LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_7_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_7_WROM;

ARCHITECTURE RTL OF L7_7_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"110100000",
  1=>"111111111",
  2=>"111010111",
  3=>"111011111",
  4=>"110111001",
  5=>"101101001",
  6=>"000000000",
  7=>"111101000",
  8=>"000000000",
  9=>"000000000",
  10=>"110000000",
  11=>"011111111",
  12=>"110110011",
  13=>"001001000",
  14=>"000000000",
  15=>"111111111",
  16=>"111111111",
  17=>"000110110",
  18=>"000000000",
  19=>"001011001",
  20=>"111000111",
  21=>"000110110",
  22=>"111111111",
  23=>"001001011",
  24=>"000000111",
  25=>"010000000",
  26=>"001001000",
  27=>"111010000",
  28=>"000000000",
  29=>"000111111",
  30=>"001001001",
  31=>"000000110",
  32=>"000000000",
  33=>"111111111",
  34=>"011111111",
  35=>"000000000",
  36=>"001111111",
  37=>"011011111",
  38=>"111111111",
  39=>"111000000",
  40=>"011111111",
  41=>"000000000",
  42=>"111111111",
  43=>"000001111",
  44=>"000000001",
  45=>"111111111",
  46=>"111111111",
  47=>"000000110",
  48=>"001001001",
  49=>"000000000",
  50=>"001001010",
  51=>"001111111",
  52=>"000011111",
  53=>"000000001",
  54=>"000111111",
  55=>"111111001",
  56=>"100110000",
  57=>"011111111",
  58=>"011111111",
  59=>"010110110",
  60=>"001000000",
  61=>"000000000",
  62=>"000000001",
  63=>"111111110",
  64=>"011111111",
  65=>"000010000",
  66=>"111111010",
  67=>"000000000",
  68=>"111110001",
  69=>"000000000",
  70=>"111000000",
  71=>"010111111",
  72=>"111100100",
  73=>"101000000",
  74=>"011111111",
  75=>"001000000",
  76=>"000100000",
  77=>"000000000",
  78=>"000000111",
  79=>"111111111",
  80=>"111111111",
  81=>"000000000",
  82=>"010010000",
  83=>"001101000",
  84=>"000000000",
  85=>"000011001",
  86=>"000000001",
  87=>"000000000",
  88=>"111111000",
  89=>"111000000",
  90=>"111101111",
  91=>"110000001",
  92=>"101111011",
  93=>"000000000",
  94=>"111111111",
  95=>"011111000",
  96=>"110010100",
  97=>"000000000",
  98=>"110110111",
  99=>"000000000",
  100=>"111011001",
  101=>"000011010",
  102=>"000000111",
  103=>"000000001",
  104=>"110110000",
  105=>"110111110",
  106=>"111111111",
  107=>"000100000",
  108=>"000000100",
  109=>"000000111",
  110=>"111111111",
  111=>"000000000",
  112=>"111111000",
  113=>"000000000",
  114=>"011011001",
  115=>"010111111",
  116=>"111000001",
  117=>"111111101",
  118=>"111110000",
  119=>"000000001",
  120=>"000111011",
  121=>"111111111",
  122=>"000000000",
  123=>"000011111",
  124=>"000011011",
  125=>"111011001",
  126=>"001011111",
  127=>"000000000",
  128=>"000110111",
  129=>"111111111",
  130=>"111111111",
  131=>"110110001",
  132=>"000000110",
  133=>"111100111",
  134=>"111110000",
  135=>"000000000",
  136=>"000000000",
  137=>"111110000",
  138=>"111000000",
  139=>"100000000",
  140=>"000000000",
  141=>"111111110",
  142=>"001000101",
  143=>"111111010",
  144=>"111111111",
  145=>"001001011",
  146=>"000000000",
  147=>"100000001",
  148=>"000100100",
  149=>"000000000",
  150=>"000000001",
  151=>"011000111",
  152=>"111111111",
  153=>"111100001",
  154=>"111000000",
  155=>"111111111",
  156=>"111101111",
  157=>"111111111",
  158=>"001011111",
  159=>"101001000",
  160=>"000000000",
  161=>"111011110",
  162=>"001001001",
  163=>"111111011",
  164=>"000000000",
  165=>"001000000",
  166=>"001001000",
  167=>"100100100",
  168=>"011111111",
  169=>"000000000",
  170=>"000000000",
  171=>"111111111",
  172=>"011111111",
  173=>"001011100",
  174=>"001000000",
  175=>"000000000",
  176=>"000100101",
  177=>"001001001",
  178=>"111111111",
  179=>"001000000",
  180=>"000000000",
  181=>"111111111",
  182=>"000000000",
  183=>"111000000",
  184=>"111111111",
  185=>"000001110",
  186=>"111110101",
  187=>"111111000",
  188=>"000000000",
  189=>"111111111",
  190=>"111100000",
  191=>"000001001",
  192=>"000011011",
  193=>"111111000",
  194=>"111111111",
  195=>"000111111",
  196=>"001111111",
  197=>"111111111",
  198=>"111111111",
  199=>"001001000",
  200=>"110100000",
  201=>"000000000",
  202=>"111111101",
  203=>"000000000",
  204=>"001011111",
  205=>"111110110",
  206=>"000000000",
  207=>"111000000",
  208=>"000000000",
  209=>"000000000",
  210=>"000000000",
  211=>"111011000",
  212=>"000111111",
  213=>"100100110",
  214=>"111111010",
  215=>"110000000",
  216=>"111111111",
  217=>"000000111",
  218=>"000000110",
  219=>"000001000",
  220=>"111111000",
  221=>"000000000",
  222=>"000000111",
  223=>"000000000",
  224=>"000000000",
  225=>"110010000",
  226=>"000000000",
  227=>"111111111",
  228=>"111111101",
  229=>"001000001",
  230=>"111111111",
  231=>"111001001",
  232=>"111010011",
  233=>"000000101",
  234=>"101101111",
  235=>"000000000",
  236=>"110000000",
  237=>"010111111",
  238=>"111110110",
  239=>"000001100",
  240=>"111111111",
  241=>"110101111",
  242=>"111111111",
  243=>"111000000",
  244=>"111000111",
  245=>"111111100",
  246=>"000001001",
  247=>"011011010",
  248=>"100000000",
  249=>"111111111",
  250=>"001001001",
  251=>"000001111",
  252=>"000111110",
  253=>"100111111",
  254=>"111111100",
  255=>"000000000",
  256=>"000000000",
  257=>"000100100",
  258=>"111111111",
  259=>"111111110",
  260=>"111100000",
  261=>"110110111",
  262=>"010000101",
  263=>"100110100",
  264=>"001001001",
  265=>"000000000",
  266=>"111001001",
  267=>"000000000",
  268=>"111101101",
  269=>"111001000",
  270=>"111000001",
  271=>"111111011",
  272=>"000000000",
  273=>"111111000",
  274=>"000000111",
  275=>"001111111",
  276=>"110111111",
  277=>"000110000",
  278=>"001000000",
  279=>"000000000",
  280=>"101011011",
  281=>"010000010",
  282=>"110111111",
  283=>"111101111",
  284=>"111111111",
  285=>"100000000",
  286=>"110111111",
  287=>"000000111",
  288=>"000000000",
  289=>"000000000",
  290=>"100110101",
  291=>"111111111",
  292=>"110000000",
  293=>"011111111",
  294=>"001001111",
  295=>"000000000",
  296=>"000001000",
  297=>"100100111",
  298=>"111101111",
  299=>"110111000",
  300=>"110100000",
  301=>"000101101",
  302=>"111101111",
  303=>"000000000",
  304=>"001001111",
  305=>"000000000",
  306=>"110111111",
  307=>"000000000",
  308=>"111100111",
  309=>"000000000",
  310=>"001001011",
  311=>"010111111",
  312=>"000000100",
  313=>"111011000",
  314=>"000000000",
  315=>"000000000",
  316=>"111111100",
  317=>"000000000",
  318=>"111101101",
  319=>"001011000",
  320=>"000000000",
  321=>"000001000",
  322=>"111111111",
  323=>"111111111",
  324=>"111111000",
  325=>"000000000",
  326=>"000111111",
  327=>"111111111",
  328=>"000000000",
  329=>"000000000",
  330=>"011001000",
  331=>"000000101",
  332=>"111111111",
  333=>"110110110",
  334=>"111001000",
  335=>"111111111",
  336=>"001011111",
  337=>"111111011",
  338=>"111111111",
  339=>"111111111",
  340=>"000000110",
  341=>"011110011",
  342=>"000000000",
  343=>"000111011",
  344=>"111111111",
  345=>"111111000",
  346=>"111111011",
  347=>"101111111",
  348=>"000000000",
  349=>"111110010",
  350=>"110111111",
  351=>"111011001",
  352=>"111111011",
  353=>"111111111",
  354=>"000110110",
  355=>"011001000",
  356=>"000111111",
  357=>"001000000",
  358=>"111011011",
  359=>"010100110",
  360=>"000111100",
  361=>"111111111",
  362=>"111111110",
  363=>"000000000",
  364=>"000000110",
  365=>"000000100",
  366=>"000000000",
  367=>"111111000",
  368=>"000000000",
  369=>"111111111",
  370=>"000000000",
  371=>"000100111",
  372=>"110000000",
  373=>"000000000",
  374=>"000000000",
  375=>"000100000",
  376=>"111111111",
  377=>"000000000",
  378=>"101001001",
  379=>"111111011",
  380=>"000000000",
  381=>"000000000",
  382=>"000000000",
  383=>"110100000",
  384=>"110110110",
  385=>"000000001",
  386=>"001001001",
  387=>"111111111",
  388=>"011111111",
  389=>"000110110",
  390=>"000000100",
  391=>"000001001",
  392=>"111111111",
  393=>"000000000",
  394=>"000001001",
  395=>"111111111",
  396=>"000000010",
  397=>"000111111",
  398=>"001001111",
  399=>"000000000",
  400=>"000000000",
  401=>"000000000",
  402=>"111111111",
  403=>"110100000",
  404=>"000000000",
  405=>"000000100",
  406=>"011011001",
  407=>"000000000",
  408=>"111111000",
  409=>"111000000",
  410=>"111111111",
  411=>"010000000",
  412=>"000000000",
  413=>"111110111",
  414=>"111111111",
  415=>"000000000",
  416=>"001001001",
  417=>"001111111",
  418=>"000000010",
  419=>"111111010",
  420=>"111000000",
  421=>"100000001",
  422=>"000100111",
  423=>"111111111",
  424=>"010010000",
  425=>"000011000",
  426=>"011011011",
  427=>"101000110",
  428=>"000000000",
  429=>"011001001",
  430=>"111010000",
  431=>"000011111",
  432=>"001000100",
  433=>"111111110",
  434=>"000000110",
  435=>"011011111",
  436=>"110111000",
  437=>"111111111",
  438=>"000000000",
  439=>"000000000",
  440=>"111111111",
  441=>"000001011",
  442=>"110100000",
  443=>"111100000",
  444=>"000000010",
  445=>"001001001",
  446=>"110000000",
  447=>"101001001",
  448=>"000000000",
  449=>"111111111",
  450=>"111111011",
  451=>"000000100",
  452=>"001001001",
  453=>"001001001",
  454=>"000000000",
  455=>"000000000",
  456=>"111111111",
  457=>"000000000",
  458=>"011000000",
  459=>"111000000",
  460=>"000000000",
  461=>"001011000",
  462=>"101000001",
  463=>"111011000",
  464=>"000000001",
  465=>"000000000",
  466=>"111111111",
  467=>"011000000",
  468=>"000000000",
  469=>"101101111",
  470=>"010011000",
  471=>"110110111",
  472=>"111111111",
  473=>"001000000",
  474=>"111011000",
  475=>"000000000",
  476=>"111110100",
  477=>"111001000",
  478=>"000001011",
  479=>"011101101",
  480=>"111111110",
  481=>"111001000",
  482=>"000000000",
  483=>"000000000",
  484=>"011111011",
  485=>"000000000",
  486=>"110110111",
  487=>"000000000",
  488=>"010111111",
  489=>"111111111",
  490=>"011101101",
  491=>"111111111",
  492=>"110111110",
  493=>"000000000",
  494=>"000000000",
  495=>"111111111",
  496=>"100100001",
  497=>"000000100",
  498=>"001001000",
  499=>"111111111",
  500=>"111111001",
  501=>"000000000",
  502=>"000000100",
  503=>"100100110",
  504=>"000000110",
  505=>"111101001",
  506=>"000111111",
  507=>"001001000",
  508=>"000000111",
  509=>"011000100",
  510=>"000000000",
  511=>"000000111",
  512=>"000000000",
  513=>"110000000",
  514=>"111111111",
  515=>"000001111",
  516=>"111111100",
  517=>"000101111",
  518=>"111010000",
  519=>"000000111",
  520=>"111111111",
  521=>"000010011",
  522=>"100101000",
  523=>"000010011",
  524=>"111111000",
  525=>"100001000",
  526=>"111001000",
  527=>"110000000",
  528=>"100111111",
  529=>"111111000",
  530=>"000111100",
  531=>"111111111",
  532=>"000110100",
  533=>"000100111",
  534=>"111000000",
  535=>"000000100",
  536=>"100100111",
  537=>"000100001",
  538=>"000000101",
  539=>"111111110",
  540=>"000000000",
  541=>"101000100",
  542=>"111011001",
  543=>"111111111",
  544=>"000001000",
  545=>"000111111",
  546=>"110110111",
  547=>"100000000",
  548=>"001000000",
  549=>"000000000",
  550=>"000111111",
  551=>"000000011",
  552=>"111111000",
  553=>"000000000",
  554=>"011111111",
  555=>"001100100",
  556=>"111111111",
  557=>"111111010",
  558=>"100100111",
  559=>"000000000",
  560=>"111111101",
  561=>"111011011",
  562=>"100000000",
  563=>"111000000",
  564=>"011001110",
  565=>"010010110",
  566=>"001000111",
  567=>"010110110",
  568=>"111000000",
  569=>"101101000",
  570=>"000000010",
  571=>"000000011",
  572=>"101000000",
  573=>"001001001",
  574=>"110010000",
  575=>"000111111",
  576=>"000000111",
  577=>"001001011",
  578=>"111111000",
  579=>"000000000",
  580=>"000000000",
  581=>"000011111",
  582=>"110000000",
  583=>"000001000",
  584=>"000000001",
  585=>"001001000",
  586=>"000000011",
  587=>"111111010",
  588=>"110000001",
  589=>"111101111",
  590=>"001001001",
  591=>"111110110",
  592=>"000000000",
  593=>"000000000",
  594=>"000000101",
  595=>"111110110",
  596=>"111111001",
  597=>"000000000",
  598=>"110110000",
  599=>"111111111",
  600=>"000000000",
  601=>"101000000",
  602=>"110110100",
  603=>"100111111",
  604=>"111001001",
  605=>"000000000",
  606=>"000110111",
  607=>"000010000",
  608=>"101000000",
  609=>"101111001",
  610=>"111111111",
  611=>"000101000",
  612=>"110010000",
  613=>"000001011",
  614=>"001111111",
  615=>"001101101",
  616=>"000000000",
  617=>"111000000",
  618=>"110111111",
  619=>"000000000",
  620=>"010000000",
  621=>"111000010",
  622=>"100001111",
  623=>"011111110",
  624=>"111111111",
  625=>"101111111",
  626=>"001001001",
  627=>"111101000",
  628=>"111000000",
  629=>"110000000",
  630=>"111100100",
  631=>"111111001",
  632=>"000001111",
  633=>"000111101",
  634=>"100100100",
  635=>"001001001",
  636=>"100110110",
  637=>"111100000",
  638=>"000001111",
  639=>"001000000",
  640=>"111101101",
  641=>"000000000",
  642=>"110110000",
  643=>"111011010",
  644=>"111111111",
  645=>"000100101",
  646=>"000110000",
  647=>"000100000",
  648=>"000000001",
  649=>"000000000",
  650=>"011011000",
  651=>"011000000",
  652=>"111010010",
  653=>"100000001",
  654=>"110001000",
  655=>"111101000",
  656=>"111111111",
  657=>"111001001",
  658=>"110110100",
  659=>"001000001",
  660=>"001001000",
  661=>"111000000",
  662=>"000011111",
  663=>"000000000",
  664=>"100100000",
  665=>"000000000",
  666=>"111101100",
  667=>"001001000",
  668=>"101110111",
  669=>"000000111",
  670=>"000000100",
  671=>"111111111",
  672=>"111111111",
  673=>"111110110",
  674=>"111110000",
  675=>"000111111",
  676=>"010000100",
  677=>"111011001",
  678=>"111111001",
  679=>"101101100",
  680=>"110000000",
  681=>"100101000",
  682=>"011111000",
  683=>"000000000",
  684=>"110110111",
  685=>"111000000",
  686=>"101001111",
  687=>"000000000",
  688=>"000000111",
  689=>"000111111",
  690=>"010011011",
  691=>"000000111",
  692=>"110111111",
  693=>"111000000",
  694=>"000110111",
  695=>"000100110",
  696=>"111101100",
  697=>"111011011",
  698=>"111000000",
  699=>"110111111",
  700=>"000000000",
  701=>"000000000",
  702=>"000111111",
  703=>"111000110",
  704=>"000111111",
  705=>"001000000",
  706=>"111111111",
  707=>"111111111",
  708=>"111111111",
  709=>"000000000",
  710=>"001000000",
  711=>"001111111",
  712=>"000000010",
  713=>"000000010",
  714=>"000000000",
  715=>"011011011",
  716=>"111111000",
  717=>"100110100",
  718=>"111000100",
  719=>"111000000",
  720=>"000000101",
  721=>"000001000",
  722=>"110000000",
  723=>"000111100",
  724=>"111010101",
  725=>"111111000",
  726=>"010000000",
  727=>"111011001",
  728=>"000000000",
  729=>"000000000",
  730=>"111110111",
  731=>"000000000",
  732=>"000000000",
  733=>"000110010",
  734=>"111111000",
  735=>"111001101",
  736=>"000000000",
  737=>"000000000",
  738=>"111111011",
  739=>"111111111",
  740=>"000100000",
  741=>"000111111",
  742=>"011111111",
  743=>"000000000",
  744=>"011000000",
  745=>"100000111",
  746=>"111101101",
  747=>"000100100",
  748=>"111111111",
  749=>"111011011",
  750=>"000000000",
  751=>"000000000",
  752=>"111111001",
  753=>"011000000",
  754=>"001111111",
  755=>"001001111",
  756=>"011000000",
  757=>"001000000",
  758=>"100110100",
  759=>"000000000",
  760=>"000000000",
  761=>"111111111",
  762=>"111111100",
  763=>"111111111",
  764=>"000000100",
  765=>"000000100",
  766=>"110110111",
  767=>"111100000",
  768=>"000100000",
  769=>"000000011",
  770=>"001000000",
  771=>"110110111",
  772=>"000000100",
  773=>"111001111",
  774=>"000100000",
  775=>"001011000",
  776=>"111110110",
  777=>"000000000",
  778=>"010111111",
  779=>"111111111",
  780=>"011000011",
  781=>"110110111",
  782=>"000000000",
  783=>"000000000",
  784=>"011000000",
  785=>"000000100",
  786=>"000000111",
  787=>"000000000",
  788=>"110100110",
  789=>"000000000",
  790=>"110111100",
  791=>"001101101",
  792=>"111110111",
  793=>"000000000",
  794=>"110111111",
  795=>"010000000",
  796=>"000000110",
  797=>"000000000",
  798=>"111000000",
  799=>"111001011",
  800=>"110111101",
  801=>"000111111",
  802=>"000000100",
  803=>"011111111",
  804=>"110111111",
  805=>"000000000",
  806=>"111000000",
  807=>"000001111",
  808=>"111111111",
  809=>"111000011",
  810=>"111111111",
  811=>"101100111",
  812=>"001011111",
  813=>"010110111",
  814=>"000000001",
  815=>"000000001",
  816=>"011011011",
  817=>"111100000",
  818=>"001001000",
  819=>"111111000",
  820=>"101111111",
  821=>"111111101",
  822=>"100111111",
  823=>"000000010",
  824=>"000000000",
  825=>"101000000",
  826=>"111000000",
  827=>"111001001",
  828=>"100000000",
  829=>"111001011",
  830=>"000000000",
  831=>"110100100",
  832=>"111111101",
  833=>"110111111",
  834=>"000000000",
  835=>"010010110",
  836=>"000000000",
  837=>"000000000",
  838=>"000000000",
  839=>"001000000",
  840=>"111001000",
  841=>"000000000",
  842=>"111001111",
  843=>"110110111",
  844=>"000000000",
  845=>"001000000",
  846=>"001001000",
  847=>"000110110",
  848=>"000110110",
  849=>"111110100",
  850=>"000000010",
  851=>"000101001",
  852=>"011011000",
  853=>"001011011",
  854=>"111111010",
  855=>"000011111",
  856=>"000111111",
  857=>"000000000",
  858=>"000000100",
  859=>"111000000",
  860=>"111111111",
  861=>"111011001",
  862=>"000000000",
  863=>"100000011",
  864=>"000000000",
  865=>"000000000",
  866=>"010010000",
  867=>"101000000",
  868=>"110111111",
  869=>"000000000",
  870=>"000000000",
  871=>"000110110",
  872=>"110111111",
  873=>"000000100",
  874=>"001111111",
  875=>"000000101",
  876=>"111110000",
  877=>"001001011",
  878=>"000110000",
  879=>"111000000",
  880=>"111111011",
  881=>"111001011",
  882=>"111111111",
  883=>"001000000",
  884=>"001011011",
  885=>"101100110",
  886=>"001001101",
  887=>"000001011",
  888=>"001101111",
  889=>"000111000",
  890=>"000000001",
  891=>"111011111",
  892=>"011000001",
  893=>"100100100",
  894=>"000111000",
  895=>"110111111",
  896=>"000111001",
  897=>"000001000",
  898=>"110110111",
  899=>"000001111",
  900=>"110111111",
  901=>"111111110",
  902=>"000100111",
  903=>"111111111",
  904=>"110000000",
  905=>"011001000",
  906=>"011001001",
  907=>"111111111",
  908=>"000111111",
  909=>"000000000",
  910=>"000000000",
  911=>"011111110",
  912=>"000000001",
  913=>"110000001",
  914=>"110111111",
  915=>"001000000",
  916=>"000100001",
  917=>"110100110",
  918=>"100110000",
  919=>"110110110",
  920=>"000001111",
  921=>"000000111",
  922=>"000000000",
  923=>"111111111",
  924=>"010010101",
  925=>"111011000",
  926=>"111111111",
  927=>"111111111",
  928=>"111000000",
  929=>"000000001",
  930=>"110100111",
  931=>"110111111",
  932=>"100111011",
  933=>"111110110",
  934=>"001000000",
  935=>"111111111",
  936=>"111111111",
  937=>"000001000",
  938=>"000000001",
  939=>"111000000",
  940=>"000101111",
  941=>"000100000",
  942=>"000000101",
  943=>"001000000",
  944=>"100000000",
  945=>"100000000",
  946=>"001001000",
  947=>"111111000",
  948=>"000111111",
  949=>"011000011",
  950=>"000000011",
  951=>"000000001",
  952=>"100111111",
  953=>"111111000",
  954=>"110000001",
  955=>"000111000",
  956=>"000010111",
  957=>"001000110",
  958=>"000000000",
  959=>"110111110",
  960=>"111111111",
  961=>"000000000",
  962=>"000000000",
  963=>"100100000",
  964=>"111111111",
  965=>"000000000",
  966=>"101111111",
  967=>"001000000",
  968=>"000000000",
  969=>"001000000",
  970=>"010001011",
  971=>"010000111",
  972=>"000000000",
  973=>"000000000",
  974=>"000000111",
  975=>"000000111",
  976=>"000011111",
  977=>"011111110",
  978=>"000000000",
  979=>"000000001",
  980=>"100001001",
  981=>"111000110",
  982=>"000000000",
  983=>"000010010",
  984=>"000000000",
  985=>"000011111",
  986=>"001000000",
  987=>"111111001",
  988=>"011111111",
  989=>"100000000",
  990=>"111000000",
  991=>"111101101",
  992=>"111101000",
  993=>"111000000",
  994=>"111100000",
  995=>"110000000",
  996=>"111111111",
  997=>"100100100",
  998=>"111111111",
  999=>"111111000",
  1000=>"111000001",
  1001=>"100101100",
  1002=>"011011111",
  1003=>"001000000",
  1004=>"000111111",
  1005=>"111001000",
  1006=>"111111111",
  1007=>"111000101",
  1008=>"111011011",
  1009=>"000100110",
  1010=>"111001000",
  1011=>"010011011",
  1012=>"000000100",
  1013=>"111111011",
  1014=>"000000000",
  1015=>"000000100",
  1016=>"000000000",
  1017=>"000110100",
  1018=>"111111001",
  1019=>"000000000",
  1020=>"000110000",
  1021=>"000110111",
  1022=>"111111111",
  1023=>"000000000",
  1024=>"111100100",
  1025=>"000000000",
  1026=>"111110000",
  1027=>"111110100",
  1028=>"111000000",
  1029=>"001000000",
  1030=>"000000111",
  1031=>"000000111",
  1032=>"111100100",
  1033=>"000001101",
  1034=>"000000110",
  1035=>"000110111",
  1036=>"110111111",
  1037=>"111111111",
  1038=>"000111111",
  1039=>"111111101",
  1040=>"000000001",
  1041=>"111011111",
  1042=>"010001000",
  1043=>"111111111",
  1044=>"000000111",
  1045=>"000000000",
  1046=>"111111000",
  1047=>"000000000",
  1048=>"111111101",
  1049=>"111111100",
  1050=>"111000110",
  1051=>"000000001",
  1052=>"000000011",
  1053=>"101111111",
  1054=>"110110100",
  1055=>"111010001",
  1056=>"111111111",
  1057=>"001001001",
  1058=>"110111000",
  1059=>"000010000",
  1060=>"110111111",
  1061=>"111111111",
  1062=>"000000000",
  1063=>"000000111",
  1064=>"001000111",
  1065=>"110111111",
  1066=>"000000111",
  1067=>"000011111",
  1068=>"011001000",
  1069=>"111111110",
  1070=>"110000001",
  1071=>"011001101",
  1072=>"111000000",
  1073=>"010000000",
  1074=>"001000110",
  1075=>"111111000",
  1076=>"001111111",
  1077=>"110100000",
  1078=>"110000000",
  1079=>"000000000",
  1080=>"111111010",
  1081=>"000000001",
  1082=>"000010111",
  1083=>"011000001",
  1084=>"111000011",
  1085=>"111111111",
  1086=>"100111000",
  1087=>"111111110",
  1088=>"011011000",
  1089=>"001001001",
  1090=>"001111111",
  1091=>"111000000",
  1092=>"100000000",
  1093=>"011101100",
  1094=>"111111111",
  1095=>"000000101",
  1096=>"011111000",
  1097=>"000000000",
  1098=>"110100111",
  1099=>"000111111",
  1100=>"110000000",
  1101=>"001011001",
  1102=>"011111111",
  1103=>"000000110",
  1104=>"000000000",
  1105=>"011011111",
  1106=>"111111001",
  1107=>"110001001",
  1108=>"000010000",
  1109=>"010000000",
  1110=>"000000011",
  1111=>"111111111",
  1112=>"111111110",
  1113=>"000000111",
  1114=>"000000111",
  1115=>"111001001",
  1116=>"111110000",
  1117=>"111111111",
  1118=>"111111111",
  1119=>"111101001",
  1120=>"001111111",
  1121=>"010000000",
  1122=>"000111111",
  1123=>"001111111",
  1124=>"101000000",
  1125=>"000000010",
  1126=>"000011111",
  1127=>"001000000",
  1128=>"111111111",
  1129=>"001000000",
  1130=>"000000000",
  1131=>"111111000",
  1132=>"000000000",
  1133=>"000000110",
  1134=>"000000000",
  1135=>"111001001",
  1136=>"000000100",
  1137=>"111011001",
  1138=>"100110111",
  1139=>"000011011",
  1140=>"000100111",
  1141=>"000000000",
  1142=>"000000000",
  1143=>"011111111",
  1144=>"000000100",
  1145=>"111111001",
  1146=>"000000000",
  1147=>"100000101",
  1148=>"111010000",
  1149=>"000001000",
  1150=>"111111110",
  1151=>"000000000",
  1152=>"101001000",
  1153=>"011000000",
  1154=>"110111111",
  1155=>"110000000",
  1156=>"000000000",
  1157=>"100111011",
  1158=>"111000001",
  1159=>"001000000",
  1160=>"011000001",
  1161=>"000011001",
  1162=>"001001101",
  1163=>"000000111",
  1164=>"000000000",
  1165=>"011111011",
  1166=>"100100110",
  1167=>"000000000",
  1168=>"000000111",
  1169=>"101000000",
  1170=>"001001000",
  1171=>"110000000",
  1172=>"000000101",
  1173=>"110111011",
  1174=>"000000001",
  1175=>"110100000",
  1176=>"001001101",
  1177=>"000010010",
  1178=>"111111111",
  1179=>"010000000",
  1180=>"111111010",
  1181=>"000000100",
  1182=>"110110111",
  1183=>"001000000",
  1184=>"000000000",
  1185=>"010000000",
  1186=>"111111100",
  1187=>"111001011",
  1188=>"101011000",
  1189=>"111111110",
  1190=>"001000000",
  1191=>"100000000",
  1192=>"111111111",
  1193=>"111000101",
  1194=>"111111000",
  1195=>"000000000",
  1196=>"011111111",
  1197=>"111110000",
  1198=>"111110110",
  1199=>"011000000",
  1200=>"111001111",
  1201=>"001001111",
  1202=>"111111110",
  1203=>"000000000",
  1204=>"000000000",
  1205=>"010110111",
  1206=>"011111110",
  1207=>"000000010",
  1208=>"111110010",
  1209=>"000000000",
  1210=>"101110000",
  1211=>"001001000",
  1212=>"000000010",
  1213=>"000000111",
  1214=>"100000100",
  1215=>"000101000",
  1216=>"111011001",
  1217=>"111111111",
  1218=>"000000111",
  1219=>"110100000",
  1220=>"011001000",
  1221=>"000000000",
  1222=>"110110111",
  1223=>"001001000",
  1224=>"111000111",
  1225=>"111110000",
  1226=>"000001101",
  1227=>"000000011",
  1228=>"111110000",
  1229=>"010111111",
  1230=>"000001000",
  1231=>"000000011",
  1232=>"111000000",
  1233=>"000000000",
  1234=>"111011001",
  1235=>"000000000",
  1236=>"110110000",
  1237=>"100011111",
  1238=>"111001111",
  1239=>"000000000",
  1240=>"110010000",
  1241=>"000000001",
  1242=>"000111111",
  1243=>"111011000",
  1244=>"000000011",
  1245=>"000000111",
  1246=>"000001000",
  1247=>"110000111",
  1248=>"000000000",
  1249=>"000111111",
  1250=>"111111111",
  1251=>"111111111",
  1252=>"000110010",
  1253=>"111001000",
  1254=>"000111011",
  1255=>"111111111",
  1256=>"111111011",
  1257=>"111101000",
  1258=>"101111111",
  1259=>"000110010",
  1260=>"111111111",
  1261=>"111100100",
  1262=>"110110111",
  1263=>"000000001",
  1264=>"000111110",
  1265=>"100000000",
  1266=>"011111110",
  1267=>"000100100",
  1268=>"111111010",
  1269=>"001001100",
  1270=>"111111000",
  1271=>"111011000",
  1272=>"000001111",
  1273=>"000011000",
  1274=>"110110000",
  1275=>"011011110",
  1276=>"011000111",
  1277=>"001011111",
  1278=>"111010000",
  1279=>"000111111",
  1280=>"000000000",
  1281=>"111111110",
  1282=>"111111111",
  1283=>"000000011",
  1284=>"000000111",
  1285=>"111111111",
  1286=>"111111100",
  1287=>"111111111",
  1288=>"000000000",
  1289=>"011010101",
  1290=>"111111111",
  1291=>"000111111",
  1292=>"100100110",
  1293=>"111111011",
  1294=>"111111011",
  1295=>"111001000",
  1296=>"110111111",
  1297=>"110110000",
  1298=>"000000110",
  1299=>"000000000",
  1300=>"000000000",
  1301=>"111000011",
  1302=>"111111111",
  1303=>"100000001",
  1304=>"111101000",
  1305=>"100110000",
  1306=>"110111000",
  1307=>"000011111",
  1308=>"000000111",
  1309=>"000000000",
  1310=>"000000000",
  1311=>"111111111",
  1312=>"111111000",
  1313=>"000000000",
  1314=>"000000001",
  1315=>"000000111",
  1316=>"111111111",
  1317=>"000000111",
  1318=>"000110110",
  1319=>"100000000",
  1320=>"000000001",
  1321=>"000000000",
  1322=>"111110000",
  1323=>"000010111",
  1324=>"111111001",
  1325=>"000000000",
  1326=>"111110111",
  1327=>"000000001",
  1328=>"101001000",
  1329=>"000001011",
  1330=>"110110101",
  1331=>"000000000",
  1332=>"000110010",
  1333=>"111111000",
  1334=>"110110111",
  1335=>"010000000",
  1336=>"000000000",
  1337=>"100000000",
  1338=>"111101001",
  1339=>"000000111",
  1340=>"000111111",
  1341=>"111000000",
  1342=>"000000000",
  1343=>"111011001",
  1344=>"000000111",
  1345=>"111111111",
  1346=>"111111111",
  1347=>"000000000",
  1348=>"000001001",
  1349=>"110001111",
  1350=>"000000000",
  1351=>"000001000",
  1352=>"111111111",
  1353=>"000000000",
  1354=>"000000000",
  1355=>"110100000",
  1356=>"000000000",
  1357=>"000000000",
  1358=>"111111000",
  1359=>"110110110",
  1360=>"110000100",
  1361=>"001000000",
  1362=>"111111011",
  1363=>"000010000",
  1364=>"110000010",
  1365=>"011011001",
  1366=>"111111111",
  1367=>"111110000",
  1368=>"111110000",
  1369=>"000000000",
  1370=>"011011001",
  1371=>"000000000",
  1372=>"111111001",
  1373=>"001001000",
  1374=>"000000001",
  1375=>"110111111",
  1376=>"011111101",
  1377=>"111000000",
  1378=>"111011001",
  1379=>"111101111",
  1380=>"000111111",
  1381=>"111111011",
  1382=>"000000000",
  1383=>"000011111",
  1384=>"111101000",
  1385=>"001101111",
  1386=>"000001001",
  1387=>"100001000",
  1388=>"110110110",
  1389=>"000111110",
  1390=>"000011111",
  1391=>"100000111",
  1392=>"011111111",
  1393=>"011000000",
  1394=>"000000000",
  1395=>"011001000",
  1396=>"111010000",
  1397=>"111111111",
  1398=>"000000101",
  1399=>"000001111",
  1400=>"111001001",
  1401=>"101000111",
  1402=>"111111111",
  1403=>"111111111",
  1404=>"111000000",
  1405=>"000100100",
  1406=>"100000000",
  1407=>"000000111",
  1408=>"010110010",
  1409=>"110110110",
  1410=>"111111011",
  1411=>"001001000",
  1412=>"111111111",
  1413=>"111111110",
  1414=>"110111000",
  1415=>"000000101",
  1416=>"000000000",
  1417=>"000010111",
  1418=>"111111111",
  1419=>"000111111",
  1420=>"111011111",
  1421=>"000110010",
  1422=>"000111111",
  1423=>"001011011",
  1424=>"111000000",
  1425=>"110000000",
  1426=>"000101101",
  1427=>"001100110",
  1428=>"000000000",
  1429=>"010011111",
  1430=>"111111011",
  1431=>"101100000",
  1432=>"001101111",
  1433=>"111011111",
  1434=>"000000111",
  1435=>"111110000",
  1436=>"111111000",
  1437=>"111111111",
  1438=>"000000010",
  1439=>"111000000",
  1440=>"000000000",
  1441=>"110000000",
  1442=>"001000000",
  1443=>"000000100",
  1444=>"000100100",
  1445=>"111001011",
  1446=>"000000100",
  1447=>"111110000",
  1448=>"111000000",
  1449=>"000100001",
  1450=>"000000000",
  1451=>"000000000",
  1452=>"000000000",
  1453=>"000000000",
  1454=>"000000001",
  1455=>"111000001",
  1456=>"000011011",
  1457=>"111111111",
  1458=>"111111000",
  1459=>"000000000",
  1460=>"101001000",
  1461=>"000000000",
  1462=>"000000000",
  1463=>"000000000",
  1464=>"111111000",
  1465=>"000000000",
  1466=>"100000001",
  1467=>"000000000",
  1468=>"000111111",
  1469=>"000011011",
  1470=>"111110100",
  1471=>"011011001",
  1472=>"111101000",
  1473=>"011110110",
  1474=>"011011111",
  1475=>"000011111",
  1476=>"111111111",
  1477=>"000000110",
  1478=>"110110111",
  1479=>"001000011",
  1480=>"110111111",
  1481=>"000000000",
  1482=>"000000101",
  1483=>"000110000",
  1484=>"000000100",
  1485=>"000010000",
  1486=>"000000001",
  1487=>"111111000",
  1488=>"111100111",
  1489=>"000000000",
  1490=>"111111001",
  1491=>"000000111",
  1492=>"001001001",
  1493=>"000000011",
  1494=>"001001010",
  1495=>"011111100",
  1496=>"111111000",
  1497=>"111011010",
  1498=>"001000011",
  1499=>"111111001",
  1500=>"111110111",
  1501=>"011000110",
  1502=>"100100000",
  1503=>"000110111",
  1504=>"001000111",
  1505=>"000000000",
  1506=>"001001111",
  1507=>"001001111",
  1508=>"000000000",
  1509=>"000010111",
  1510=>"100100101",
  1511=>"100001001",
  1512=>"000000111",
  1513=>"110011001",
  1514=>"000000000",
  1515=>"000111011",
  1516=>"111111111",
  1517=>"000001000",
  1518=>"000000111",
  1519=>"111111111",
  1520=>"101000000",
  1521=>"111111110",
  1522=>"010110111",
  1523=>"010010010",
  1524=>"111111110",
  1525=>"010110100",
  1526=>"111000000",
  1527=>"111110100",
  1528=>"111111000",
  1529=>"100000100",
  1530=>"110000000",
  1531=>"000000000",
  1532=>"110000011",
  1533=>"000100000",
  1534=>"000110111",
  1535=>"111111111",
  1536=>"100100000",
  1537=>"000000000",
  1538=>"000000100",
  1539=>"000000000",
  1540=>"101101100",
  1541=>"011100000",
  1542=>"111111000",
  1543=>"100100000",
  1544=>"000111111",
  1545=>"000000000",
  1546=>"111111111",
  1547=>"111111111",
  1548=>"111000100",
  1549=>"000000000",
  1550=>"111111000",
  1551=>"111000100",
  1552=>"111111001",
  1553=>"000000000",
  1554=>"000000111",
  1555=>"000000001",
  1556=>"111111111",
  1557=>"111111111",
  1558=>"111111001",
  1559=>"110100100",
  1560=>"100000111",
  1561=>"100000000",
  1562=>"111110110",
  1563=>"010000001",
  1564=>"000111111",
  1565=>"111111001",
  1566=>"110111001",
  1567=>"000001001",
  1568=>"111111000",
  1569=>"000000000",
  1570=>"000000000",
  1571=>"000000000",
  1572=>"111111101",
  1573=>"111111000",
  1574=>"000000000",
  1575=>"111111111",
  1576=>"000000000",
  1577=>"110000110",
  1578=>"000000000",
  1579=>"100111101",
  1580=>"000000001",
  1581=>"100110000",
  1582=>"000000111",
  1583=>"111011000",
  1584=>"011000000",
  1585=>"111000000",
  1586=>"011111110",
  1587=>"111111111",
  1588=>"111010000",
  1589=>"000001000",
  1590=>"111100000",
  1591=>"000000000",
  1592=>"011111001",
  1593=>"111111111",
  1594=>"111000000",
  1595=>"000000000",
  1596=>"101101111",
  1597=>"100000000",
  1598=>"111111000",
  1599=>"000000000",
  1600=>"110110111",
  1601=>"010000000",
  1602=>"110110111",
  1603=>"000010110",
  1604=>"111111101",
  1605=>"111111011",
  1606=>"000000101",
  1607=>"000000000",
  1608=>"110110111",
  1609=>"101001101",
  1610=>"111110000",
  1611=>"000100100",
  1612=>"000110111",
  1613=>"100101100",
  1614=>"000000110",
  1615=>"111111000",
  1616=>"101101000",
  1617=>"000001111",
  1618=>"111110111",
  1619=>"110111000",
  1620=>"111001000",
  1621=>"000000111",
  1622=>"110110000",
  1623=>"000101111",
  1624=>"000000000",
  1625=>"101000111",
  1626=>"100111000",
  1627=>"000000000",
  1628=>"111100000",
  1629=>"100111111",
  1630=>"000000011",
  1631=>"011011000",
  1632=>"000000000",
  1633=>"111000000",
  1634=>"100011000",
  1635=>"000000000",
  1636=>"111111111",
  1637=>"111101101",
  1638=>"000000000",
  1639=>"111111000",
  1640=>"000111111",
  1641=>"000000001",
  1642=>"000000100",
  1643=>"100111110",
  1644=>"111100000",
  1645=>"001000000",
  1646=>"000000000",
  1647=>"111111000",
  1648=>"000000000",
  1649=>"000000000",
  1650=>"111000000",
  1651=>"000000111",
  1652=>"000000000",
  1653=>"100111111",
  1654=>"111110111",
  1655=>"111000000",
  1656=>"111110111",
  1657=>"000111111",
  1658=>"111111111",
  1659=>"000000000",
  1660=>"110110111",
  1661=>"111101000",
  1662=>"111011000",
  1663=>"110111111",
  1664=>"000001111",
  1665=>"000000000",
  1666=>"110000000",
  1667=>"011000000",
  1668=>"001000011",
  1669=>"000000001",
  1670=>"111110000",
  1671=>"100100111",
  1672=>"000000000",
  1673=>"111111111",
  1674=>"000000001",
  1675=>"000111010",
  1676=>"000000000",
  1677=>"000000001",
  1678=>"000010111",
  1679=>"111000000",
  1680=>"000101111",
  1681=>"000000000",
  1682=>"000000000",
  1683=>"000010000",
  1684=>"000000110",
  1685=>"000000110",
  1686=>"000100111",
  1687=>"000000100",
  1688=>"000000110",
  1689=>"100000011",
  1690=>"000001000",
  1691=>"000000000",
  1692=>"111111110",
  1693=>"000000100",
  1694=>"011111000",
  1695=>"000000100",
  1696=>"000010111",
  1697=>"000010000",
  1698=>"000000000",
  1699=>"110100000",
  1700=>"100001110",
  1701=>"000011011",
  1702=>"001101111",
  1703=>"000100000",
  1704=>"000000000",
  1705=>"000000111",
  1706=>"000010000",
  1707=>"111001000",
  1708=>"100111111",
  1709=>"000000001",
  1710=>"000000000",
  1711=>"111000111",
  1712=>"111111000",
  1713=>"001000000",
  1714=>"111111111",
  1715=>"010111111",
  1716=>"111101100",
  1717=>"001001111",
  1718=>"111111111",
  1719=>"000000010",
  1720=>"000000000",
  1721=>"111100111",
  1722=>"100101001",
  1723=>"111001011",
  1724=>"100000101",
  1725=>"110111100",
  1726=>"000000000",
  1727=>"111100100",
  1728=>"000000111",
  1729=>"100111111",
  1730=>"111100101",
  1731=>"110111111",
  1732=>"111111111",
  1733=>"000101111",
  1734=>"000000000",
  1735=>"111111011",
  1736=>"111111111",
  1737=>"000001111",
  1738=>"111110100",
  1739=>"000010111",
  1740=>"001010110",
  1741=>"110001000",
  1742=>"110000000",
  1743=>"000001000",
  1744=>"110000000",
  1745=>"000000011",
  1746=>"111000000",
  1747=>"111011001",
  1748=>"111111111",
  1749=>"000000000",
  1750=>"000000000",
  1751=>"010000000",
  1752=>"000000011",
  1753=>"000000010",
  1754=>"111111111",
  1755=>"011001100",
  1756=>"111111111",
  1757=>"111111111",
  1758=>"011111000",
  1759=>"111111111",
  1760=>"000000111",
  1761=>"000000000",
  1762=>"110011010",
  1763=>"110111000",
  1764=>"111111111",
  1765=>"010010000",
  1766=>"110000000",
  1767=>"011000110",
  1768=>"000000001",
  1769=>"110111001",
  1770=>"111011000",
  1771=>"000000100",
  1772=>"111111111",
  1773=>"100000000",
  1774=>"000010010",
  1775=>"111001111",
  1776=>"000000111",
  1777=>"000000011",
  1778=>"000000000",
  1779=>"111111100",
  1780=>"000000000",
  1781=>"000010000",
  1782=>"111001111",
  1783=>"100111111",
  1784=>"100101101",
  1785=>"000000111",
  1786=>"000111111",
  1787=>"111111000",
  1788=>"000000000",
  1789=>"000001011",
  1790=>"000000000",
  1791=>"000000000",
  1792=>"100000000",
  1793=>"111111011",
  1794=>"000000111",
  1795=>"000000101",
  1796=>"100011011",
  1797=>"000000010",
  1798=>"000000000",
  1799=>"000000000",
  1800=>"100111000",
  1801=>"000101111",
  1802=>"011001000",
  1803=>"011011001",
  1804=>"000000100",
  1805=>"000010111",
  1806=>"011010010",
  1807=>"100100111",
  1808=>"111101001",
  1809=>"111111111",
  1810=>"111111111",
  1811=>"100101111",
  1812=>"111111110",
  1813=>"000000100",
  1814=>"000010000",
  1815=>"000001001",
  1816=>"000111111",
  1817=>"000101111",
  1818=>"111111111",
  1819=>"100000011",
  1820=>"110111111",
  1821=>"110110110",
  1822=>"000110110",
  1823=>"000000111",
  1824=>"011011011",
  1825=>"111111111",
  1826=>"000110000",
  1827=>"001011000",
  1828=>"111011011",
  1829=>"000000000",
  1830=>"011001011",
  1831=>"111110000",
  1832=>"101001111",
  1833=>"111111000",
  1834=>"000000010",
  1835=>"111111111",
  1836=>"000000111",
  1837=>"001001011",
  1838=>"111000111",
  1839=>"110000000",
  1840=>"000111110",
  1841=>"110111001",
  1842=>"000000000",
  1843=>"010000011",
  1844=>"111111000",
  1845=>"011111111",
  1846=>"000010011",
  1847=>"000000110",
  1848=>"000000000",
  1849=>"000110111",
  1850=>"001111111",
  1851=>"111000000",
  1852=>"001000000",
  1853=>"111111000",
  1854=>"000000100",
  1855=>"010011111",
  1856=>"010111111",
  1857=>"001011111",
  1858=>"101001101",
  1859=>"000000111",
  1860=>"000110000",
  1861=>"001000110",
  1862=>"000000100",
  1863=>"000111001",
  1864=>"100111111",
  1865=>"000000001",
  1866=>"000000111",
  1867=>"110111011",
  1868=>"000000001",
  1869=>"001011111",
  1870=>"000001001",
  1871=>"100111111",
  1872=>"011111110",
  1873=>"000000100",
  1874=>"111001000",
  1875=>"000000000",
  1876=>"111111111",
  1877=>"001001001",
  1878=>"000111111",
  1879=>"111111111",
  1880=>"000000011",
  1881=>"001001111",
  1882=>"000001111",
  1883=>"111000000",
  1884=>"111000010",
  1885=>"111111111",
  1886=>"110111111",
  1887=>"000000100",
  1888=>"000000001",
  1889=>"111111111",
  1890=>"111111111",
  1891=>"001000110",
  1892=>"001001001",
  1893=>"000000000",
  1894=>"111111111",
  1895=>"111001001",
  1896=>"111001001",
  1897=>"111010000",
  1898=>"000000111",
  1899=>"010111111",
  1900=>"111110000",
  1901=>"111111000",
  1902=>"000111111",
  1903=>"000000000",
  1904=>"000000001",
  1905=>"000100111",
  1906=>"111010001",
  1907=>"000000100",
  1908=>"000000000",
  1909=>"000111010",
  1910=>"111111111",
  1911=>"000001111",
  1912=>"100000101",
  1913=>"111111111",
  1914=>"000101101",
  1915=>"111011010",
  1916=>"000000101",
  1917=>"000000000",
  1918=>"000001111",
  1919=>"000000111",
  1920=>"111000000",
  1921=>"000000000",
  1922=>"110111110",
  1923=>"111011111",
  1924=>"110100100",
  1925=>"111111111",
  1926=>"111100100",
  1927=>"111011111",
  1928=>"111000000",
  1929=>"110110111",
  1930=>"000000010",
  1931=>"000000000",
  1932=>"100000001",
  1933=>"001001000",
  1934=>"111000000",
  1935=>"000100101",
  1936=>"000000000",
  1937=>"111111000",
  1938=>"101111111",
  1939=>"100110000",
  1940=>"011000000",
  1941=>"000000000",
  1942=>"100110111",
  1943=>"000111000",
  1944=>"000000011",
  1945=>"000000000",
  1946=>"000000000",
  1947=>"110111111",
  1948=>"111111000",
  1949=>"111111111",
  1950=>"100100000",
  1951=>"110111111",
  1952=>"000000000",
  1953=>"011011001",
  1954=>"111111000",
  1955=>"000000000",
  1956=>"111111000",
  1957=>"000000000",
  1958=>"111000111",
  1959=>"010111010",
  1960=>"110000000",
  1961=>"000000000",
  1962=>"111111110",
  1963=>"000000000",
  1964=>"111000000",
  1965=>"000000000",
  1966=>"111101000",
  1967=>"100000001",
  1968=>"011111111",
  1969=>"000110111",
  1970=>"000000011",
  1971=>"111000111",
  1972=>"000000000",
  1973=>"000001011",
  1974=>"001111000",
  1975=>"010010000",
  1976=>"000000000",
  1977=>"001111010",
  1978=>"111000110",
  1979=>"111111111",
  1980=>"010000000",
  1981=>"111000100",
  1982=>"000000000",
  1983=>"000001001",
  1984=>"000000000",
  1985=>"111100111",
  1986=>"000000000",
  1987=>"000000000",
  1988=>"111111000",
  1989=>"000010100",
  1990=>"111111010",
  1991=>"110110110",
  1992=>"100111111",
  1993=>"000001111",
  1994=>"000000000",
  1995=>"001000111",
  1996=>"111010100",
  1997=>"011010111",
  1998=>"111000000",
  1999=>"000110111",
  2000=>"000010000",
  2001=>"111000100",
  2002=>"111111111",
  2003=>"000000101",
  2004=>"111111000",
  2005=>"000000000",
  2006=>"000000110",
  2007=>"110111111",
  2008=>"000000000",
  2009=>"001001111",
  2010=>"111111111",
  2011=>"000001000",
  2012=>"010110111",
  2013=>"000011111",
  2014=>"111111111",
  2015=>"101111111",
  2016=>"111010110",
  2017=>"110111111",
  2018=>"111010011",
  2019=>"000000000",
  2020=>"000000001",
  2021=>"111111111",
  2022=>"000000001",
  2023=>"111101111",
  2024=>"111100000",
  2025=>"111111000",
  2026=>"010000000",
  2027=>"000000100",
  2028=>"000100110",
  2029=>"000000100",
  2030=>"111111111",
  2031=>"111111111",
  2032=>"000111111",
  2033=>"000000010",
  2034=>"011011001",
  2035=>"110000000",
  2036=>"111000000",
  2037=>"111001001",
  2038=>"000100101",
  2039=>"110110000",
  2040=>"111111111",
  2041=>"000000000",
  2042=>"101000000",
  2043=>"111000000",
  2044=>"010110011",
  2045=>"001001001",
  2046=>"101000000",
  2047=>"000111111",
  2048=>"111111111",
  2049=>"000000000",
  2050=>"111111111",
  2051=>"000000000",
  2052=>"111111111",
  2053=>"011011010",
  2054=>"111111111",
  2055=>"111001001",
  2056=>"000000000",
  2057=>"110010000",
  2058=>"000000000",
  2059=>"000000000",
  2060=>"000010000",
  2061=>"000100100",
  2062=>"000000001",
  2063=>"111111111",
  2064=>"111111000",
  2065=>"000011011",
  2066=>"000001001",
  2067=>"111111111",
  2068=>"000000000",
  2069=>"111000000",
  2070=>"111111111",
  2071=>"000000001",
  2072=>"010010100",
  2073=>"010110000",
  2074=>"111111100",
  2075=>"111011000",
  2076=>"000000000",
  2077=>"011001100",
  2078=>"001101111",
  2079=>"000000001",
  2080=>"000000000",
  2081=>"000110111",
  2082=>"100100000",
  2083=>"001000111",
  2084=>"000000010",
  2085=>"000001000",
  2086=>"000000110",
  2087=>"111000000",
  2088=>"000000000",
  2089=>"010111011",
  2090=>"111111111",
  2091=>"100110110",
  2092=>"000000000",
  2093=>"111111111",
  2094=>"111100111",
  2095=>"111111110",
  2096=>"111111111",
  2097=>"000000000",
  2098=>"000100011",
  2099=>"000000000",
  2100=>"000111111",
  2101=>"011011011",
  2102=>"000101110",
  2103=>"111111111",
  2104=>"111100000",
  2105=>"101100000",
  2106=>"111110110",
  2107=>"101111111",
  2108=>"000101111",
  2109=>"111111011",
  2110=>"110110000",
  2111=>"111011000",
  2112=>"000010000",
  2113=>"000000000",
  2114=>"100100111",
  2115=>"110111111",
  2116=>"000000110",
  2117=>"111111111",
  2118=>"111111000",
  2119=>"111111111",
  2120=>"111111111",
  2121=>"000000111",
  2122=>"111111111",
  2123=>"001000111",
  2124=>"100001111",
  2125=>"000000111",
  2126=>"001000000",
  2127=>"000000100",
  2128=>"111111000",
  2129=>"111000011",
  2130=>"111101100",
  2131=>"111111111",
  2132=>"000000010",
  2133=>"000000000",
  2134=>"000100000",
  2135=>"000000000",
  2136=>"000000110",
  2137=>"000101111",
  2138=>"111101001",
  2139=>"011001000",
  2140=>"111110000",
  2141=>"011111111",
  2142=>"000000100",
  2143=>"100100110",
  2144=>"111000000",
  2145=>"100100111",
  2146=>"111111111",
  2147=>"111011010",
  2148=>"100100000",
  2149=>"000000000",
  2150=>"101111110",
  2151=>"000100111",
  2152=>"001000000",
  2153=>"111111000",
  2154=>"000000000",
  2155=>"000000000",
  2156=>"000001000",
  2157=>"111111111",
  2158=>"111111111",
  2159=>"011010010",
  2160=>"100000000",
  2161=>"111111111",
  2162=>"111100111",
  2163=>"000110111",
  2164=>"000000000",
  2165=>"011000000",
  2166=>"100000000",
  2167=>"000111111",
  2168=>"001000011",
  2169=>"000111111",
  2170=>"001000000",
  2171=>"011001001",
  2172=>"000000000",
  2173=>"000000011",
  2174=>"000000111",
  2175=>"000000000",
  2176=>"000000000",
  2177=>"111110111",
  2178=>"000000000",
  2179=>"001101111",
  2180=>"110110000",
  2181=>"000000000",
  2182=>"111111111",
  2183=>"000000000",
  2184=>"000000000",
  2185=>"000000000",
  2186=>"000000000",
  2187=>"111101111",
  2188=>"000000000",
  2189=>"111110000",
  2190=>"110011011",
  2191=>"000000100",
  2192=>"111111111",
  2193=>"010010111",
  2194=>"000000000",
  2195=>"111111111",
  2196=>"000100100",
  2197=>"000100111",
  2198=>"111001000",
  2199=>"111100000",
  2200=>"111111111",
  2201=>"000000000",
  2202=>"000000000",
  2203=>"111111111",
  2204=>"111111111",
  2205=>"111110011",
  2206=>"011011111",
  2207=>"000000110",
  2208=>"110110110",
  2209=>"000100110",
  2210=>"111111000",
  2211=>"111111000",
  2212=>"000000000",
  2213=>"111111001",
  2214=>"111111111",
  2215=>"000100110",
  2216=>"101101111",
  2217=>"000000111",
  2218=>"100000000",
  2219=>"000000010",
  2220=>"111011000",
  2221=>"000001001",
  2222=>"111111111",
  2223=>"001111000",
  2224=>"000011000",
  2225=>"011011101",
  2226=>"110100100",
  2227=>"000000000",
  2228=>"000011011",
  2229=>"000000000",
  2230=>"111101111",
  2231=>"111110111",
  2232=>"110111101",
  2233=>"101101111",
  2234=>"000111100",
  2235=>"101101101",
  2236=>"000000001",
  2237=>"001001001",
  2238=>"000000011",
  2239=>"111111100",
  2240=>"111111000",
  2241=>"001111111",
  2242=>"000000000",
  2243=>"000110111",
  2244=>"000000000",
  2245=>"000000010",
  2246=>"111111111",
  2247=>"011110000",
  2248=>"000100000",
  2249=>"000000001",
  2250=>"110111111",
  2251=>"011111111",
  2252=>"000000000",
  2253=>"000110000",
  2254=>"000000000",
  2255=>"000000000",
  2256=>"000000000",
  2257=>"111110110",
  2258=>"001000000",
  2259=>"111111111",
  2260=>"000000000",
  2261=>"111011001",
  2262=>"001000000",
  2263=>"000000011",
  2264=>"111010000",
  2265=>"111000000",
  2266=>"000000000",
  2267=>"000001000",
  2268=>"001001001",
  2269=>"111111110",
  2270=>"000000111",
  2271=>"011000000",
  2272=>"000000000",
  2273=>"111111101",
  2274=>"111111000",
  2275=>"001001000",
  2276=>"100000000",
  2277=>"011011111",
  2278=>"000000110",
  2279=>"110111100",
  2280=>"111001000",
  2281=>"111101000",
  2282=>"111111001",
  2283=>"000111111",
  2284=>"001111000",
  2285=>"100000000",
  2286=>"000000000",
  2287=>"111101101",
  2288=>"111110000",
  2289=>"111111000",
  2290=>"111101100",
  2291=>"000000000",
  2292=>"111111111",
  2293=>"001001011",
  2294=>"111111110",
  2295=>"111100000",
  2296=>"000000111",
  2297=>"010000000",
  2298=>"000000000",
  2299=>"111011010",
  2300=>"000001011",
  2301=>"100010010",
  2302=>"001000000",
  2303=>"110001011",
  2304=>"111111111",
  2305=>"100100110",
  2306=>"000000100",
  2307=>"000000000",
  2308=>"100110111",
  2309=>"110000000",
  2310=>"111111111",
  2311=>"100100101",
  2312=>"000000001",
  2313=>"101001001",
  2314=>"001001001",
  2315=>"111001000",
  2316=>"111111111",
  2317=>"000100101",
  2318=>"101001000",
  2319=>"001111111",
  2320=>"000010110",
  2321=>"001001000",
  2322=>"001000000",
  2323=>"001001001",
  2324=>"100110111",
  2325=>"000111111",
  2326=>"001000101",
  2327=>"000000100",
  2328=>"000000000",
  2329=>"001000101",
  2330=>"000100111",
  2331=>"000000000",
  2332=>"001011010",
  2333=>"000000000",
  2334=>"111111111",
  2335=>"000001111",
  2336=>"000000011",
  2337=>"101111111",
  2338=>"101001000",
  2339=>"110111111",
  2340=>"000110101",
  2341=>"111111110",
  2342=>"000000100",
  2343=>"000100100",
  2344=>"000000000",
  2345=>"000000000",
  2346=>"000000101",
  2347=>"000000000",
  2348=>"011001111",
  2349=>"111111111",
  2350=>"000111000",
  2351=>"000111111",
  2352=>"111111111",
  2353=>"000000000",
  2354=>"111111111",
  2355=>"000000000",
  2356=>"001000000",
  2357=>"111111111",
  2358=>"000100100",
  2359=>"101101000",
  2360=>"111111111",
  2361=>"111001111",
  2362=>"000000001",
  2363=>"111111111",
  2364=>"100110100",
  2365=>"111111000",
  2366=>"000100100",
  2367=>"111111111",
  2368=>"000000100",
  2369=>"011000000",
  2370=>"000000000",
  2371=>"001000000",
  2372=>"100000111",
  2373=>"011111000",
  2374=>"111111111",
  2375=>"111111111",
  2376=>"000011111",
  2377=>"110010000",
  2378=>"011001101",
  2379=>"100000100",
  2380=>"000000000",
  2381=>"111111111",
  2382=>"000000101",
  2383=>"111111111",
  2384=>"100100100",
  2385=>"100101111",
  2386=>"000000000",
  2387=>"111111111",
  2388=>"000101101",
  2389=>"000001011",
  2390=>"100111100",
  2391=>"100000000",
  2392=>"000000000",
  2393=>"000000000",
  2394=>"111110001",
  2395=>"000110111",
  2396=>"111111111",
  2397=>"111110000",
  2398=>"111101000",
  2399=>"001011011",
  2400=>"111111111",
  2401=>"111111111",
  2402=>"100010011",
  2403=>"000111111",
  2404=>"000000000",
  2405=>"000000100",
  2406=>"111111000",
  2407=>"111111110",
  2408=>"101001111",
  2409=>"000011000",
  2410=>"000110000",
  2411=>"110100000",
  2412=>"000011001",
  2413=>"101000111",
  2414=>"111111111",
  2415=>"010111100",
  2416=>"111111000",
  2417=>"000000000",
  2418=>"111111111",
  2419=>"011011111",
  2420=>"111111101",
  2421=>"111111111",
  2422=>"011000000",
  2423=>"000011001",
  2424=>"101001000",
  2425=>"001111111",
  2426=>"110111111",
  2427=>"101100100",
  2428=>"011000110",
  2429=>"111111111",
  2430=>"111111111",
  2431=>"111101000",
  2432=>"111110000",
  2433=>"010110011",
  2434=>"111111111",
  2435=>"000000000",
  2436=>"111000000",
  2437=>"001000001",
  2438=>"100000000",
  2439=>"001001000",
  2440=>"000000000",
  2441=>"001001000",
  2442=>"001000000",
  2443=>"001111101",
  2444=>"111111111",
  2445=>"000000000",
  2446=>"001001111",
  2447=>"111111000",
  2448=>"111110000",
  2449=>"110000000",
  2450=>"000000000",
  2451=>"011111001",
  2452=>"111001000",
  2453=>"000000111",
  2454=>"100000001",
  2455=>"000000000",
  2456=>"111100111",
  2457=>"111110010",
  2458=>"111111111",
  2459=>"000101111",
  2460=>"111111110",
  2461=>"111111000",
  2462=>"000000000",
  2463=>"010010000",
  2464=>"001000000",
  2465=>"100110110",
  2466=>"000001001",
  2467=>"111111111",
  2468=>"111111001",
  2469=>"000001110",
  2470=>"011011000",
  2471=>"000100000",
  2472=>"001000110",
  2473=>"111111101",
  2474=>"000000000",
  2475=>"000000101",
  2476=>"110111111",
  2477=>"000000000",
  2478=>"111011011",
  2479=>"111111111",
  2480=>"000000100",
  2481=>"110111110",
  2482=>"000000000",
  2483=>"111111111",
  2484=>"000000000",
  2485=>"111111111",
  2486=>"001000000",
  2487=>"000000000",
  2488=>"111111110",
  2489=>"111111111",
  2490=>"000111111",
  2491=>"000000000",
  2492=>"000000111",
  2493=>"000000000",
  2494=>"001111111",
  2495=>"000011111",
  2496=>"101101000",
  2497=>"001011011",
  2498=>"000000000",
  2499=>"000111111",
  2500=>"111100111",
  2501=>"001001001",
  2502=>"111111111",
  2503=>"111111111",
  2504=>"110001111",
  2505=>"000010111",
  2506=>"111111000",
  2507=>"000000101",
  2508=>"110000000",
  2509=>"111111000",
  2510=>"111111100",
  2511=>"111111001",
  2512=>"000000111",
  2513=>"001111111",
  2514=>"000000011",
  2515=>"111111111",
  2516=>"111111111",
  2517=>"000000000",
  2518=>"000011011",
  2519=>"000000000",
  2520=>"100100000",
  2521=>"100111111",
  2522=>"000100101",
  2523=>"111111000",
  2524=>"000000000",
  2525=>"100100101",
  2526=>"000001111",
  2527=>"111111111",
  2528=>"000000000",
  2529=>"000111010",
  2530=>"111111111",
  2531=>"111111111",
  2532=>"110110111",
  2533=>"000110011",
  2534=>"001000000",
  2535=>"001000111",
  2536=>"111111000",
  2537=>"000100111",
  2538=>"000000100",
  2539=>"000001111",
  2540=>"000000000",
  2541=>"000011011",
  2542=>"010010000",
  2543=>"111111111",
  2544=>"000001111",
  2545=>"110000000",
  2546=>"111111111",
  2547=>"000000000",
  2548=>"001001110",
  2549=>"111001000",
  2550=>"000000100",
  2551=>"000000111",
  2552=>"001111111",
  2553=>"000000100",
  2554=>"000011000",
  2555=>"111111000",
  2556=>"000000000",
  2557=>"111111000",
  2558=>"111111111",
  2559=>"000000000",
  2560=>"111110111",
  2561=>"111111111",
  2562=>"011001111",
  2563=>"110110110",
  2564=>"100101001",
  2565=>"011000100",
  2566=>"000000000",
  2567=>"111111111",
  2568=>"011011111",
  2569=>"000000100",
  2570=>"011000000",
  2571=>"111111111",
  2572=>"100010010",
  2573=>"000000110",
  2574=>"001000110",
  2575=>"000010010",
  2576=>"101101001",
  2577=>"000000000",
  2578=>"000000010",
  2579=>"000000000",
  2580=>"111100000",
  2581=>"111011000",
  2582=>"111111111",
  2583=>"000000100",
  2584=>"111000000",
  2585=>"100000100",
  2586=>"111100100",
  2587=>"000000000",
  2588=>"111111111",
  2589=>"000000001",
  2590=>"101101101",
  2591=>"110000111",
  2592=>"010110110",
  2593=>"000000000",
  2594=>"110110110",
  2595=>"111111111",
  2596=>"111111111",
  2597=>"001111111",
  2598=>"011000000",
  2599=>"111111101",
  2600=>"000000111",
  2601=>"001001111",
  2602=>"001100111",
  2603=>"000000000",
  2604=>"000000000",
  2605=>"010011001",
  2606=>"011011111",
  2607=>"000100100",
  2608=>"000000100",
  2609=>"000000001",
  2610=>"000100110",
  2611=>"111111111",
  2612=>"000011011",
  2613=>"101101101",
  2614=>"011000000",
  2615=>"111111111",
  2616=>"111000001",
  2617=>"000000000",
  2618=>"111000000",
  2619=>"111111111",
  2620=>"111111111",
  2621=>"000000000",
  2622=>"110110100",
  2623=>"010011111",
  2624=>"000110111",
  2625=>"000000001",
  2626=>"111110110",
  2627=>"011000000",
  2628=>"111001000",
  2629=>"000000000",
  2630=>"000000001",
  2631=>"111111111",
  2632=>"000000000",
  2633=>"001100100",
  2634=>"011011111",
  2635=>"111111100",
  2636=>"101000000",
  2637=>"111111100",
  2638=>"001001011",
  2639=>"111000000",
  2640=>"000000000",
  2641=>"000000111",
  2642=>"110111111",
  2643=>"100000000",
  2644=>"110111100",
  2645=>"000000100",
  2646=>"000000000",
  2647=>"000000000",
  2648=>"000100100",
  2649=>"111001000",
  2650=>"101101101",
  2651=>"111111111",
  2652=>"111111111",
  2653=>"000000000",
  2654=>"111111111",
  2655=>"111011111",
  2656=>"110110111",
  2657=>"100111111",
  2658=>"011111010",
  2659=>"111111111",
  2660=>"001001001",
  2661=>"010010000",
  2662=>"111100100",
  2663=>"111101000",
  2664=>"110000110",
  2665=>"010011111",
  2666=>"101001111",
  2667=>"111111111",
  2668=>"111111111",
  2669=>"110111101",
  2670=>"111100111",
  2671=>"000000000",
  2672=>"010000000",
  2673=>"111101101",
  2674=>"101101101",
  2675=>"111111111",
  2676=>"111110100",
  2677=>"110100100",
  2678=>"000000000",
  2679=>"111111111",
  2680=>"111111111",
  2681=>"110110000",
  2682=>"101101001",
  2683=>"111111111",
  2684=>"111111111",
  2685=>"101000000",
  2686=>"110100011",
  2687=>"110111111",
  2688=>"000000000",
  2689=>"100111101",
  2690=>"000001111",
  2691=>"000000000",
  2692=>"000000100",
  2693=>"000000001",
  2694=>"110110000",
  2695=>"111110111",
  2696=>"000000100",
  2697=>"111011011",
  2698=>"111111111",
  2699=>"110110100",
  2700=>"000000001",
  2701=>"111001011",
  2702=>"111101101",
  2703=>"011101100",
  2704=>"010111111",
  2705=>"000010000",
  2706=>"010110111",
  2707=>"000000000",
  2708=>"000000000",
  2709=>"000100110",
  2710=>"000000000",
  2711=>"001111111",
  2712=>"111111111",
  2713=>"001001111",
  2714=>"100111000",
  2715=>"000000000",
  2716=>"000000110",
  2717=>"110100100",
  2718=>"101001100",
  2719=>"111111111",
  2720=>"110111111",
  2721=>"111011111",
  2722=>"111111111",
  2723=>"111111111",
  2724=>"111101111",
  2725=>"110111111",
  2726=>"110110111",
  2727=>"000111111",
  2728=>"111111111",
  2729=>"000110000",
  2730=>"001000000",
  2731=>"110000110",
  2732=>"001001000",
  2733=>"110100101",
  2734=>"111111111",
  2735=>"110110000",
  2736=>"000000110",
  2737=>"001000000",
  2738=>"111111111",
  2739=>"111111111",
  2740=>"110100111",
  2741=>"111111111",
  2742=>"000000000",
  2743=>"000000001",
  2744=>"000100000",
  2745=>"000000100",
  2746=>"101100000",
  2747=>"101110111",
  2748=>"111000111",
  2749=>"000000000",
  2750=>"111111100",
  2751=>"111111111",
  2752=>"111111111",
  2753=>"000000000",
  2754=>"111111111",
  2755=>"000100111",
  2756=>"000000000",
  2757=>"100111111",
  2758=>"000000001",
  2759=>"111111111",
  2760=>"101000000",
  2761=>"000001111",
  2762=>"000000100",
  2763=>"111111110",
  2764=>"000000111",
  2765=>"000000000",
  2766=>"000000111",
  2767=>"000000110",
  2768=>"000001000",
  2769=>"000000000",
  2770=>"110000000",
  2771=>"111111111",
  2772=>"111111000",
  2773=>"000011111",
  2774=>"111000000",
  2775=>"110110000",
  2776=>"110110111",
  2777=>"101000000",
  2778=>"000000000",
  2779=>"110000000",
  2780=>"111111111",
  2781=>"000110100",
  2782=>"000000000",
  2783=>"000110111",
  2784=>"000000000",
  2785=>"001001000",
  2786=>"001000000",
  2787=>"110111011",
  2788=>"111111111",
  2789=>"001001000",
  2790=>"111000000",
  2791=>"111111100",
  2792=>"111110001",
  2793=>"111111111",
  2794=>"000001111",
  2795=>"101101001",
  2796=>"111111110",
  2797=>"111111111",
  2798=>"000000000",
  2799=>"111111111",
  2800=>"000000001",
  2801=>"101111001",
  2802=>"000000111",
  2803=>"111111011",
  2804=>"010001111",
  2805=>"111111111",
  2806=>"011111110",
  2807=>"111111000",
  2808=>"110000110",
  2809=>"000010010",
  2810=>"000000111",
  2811=>"111111111",
  2812=>"100111011",
  2813=>"010010111",
  2814=>"100000100",
  2815=>"111111111",
  2816=>"110000000",
  2817=>"000000101",
  2818=>"000000000",
  2819=>"010110100",
  2820=>"111111001",
  2821=>"111111010",
  2822=>"111111000",
  2823=>"100100100",
  2824=>"100000000",
  2825=>"111111111",
  2826=>"000000000",
  2827=>"000000000",
  2828=>"111111111",
  2829=>"011111111",
  2830=>"110111101",
  2831=>"110111100",
  2832=>"100100101",
  2833=>"011011000",
  2834=>"000000000",
  2835=>"111111101",
  2836=>"111111101",
  2837=>"111000000",
  2838=>"011111000",
  2839=>"000000000",
  2840=>"110111110",
  2841=>"101001001",
  2842=>"110100000",
  2843=>"000001011",
  2844=>"111111010",
  2845=>"000000111",
  2846=>"111111111",
  2847=>"000000000",
  2848=>"011101111",
  2849=>"111111111",
  2850=>"001000111",
  2851=>"111000000",
  2852=>"001011111",
  2853=>"000000001",
  2854=>"111111110",
  2855=>"111011101",
  2856=>"001000010",
  2857=>"000000000",
  2858=>"000000111",
  2859=>"111111100",
  2860=>"000001001",
  2861=>"111111111",
  2862=>"111100111",
  2863=>"100100111",
  2864=>"000000000",
  2865=>"001001111",
  2866=>"000000010",
  2867=>"000000100",
  2868=>"111101000",
  2869=>"010011000",
  2870=>"110110111",
  2871=>"000000111",
  2872=>"111111100",
  2873=>"111111111",
  2874=>"100100100",
  2875=>"000100111",
  2876=>"001001001",
  2877=>"110111000",
  2878=>"110110110",
  2879=>"111111011",
  2880=>"000000000",
  2881=>"111111111",
  2882=>"000000001",
  2883=>"111111111",
  2884=>"010110111",
  2885=>"111111111",
  2886=>"000000001",
  2887=>"101001001",
  2888=>"000110011",
  2889=>"000000000",
  2890=>"000111100",
  2891=>"010000000",
  2892=>"011111111",
  2893=>"000000000",
  2894=>"100100111",
  2895=>"000001001",
  2896=>"001010110",
  2897=>"111111111",
  2898=>"000110000",
  2899=>"000000000",
  2900=>"000000111",
  2901=>"011011000",
  2902=>"000000111",
  2903=>"000100100",
  2904=>"000000001",
  2905=>"001000001",
  2906=>"010010111",
  2907=>"101101100",
  2908=>"111111111",
  2909=>"111111111",
  2910=>"111111111",
  2911=>"011001001",
  2912=>"011111001",
  2913=>"000000000",
  2914=>"000000000",
  2915=>"000000000",
  2916=>"000011010",
  2917=>"111111111",
  2918=>"000000000",
  2919=>"011111110",
  2920=>"011101001",
  2921=>"111000000",
  2922=>"000000111",
  2923=>"011011011",
  2924=>"001000000",
  2925=>"101000001",
  2926=>"111111111",
  2927=>"110010011",
  2928=>"111111000",
  2929=>"110110111",
  2930=>"100110110",
  2931=>"101001111",
  2932=>"100000000",
  2933=>"000000001",
  2934=>"101110111",
  2935=>"001011011",
  2936=>"000000110",
  2937=>"110111111",
  2938=>"110110100",
  2939=>"101101101",
  2940=>"111111011",
  2941=>"000000000",
  2942=>"000000000",
  2943=>"000000000",
  2944=>"001011000",
  2945=>"000000000",
  2946=>"001001100",
  2947=>"000000000",
  2948=>"000000000",
  2949=>"001001001",
  2950=>"001011111",
  2951=>"101100100",
  2952=>"111101111",
  2953=>"111101101",
  2954=>"111000111",
  2955=>"001001000",
  2956=>"111111111",
  2957=>"111111111",
  2958=>"001000000",
  2959=>"111111010",
  2960=>"000010010",
  2961=>"010000000",
  2962=>"010000000",
  2963=>"110110110",
  2964=>"000000000",
  2965=>"000000000",
  2966=>"111101000",
  2967=>"111111101",
  2968=>"111111001",
  2969=>"111111111",
  2970=>"000010000",
  2971=>"000100100",
  2972=>"000000010",
  2973=>"000010011",
  2974=>"000010110",
  2975=>"000000001",
  2976=>"000111111",
  2977=>"111111111",
  2978=>"111001000",
  2979=>"111001111",
  2980=>"111111111",
  2981=>"100000100",
  2982=>"000000000",
  2983=>"110110111",
  2984=>"000000000",
  2985=>"001011111",
  2986=>"111111111",
  2987=>"011010000",
  2988=>"000000001",
  2989=>"111101111",
  2990=>"001000000",
  2991=>"110110110",
  2992=>"111111111",
  2993=>"111111010",
  2994=>"000001000",
  2995=>"000111100",
  2996=>"111111111",
  2997=>"100100000",
  2998=>"111001011",
  2999=>"000000000",
  3000=>"111110000",
  3001=>"111111111",
  3002=>"000100011",
  3003=>"001011111",
  3004=>"111111111",
  3005=>"000001100",
  3006=>"110111111",
  3007=>"101101111",
  3008=>"111001011",
  3009=>"001011000",
  3010=>"111111111",
  3011=>"000000000",
  3012=>"111000000",
  3013=>"100101111",
  3014=>"110111110",
  3015=>"111111110",
  3016=>"110100111",
  3017=>"000000110",
  3018=>"110000000",
  3019=>"000011000",
  3020=>"110000001",
  3021=>"111111001",
  3022=>"001110110",
  3023=>"000000000",
  3024=>"000000000",
  3025=>"111101101",
  3026=>"000000000",
  3027=>"000110110",
  3028=>"111111101",
  3029=>"000000011",
  3030=>"110101001",
  3031=>"000000000",
  3032=>"011000100",
  3033=>"000000001",
  3034=>"111000000",
  3035=>"000000000",
  3036=>"110000111",
  3037=>"110111000",
  3038=>"100100000",
  3039=>"100100101",
  3040=>"001000111",
  3041=>"000000001",
  3042=>"111111111",
  3043=>"001000111",
  3044=>"110000000",
  3045=>"111111111",
  3046=>"111011111",
  3047=>"001000000",
  3048=>"000000000",
  3049=>"101100111",
  3050=>"000100110",
  3051=>"111001000",
  3052=>"000000000",
  3053=>"000010010",
  3054=>"000000000",
  3055=>"000000000",
  3056=>"100110111",
  3057=>"111111111",
  3058=>"111100100",
  3059=>"101111111",
  3060=>"110011111",
  3061=>"000001011",
  3062=>"000000111",
  3063=>"111111111",
  3064=>"001001111",
  3065=>"101100110",
  3066=>"111111111",
  3067=>"111111011",
  3068=>"000000100",
  3069=>"100100111",
  3070=>"001001100",
  3071=>"010010111",
  3072=>"000001111",
  3073=>"100000001",
  3074=>"000000100",
  3075=>"111111111",
  3076=>"111111000",
  3077=>"111100000",
  3078=>"000000111",
  3079=>"000001111",
  3080=>"011111110",
  3081=>"111011000",
  3082=>"001100111",
  3083=>"111000000",
  3084=>"110000000",
  3085=>"000000111",
  3086=>"000001101",
  3087=>"000100110",
  3088=>"000000001",
  3089=>"011000111",
  3090=>"000001000",
  3091=>"111111110",
  3092=>"101111111",
  3093=>"110000111",
  3094=>"000000000",
  3095=>"011011111",
  3096=>"111111111",
  3097=>"011111111",
  3098=>"000000000",
  3099=>"111111000",
  3100=>"111000001",
  3101=>"000000011",
  3102=>"000110000",
  3103=>"000010111",
  3104=>"000111111",
  3105=>"111111110",
  3106=>"011011000",
  3107=>"000001000",
  3108=>"000011111",
  3109=>"111111001",
  3110=>"111111111",
  3111=>"000000111",
  3112=>"000000111",
  3113=>"000000000",
  3114=>"111111111",
  3115=>"110111111",
  3116=>"000000101",
  3117=>"110111101",
  3118=>"000000100",
  3119=>"010110000",
  3120=>"000001001",
  3121=>"000000000",
  3122=>"000001001",
  3123=>"101000000",
  3124=>"111111110",
  3125=>"111111100",
  3126=>"001001111",
  3127=>"000110110",
  3128=>"000000110",
  3129=>"111000000",
  3130=>"111000101",
  3131=>"111001001",
  3132=>"111111001",
  3133=>"111100100",
  3134=>"111101011",
  3135=>"111000111",
  3136=>"111111000",
  3137=>"000000111",
  3138=>"000000000",
  3139=>"011000101",
  3140=>"000011110",
  3141=>"000000001",
  3142=>"111111111",
  3143=>"111111111",
  3144=>"001000000",
  3145=>"111111111",
  3146=>"000100111",
  3147=>"111111110",
  3148=>"000001001",
  3149=>"111111111",
  3150=>"011000001",
  3151=>"111010010",
  3152=>"000000000",
  3153=>"111000000",
  3154=>"111000000",
  3155=>"001001111",
  3156=>"001000111",
  3157=>"000000000",
  3158=>"000000000",
  3159=>"101101111",
  3160=>"000011001",
  3161=>"111111000",
  3162=>"001000111",
  3163=>"001000111",
  3164=>"000111000",
  3165=>"101001000",
  3166=>"111111111",
  3167=>"101100000",
  3168=>"000000000",
  3169=>"111110110",
  3170=>"111000000",
  3171=>"100100000",
  3172=>"000000000",
  3173=>"000111111",
  3174=>"000000000",
  3175=>"000000111",
  3176=>"111111111",
  3177=>"000000100",
  3178=>"111111111",
  3179=>"111111000",
  3180=>"111110000",
  3181=>"000000000",
  3182=>"111111111",
  3183=>"110111011",
  3184=>"110111111",
  3185=>"111111000",
  3186=>"000111111",
  3187=>"111011000",
  3188=>"110100100",
  3189=>"001000000",
  3190=>"100000000",
  3191=>"000000110",
  3192=>"111011001",
  3193=>"001101111",
  3194=>"000000000",
  3195=>"111111101",
  3196=>"110100100",
  3197=>"000000111",
  3198=>"000111111",
  3199=>"111000000",
  3200=>"000000000",
  3201=>"000000001",
  3202=>"111111111",
  3203=>"000000110",
  3204=>"000000111",
  3205=>"111101100",
  3206=>"011000000",
  3207=>"111111000",
  3208=>"101111111",
  3209=>"000000001",
  3210=>"000000110",
  3211=>"000000000",
  3212=>"001010111",
  3213=>"110111111",
  3214=>"111111000",
  3215=>"000110100",
  3216=>"000010110",
  3217=>"000011111",
  3218=>"001000000",
  3219=>"100110000",
  3220=>"010000101",
  3221=>"111101100",
  3222=>"100110110",
  3223=>"111000000",
  3224=>"111001000",
  3225=>"111111111",
  3226=>"111000000",
  3227=>"111000000",
  3228=>"000000110",
  3229=>"000000011",
  3230=>"000000001",
  3231=>"001111111",
  3232=>"011010000",
  3233=>"111010110",
  3234=>"111000000",
  3235=>"100111111",
  3236=>"000000000",
  3237=>"000000000",
  3238=>"000110111",
  3239=>"011011011",
  3240=>"000100111",
  3241=>"000010111",
  3242=>"000111010",
  3243=>"000000000",
  3244=>"000000000",
  3245=>"000000111",
  3246=>"001100100",
  3247=>"000011111",
  3248=>"000001001",
  3249=>"110111110",
  3250=>"111111111",
  3251=>"000111100",
  3252=>"111101000",
  3253=>"000000000",
  3254=>"000000111",
  3255=>"000111101",
  3256=>"001111111",
  3257=>"001101000",
  3258=>"000000000",
  3259=>"000000000",
  3260=>"110111111",
  3261=>"000110111",
  3262=>"000111111",
  3263=>"000111111",
  3264=>"011111111",
  3265=>"000111111",
  3266=>"111000000",
  3267=>"110110001",
  3268=>"111111111",
  3269=>"111011000",
  3270=>"111000000",
  3271=>"000011111",
  3272=>"000000111",
  3273=>"001000000",
  3274=>"001001111",
  3275=>"111111000",
  3276=>"111111000",
  3277=>"000000000",
  3278=>"100111111",
  3279=>"111111111",
  3280=>"111111111",
  3281=>"110110011",
  3282=>"000000111",
  3283=>"000000000",
  3284=>"000000111",
  3285=>"110100100",
  3286=>"000000000",
  3287=>"111110000",
  3288=>"000001000",
  3289=>"000000110",
  3290=>"000000000",
  3291=>"010111111",
  3292=>"111111111",
  3293=>"101111110",
  3294=>"000000000",
  3295=>"111111000",
  3296=>"111000111",
  3297=>"000000101",
  3298=>"000000000",
  3299=>"100000000",
  3300=>"000000000",
  3301=>"111111111",
  3302=>"001000001",
  3303=>"100111011",
  3304=>"111111111",
  3305=>"000001011",
  3306=>"111011000",
  3307=>"111111111",
  3308=>"011000000",
  3309=>"000110111",
  3310=>"000111000",
  3311=>"001000000",
  3312=>"100110000",
  3313=>"110000000",
  3314=>"000011011",
  3315=>"000000111",
  3316=>"001001001",
  3317=>"111111000",
  3318=>"011011001",
  3319=>"111111000",
  3320=>"110111111",
  3321=>"010000000",
  3322=>"111101111",
  3323=>"111100000",
  3324=>"000001111",
  3325=>"000000001",
  3326=>"000000000",
  3327=>"000000101",
  3328=>"000100110",
  3329=>"111110111",
  3330=>"111101111",
  3331=>"110111111",
  3332=>"111111000",
  3333=>"111000000",
  3334=>"100111111",
  3335=>"100000000",
  3336=>"000000000",
  3337=>"000100111",
  3338=>"111001111",
  3339=>"110110111",
  3340=>"001000101",
  3341=>"000000111",
  3342=>"111000000",
  3343=>"111111101",
  3344=>"001111111",
  3345=>"111111000",
  3346=>"111000000",
  3347=>"000000000",
  3348=>"100000001",
  3349=>"111101000",
  3350=>"000000100",
  3351=>"000000111",
  3352=>"000011110",
  3353=>"111111000",
  3354=>"111111111",
  3355=>"100100110",
  3356=>"011011111",
  3357=>"111111100",
  3358=>"000000010",
  3359=>"111000001",
  3360=>"000100110",
  3361=>"000000100",
  3362=>"010110000",
  3363=>"000000000",
  3364=>"000110111",
  3365=>"111101111",
  3366=>"100111111",
  3367=>"000000000",
  3368=>"000000000",
  3369=>"000000000",
  3370=>"110110111",
  3371=>"111000000",
  3372=>"000000110",
  3373=>"111111000",
  3374=>"101111001",
  3375=>"000000001",
  3376=>"110000000",
  3377=>"100110100",
  3378=>"111111110",
  3379=>"110111000",
  3380=>"111101001",
  3381=>"000000101",
  3382=>"011000000",
  3383=>"111111111",
  3384=>"110111000",
  3385=>"111000101",
  3386=>"000000010",
  3387=>"111111000",
  3388=>"110100111",
  3389=>"000000111",
  3390=>"011111111",
  3391=>"111000000",
  3392=>"000000000",
  3393=>"111111111",
  3394=>"000000111",
  3395=>"000000000",
  3396=>"111111110",
  3397=>"111111100",
  3398=>"111111111",
  3399=>"000000101",
  3400=>"010000000",
  3401=>"111001011",
  3402=>"111000000",
  3403=>"000000000",
  3404=>"000110111",
  3405=>"111111001",
  3406=>"000000100",
  3407=>"111111000",
  3408=>"000000111",
  3409=>"000100111",
  3410=>"111111111",
  3411=>"111000000",
  3412=>"000111000",
  3413=>"011011011",
  3414=>"000000000",
  3415=>"111111000",
  3416=>"001000000",
  3417=>"000000000",
  3418=>"110111000",
  3419=>"001000001",
  3420=>"000000000",
  3421=>"001000000",
  3422=>"111001000",
  3423=>"000001001",
  3424=>"111011010",
  3425=>"000000011",
  3426=>"001111001",
  3427=>"111101111",
  3428=>"000000110",
  3429=>"000000001",
  3430=>"000001111",
  3431=>"111111111",
  3432=>"000000110",
  3433=>"111110110",
  3434=>"000000010",
  3435=>"011000000",
  3436=>"000000000",
  3437=>"011000100",
  3438=>"001111111",
  3439=>"000000000",
  3440=>"101000000",
  3441=>"000000000",
  3442=>"000000000",
  3443=>"000011011",
  3444=>"000011111",
  3445=>"010011000",
  3446=>"101111111",
  3447=>"011000010",
  3448=>"001000111",
  3449=>"111000000",
  3450=>"111111111",
  3451=>"011000010",
  3452=>"111111000",
  3453=>"111001000",
  3454=>"111111111",
  3455=>"111111111",
  3456=>"001000000",
  3457=>"000011011",
  3458=>"000000000",
  3459=>"101101100",
  3460=>"000000000",
  3461=>"100111111",
  3462=>"111111110",
  3463=>"000000000",
  3464=>"001000000",
  3465=>"100111111",
  3466=>"111111000",
  3467=>"110111111",
  3468=>"111000000",
  3469=>"000110100",
  3470=>"101010000",
  3471=>"000000000",
  3472=>"000000010",
  3473=>"000000000",
  3474=>"000010111",
  3475=>"001100110",
  3476=>"000000000",
  3477=>"000010000",
  3478=>"000001111",
  3479=>"000000100",
  3480=>"100111111",
  3481=>"000000000",
  3482=>"111111111",
  3483=>"111111111",
  3484=>"000010111",
  3485=>"001111111",
  3486=>"000000000",
  3487=>"000000000",
  3488=>"100111100",
  3489=>"001010000",
  3490=>"111111000",
  3491=>"011111011",
  3492=>"111111001",
  3493=>"000111111",
  3494=>"111100111",
  3495=>"111111111",
  3496=>"111111111",
  3497=>"000000000",
  3498=>"001000011",
  3499=>"100110110",
  3500=>"000000000",
  3501=>"010111011",
  3502=>"111001000",
  3503=>"000000110",
  3504=>"101111111",
  3505=>"111001011",
  3506=>"110111111",
  3507=>"111111000",
  3508=>"000000000",
  3509=>"000000111",
  3510=>"000100110",
  3511=>"000000000",
  3512=>"000000001",
  3513=>"000000000",
  3514=>"000100000",
  3515=>"000000111",
  3516=>"010010011",
  3517=>"111110000",
  3518=>"111000011",
  3519=>"100100111",
  3520=>"000110110",
  3521=>"111011010",
  3522=>"111111111",
  3523=>"000100110",
  3524=>"101000100",
  3525=>"111111111",
  3526=>"011011000",
  3527=>"110110111",
  3528=>"110111111",
  3529=>"000000000",
  3530=>"000001111",
  3531=>"110000000",
  3532=>"111000000",
  3533=>"000000111",
  3534=>"010000000",
  3535=>"000100100",
  3536=>"000000000",
  3537=>"111111111",
  3538=>"000000000",
  3539=>"111110110",
  3540=>"101000000",
  3541=>"000000000",
  3542=>"000000000",
  3543=>"110100000",
  3544=>"000000000",
  3545=>"111000000",
  3546=>"111000000",
  3547=>"111111111",
  3548=>"000000010",
  3549=>"010000111",
  3550=>"010110000",
  3551=>"001011111",
  3552=>"111111011",
  3553=>"000101111",
  3554=>"000000000",
  3555=>"000000111",
  3556=>"000000011",
  3557=>"111111111",
  3558=>"111111111",
  3559=>"111000000",
  3560=>"000000111",
  3561=>"011111111",
  3562=>"111111011",
  3563=>"000000000",
  3564=>"000000111",
  3565=>"000000011",
  3566=>"111000000",
  3567=>"111011011",
  3568=>"010110110",
  3569=>"111000000",
  3570=>"000000000",
  3571=>"000110110",
  3572=>"111111111",
  3573=>"000000111",
  3574=>"000000000",
  3575=>"110011111",
  3576=>"000101000",
  3577=>"011001011",
  3578=>"111111110",
  3579=>"111110010",
  3580=>"111111100",
  3581=>"000100111",
  3582=>"111011111",
  3583=>"000000000",
  3584=>"000000000",
  3585=>"110111111",
  3586=>"000000111",
  3587=>"000000011",
  3588=>"101001001",
  3589=>"111111000",
  3590=>"000000000",
  3591=>"111111111",
  3592=>"000000000",
  3593=>"110111011",
  3594=>"111000000",
  3595=>"111111111",
  3596=>"000000000",
  3597=>"001111111",
  3598=>"011111100",
  3599=>"001001111",
  3600=>"000111111",
  3601=>"000111111",
  3602=>"011001001",
  3603=>"100111000",
  3604=>"111111000",
  3605=>"000111111",
  3606=>"000000001",
  3607=>"000011011",
  3608=>"011111111",
  3609=>"011011011",
  3610=>"111111111",
  3611=>"111111000",
  3612=>"111000000",
  3613=>"000111111",
  3614=>"000000101",
  3615=>"110110000",
  3616=>"010110000",
  3617=>"000000111",
  3618=>"110111111",
  3619=>"000000000",
  3620=>"111111001",
  3621=>"100100111",
  3622=>"011111111",
  3623=>"111111111",
  3624=>"110001001",
  3625=>"111000000",
  3626=>"100111111",
  3627=>"000000101",
  3628=>"111111111",
  3629=>"000111111",
  3630=>"111000000",
  3631=>"000011010",
  3632=>"111100000",
  3633=>"000000000",
  3634=>"011111100",
  3635=>"000000011",
  3636=>"111001000",
  3637=>"000110100",
  3638=>"000000001",
  3639=>"000000000",
  3640=>"111111110",
  3641=>"110111111",
  3642=>"000000000",
  3643=>"011011000",
  3644=>"000000011",
  3645=>"111000000",
  3646=>"000000000",
  3647=>"111011100",
  3648=>"111111001",
  3649=>"111101101",
  3650=>"111111111",
  3651=>"000000111",
  3652=>"010010111",
  3653=>"100100100",
  3654=>"111111111",
  3655=>"110000000",
  3656=>"111111001",
  3657=>"111111100",
  3658=>"111000000",
  3659=>"100000010",
  3660=>"000000000",
  3661=>"110111100",
  3662=>"011011000",
  3663=>"000110111",
  3664=>"000011000",
  3665=>"000000000",
  3666=>"000000110",
  3667=>"000000100",
  3668=>"111000000",
  3669=>"000000000",
  3670=>"100000000",
  3671=>"111111111",
  3672=>"111011111",
  3673=>"111101111",
  3674=>"111111111",
  3675=>"001000000",
  3676=>"111001111",
  3677=>"011011011",
  3678=>"110110000",
  3679=>"111100110",
  3680=>"000000000",
  3681=>"111100000",
  3682=>"010010111",
  3683=>"111111101",
  3684=>"110110011",
  3685=>"000000000",
  3686=>"000000000",
  3687=>"000000000",
  3688=>"011011111",
  3689=>"000000000",
  3690=>"111111111",
  3691=>"001001000",
  3692=>"000000011",
  3693=>"011111111",
  3694=>"000000111",
  3695=>"000000000",
  3696=>"100000000",
  3697=>"000000000",
  3698=>"111111111",
  3699=>"111111000",
  3700=>"000000000",
  3701=>"001001001",
  3702=>"000000001",
  3703=>"111111011",
  3704=>"110110111",
  3705=>"000000100",
  3706=>"000000000",
  3707=>"110010000",
  3708=>"110000000",
  3709=>"000000000",
  3710=>"111000000",
  3711=>"000111111",
  3712=>"000000111",
  3713=>"000000000",
  3714=>"111111111",
  3715=>"000000001",
  3716=>"011111011",
  3717=>"000000000",
  3718=>"111011111",
  3719=>"000111111",
  3720=>"111111111",
  3721=>"101000111",
  3722=>"000000000",
  3723=>"000101111",
  3724=>"111011000",
  3725=>"000110110",
  3726=>"111111111",
  3727=>"000000000",
  3728=>"000000111",
  3729=>"100000000",
  3730=>"111111000",
  3731=>"111011111",
  3732=>"000001001",
  3733=>"100000111",
  3734=>"000111111",
  3735=>"111000100",
  3736=>"000000000",
  3737=>"111111111",
  3738=>"000000110",
  3739=>"000001001",
  3740=>"000000111",
  3741=>"111111010",
  3742=>"100000000",
  3743=>"110111111",
  3744=>"100100111",
  3745=>"111111000",
  3746=>"000000001",
  3747=>"000000000",
  3748=>"000010000",
  3749=>"111111111",
  3750=>"111111111",
  3751=>"010100000",
  3752=>"111000000",
  3753=>"000000111",
  3754=>"111110000",
  3755=>"000000000",
  3756=>"111011000",
  3757=>"110000111",
  3758=>"110111111",
  3759=>"111111111",
  3760=>"111111000",
  3761=>"111110100",
  3762=>"111111110",
  3763=>"000011111",
  3764=>"111000000",
  3765=>"111000101",
  3766=>"000000000",
  3767=>"000000000",
  3768=>"000010111",
  3769=>"111111111",
  3770=>"000000000",
  3771=>"000000001",
  3772=>"000000000",
  3773=>"001011011",
  3774=>"111000111",
  3775=>"000000000",
  3776=>"111111000",
  3777=>"111110000",
  3778=>"111111111",
  3779=>"111111000",
  3780=>"000000010",
  3781=>"000111111",
  3782=>"111100100",
  3783=>"111111111",
  3784=>"111111111",
  3785=>"000000000",
  3786=>"111111100",
  3787=>"111111111",
  3788=>"101000000",
  3789=>"111111111",
  3790=>"011011111",
  3791=>"010000000",
  3792=>"111111111",
  3793=>"000000000",
  3794=>"100111101",
  3795=>"010110010",
  3796=>"000000000",
  3797=>"110111110",
  3798=>"001000000",
  3799=>"001000011",
  3800=>"111111111",
  3801=>"110000001",
  3802=>"111111111",
  3803=>"111100000",
  3804=>"111111111",
  3805=>"111111110",
  3806=>"000111010",
  3807=>"000111111",
  3808=>"111111111",
  3809=>"001111111",
  3810=>"000000000",
  3811=>"001101000",
  3812=>"111111111",
  3813=>"100100000",
  3814=>"000000110",
  3815=>"000100000",
  3816=>"111111011",
  3817=>"000010110",
  3818=>"111111011",
  3819=>"100111110",
  3820=>"000000101",
  3821=>"000000000",
  3822=>"000000101",
  3823=>"000001001",
  3824=>"000000000",
  3825=>"000000111",
  3826=>"011000000",
  3827=>"000001111",
  3828=>"111111111",
  3829=>"110110001",
  3830=>"000111111",
  3831=>"111000100",
  3832=>"111111000",
  3833=>"000000000",
  3834=>"000000000",
  3835=>"011111111",
  3836=>"000110110",
  3837=>"101111101",
  3838=>"000000000",
  3839=>"000000001",
  3840=>"001011000",
  3841=>"000100111",
  3842=>"001000000",
  3843=>"000000001",
  3844=>"111001000",
  3845=>"111111111",
  3846=>"000110111",
  3847=>"000000000",
  3848=>"000000001",
  3849=>"100101000",
  3850=>"111111111",
  3851=>"111111111",
  3852=>"111101000",
  3853=>"100000000",
  3854=>"001000000",
  3855=>"000011001",
  3856=>"000110100",
  3857=>"000110111",
  3858=>"111111100",
  3859=>"000000100",
  3860=>"111111000",
  3861=>"000000110",
  3862=>"111111110",
  3863=>"110101111",
  3864=>"110111111",
  3865=>"110100100",
  3866=>"110111010",
  3867=>"111111111",
  3868=>"111111110",
  3869=>"111111110",
  3870=>"000000000",
  3871=>"010111111",
  3872=>"000110110",
  3873=>"001000111",
  3874=>"000000000",
  3875=>"000000000",
  3876=>"110000000",
  3877=>"000000100",
  3878=>"011111000",
  3879=>"111111111",
  3880=>"110110110",
  3881=>"000000111",
  3882=>"110111111",
  3883=>"111000100",
  3884=>"111111111",
  3885=>"010111001",
  3886=>"001000111",
  3887=>"000000000",
  3888=>"010110111",
  3889=>"000000001",
  3890=>"000111111",
  3891=>"000000000",
  3892=>"000000101",
  3893=>"000000000",
  3894=>"011111111",
  3895=>"111001000",
  3896=>"111101111",
  3897=>"101000000",
  3898=>"010000000",
  3899=>"111101000",
  3900=>"111111110",
  3901=>"000000111",
  3902=>"000000000",
  3903=>"111111000",
  3904=>"000000111",
  3905=>"000101111",
  3906=>"000000100",
  3907=>"111011000",
  3908=>"001001000",
  3909=>"110100100",
  3910=>"110111111",
  3911=>"111111111",
  3912=>"111000000",
  3913=>"100101001",
  3914=>"110111111",
  3915=>"000000100",
  3916=>"000000000",
  3917=>"000000000",
  3918=>"111111111",
  3919=>"110111111",
  3920=>"100111011",
  3921=>"111111000",
  3922=>"111010000",
  3923=>"000000000",
  3924=>"000000110",
  3925=>"011011001",
  3926=>"111111101",
  3927=>"000100000",
  3928=>"000000111",
  3929=>"000001001",
  3930=>"000000011",
  3931=>"001000000",
  3932=>"000111111",
  3933=>"111111111",
  3934=>"111100000",
  3935=>"111011111",
  3936=>"000111110",
  3937=>"001001001",
  3938=>"000111000",
  3939=>"111111111",
  3940=>"011111111",
  3941=>"000000000",
  3942=>"111111111",
  3943=>"000001111",
  3944=>"000000000",
  3945=>"000000111",
  3946=>"111111000",
  3947=>"111111110",
  3948=>"111011010",
  3949=>"000001001",
  3950=>"000000000",
  3951=>"100111101",
  3952=>"000000000",
  3953=>"110111111",
  3954=>"000000111",
  3955=>"000000000",
  3956=>"100111111",
  3957=>"111101000",
  3958=>"011000000",
  3959=>"000010000",
  3960=>"110000000",
  3961=>"000100111",
  3962=>"111111000",
  3963=>"111111111",
  3964=>"100111111",
  3965=>"111111111",
  3966=>"000000000",
  3967=>"000011111",
  3968=>"011111111",
  3969=>"111111111",
  3970=>"001001011",
  3971=>"111101000",
  3972=>"111111111",
  3973=>"000000111",
  3974=>"011000000",
  3975=>"111111110",
  3976=>"111000000",
  3977=>"111000100",
  3978=>"111000000",
  3979=>"111111001",
  3980=>"111111111",
  3981=>"001000000",
  3982=>"000000000",
  3983=>"000011000",
  3984=>"000000000",
  3985=>"100100101",
  3986=>"000000111",
  3987=>"011110010",
  3988=>"111111111",
  3989=>"000000001",
  3990=>"000000001",
  3991=>"000000000",
  3992=>"000000111",
  3993=>"111110010",
  3994=>"111111110",
  3995=>"110111111",
  3996=>"110010000",
  3997=>"000100100",
  3998=>"110010111",
  3999=>"000000000",
  4000=>"000111111",
  4001=>"111111110",
  4002=>"000000000",
  4003=>"111111111",
  4004=>"100000001",
  4005=>"100111000",
  4006=>"111101001",
  4007=>"111100000",
  4008=>"000000000",
  4009=>"011000000",
  4010=>"000000000",
  4011=>"110111100",
  4012=>"000000000",
  4013=>"110100110",
  4014=>"000000000",
  4015=>"010111111",
  4016=>"111100000",
  4017=>"001000000",
  4018=>"000000000",
  4019=>"000000111",
  4020=>"000000000",
  4021=>"000000000",
  4022=>"111101111",
  4023=>"000010111",
  4024=>"011010000",
  4025=>"111011000",
  4026=>"000000000",
  4027=>"000000111",
  4028=>"000000111",
  4029=>"111111111",
  4030=>"000111111",
  4031=>"001010000",
  4032=>"000000000",
  4033=>"000110110",
  4034=>"001000000",
  4035=>"000111111",
  4036=>"111111111",
  4037=>"011001000",
  4038=>"011000001",
  4039=>"000000000",
  4040=>"011000000",
  4041=>"010000110",
  4042=>"101000000",
  4043=>"000001111",
  4044=>"011000000",
  4045=>"111000111",
  4046=>"101111011",
  4047=>"100100111",
  4048=>"001000000",
  4049=>"110111111",
  4050=>"000000000",
  4051=>"000000000",
  4052=>"001001000",
  4053=>"101000000",
  4054=>"000000111",
  4055=>"000000000",
  4056=>"111000000",
  4057=>"111000000",
  4058=>"000010000",
  4059=>"100000001",
  4060=>"000100111",
  4061=>"111111111",
  4062=>"000000111",
  4063=>"011111001",
  4064=>"111111111",
  4065=>"100110111",
  4066=>"000000000",
  4067=>"000001001",
  4068=>"110010000",
  4069=>"001111111",
  4070=>"111001000",
  4071=>"000000000",
  4072=>"000000111",
  4073=>"111011110",
  4074=>"100000100",
  4075=>"000000001",
  4076=>"000111101",
  4077=>"000000001",
  4078=>"011111001",
  4079=>"001011111",
  4080=>"010011000",
  4081=>"000010010",
  4082=>"111000100",
  4083=>"001111000",
  4084=>"111001111",
  4085=>"101001001",
  4086=>"000000000",
  4087=>"100111011",
  4088=>"000000101",
  4089=>"100111001",
  4090=>"111111110",
  4091=>"000000111",
  4092=>"111111111",
  4093=>"000000000",
  4094=>"111000000",
  4095=>"111001000",
  4096=>"011001001",
  4097=>"111111001",
  4098=>"001000000",
  4099=>"011011111",
  4100=>"000000000",
  4101=>"000100110",
  4102=>"000000001",
  4103=>"101000000",
  4104=>"111111111",
  4105=>"000111010",
  4106=>"111111111",
  4107=>"110110111",
  4108=>"111011000",
  4109=>"111000000",
  4110=>"100000001",
  4111=>"111111111",
  4112=>"111111111",
  4113=>"000101111",
  4114=>"000000000",
  4115=>"100000000",
  4116=>"111111111",
  4117=>"111111000",
  4118=>"000000111",
  4119=>"111110010",
  4120=>"111011110",
  4121=>"011111111",
  4122=>"100111111",
  4123=>"100000001",
  4124=>"011000000",
  4125=>"000000100",
  4126=>"111111011",
  4127=>"010000110",
  4128=>"011111111",
  4129=>"111111011",
  4130=>"010000000",
  4131=>"000000111",
  4132=>"000000000",
  4133=>"000000000",
  4134=>"111111111",
  4135=>"000000000",
  4136=>"000111111",
  4137=>"101111111",
  4138=>"000000000",
  4139=>"000000000",
  4140=>"110110111",
  4141=>"111111001",
  4142=>"000100100",
  4143=>"000100100",
  4144=>"111101000",
  4145=>"110100000",
  4146=>"111111011",
  4147=>"000000000",
  4148=>"011111110",
  4149=>"111111111",
  4150=>"111001111",
  4151=>"111111111",
  4152=>"010011001",
  4153=>"101000100",
  4154=>"111101111",
  4155=>"111111110",
  4156=>"111111111",
  4157=>"000000000",
  4158=>"001011011",
  4159=>"000000000",
  4160=>"111111111",
  4161=>"100000000",
  4162=>"110010011",
  4163=>"110110111",
  4164=>"000000000",
  4165=>"001000111",
  4166=>"111111111",
  4167=>"111110100",
  4168=>"110010011",
  4169=>"111000111",
  4170=>"011111111",
  4171=>"100000110",
  4172=>"000000001",
  4173=>"111111111",
  4174=>"000111111",
  4175=>"011011001",
  4176=>"100100111",
  4177=>"011001011",
  4178=>"111111111",
  4179=>"000110110",
  4180=>"000000000",
  4181=>"000000000",
  4182=>"001000100",
  4183=>"000000000",
  4184=>"110110000",
  4185=>"111001101",
  4186=>"000110000",
  4187=>"111111100",
  4188=>"111111001",
  4189=>"001111111",
  4190=>"110110111",
  4191=>"100110011",
  4192=>"000101111",
  4193=>"111111111",
  4194=>"111011001",
  4195=>"000000000",
  4196=>"111111100",
  4197=>"111010110",
  4198=>"000000000",
  4199=>"111111111",
  4200=>"100100000",
  4201=>"000000000",
  4202=>"000000111",
  4203=>"111000000",
  4204=>"000000000",
  4205=>"111111111",
  4206=>"000000000",
  4207=>"111111111",
  4208=>"101111001",
  4209=>"000000000",
  4210=>"111111000",
  4211=>"000000000",
  4212=>"111011000",
  4213=>"000111111",
  4214=>"000000110",
  4215=>"111101000",
  4216=>"000000000",
  4217=>"100000101",
  4218=>"100100000",
  4219=>"111111111",
  4220=>"111111111",
  4221=>"000111111",
  4222=>"111111111",
  4223=>"010000000",
  4224=>"000000111",
  4225=>"111111111",
  4226=>"100000111",
  4227=>"011011011",
  4228=>"100100000",
  4229=>"000000000",
  4230=>"100111111",
  4231=>"111111000",
  4232=>"000100111",
  4233=>"000001111",
  4234=>"001000010",
  4235=>"000000000",
  4236=>"000000000",
  4237=>"000000000",
  4238=>"000001111",
  4239=>"111111011",
  4240=>"111111111",
  4241=>"000000000",
  4242=>"000000111",
  4243=>"111001001",
  4244=>"101000000",
  4245=>"000011001",
  4246=>"100100000",
  4247=>"111000000",
  4248=>"111111111",
  4249=>"111111111",
  4250=>"100000111",
  4251=>"111000000",
  4252=>"000000000",
  4253=>"000000000",
  4254=>"101100000",
  4255=>"000000111",
  4256=>"000000000",
  4257=>"111111111",
  4258=>"000000000",
  4259=>"111111111",
  4260=>"111011000",
  4261=>"111111000",
  4262=>"111111001",
  4263=>"111111111",
  4264=>"111111110",
  4265=>"111110010",
  4266=>"000001111",
  4267=>"111111111",
  4268=>"111101001",
  4269=>"011000000",
  4270=>"000000110",
  4271=>"001011111",
  4272=>"111100111",
  4273=>"111111111",
  4274=>"111111111",
  4275=>"000000000",
  4276=>"000001001",
  4277=>"000110010",
  4278=>"001111111",
  4279=>"000000001",
  4280=>"011001100",
  4281=>"111111000",
  4282=>"011111100",
  4283=>"000111111",
  4284=>"111111111",
  4285=>"000000000",
  4286=>"000000010",
  4287=>"111111110",
  4288=>"001000000",
  4289=>"101001001",
  4290=>"000001000",
  4291=>"111111010",
  4292=>"101111111",
  4293=>"000000000",
  4294=>"111111001",
  4295=>"111111011",
  4296=>"111111111",
  4297=>"111111111",
  4298=>"111111110",
  4299=>"011000001",
  4300=>"001000000",
  4301=>"010010000",
  4302=>"110111111",
  4303=>"111000000",
  4304=>"000000000",
  4305=>"000000001",
  4306=>"111111110",
  4307=>"000000111",
  4308=>"000000111",
  4309=>"111111111",
  4310=>"111111111",
  4311=>"111100000",
  4312=>"111111001",
  4313=>"011111000",
  4314=>"111111111",
  4315=>"000000110",
  4316=>"000111101",
  4317=>"111111111",
  4318=>"000000000",
  4319=>"111011111",
  4320=>"011010000",
  4321=>"111000000",
  4322=>"111111111",
  4323=>"111111111",
  4324=>"100100001",
  4325=>"111111111",
  4326=>"111111111",
  4327=>"111011001",
  4328=>"011011000",
  4329=>"011011000",
  4330=>"001000000",
  4331=>"000000000",
  4332=>"111111110",
  4333=>"110111111",
  4334=>"001100000",
  4335=>"011010000",
  4336=>"100100110",
  4337=>"010000000",
  4338=>"111111100",
  4339=>"000000000",
  4340=>"000000000",
  4341=>"000100111",
  4342=>"000000000",
  4343=>"111001011",
  4344=>"001000000",
  4345=>"111111111",
  4346=>"001000000",
  4347=>"001001000",
  4348=>"010111101",
  4349=>"110100100",
  4350=>"000000000",
  4351=>"000110111",
  4352=>"011011011",
  4353=>"111100100",
  4354=>"000000000",
  4355=>"000101111",
  4356=>"111111001",
  4357=>"000000000",
  4358=>"000000000",
  4359=>"111111111",
  4360=>"000011111",
  4361=>"000110111",
  4362=>"000000000",
  4363=>"000000001",
  4364=>"001101111",
  4365=>"011111011",
  4366=>"000000000",
  4367=>"111111111",
  4368=>"000000100",
  4369=>"001111001",
  4370=>"111111111",
  4371=>"000010111",
  4372=>"111111111",
  4373=>"000111111",
  4374=>"100100100",
  4375=>"001111110",
  4376=>"000000000",
  4377=>"000011111",
  4378=>"000000000",
  4379=>"000000000",
  4380=>"111111000",
  4381=>"111011000",
  4382=>"111111111",
  4383=>"000100000",
  4384=>"000000000",
  4385=>"100011111",
  4386=>"000000000",
  4387=>"011111011",
  4388=>"000000000",
  4389=>"111111111",
  4390=>"000000000",
  4391=>"011000011",
  4392=>"000011111",
  4393=>"111111111",
  4394=>"111000000",
  4395=>"111111111",
  4396=>"000111111",
  4397=>"000000001",
  4398=>"000000000",
  4399=>"111110110",
  4400=>"000000000",
  4401=>"111111111",
  4402=>"111111111",
  4403=>"000000110",
  4404=>"111001111",
  4405=>"000000110",
  4406=>"001000000",
  4407=>"000010000",
  4408=>"110100100",
  4409=>"111100111",
  4410=>"100111111",
  4411=>"111000100",
  4412=>"111111110",
  4413=>"000000111",
  4414=>"010001001",
  4415=>"011011111",
  4416=>"000000000",
  4417=>"111111111",
  4418=>"011000100",
  4419=>"111111111",
  4420=>"111000000",
  4421=>"100000000",
  4422=>"111111111",
  4423=>"000000000",
  4424=>"001000000",
  4425=>"000010001",
  4426=>"111111111",
  4427=>"000000000",
  4428=>"111111111",
  4429=>"000111111",
  4430=>"111111111",
  4431=>"011011000",
  4432=>"010011011",
  4433=>"000000000",
  4434=>"000000111",
  4435=>"000000000",
  4436=>"000000000",
  4437=>"011011001",
  4438=>"001000000",
  4439=>"110110110",
  4440=>"110100000",
  4441=>"011111011",
  4442=>"000111111",
  4443=>"111111111",
  4444=>"000000000",
  4445=>"000000010",
  4446=>"011111100",
  4447=>"111111111",
  4448=>"001000000",
  4449=>"110100000",
  4450=>"111111101",
  4451=>"111100101",
  4452=>"000000101",
  4453=>"011001111",
  4454=>"111000000",
  4455=>"110111111",
  4456=>"000000000",
  4457=>"000010000",
  4458=>"111111111",
  4459=>"011111111",
  4460=>"000100100",
  4461=>"011111111",
  4462=>"110111111",
  4463=>"111011000",
  4464=>"111111000",
  4465=>"111111111",
  4466=>"111100000",
  4467=>"001011011",
  4468=>"111111111",
  4469=>"111011000",
  4470=>"000000000",
  4471=>"000000100",
  4472=>"111101000",
  4473=>"111111000",
  4474=>"000000000",
  4475=>"110000001",
  4476=>"111111011",
  4477=>"000000000",
  4478=>"000000000",
  4479=>"111111110",
  4480=>"000100111",
  4481=>"000000100",
  4482=>"100000000",
  4483=>"111000111",
  4484=>"000001011",
  4485=>"000000111",
  4486=>"111100000",
  4487=>"000000011",
  4488=>"001111111",
  4489=>"000000000",
  4490=>"000100100",
  4491=>"111111110",
  4492=>"001000111",
  4493=>"011111111",
  4494=>"111111111",
  4495=>"000000000",
  4496=>"111111111",
  4497=>"111111111",
  4498=>"001000010",
  4499=>"111001001",
  4500=>"000000000",
  4501=>"010010000",
  4502=>"100000100",
  4503=>"000000000",
  4504=>"000000000",
  4505=>"000000001",
  4506=>"111111111",
  4507=>"110010000",
  4508=>"000000000",
  4509=>"000000000",
  4510=>"000000000",
  4511=>"000000000",
  4512=>"000010111",
  4513=>"110000000",
  4514=>"000100100",
  4515=>"001000000",
  4516=>"111111111",
  4517=>"000000000",
  4518=>"111001000",
  4519=>"110110111",
  4520=>"111111111",
  4521=>"111101111",
  4522=>"100100110",
  4523=>"111011000",
  4524=>"000000000",
  4525=>"001001001",
  4526=>"111111111",
  4527=>"011111111",
  4528=>"000111111",
  4529=>"111111111",
  4530=>"111111111",
  4531=>"000100111",
  4532=>"100001000",
  4533=>"111111111",
  4534=>"111111011",
  4535=>"111111111",
  4536=>"001010000",
  4537=>"101111111",
  4538=>"000001001",
  4539=>"111001111",
  4540=>"000000000",
  4541=>"100100111",
  4542=>"000000001",
  4543=>"100100100",
  4544=>"001000000",
  4545=>"111111111",
  4546=>"000000000",
  4547=>"111111111",
  4548=>"100000100",
  4549=>"011011011",
  4550=>"000000000",
  4551=>"000000011",
  4552=>"111111111",
  4553=>"011011000",
  4554=>"111111000",
  4555=>"000000000",
  4556=>"111010001",
  4557=>"111111111",
  4558=>"000000101",
  4559=>"000111011",
  4560=>"111101000",
  4561=>"000000000",
  4562=>"010010010",
  4563=>"111111110",
  4564=>"111111111",
  4565=>"111111101",
  4566=>"000111111",
  4567=>"001000000",
  4568=>"101101101",
  4569=>"100111110",
  4570=>"000000001",
  4571=>"111111111",
  4572=>"000000000",
  4573=>"111010000",
  4574=>"010000000",
  4575=>"101000110",
  4576=>"111111111",
  4577=>"111101101",
  4578=>"000111111",
  4579=>"111100101",
  4580=>"001111111",
  4581=>"100000000",
  4582=>"000000001",
  4583=>"000000000",
  4584=>"100000000",
  4585=>"001000000",
  4586=>"111111001",
  4587=>"001000100",
  4588=>"000000000",
  4589=>"000000010",
  4590=>"000000111",
  4591=>"000000000",
  4592=>"010110110",
  4593=>"111111111",
  4594=>"111111111",
  4595=>"110110000",
  4596=>"010100100",
  4597=>"000000011",
  4598=>"000000000",
  4599=>"001001000",
  4600=>"110000000",
  4601=>"111101000",
  4602=>"100110111",
  4603=>"000000001",
  4604=>"000000000",
  4605=>"111001000",
  4606=>"111101111",
  4607=>"111000111",
  4608=>"110110000",
  4609=>"000000000",
  4610=>"000000111",
  4611=>"001111111",
  4612=>"101101111",
  4613=>"111111110",
  4614=>"111111111",
  4615=>"111000000",
  4616=>"000000111",
  4617=>"111111011",
  4618=>"111111111",
  4619=>"000111111",
  4620=>"000000000",
  4621=>"100100111",
  4622=>"011011000",
  4623=>"000000000",
  4624=>"111001111",
  4625=>"000000111",
  4626=>"011001000",
  4627=>"111111110",
  4628=>"100000011",
  4629=>"111111111",
  4630=>"001001011",
  4631=>"110100100",
  4632=>"001001111",
  4633=>"110110100",
  4634=>"000000000",
  4635=>"000000011",
  4636=>"000000000",
  4637=>"111000000",
  4638=>"001001001",
  4639=>"000000000",
  4640=>"111001000",
  4641=>"111111111",
  4642=>"000000010",
  4643=>"111111011",
  4644=>"000000000",
  4645=>"100000001",
  4646=>"000001000",
  4647=>"000000001",
  4648=>"010111001",
  4649=>"001001000",
  4650=>"111111111",
  4651=>"111111111",
  4652=>"100110100",
  4653=>"111111011",
  4654=>"001001001",
  4655=>"001000000",
  4656=>"000000000",
  4657=>"000000000",
  4658=>"100110110",
  4659=>"100010111",
  4660=>"000100111",
  4661=>"111010110",
  4662=>"000000000",
  4663=>"110101000",
  4664=>"000000000",
  4665=>"100100000",
  4666=>"111111000",
  4667=>"000000111",
  4668=>"101000000",
  4669=>"000000000",
  4670=>"100111011",
  4671=>"111111111",
  4672=>"000111111",
  4673=>"111001100",
  4674=>"000111111",
  4675=>"001000000",
  4676=>"011110010",
  4677=>"100001111",
  4678=>"111111010",
  4679=>"111111000",
  4680=>"110100110",
  4681=>"111100111",
  4682=>"001110111",
  4683=>"000111111",
  4684=>"010010000",
  4685=>"111111000",
  4686=>"111001000",
  4687=>"000100101",
  4688=>"111111111",
  4689=>"000000001",
  4690=>"000000000",
  4691=>"111111010",
  4692=>"000000000",
  4693=>"110100100",
  4694=>"111110110",
  4695=>"000000000",
  4696=>"111111111",
  4697=>"000000000",
  4698=>"111111101",
  4699=>"111110110",
  4700=>"001001000",
  4701=>"000000001",
  4702=>"001000000",
  4703=>"001001000",
  4704=>"001001111",
  4705=>"000000000",
  4706=>"000111111",
  4707=>"111100100",
  4708=>"001111110",
  4709=>"000001011",
  4710=>"100000100",
  4711=>"111111111",
  4712=>"111111111",
  4713=>"000000100",
  4714=>"000000000",
  4715=>"000001011",
  4716=>"111110110",
  4717=>"100000000",
  4718=>"111110111",
  4719=>"100111101",
  4720=>"000000000",
  4721=>"000000000",
  4722=>"011010011",
  4723=>"111010111",
  4724=>"000000000",
  4725=>"001001001",
  4726=>"111000100",
  4727=>"000000000",
  4728=>"000110111",
  4729=>"000000000",
  4730=>"001101110",
  4731=>"000000000",
  4732=>"110100100",
  4733=>"001000000",
  4734=>"111111111",
  4735=>"111111111",
  4736=>"111111111",
  4737=>"100100100",
  4738=>"111111110",
  4739=>"010000011",
  4740=>"000000000",
  4741=>"111000000",
  4742=>"111111111",
  4743=>"111111111",
  4744=>"111111111",
  4745=>"000000000",
  4746=>"100111111",
  4747=>"000000000",
  4748=>"000000000",
  4749=>"001111111",
  4750=>"001011111",
  4751=>"111111000",
  4752=>"000000000",
  4753=>"111111111",
  4754=>"100100111",
  4755=>"001001000",
  4756=>"000000000",
  4757=>"000010111",
  4758=>"011001000",
  4759=>"111111000",
  4760=>"000000111",
  4761=>"111111110",
  4762=>"000000000",
  4763=>"000000001",
  4764=>"000111111",
  4765=>"001000110",
  4766=>"001001000",
  4767=>"000000001",
  4768=>"101101111",
  4769=>"111111111",
  4770=>"111111000",
  4771=>"111111111",
  4772=>"000000001",
  4773=>"000000000",
  4774=>"000000000",
  4775=>"010111111",
  4776=>"111111111",
  4777=>"000000000",
  4778=>"000000000",
  4779=>"001000100",
  4780=>"101111011",
  4781=>"111001111",
  4782=>"000000000",
  4783=>"111111000",
  4784=>"000010000",
  4785=>"111101001",
  4786=>"111111110",
  4787=>"000111110",
  4788=>"001001111",
  4789=>"111111100",
  4790=>"111100000",
  4791=>"001111111",
  4792=>"111111111",
  4793=>"000000111",
  4794=>"111111111",
  4795=>"001000001",
  4796=>"000010110",
  4797=>"111111001",
  4798=>"000110110",
  4799=>"000000100",
  4800=>"111111111",
  4801=>"011111000",
  4802=>"111101101",
  4803=>"110111111",
  4804=>"000110110",
  4805=>"000000000",
  4806=>"000000000",
  4807=>"001000000",
  4808=>"001011011",
  4809=>"111000000",
  4810=>"000100000",
  4811=>"001000000",
  4812=>"100111000",
  4813=>"111111001",
  4814=>"111111111",
  4815=>"111111111",
  4816=>"111000000",
  4817=>"001001111",
  4818=>"111111110",
  4819=>"001100110",
  4820=>"111001000",
  4821=>"001000001",
  4822=>"000001111",
  4823=>"110000000",
  4824=>"000000000",
  4825=>"101011000",
  4826=>"110100111",
  4827=>"000000000",
  4828=>"111101111",
  4829=>"111111000",
  4830=>"000000001",
  4831=>"100000000",
  4832=>"000000000",
  4833=>"000011111",
  4834=>"001000000",
  4835=>"111111111",
  4836=>"000001000",
  4837=>"000000000",
  4838=>"111111110",
  4839=>"110101001",
  4840=>"111111111",
  4841=>"100110111",
  4842=>"000000110",
  4843=>"000000000",
  4844=>"001000000",
  4845=>"001000000",
  4846=>"000000000",
  4847=>"111011000",
  4848=>"011000000",
  4849=>"100000000",
  4850=>"011111111",
  4851=>"101000000",
  4852=>"000111111",
  4853=>"101100100",
  4854=>"001001101",
  4855=>"000000110",
  4856=>"000000000",
  4857=>"100100111",
  4858=>"111100110",
  4859=>"101111111",
  4860=>"111010000",
  4861=>"001001011",
  4862=>"111111111",
  4863=>"000000111",
  4864=>"000000000",
  4865=>"001111011",
  4866=>"000000001",
  4867=>"101101111",
  4868=>"110010011",
  4869=>"000111111",
  4870=>"000000111",
  4871=>"100110010",
  4872=>"100100000",
  4873=>"000000100",
  4874=>"110000100",
  4875=>"111111001",
  4876=>"000000100",
  4877=>"100000000",
  4878=>"111111000",
  4879=>"111111111",
  4880=>"000010001",
  4881=>"110111111",
  4882=>"110100000",
  4883=>"111101100",
  4884=>"011001111",
  4885=>"000110100",
  4886=>"011011011",
  4887=>"000000111",
  4888=>"111111111",
  4889=>"111111111",
  4890=>"111111000",
  4891=>"001001001",
  4892=>"001001001",
  4893=>"000000101",
  4894=>"111111100",
  4895=>"111110000",
  4896=>"111000111",
  4897=>"000101001",
  4898=>"111111111",
  4899=>"110111010",
  4900=>"111111111",
  4901=>"000000000",
  4902=>"100100000",
  4903=>"011000000",
  4904=>"000100111",
  4905=>"110111000",
  4906=>"101011000",
  4907=>"111111111",
  4908=>"110110010",
  4909=>"111111011",
  4910=>"101110000",
  4911=>"000000000",
  4912=>"011011000",
  4913=>"111111000",
  4914=>"011000000",
  4915=>"000000000",
  4916=>"000000000",
  4917=>"101111010",
  4918=>"000000000",
  4919=>"101111111",
  4920=>"110111100",
  4921=>"001000000",
  4922=>"011000000",
  4923=>"001010001",
  4924=>"111011111",
  4925=>"100100000",
  4926=>"111111100",
  4927=>"111010000",
  4928=>"000000000",
  4929=>"000000111",
  4930=>"001001000",
  4931=>"000000000",
  4932=>"111010110",
  4933=>"110111111",
  4934=>"001101111",
  4935=>"000000000",
  4936=>"011010011",
  4937=>"000000000",
  4938=>"001001000",
  4939=>"000000000",
  4940=>"111111101",
  4941=>"111111111",
  4942=>"000000111",
  4943=>"100100100",
  4944=>"111110000",
  4945=>"000000001",
  4946=>"100000000",
  4947=>"000000000",
  4948=>"111100000",
  4949=>"001001011",
  4950=>"111111111",
  4951=>"111011011",
  4952=>"001011011",
  4953=>"000100000",
  4954=>"101000111",
  4955=>"111110111",
  4956=>"111001111",
  4957=>"111111111",
  4958=>"111000000",
  4959=>"000001001",
  4960=>"000000001",
  4961=>"001001001",
  4962=>"000000000",
  4963=>"111111111",
  4964=>"110110010",
  4965=>"000000000",
  4966=>"111111001",
  4967=>"000000000",
  4968=>"001000001",
  4969=>"000100111",
  4970=>"101111000",
  4971=>"111111111",
  4972=>"101111010",
  4973=>"111000000",
  4974=>"111111111",
  4975=>"111111100",
  4976=>"101000010",
  4977=>"000000000",
  4978=>"110110111",
  4979=>"011011111",
  4980=>"000000000",
  4981=>"000000000",
  4982=>"101000001",
  4983=>"001000000",
  4984=>"000000000",
  4985=>"000000000",
  4986=>"111001001",
  4987=>"111111111",
  4988=>"111111111",
  4989=>"000000000",
  4990=>"111101111",
  4991=>"000000000",
  4992=>"110000000",
  4993=>"111111010",
  4994=>"111111111",
  4995=>"100110111",
  4996=>"000000000",
  4997=>"110110000",
  4998=>"011000000",
  4999=>"100100100",
  5000=>"111000000",
  5001=>"111100000",
  5002=>"001100000",
  5003=>"101001000",
  5004=>"001000000",
  5005=>"100011001",
  5006=>"111001000",
  5007=>"001111111",
  5008=>"010011001",
  5009=>"011111111",
  5010=>"111111000",
  5011=>"110111111",
  5012=>"000000000",
  5013=>"000000000",
  5014=>"000000011",
  5015=>"100000011",
  5016=>"110111111",
  5017=>"000000000",
  5018=>"111100110",
  5019=>"000000000",
  5020=>"000000100",
  5021=>"001111111",
  5022=>"001111001",
  5023=>"111111001",
  5024=>"111111111",
  5025=>"000001001",
  5026=>"111111011",
  5027=>"111001000",
  5028=>"111111010",
  5029=>"000111111",
  5030=>"100010010",
  5031=>"111111111",
  5032=>"000000101",
  5033=>"110110000",
  5034=>"000000000",
  5035=>"110100111",
  5036=>"000000000",
  5037=>"000000011",
  5038=>"111111110",
  5039=>"111111111",
  5040=>"000000000",
  5041=>"111111111",
  5042=>"111111111",
  5043=>"111111111",
  5044=>"000000110",
  5045=>"111111010",
  5046=>"111111000",
  5047=>"001001100",
  5048=>"111111101",
  5049=>"000111111",
  5050=>"000000000",
  5051=>"110110111",
  5052=>"001111111",
  5053=>"111111111",
  5054=>"001000000",
  5055=>"111010010",
  5056=>"000111111",
  5057=>"000000000",
  5058=>"111111111",
  5059=>"110100000",
  5060=>"000010000",
  5061=>"100110110",
  5062=>"110110010",
  5063=>"000000001",
  5064=>"101000000",
  5065=>"000000000",
  5066=>"110111011",
  5067=>"111111000",
  5068=>"000000000",
  5069=>"000000001",
  5070=>"000000000",
  5071=>"110111111",
  5072=>"001001011",
  5073=>"001100101",
  5074=>"111110111",
  5075=>"111111111",
  5076=>"000000000",
  5077=>"000000000",
  5078=>"000000000",
  5079=>"110110110",
  5080=>"000000001",
  5081=>"001100111",
  5082=>"000000000",
  5083=>"000000000",
  5084=>"000000000",
  5085=>"000000111",
  5086=>"000000000",
  5087=>"001001001",
  5088=>"000100110",
  5089=>"000000000",
  5090=>"011111111",
  5091=>"000000000",
  5092=>"000101111",
  5093=>"001001111",
  5094=>"111010110",
  5095=>"111111111",
  5096=>"000101001",
  5097=>"000100111",
  5098=>"111110111",
  5099=>"111111111",
  5100=>"011000110",
  5101=>"111111001",
  5102=>"111111011",
  5103=>"101111011",
  5104=>"111111001",
  5105=>"011001000",
  5106=>"110110111",
  5107=>"010000000",
  5108=>"111111111",
  5109=>"011000000",
  5110=>"110111111",
  5111=>"111111111",
  5112=>"111111111",
  5113=>"110110110",
  5114=>"111111011",
  5115=>"111110111",
  5116=>"111111111",
  5117=>"111111010",
  5118=>"001111111",
  5119=>"000000110",
  5120=>"111110110",
  5121=>"011000000",
  5122=>"000000111",
  5123=>"111110000",
  5124=>"100100100",
  5125=>"000000001",
  5126=>"000000000",
  5127=>"111100111",
  5128=>"000000010",
  5129=>"000011000",
  5130=>"110100000",
  5131=>"110000000",
  5132=>"000000000",
  5133=>"001001111",
  5134=>"111100100",
  5135=>"000110111",
  5136=>"110000111",
  5137=>"000000000",
  5138=>"010111100",
  5139=>"110111111",
  5140=>"101100000",
  5141=>"000000111",
  5142=>"000001001",
  5143=>"000000100",
  5144=>"100110110",
  5145=>"000000001",
  5146=>"000110111",
  5147=>"111011110",
  5148=>"000000000",
  5149=>"111111111",
  5150=>"111111111",
  5151=>"111111111",
  5152=>"111111000",
  5153=>"111111111",
  5154=>"000100111",
  5155=>"111100100",
  5156=>"000000000",
  5157=>"000000000",
  5158=>"000110111",
  5159=>"100101000",
  5160=>"000000001",
  5161=>"111101001",
  5162=>"111111111",
  5163=>"000000110",
  5164=>"000000000",
  5165=>"000000000",
  5166=>"111111001",
  5167=>"001000000",
  5168=>"000000000",
  5169=>"000000000",
  5170=>"100100000",
  5171=>"000111110",
  5172=>"000000000",
  5173=>"000000000",
  5174=>"001001100",
  5175=>"000000101",
  5176=>"001000000",
  5177=>"011001001",
  5178=>"110000000",
  5179=>"000000000",
  5180=>"111000111",
  5181=>"111101111",
  5182=>"001101111",
  5183=>"000000000",
  5184=>"000000001",
  5185=>"011001000",
  5186=>"110000000",
  5187=>"000000000",
  5188=>"010000000",
  5189=>"111110111",
  5190=>"111000111",
  5191=>"111000000",
  5192=>"110110110",
  5193=>"111111100",
  5194=>"101000111",
  5195=>"111101100",
  5196=>"111011000",
  5197=>"000000000",
  5198=>"000000000",
  5199=>"111111111",
  5200=>"001000000",
  5201=>"001000001",
  5202=>"000000111",
  5203=>"100000000",
  5204=>"000000111",
  5205=>"000000000",
  5206=>"000000001",
  5207=>"011011011",
  5208=>"111001000",
  5209=>"111100000",
  5210=>"111111111",
  5211=>"111100001",
  5212=>"000000000",
  5213=>"111111111",
  5214=>"110111111",
  5215=>"111111111",
  5216=>"111100000",
  5217=>"000000000",
  5218=>"000000111",
  5219=>"000100111",
  5220=>"000000000",
  5221=>"111111110",
  5222=>"011011111",
  5223=>"000000000",
  5224=>"000111111",
  5225=>"001000000",
  5226=>"111000000",
  5227=>"000111111",
  5228=>"101001011",
  5229=>"110110110",
  5230=>"111001000",
  5231=>"000000001",
  5232=>"111111111",
  5233=>"000000000",
  5234=>"111111001",
  5235=>"011111110",
  5236=>"000000000",
  5237=>"000000000",
  5238=>"101111000",
  5239=>"011011100",
  5240=>"111010110",
  5241=>"000000000",
  5242=>"000010000",
  5243=>"110010011",
  5244=>"110100100",
  5245=>"111111111",
  5246=>"000000000",
  5247=>"110010000",
  5248=>"000000011",
  5249=>"000000000",
  5250=>"111111111",
  5251=>"111000000",
  5252=>"111111111",
  5253=>"111111001",
  5254=>"100110110",
  5255=>"011011010",
  5256=>"000000100",
  5257=>"000011001",
  5258=>"111000000",
  5259=>"101111100",
  5260=>"101001111",
  5261=>"000000111",
  5262=>"001101001",
  5263=>"000111110",
  5264=>"000000011",
  5265=>"111100000",
  5266=>"011111111",
  5267=>"110111010",
  5268=>"011111111",
  5269=>"000110111",
  5270=>"000110110",
  5271=>"010000111",
  5272=>"100100000",
  5273=>"101100101",
  5274=>"100111111",
  5275=>"000000000",
  5276=>"110101101",
  5277=>"011011011",
  5278=>"111111011",
  5279=>"111111111",
  5280=>"111001001",
  5281=>"111000000",
  5282=>"000011000",
  5283=>"111000000",
  5284=>"000010000",
  5285=>"110110000",
  5286=>"000000000",
  5287=>"111111001",
  5288=>"001001111",
  5289=>"000000000",
  5290=>"111111000",
  5291=>"011001000",
  5292=>"111111011",
  5293=>"011001101",
  5294=>"111101111",
  5295=>"110110000",
  5296=>"000110110",
  5297=>"110110100",
  5298=>"110111111",
  5299=>"000000101",
  5300=>"010111100",
  5301=>"111111000",
  5302=>"000000000",
  5303=>"011001111",
  5304=>"111101100",
  5305=>"111111111",
  5306=>"010111111",
  5307=>"111100000",
  5308=>"110110111",
  5309=>"101100000",
  5310=>"111001001",
  5311=>"000000000",
  5312=>"110011111",
  5313=>"111011001",
  5314=>"111001001",
  5315=>"010111111",
  5316=>"000111000",
  5317=>"000111111",
  5318=>"000001001",
  5319=>"111111111",
  5320=>"000000000",
  5321=>"000000001",
  5322=>"011011011",
  5323=>"111111111",
  5324=>"110110100",
  5325=>"000111001",
  5326=>"110110101",
  5327=>"000000000",
  5328=>"000011111",
  5329=>"000000111",
  5330=>"000110110",
  5331=>"100000000",
  5332=>"000000100",
  5333=>"100110110",
  5334=>"000000000",
  5335=>"110111111",
  5336=>"111001000",
  5337=>"111101101",
  5338=>"001001001",
  5339=>"111100100",
  5340=>"111001101",
  5341=>"000110110",
  5342=>"000111110",
  5343=>"111111111",
  5344=>"111111111",
  5345=>"000111111",
  5346=>"000000000",
  5347=>"111101000",
  5348=>"110100100",
  5349=>"110100100",
  5350=>"100100111",
  5351=>"111111111",
  5352=>"001011011",
  5353=>"010000010",
  5354=>"100100111",
  5355=>"110110111",
  5356=>"001011001",
  5357=>"000000000",
  5358=>"000110110",
  5359=>"000000111",
  5360=>"000000000",
  5361=>"000000000",
  5362=>"110100000",
  5363=>"001000000",
  5364=>"111111111",
  5365=>"111111111",
  5366=>"111111110",
  5367=>"001000000",
  5368=>"111111111",
  5369=>"000111111",
  5370=>"000000000",
  5371=>"000001111",
  5372=>"111001011",
  5373=>"001001111",
  5374=>"000000000",
  5375=>"110110110",
  5376=>"111000000",
  5377=>"001000000",
  5378=>"100000000",
  5379=>"001000000",
  5380=>"110110101",
  5381=>"011011001",
  5382=>"111111111",
  5383=>"111010000",
  5384=>"111101001",
  5385=>"000100110",
  5386=>"111111111",
  5387=>"111111110",
  5388=>"111111001",
  5389=>"111111111",
  5390=>"100000000",
  5391=>"000010010",
  5392=>"111111111",
  5393=>"011011001",
  5394=>"011000000",
  5395=>"000000000",
  5396=>"000110111",
  5397=>"000000111",
  5398=>"110111111",
  5399=>"100000111",
  5400=>"100001111",
  5401=>"000000000",
  5402=>"111111110",
  5403=>"100000100",
  5404=>"000001000",
  5405=>"000000000",
  5406=>"111111111",
  5407=>"010111111",
  5408=>"000000001",
  5409=>"111001001",
  5410=>"111111111",
  5411=>"100101111",
  5412=>"111111111",
  5413=>"111111111",
  5414=>"111111011",
  5415=>"111110110",
  5416=>"111010111",
  5417=>"110000100",
  5418=>"111001111",
  5419=>"111100111",
  5420=>"111111111",
  5421=>"000000011",
  5422=>"000000000",
  5423=>"000100110",
  5424=>"000001010",
  5425=>"000000000",
  5426=>"000000000",
  5427=>"000000000",
  5428=>"000000100",
  5429=>"111111111",
  5430=>"000100000",
  5431=>"111111111",
  5432=>"000011000",
  5433=>"110000111",
  5434=>"000000000",
  5435=>"000000000",
  5436=>"111111111",
  5437=>"000000110",
  5438=>"000000000",
  5439=>"110111111",
  5440=>"000000000",
  5441=>"000000000",
  5442=>"110000000",
  5443=>"011111010",
  5444=>"000000111",
  5445=>"000000000",
  5446=>"000000000",
  5447=>"111111001",
  5448=>"111111000",
  5449=>"110000000",
  5450=>"000000000",
  5451=>"000000000",
  5452=>"000000000",
  5453=>"111101000",
  5454=>"111100111",
  5455=>"100100001",
  5456=>"100100100",
  5457=>"101100111",
  5458=>"100000000",
  5459=>"000000010",
  5460=>"000000000",
  5461=>"011001001",
  5462=>"111000000",
  5463=>"111111111",
  5464=>"111000000",
  5465=>"000000000",
  5466=>"000000000",
  5467=>"101100100",
  5468=>"000000111",
  5469=>"000001111",
  5470=>"111000000",
  5471=>"111101111",
  5472=>"111111000",
  5473=>"110111111",
  5474=>"111111111",
  5475=>"111000000",
  5476=>"000011111",
  5477=>"000011111",
  5478=>"111111001",
  5479=>"001101101",
  5480=>"000000001",
  5481=>"000000100",
  5482=>"111111110",
  5483=>"110000111",
  5484=>"110011111",
  5485=>"111011000",
  5486=>"100000000",
  5487=>"000000000",
  5488=>"011000000",
  5489=>"000001010",
  5490=>"010010000",
  5491=>"000000000",
  5492=>"100110111",
  5493=>"111111111",
  5494=>"000000111",
  5495=>"110111111",
  5496=>"111100000",
  5497=>"000010011",
  5498=>"111111111",
  5499=>"000001011",
  5500=>"001101111",
  5501=>"100100111",
  5502=>"111111111",
  5503=>"111000000",
  5504=>"000000100",
  5505=>"000000000",
  5506=>"111111111",
  5507=>"111111011",
  5508=>"000000000",
  5509=>"111111101",
  5510=>"111111110",
  5511=>"000000011",
  5512=>"010111111",
  5513=>"000000000",
  5514=>"110000000",
  5515=>"000011000",
  5516=>"111111001",
  5517=>"111111000",
  5518=>"100000000",
  5519=>"110111000",
  5520=>"000000000",
  5521=>"100100100",
  5522=>"100110000",
  5523=>"111111111",
  5524=>"111101100",
  5525=>"000000000",
  5526=>"111111111",
  5527=>"111110100",
  5528=>"000000111",
  5529=>"111010000",
  5530=>"100000000",
  5531=>"111111100",
  5532=>"100100110",
  5533=>"000001000",
  5534=>"000001000",
  5535=>"000000000",
  5536=>"100110110",
  5537=>"000000111",
  5538=>"001000001",
  5539=>"111111111",
  5540=>"100101101",
  5541=>"100111010",
  5542=>"000000111",
  5543=>"010000000",
  5544=>"000000101",
  5545=>"000111111",
  5546=>"111111100",
  5547=>"011000100",
  5548=>"000000000",
  5549=>"111111011",
  5550=>"111111111",
  5551=>"000000000",
  5552=>"000000001",
  5553=>"111111000",
  5554=>"000110010",
  5555=>"110111111",
  5556=>"101101000",
  5557=>"111100001",
  5558=>"101101111",
  5559=>"000000110",
  5560=>"011111000",
  5561=>"000111111",
  5562=>"111111111",
  5563=>"111100111",
  5564=>"000111111",
  5565=>"111111111",
  5566=>"000111111",
  5567=>"101100001",
  5568=>"001101000",
  5569=>"111111111",
  5570=>"100000000",
  5571=>"000111111",
  5572=>"001000000",
  5573=>"100000000",
  5574=>"010000000",
  5575=>"000000111",
  5576=>"111100100",
  5577=>"100110110",
  5578=>"000000000",
  5579=>"111111111",
  5580=>"000000000",
  5581=>"000000000",
  5582=>"111110000",
  5583=>"111111111",
  5584=>"000000000",
  5585=>"000000111",
  5586=>"001000000",
  5587=>"111000000",
  5588=>"111110111",
  5589=>"111101100",
  5590=>"000111000",
  5591=>"001001011",
  5592=>"111100100",
  5593=>"111000101",
  5594=>"000000111",
  5595=>"000000000",
  5596=>"011111101",
  5597=>"111111101",
  5598=>"000000111",
  5599=>"111111000",
  5600=>"001000111",
  5601=>"111000000",
  5602=>"000110111",
  5603=>"111111000",
  5604=>"111110000",
  5605=>"000000000",
  5606=>"000000000",
  5607=>"000000000",
  5608=>"101000000",
  5609=>"111001001",
  5610=>"011000001",
  5611=>"000000000",
  5612=>"000000100",
  5613=>"000110011",
  5614=>"000000011",
  5615=>"000000000",
  5616=>"000000000",
  5617=>"111111111",
  5618=>"111111111",
  5619=>"111111000",
  5620=>"111111000",
  5621=>"111100000",
  5622=>"000000010",
  5623=>"100110011",
  5624=>"000000111",
  5625=>"110110100",
  5626=>"000110110",
  5627=>"000111111",
  5628=>"011011011",
  5629=>"110000000",
  5630=>"111111111",
  5631=>"000110100",
  5632=>"100000000",
  5633=>"000000111",
  5634=>"111000111",
  5635=>"110001000",
  5636=>"111111111",
  5637=>"010001001",
  5638=>"111111110",
  5639=>"000001001",
  5640=>"001001111",
  5641=>"011011111",
  5642=>"100110111",
  5643=>"111111111",
  5644=>"110111110",
  5645=>"000000000",
  5646=>"000000000",
  5647=>"101101101",
  5648=>"000110111",
  5649=>"111011000",
  5650=>"010110010",
  5651=>"111111011",
  5652=>"000000000",
  5653=>"100000100",
  5654=>"000111110",
  5655=>"001001001",
  5656=>"000000000",
  5657=>"100100000",
  5658=>"000101011",
  5659=>"011011011",
  5660=>"111111000",
  5661=>"000010111",
  5662=>"000000001",
  5663=>"000000110",
  5664=>"111111111",
  5665=>"000110111",
  5666=>"101100000",
  5667=>"000000111",
  5668=>"111111000",
  5669=>"111101101",
  5670=>"110000001",
  5671=>"000010010",
  5672=>"110111110",
  5673=>"100100111",
  5674=>"111111111",
  5675=>"111111000",
  5676=>"001011111",
  5677=>"000110110",
  5678=>"000000100",
  5679=>"000000001",
  5680=>"101111101",
  5681=>"111100000",
  5682=>"111111111",
  5683=>"100110010",
  5684=>"100000100",
  5685=>"001001001",
  5686=>"101001001",
  5687=>"000000000",
  5688=>"100000111",
  5689=>"000000000",
  5690=>"111111111",
  5691=>"001001111",
  5692=>"101101111",
  5693=>"111001001",
  5694=>"001011111",
  5695=>"001111111",
  5696=>"110110111",
  5697=>"000000110",
  5698=>"000000101",
  5699=>"000110111",
  5700=>"111000001",
  5701=>"001001001",
  5702=>"011111111",
  5703=>"110000010",
  5704=>"001001011",
  5705=>"000000100",
  5706=>"000011011",
  5707=>"000000000",
  5708=>"101000101",
  5709=>"000000100",
  5710=>"000000001",
  5711=>"111111110",
  5712=>"000000000",
  5713=>"000000000",
  5714=>"111111111",
  5715=>"000000000",
  5716=>"000101111",
  5717=>"111111110",
  5718=>"101101100",
  5719=>"001001101",
  5720=>"101000000",
  5721=>"001101111",
  5722=>"000010000",
  5723=>"100100100",
  5724=>"000000000",
  5725=>"111111101",
  5726=>"000010000",
  5727=>"010000110",
  5728=>"010000010",
  5729=>"111111011",
  5730=>"111011011",
  5731=>"101001001",
  5732=>"110010000",
  5733=>"111000000",
  5734=>"010000000",
  5735=>"001000001",
  5736=>"111111111",
  5737=>"000000101",
  5738=>"000011111",
  5739=>"000000010",
  5740=>"000100100",
  5741=>"111111110",
  5742=>"111101001",
  5743=>"000000000",
  5744=>"000000001",
  5745=>"000000111",
  5746=>"100000101",
  5747=>"000000000",
  5748=>"111111010",
  5749=>"110100100",
  5750=>"111111111",
  5751=>"001000101",
  5752=>"111110000",
  5753=>"000011011",
  5754=>"010000000",
  5755=>"001001001",
  5756=>"001111101",
  5757=>"001000111",
  5758=>"110100110",
  5759=>"000110111",
  5760=>"111101000",
  5761=>"100000111",
  5762=>"100111100",
  5763=>"000011001",
  5764=>"111101000",
  5765=>"110111110",
  5766=>"111001011",
  5767=>"000000000",
  5768=>"000000000",
  5769=>"001011111",
  5770=>"101111111",
  5771=>"001011111",
  5772=>"111111101",
  5773=>"101111111",
  5774=>"110111011",
  5775=>"111111100",
  5776=>"000001101",
  5777=>"000000100",
  5778=>"111100000",
  5779=>"111000110",
  5780=>"101000100",
  5781=>"101001111",
  5782=>"000000100",
  5783=>"001001100",
  5784=>"001001001",
  5785=>"001000101",
  5786=>"111010111",
  5787=>"111111111",
  5788=>"011000111",
  5789=>"110000000",
  5790=>"110110010",
  5791=>"101000101",
  5792=>"000010111",
  5793=>"001001111",
  5794=>"101111111",
  5795=>"111010111",
  5796=>"000110011",
  5797=>"000000001",
  5798=>"111111111",
  5799=>"100100100",
  5800=>"000111011",
  5801=>"111111111",
  5802=>"001001001",
  5803=>"000000100",
  5804=>"011111111",
  5805=>"010011011",
  5806=>"111111010",
  5807=>"000000000",
  5808=>"011111111",
  5809=>"011001101",
  5810=>"110111110",
  5811=>"111111111",
  5812=>"110010011",
  5813=>"000100100",
  5814=>"101111111",
  5815=>"111111111",
  5816=>"000000000",
  5817=>"010111111",
  5818=>"000001000",
  5819=>"111111111",
  5820=>"111111111",
  5821=>"000000000",
  5822=>"000000100",
  5823=>"000100100",
  5824=>"111111111",
  5825=>"001000101",
  5826=>"000101111",
  5827=>"111111111",
  5828=>"000000001",
  5829=>"000000100",
  5830=>"111110000",
  5831=>"000000100",
  5832=>"111111111",
  5833=>"001001111",
  5834=>"101111111",
  5835=>"100000101",
  5836=>"011010000",
  5837=>"000000100",
  5838=>"000000010",
  5839=>"011011111",
  5840=>"100000000",
  5841=>"000001001",
  5842=>"000000000",
  5843=>"101001111",
  5844=>"100100101",
  5845=>"111111011",
  5846=>"000000000",
  5847=>"000101001",
  5848=>"000000111",
  5849=>"110101000",
  5850=>"000000000",
  5851=>"000001011",
  5852=>"111111011",
  5853=>"000000111",
  5854=>"000000100",
  5855=>"001000101",
  5856=>"111111010",
  5857=>"010010010",
  5858=>"011111000",
  5859=>"000011111",
  5860=>"101000110",
  5861=>"001111011",
  5862=>"110111010",
  5863=>"101111111",
  5864=>"000101000",
  5865=>"111110100",
  5866=>"110100100",
  5867=>"000000101",
  5868=>"111110000",
  5869=>"011001000",
  5870=>"000000001",
  5871=>"111111111",
  5872=>"001000000",
  5873=>"000000110",
  5874=>"010010000",
  5875=>"000000100",
  5876=>"011001111",
  5877=>"000000100",
  5878=>"111001011",
  5879=>"111111000",
  5880=>"111101000",
  5881=>"111111111",
  5882=>"001111111",
  5883=>"100000000",
  5884=>"001001101",
  5885=>"011001010",
  5886=>"011011001",
  5887=>"000000101",
  5888=>"100110111",
  5889=>"100100101",
  5890=>"000110111",
  5891=>"100110000",
  5892=>"111000101",
  5893=>"110111101",
  5894=>"000010111",
  5895=>"111010001",
  5896=>"111011000",
  5897=>"000000000",
  5898=>"001000101",
  5899=>"011001111",
  5900=>"000000001",
  5901=>"000110000",
  5902=>"111111111",
  5903=>"100100110",
  5904=>"111000100",
  5905=>"101110101",
  5906=>"000001001",
  5907=>"111111111",
  5908=>"111111011",
  5909=>"111111111",
  5910=>"100100110",
  5911=>"101001110",
  5912=>"001001001",
  5913=>"000000000",
  5914=>"000000011",
  5915=>"000011111",
  5916=>"000000111",
  5917=>"101000101",
  5918=>"000110000",
  5919=>"000000110",
  5920=>"000000000",
  5921=>"000000000",
  5922=>"000000000",
  5923=>"100111001",
  5924=>"001111110",
  5925=>"000000000",
  5926=>"001000101",
  5927=>"111011000",
  5928=>"110000100",
  5929=>"101001111",
  5930=>"000011100",
  5931=>"000000000",
  5932=>"011011111",
  5933=>"000000100",
  5934=>"111111000",
  5935=>"000000111",
  5936=>"000000000",
  5937=>"110011000",
  5938=>"101100100",
  5939=>"100111011",
  5940=>"100000000",
  5941=>"000000100",
  5942=>"000010100",
  5943=>"000111111",
  5944=>"010010000",
  5945=>"000000100",
  5946=>"001000101",
  5947=>"110111100",
  5948=>"100100000",
  5949=>"111110000",
  5950=>"001000111",
  5951=>"111001111",
  5952=>"000000000",
  5953=>"111110001",
  5954=>"000001011",
  5955=>"000000000",
  5956=>"000001111",
  5957=>"100111111",
  5958=>"001010000",
  5959=>"110111000",
  5960=>"101111111",
  5961=>"011000111",
  5962=>"000000000",
  5963=>"100101111",
  5964=>"110111000",
  5965=>"000000001",
  5966=>"111011111",
  5967=>"001001001",
  5968=>"001001011",
  5969=>"000000000",
  5970=>"101101101",
  5971=>"111111111",
  5972=>"101000111",
  5973=>"011111111",
  5974=>"101001101",
  5975=>"111111101",
  5976=>"110101001",
  5977=>"001101111",
  5978=>"111110111",
  5979=>"000101111",
  5980=>"110111111",
  5981=>"000000111",
  5982=>"110010010",
  5983=>"001000110",
  5984=>"111001001",
  5985=>"101101101",
  5986=>"000000111",
  5987=>"111111001",
  5988=>"001100000",
  5989=>"000000001",
  5990=>"000000000",
  5991=>"111111010",
  5992=>"001001011",
  5993=>"010110110",
  5994=>"111100100",
  5995=>"110110100",
  5996=>"010001011",
  5997=>"000111000",
  5998=>"101101111",
  5999=>"000001101",
  6000=>"111100111",
  6001=>"001111111",
  6002=>"000000100",
  6003=>"111111110",
  6004=>"111111101",
  6005=>"111101110",
  6006=>"000100100",
  6007=>"000010011",
  6008=>"101101101",
  6009=>"100000111",
  6010=>"000000101",
  6011=>"100000100",
  6012=>"011111111",
  6013=>"111010000",
  6014=>"111111011",
  6015=>"000000101",
  6016=>"111111001",
  6017=>"110111111",
  6018=>"000000000",
  6019=>"000000001",
  6020=>"111001000",
  6021=>"000000000",
  6022=>"000000100",
  6023=>"101110001",
  6024=>"111111111",
  6025=>"011111111",
  6026=>"011000111",
  6027=>"000000000",
  6028=>"001001111",
  6029=>"100100000",
  6030=>"001011001",
  6031=>"000000000",
  6032=>"111111111",
  6033=>"000000001",
  6034=>"000110000",
  6035=>"011001100",
  6036=>"000000010",
  6037=>"000000000",
  6038=>"111011011",
  6039=>"000000000",
  6040=>"111110111",
  6041=>"011111111",
  6042=>"101000000",
  6043=>"111111010",
  6044=>"000000000",
  6045=>"111111111",
  6046=>"000000100",
  6047=>"000000000",
  6048=>"000000111",
  6049=>"000000000",
  6050=>"000111111",
  6051=>"000000001",
  6052=>"010011010",
  6053=>"101101101",
  6054=>"111111001",
  6055=>"000100100",
  6056=>"000101000",
  6057=>"000000111",
  6058=>"111111010",
  6059=>"000110110",
  6060=>"111111111",
  6061=>"001010001",
  6062=>"000011111",
  6063=>"000101110",
  6064=>"111111111",
  6065=>"101110111",
  6066=>"100000101",
  6067=>"000000000",
  6068=>"001000000",
  6069=>"000001111",
  6070=>"110111010",
  6071=>"000111111",
  6072=>"000000011",
  6073=>"111101000",
  6074=>"101101111",
  6075=>"110110110",
  6076=>"000000000",
  6077=>"011000000",
  6078=>"110100110",
  6079=>"100100100",
  6080=>"000000000",
  6081=>"111111111",
  6082=>"000000111",
  6083=>"111111111",
  6084=>"101000000",
  6085=>"001111011",
  6086=>"000000111",
  6087=>"000110111",
  6088=>"000000100",
  6089=>"111111010",
  6090=>"000000001",
  6091=>"010111111",
  6092=>"010000000",
  6093=>"000000000",
  6094=>"001000000",
  6095=>"000000011",
  6096=>"000000000",
  6097=>"100111100",
  6098=>"111110110",
  6099=>"101111111",
  6100=>"110000000",
  6101=>"000000000",
  6102=>"000000010",
  6103=>"111111011",
  6104=>"000101010",
  6105=>"000000000",
  6106=>"101100100",
  6107=>"001001011",
  6108=>"011000000",
  6109=>"100100000",
  6110=>"111000111",
  6111=>"100100100",
  6112=>"000001001",
  6113=>"100100111",
  6114=>"000000000",
  6115=>"000000100",
  6116=>"000000101",
  6117=>"000100100",
  6118=>"001000001",
  6119=>"000000111",
  6120=>"000000000",
  6121=>"000000100",
  6122=>"001000000",
  6123=>"001100111",
  6124=>"000000111",
  6125=>"010011100",
  6126=>"001001011",
  6127=>"101001000",
  6128=>"111111000",
  6129=>"000000111",
  6130=>"001001101",
  6131=>"000000101",
  6132=>"110110010",
  6133=>"000000000",
  6134=>"011001001",
  6135=>"111011111",
  6136=>"111111110",
  6137=>"001001101",
  6138=>"110110000",
  6139=>"111111110",
  6140=>"100100000",
  6141=>"000000011",
  6142=>"000000001",
  6143=>"001101111",
  6144=>"111111111",
  6145=>"001001000",
  6146=>"001101101",
  6147=>"001111111",
  6148=>"111111010",
  6149=>"010010010",
  6150=>"000000000",
  6151=>"000000001",
  6152=>"111111011",
  6153=>"100000000",
  6154=>"000000000",
  6155=>"000000110",
  6156=>"000000010",
  6157=>"011011010",
  6158=>"000000000",
  6159=>"000000000",
  6160=>"111111111",
  6161=>"100000011",
  6162=>"000110111",
  6163=>"111111111",
  6164=>"000000000",
  6165=>"111111000",
  6166=>"001001001",
  6167=>"001000100",
  6168=>"001001001",
  6169=>"111111010",
  6170=>"011000111",
  6171=>"000100110",
  6172=>"000000001",
  6173=>"000100100",
  6174=>"011111111",
  6175=>"000111111",
  6176=>"100000000",
  6177=>"111111110",
  6178=>"100000000",
  6179=>"111111111",
  6180=>"111111101",
  6181=>"000000000",
  6182=>"000000111",
  6183=>"000111111",
  6184=>"011011010",
  6185=>"000000000",
  6186=>"000000000",
  6187=>"000000000",
  6188=>"100000000",
  6189=>"111111011",
  6190=>"010010000",
  6191=>"111000000",
  6192=>"111111001",
  6193=>"000000000",
  6194=>"010000000",
  6195=>"000000000",
  6196=>"111010110",
  6197=>"111101111",
  6198=>"111100111",
  6199=>"011110001",
  6200=>"000111101",
  6201=>"000000000",
  6202=>"000000000",
  6203=>"111111010",
  6204=>"000001001",
  6205=>"111101111",
  6206=>"100000000",
  6207=>"000000000",
  6208=>"110000000",
  6209=>"111111111",
  6210=>"011000110",
  6211=>"001011011",
  6212=>"000000000",
  6213=>"000000000",
  6214=>"000000000",
  6215=>"000000000",
  6216=>"000000100",
  6217=>"000000101",
  6218=>"000111110",
  6219=>"001011000",
  6220=>"011111111",
  6221=>"111111111",
  6222=>"010000000",
  6223=>"111111010",
  6224=>"111110000",
  6225=>"111111000",
  6226=>"111000001",
  6227=>"000000000",
  6228=>"010011111",
  6229=>"000011110",
  6230=>"000100010",
  6231=>"111111111",
  6232=>"100111111",
  6233=>"111101111",
  6234=>"000000001",
  6235=>"011110110",
  6236=>"000000000",
  6237=>"101111111",
  6238=>"000010000",
  6239=>"100000001",
  6240=>"100111111",
  6241=>"100000000",
  6242=>"111101000",
  6243=>"001001001",
  6244=>"011011101",
  6245=>"111111111",
  6246=>"000000110",
  6247=>"000101111",
  6248=>"001111111",
  6249=>"111111000",
  6250=>"001001100",
  6251=>"100101010",
  6252=>"000000110",
  6253=>"000000000",
  6254=>"110110100",
  6255=>"111111111",
  6256=>"000000000",
  6257=>"000110111",
  6258=>"111110111",
  6259=>"000000001",
  6260=>"101001111",
  6261=>"110111111",
  6262=>"110000000",
  6263=>"111111010",
  6264=>"000000000",
  6265=>"000000100",
  6266=>"001000001",
  6267=>"000110110",
  6268=>"111111111",
  6269=>"111111111",
  6270=>"010000001",
  6271=>"110111110",
  6272=>"111111111",
  6273=>"111111111",
  6274=>"000000100",
  6275=>"000000100",
  6276=>"111111111",
  6277=>"000000000",
  6278=>"101000000",
  6279=>"010111111",
  6280=>"100111111",
  6281=>"111111010",
  6282=>"111111000",
  6283=>"000000000",
  6284=>"111111111",
  6285=>"111111110",
  6286=>"010111111",
  6287=>"000000000",
  6288=>"110010000",
  6289=>"110111111",
  6290=>"111010000",
  6291=>"000000000",
  6292=>"111111011",
  6293=>"010100100",
  6294=>"000001001",
  6295=>"111111011",
  6296=>"111111101",
  6297=>"101101101",
  6298=>"000000000",
  6299=>"111111111",
  6300=>"111101000",
  6301=>"001000000",
  6302=>"111111111",
  6303=>"011001000",
  6304=>"000000000",
  6305=>"000000000",
  6306=>"000000100",
  6307=>"111111111",
  6308=>"111111111",
  6309=>"011011000",
  6310=>"111111111",
  6311=>"010111111",
  6312=>"011111111",
  6313=>"111111111",
  6314=>"111100100",
  6315=>"111111111",
  6316=>"111111011",
  6317=>"110110110",
  6318=>"100001001",
  6319=>"111011000",
  6320=>"000000000",
  6321=>"111111111",
  6322=>"111111111",
  6323=>"000000111",
  6324=>"111111111",
  6325=>"111001000",
  6326=>"111111111",
  6327=>"101111011",
  6328=>"000000001",
  6329=>"101001001",
  6330=>"101111000",
  6331=>"110000011",
  6332=>"111111000",
  6333=>"110110000",
  6334=>"001111111",
  6335=>"111111111",
  6336=>"000010000",
  6337=>"000000101",
  6338=>"000001001",
  6339=>"100000100",
  6340=>"110100110",
  6341=>"111111111",
  6342=>"111011000",
  6343=>"011110100",
  6344=>"000000001",
  6345=>"000000000",
  6346=>"111010110",
  6347=>"000000100",
  6348=>"011001000",
  6349=>"100111111",
  6350=>"111111111",
  6351=>"000111111",
  6352=>"001000100",
  6353=>"111100100",
  6354=>"011111110",
  6355=>"001000000",
  6356=>"111110100",
  6357=>"000000000",
  6358=>"111111111",
  6359=>"010111111",
  6360=>"001011001",
  6361=>"111111111",
  6362=>"000000000",
  6363=>"000000010",
  6364=>"111111111",
  6365=>"111000000",
  6366=>"111111111",
  6367=>"110110110",
  6368=>"000000010",
  6369=>"000000000",
  6370=>"101101001",
  6371=>"111111011",
  6372=>"111000000",
  6373=>"110111100",
  6374=>"111111111",
  6375=>"100111101",
  6376=>"111111000",
  6377=>"000000111",
  6378=>"111111101",
  6379=>"111001001",
  6380=>"111010000",
  6381=>"111110110",
  6382=>"111001000",
  6383=>"001000000",
  6384=>"000000000",
  6385=>"111000111",
  6386=>"000010110",
  6387=>"110010110",
  6388=>"000000000",
  6389=>"001001001",
  6390=>"011011100",
  6391=>"110000000",
  6392=>"000000000",
  6393=>"100100111",
  6394=>"000000000",
  6395=>"111111111",
  6396=>"100100000",
  6397=>"001001011",
  6398=>"000011011",
  6399=>"101111111",
  6400=>"110111111",
  6401=>"000000011",
  6402=>"101001000",
  6403=>"111111100",
  6404=>"111111111",
  6405=>"001011111",
  6406=>"011111111",
  6407=>"000000001",
  6408=>"111111111",
  6409=>"111111111",
  6410=>"000000001",
  6411=>"000000000",
  6412=>"001001111",
  6413=>"000000000",
  6414=>"111111001",
  6415=>"000000000",
  6416=>"000000000",
  6417=>"000000000",
  6418=>"111111110",
  6419=>"001000000",
  6420=>"000110111",
  6421=>"011000000",
  6422=>"011010000",
  6423=>"001001000",
  6424=>"010000000",
  6425=>"111000000",
  6426=>"000000111",
  6427=>"001000100",
  6428=>"000000000",
  6429=>"000001110",
  6430=>"000000111",
  6431=>"000000000",
  6432=>"000110110",
  6433=>"011000000",
  6434=>"010010110",
  6435=>"111010000",
  6436=>"001101101",
  6437=>"000100100",
  6438=>"111000000",
  6439=>"111111110",
  6440=>"111111100",
  6441=>"111111111",
  6442=>"010000010",
  6443=>"011011111",
  6444=>"000100111",
  6445=>"100110100",
  6446=>"000000111",
  6447=>"001111101",
  6448=>"000010010",
  6449=>"000000100",
  6450=>"000000101",
  6451=>"011011100",
  6452=>"000000001",
  6453=>"111111111",
  6454=>"111111000",
  6455=>"111010000",
  6456=>"110111111",
  6457=>"111100000",
  6458=>"000000000",
  6459=>"001000000",
  6460=>"110110110",
  6461=>"110110100",
  6462=>"111111000",
  6463=>"000000010",
  6464=>"111011001",
  6465=>"000001000",
  6466=>"000011111",
  6467=>"001001001",
  6468=>"100110100",
  6469=>"000010000",
  6470=>"100000000",
  6471=>"000000100",
  6472=>"100000000",
  6473=>"000000000",
  6474=>"000000000",
  6475=>"111010110",
  6476=>"000000000",
  6477=>"000000000",
  6478=>"000011111",
  6479=>"000000000",
  6480=>"110110111",
  6481=>"001101111",
  6482=>"001111111",
  6483=>"000000111",
  6484=>"000100111",
  6485=>"011111111",
  6486=>"000000111",
  6487=>"111111111",
  6488=>"110100000",
  6489=>"111101000",
  6490=>"000000000",
  6491=>"000011111",
  6492=>"111000000",
  6493=>"000000101",
  6494=>"001000100",
  6495=>"000100110",
  6496=>"000100111",
  6497=>"010000000",
  6498=>"110011011",
  6499=>"000000000",
  6500=>"100100110",
  6501=>"000000111",
  6502=>"000000111",
  6503=>"000000000",
  6504=>"110110110",
  6505=>"000101101",
  6506=>"001001000",
  6507=>"111100100",
  6508=>"001011000",
  6509=>"110110000",
  6510=>"000000000",
  6511=>"111011011",
  6512=>"111101100",
  6513=>"100111111",
  6514=>"000000111",
  6515=>"111111010",
  6516=>"111111111",
  6517=>"001001001",
  6518=>"000010111",
  6519=>"111111111",
  6520=>"111111111",
  6521=>"000000000",
  6522=>"000000000",
  6523=>"100000001",
  6524=>"100100110",
  6525=>"111100111",
  6526=>"000000000",
  6527=>"111111111",
  6528=>"000100100",
  6529=>"111001101",
  6530=>"001011011",
  6531=>"000000000",
  6532=>"111111111",
  6533=>"000001001",
  6534=>"000000110",
  6535=>"111110110",
  6536=>"000000000",
  6537=>"111111111",
  6538=>"111011000",
  6539=>"001001111",
  6540=>"101101101",
  6541=>"111111111",
  6542=>"000001011",
  6543=>"111111000",
  6544=>"111111111",
  6545=>"111111111",
  6546=>"110110110",
  6547=>"011111111",
  6548=>"000000000",
  6549=>"000010000",
  6550=>"111111111",
  6551=>"101111111",
  6552=>"011000011",
  6553=>"001011011",
  6554=>"000000100",
  6555=>"000000000",
  6556=>"100100000",
  6557=>"000110111",
  6558=>"000000000",
  6559=>"001000111",
  6560=>"001011111",
  6561=>"000011011",
  6562=>"000010000",
  6563=>"000000000",
  6564=>"000001001",
  6565=>"111111111",
  6566=>"111000111",
  6567=>"000010110",
  6568=>"101001000",
  6569=>"000100110",
  6570=>"000000000",
  6571=>"110100100",
  6572=>"101000000",
  6573=>"000000011",
  6574=>"111111001",
  6575=>"000000000",
  6576=>"111111000",
  6577=>"000000000",
  6578=>"111101000",
  6579=>"000000110",
  6580=>"000100110",
  6581=>"000000111",
  6582=>"000000000",
  6583=>"111001101",
  6584=>"011011000",
  6585=>"111000000",
  6586=>"100101111",
  6587=>"101100111",
  6588=>"111111000",
  6589=>"111101101",
  6590=>"010000000",
  6591=>"110100110",
  6592=>"000000000",
  6593=>"110000000",
  6594=>"000000000",
  6595=>"100100000",
  6596=>"000000000",
  6597=>"111111001",
  6598=>"010010111",
  6599=>"111111111",
  6600=>"111111111",
  6601=>"011111100",
  6602=>"111101000",
  6603=>"111000000",
  6604=>"000110111",
  6605=>"111111111",
  6606=>"000010110",
  6607=>"000000000",
  6608=>"001001001",
  6609=>"000000000",
  6610=>"000000001",
  6611=>"000100000",
  6612=>"000100111",
  6613=>"000111111",
  6614=>"000000000",
  6615=>"000001001",
  6616=>"110111001",
  6617=>"000000111",
  6618=>"000000000",
  6619=>"000000110",
  6620=>"111011000",
  6621=>"111111110",
  6622=>"111111110",
  6623=>"001101001",
  6624=>"111000000",
  6625=>"100111111",
  6626=>"000000000",
  6627=>"010000010",
  6628=>"001111101",
  6629=>"011011011",
  6630=>"011000001",
  6631=>"100110110",
  6632=>"110010000",
  6633=>"111111011",
  6634=>"001100101",
  6635=>"111011000",
  6636=>"001111111",
  6637=>"000000110",
  6638=>"111001000",
  6639=>"100000100",
  6640=>"110111110",
  6641=>"010110110",
  6642=>"000000000",
  6643=>"000000010",
  6644=>"000001100",
  6645=>"111000000",
  6646=>"111111111",
  6647=>"110110110",
  6648=>"110110000",
  6649=>"101101101",
  6650=>"111111001",
  6651=>"000000000",
  6652=>"101001111",
  6653=>"001101001",
  6654=>"001001010",
  6655=>"000110110",
  6656=>"111000010",
  6657=>"111000001",
  6658=>"101101111",
  6659=>"100110111",
  6660=>"111111111",
  6661=>"101101101",
  6662=>"001001001",
  6663=>"101101101",
  6664=>"000111111",
  6665=>"000000001",
  6666=>"110101000",
  6667=>"111111011",
  6668=>"111111111",
  6669=>"100101001",
  6670=>"111101101",
  6671=>"010110010",
  6672=>"111111111",
  6673=>"011011010",
  6674=>"011011110",
  6675=>"110111101",
  6676=>"011100100",
  6677=>"001000100",
  6678=>"000000000",
  6679=>"111111111",
  6680=>"111111111",
  6681=>"011010000",
  6682=>"010011001",
  6683=>"011111111",
  6684=>"101111111",
  6685=>"100000000",
  6686=>"001001111",
  6687=>"000000110",
  6688=>"000000000",
  6689=>"011011111",
  6690=>"110100111",
  6691=>"111110111",
  6692=>"000000000",
  6693=>"110111111",
  6694=>"000000000",
  6695=>"000010011",
  6696=>"101010010",
  6697=>"011010010",
  6698=>"011111111",
  6699=>"010011001",
  6700=>"100000000",
  6701=>"100110111",
  6702=>"000000001",
  6703=>"101100100",
  6704=>"001011011",
  6705=>"000000000",
  6706=>"111011001",
  6707=>"101111101",
  6708=>"000001111",
  6709=>"111111111",
  6710=>"001111111",
  6711=>"000000111",
  6712=>"101101000",
  6713=>"011001001",
  6714=>"000001111",
  6715=>"001000000",
  6716=>"100100111",
  6717=>"111111111",
  6718=>"110110110",
  6719=>"101000000",
  6720=>"101101001",
  6721=>"100101101",
  6722=>"000000010",
  6723=>"111101111",
  6724=>"110110110",
  6725=>"010011011",
  6726=>"000000100",
  6727=>"010000110",
  6728=>"111111111",
  6729=>"101101111",
  6730=>"000000001",
  6731=>"000010000",
  6732=>"110110110",
  6733=>"000010000",
  6734=>"111000011",
  6735=>"001000111",
  6736=>"011000010",
  6737=>"001001111",
  6738=>"010010010",
  6739=>"111110110",
  6740=>"001001000",
  6741=>"010010011",
  6742=>"001001001",
  6743=>"000101000",
  6744=>"001011000",
  6745=>"101100110",
  6746=>"100110111",
  6747=>"111111011",
  6748=>"100000000",
  6749=>"110111101",
  6750=>"001000000",
  6751=>"100000100",
  6752=>"001000110",
  6753=>"110110111",
  6754=>"000000101",
  6755=>"001101111",
  6756=>"111110111",
  6757=>"101111000",
  6758=>"111111110",
  6759=>"110100000",
  6760=>"111111111",
  6761=>"000000101",
  6762=>"110111100",
  6763=>"101101100",
  6764=>"011010110",
  6765=>"101000000",
  6766=>"111100111",
  6767=>"010010110",
  6768=>"000001000",
  6769=>"110110010",
  6770=>"011111001",
  6771=>"001000000",
  6772=>"000101101",
  6773=>"101111010",
  6774=>"110110000",
  6775=>"000000000",
  6776=>"010111111",
  6777=>"010111101",
  6778=>"101001000",
  6779=>"000000110",
  6780=>"111111111",
  6781=>"011111111",
  6782=>"011000000",
  6783=>"011011010",
  6784=>"010010010",
  6785=>"011001001",
  6786=>"001000000",
  6787=>"000010001",
  6788=>"101101101",
  6789=>"110110111",
  6790=>"011011110",
  6791=>"100101001",
  6792=>"000000000",
  6793=>"001101111",
  6794=>"001001101",
  6795=>"111111101",
  6796=>"001000000",
  6797=>"111111110",
  6798=>"110110010",
  6799=>"001011000",
  6800=>"000000011",
  6801=>"110110110",
  6802=>"100000000",
  6803=>"011001011",
  6804=>"100101101",
  6805=>"010011010",
  6806=>"000010110",
  6807=>"111111111",
  6808=>"001000000",
  6809=>"110111111",
  6810=>"111111011",
  6811=>"101101101",
  6812=>"000110100",
  6813=>"101001000",
  6814=>"000100100",
  6815=>"000101111",
  6816=>"000000000",
  6817=>"101100101",
  6818=>"001101111",
  6819=>"000000010",
  6820=>"001001001",
  6821=>"011111010",
  6822=>"110110110",
  6823=>"011111011",
  6824=>"111000110",
  6825=>"010010011",
  6826=>"001001000",
  6827=>"000110111",
  6828=>"111110010",
  6829=>"111001111",
  6830=>"101101111",
  6831=>"100001000",
  6832=>"000000000",
  6833=>"010011011",
  6834=>"010010010",
  6835=>"000001011",
  6836=>"111011000",
  6837=>"001000000",
  6838=>"010010010",
  6839=>"111111000",
  6840=>"101001011",
  6841=>"101000010",
  6842=>"001000101",
  6843=>"011000000",
  6844=>"100111111",
  6845=>"010000000",
  6846=>"110110110",
  6847=>"000000000",
  6848=>"111011000",
  6849=>"111011110",
  6850=>"111111110",
  6851=>"010010000",
  6852=>"000110111",
  6853=>"000000101",
  6854=>"000100100",
  6855=>"101101101",
  6856=>"000101101",
  6857=>"001101101",
  6858=>"000010000",
  6859=>"000000000",
  6860=>"111111111",
  6861=>"010010011",
  6862=>"001001001",
  6863=>"111111000",
  6864=>"111011010",
  6865=>"111111110",
  6866=>"001111111",
  6867=>"001001001",
  6868=>"010011010",
  6869=>"111111110",
  6870=>"101101001",
  6871=>"111011110",
  6872=>"000100100",
  6873=>"011011111",
  6874=>"111100000",
  6875=>"011010000",
  6876=>"000000000",
  6877=>"000000000",
  6878=>"010010010",
  6879=>"001001011",
  6880=>"101101111",
  6881=>"000000001",
  6882=>"101101101",
  6883=>"111000000",
  6884=>"000000010",
  6885=>"000111100",
  6886=>"000000111",
  6887=>"010000001",
  6888=>"111111111",
  6889=>"010010010",
  6890=>"111101101",
  6891=>"111110010",
  6892=>"001000011",
  6893=>"000000000",
  6894=>"110011011",
  6895=>"000000101",
  6896=>"000000000",
  6897=>"001111111",
  6898=>"001000101",
  6899=>"000001111",
  6900=>"000010000",
  6901=>"001001001",
  6902=>"001111011",
  6903=>"000101101",
  6904=>"110010011",
  6905=>"011111010",
  6906=>"010010010",
  6907=>"101111111",
  6908=>"001000000",
  6909=>"001001001",
  6910=>"011011000",
  6911=>"110110111",
  6912=>"011011001",
  6913=>"101101111",
  6914=>"000000010",
  6915=>"010000000",
  6916=>"000000000",
  6917=>"110111111",
  6918=>"000100111",
  6919=>"000111111",
  6920=>"001000000",
  6921=>"000000111",
  6922=>"101101101",
  6923=>"111011000",
  6924=>"110000000",
  6925=>"000000111",
  6926=>"110110111",
  6927=>"101111111",
  6928=>"111111111",
  6929=>"000000101",
  6930=>"000000010",
  6931=>"101001001",
  6932=>"101001001",
  6933=>"000111001",
  6934=>"111111111",
  6935=>"101101101",
  6936=>"000010010",
  6937=>"100000000",
  6938=>"010111101",
  6939=>"000001101",
  6940=>"101011011",
  6941=>"000000001",
  6942=>"001001001",
  6943=>"000000000",
  6944=>"110011001",
  6945=>"111111111",
  6946=>"101111101",
  6947=>"101111000",
  6948=>"100000000",
  6949=>"000000111",
  6950=>"000000010",
  6951=>"000001011",
  6952=>"101101011",
  6953=>"011000101",
  6954=>"000011110",
  6955=>"100100100",
  6956=>"110110110",
  6957=>"001001000",
  6958=>"011011111",
  6959=>"011011011",
  6960=>"010010100",
  6961=>"000010010",
  6962=>"100100100",
  6963=>"110000000",
  6964=>"010111111",
  6965=>"000010001",
  6966=>"000000000",
  6967=>"000001001",
  6968=>"001111001",
  6969=>"100101111",
  6970=>"001001100",
  6971=>"001000100",
  6972=>"000000100",
  6973=>"000000000",
  6974=>"000010011",
  6975=>"010010110",
  6976=>"000000000",
  6977=>"100101101",
  6978=>"011111011",
  6979=>"101100100",
  6980=>"101011000",
  6981=>"000000101",
  6982=>"001101011",
  6983=>"101101111",
  6984=>"010000000",
  6985=>"000001001",
  6986=>"101101001",
  6987=>"100100100",
  6988=>"001011111",
  6989=>"011011000",
  6990=>"001100101",
  6991=>"010011011",
  6992=>"100111101",
  6993=>"111111000",
  6994=>"101000001",
  6995=>"010010000",
  6996=>"010000000",
  6997=>"010011001",
  6998=>"111111111",
  6999=>"110111010",
  7000=>"001001001",
  7001=>"111011010",
  7002=>"010010001",
  7003=>"111111001",
  7004=>"001001001",
  7005=>"000000000",
  7006=>"110010010",
  7007=>"000100001",
  7008=>"111010000",
  7009=>"100100110",
  7010=>"110110100",
  7011=>"100100111",
  7012=>"100111110",
  7013=>"000001011",
  7014=>"111111111",
  7015=>"101111111",
  7016=>"111011011",
  7017=>"010110010",
  7018=>"111111011",
  7019=>"101101111",
  7020=>"000111000",
  7021=>"000110001",
  7022=>"011110010",
  7023=>"000000101",
  7024=>"011010111",
  7025=>"011111111",
  7026=>"000010000",
  7027=>"010010010",
  7028=>"001011011",
  7029=>"110110110",
  7030=>"101101100",
  7031=>"011111100",
  7032=>"011000000",
  7033=>"000000000",
  7034=>"000000110",
  7035=>"111110111",
  7036=>"000010000",
  7037=>"111000000",
  7038=>"000000111",
  7039=>"000000010",
  7040=>"110110111",
  7041=>"001001011",
  7042=>"111111111",
  7043=>"000000001",
  7044=>"010111111",
  7045=>"101100111",
  7046=>"101001000",
  7047=>"010110110",
  7048=>"100000000",
  7049=>"001000000",
  7050=>"111110000",
  7051=>"100101111",
  7052=>"101100111",
  7053=>"000000000",
  7054=>"110111111",
  7055=>"110111011",
  7056=>"010011000",
  7057=>"111110110",
  7058=>"110110000",
  7059=>"000000001",
  7060=>"100100111",
  7061=>"000010000",
  7062=>"011001010",
  7063=>"001001011",
  7064=>"111110111",
  7065=>"000000101",
  7066=>"000000100",
  7067=>"100101110",
  7068=>"010000000",
  7069=>"000000011",
  7070=>"000000101",
  7071=>"010000100",
  7072=>"010011001",
  7073=>"000100100",
  7074=>"011010110",
  7075=>"001111111",
  7076=>"000100110",
  7077=>"000010111",
  7078=>"100100101",
  7079=>"110110110",
  7080=>"101101100",
  7081=>"000100101",
  7082=>"111010000",
  7083=>"111111110",
  7084=>"000000011",
  7085=>"010010010",
  7086=>"101101000",
  7087=>"001000100",
  7088=>"101100000",
  7089=>"000010010",
  7090=>"111001011",
  7091=>"000010010",
  7092=>"111111001",
  7093=>"110100100",
  7094=>"111111100",
  7095=>"011001001",
  7096=>"000011111",
  7097=>"000000110",
  7098=>"011001001",
  7099=>"000010010",
  7100=>"000000000",
  7101=>"110110110",
  7102=>"111101101",
  7103=>"111101101",
  7104=>"000001011",
  7105=>"010010110",
  7106=>"000000001",
  7107=>"010000000",
  7108=>"100000000",
  7109=>"001000010",
  7110=>"000010000",
  7111=>"100101110",
  7112=>"001101100",
  7113=>"000001011",
  7114=>"001001001",
  7115=>"000000000",
  7116=>"110110000",
  7117=>"100110110",
  7118=>"001001001",
  7119=>"010010111",
  7120=>"101001001",
  7121=>"000000001",
  7122=>"111111111",
  7123=>"010111111",
  7124=>"000000000",
  7125=>"011011111",
  7126=>"000010010",
  7127=>"100001001",
  7128=>"000000000",
  7129=>"011010100",
  7130=>"000001000",
  7131=>"011000000",
  7132=>"001111100",
  7133=>"010111111",
  7134=>"011110100",
  7135=>"001001001",
  7136=>"001101100",
  7137=>"111001111",
  7138=>"000010111",
  7139=>"100100101",
  7140=>"111111000",
  7141=>"111110111",
  7142=>"110110110",
  7143=>"000000000",
  7144=>"001001001",
  7145=>"011111001",
  7146=>"000000011",
  7147=>"111011111",
  7148=>"000000101",
  7149=>"111111101",
  7150=>"101111101",
  7151=>"000000100",
  7152=>"111101000",
  7153=>"010010010",
  7154=>"101101111",
  7155=>"000000001",
  7156=>"011101001",
  7157=>"000000000",
  7158=>"110110110",
  7159=>"111111001",
  7160=>"111111101",
  7161=>"000000000",
  7162=>"101101011",
  7163=>"000000000",
  7164=>"000100000",
  7165=>"000101001",
  7166=>"000000010",
  7167=>"000000000",
  7168=>"111001001",
  7169=>"000000000",
  7170=>"000000000",
  7171=>"000001001",
  7172=>"001001001",
  7173=>"111111111",
  7174=>"011011011",
  7175=>"111111111",
  7176=>"000111000",
  7177=>"001001111",
  7178=>"111101111",
  7179=>"011111111",
  7180=>"110111110",
  7181=>"111111111",
  7182=>"000000111",
  7183=>"011111111",
  7184=>"000100100",
  7185=>"000001111",
  7186=>"000000001",
  7187=>"000000000",
  7188=>"111111111",
  7189=>"000000000",
  7190=>"000100000",
  7191=>"000010111",
  7192=>"111001000",
  7193=>"100000000",
  7194=>"110111111",
  7195=>"000000111",
  7196=>"000000000",
  7197=>"001101100",
  7198=>"100110110",
  7199=>"111111000",
  7200=>"001011010",
  7201=>"000000111",
  7202=>"101001001",
  7203=>"000000101",
  7204=>"111110000",
  7205=>"110111110",
  7206=>"111111011",
  7207=>"101111001",
  7208=>"100101111",
  7209=>"011001011",
  7210=>"111111111",
  7211=>"111111111",
  7212=>"000000000",
  7213=>"000000001",
  7214=>"000000000",
  7215=>"111111111",
  7216=>"000000000",
  7217=>"100110000",
  7218=>"111110010",
  7219=>"100101100",
  7220=>"000001001",
  7221=>"100010000",
  7222=>"001111111",
  7223=>"000000000",
  7224=>"111101011",
  7225=>"001111000",
  7226=>"000000000",
  7227=>"011111111",
  7228=>"111111111",
  7229=>"111000000",
  7230=>"000101111",
  7231=>"111001000",
  7232=>"011001110",
  7233=>"000010010",
  7234=>"110111110",
  7235=>"111111111",
  7236=>"000000000",
  7237=>"111111111",
  7238=>"011011110",
  7239=>"000000000",
  7240=>"111111011",
  7241=>"111111111",
  7242=>"110111111",
  7243=>"111111101",
  7244=>"000000000",
  7245=>"000001100",
  7246=>"111101100",
  7247=>"000000000",
  7248=>"011011111",
  7249=>"000000111",
  7250=>"000101000",
  7251=>"000100100",
  7252=>"101111100",
  7253=>"100111100",
  7254=>"111111100",
  7255=>"111111111",
  7256=>"000011111",
  7257=>"000001111",
  7258=>"111111111",
  7259=>"001011001",
  7260=>"000000000",
  7261=>"011111111",
  7262=>"000000100",
  7263=>"000000011",
  7264=>"111001001",
  7265=>"111111011",
  7266=>"000000000",
  7267=>"111111000",
  7268=>"000000111",
  7269=>"111100101",
  7270=>"111111111",
  7271=>"011111111",
  7272=>"000000000",
  7273=>"000111111",
  7274=>"001000000",
  7275=>"000011000",
  7276=>"000000100",
  7277=>"111111111",
  7278=>"111111111",
  7279=>"111001001",
  7280=>"000000000",
  7281=>"000000000",
  7282=>"001000000",
  7283=>"111000110",
  7284=>"000000000",
  7285=>"000100110",
  7286=>"111111110",
  7287=>"111111111",
  7288=>"111111111",
  7289=>"000000000",
  7290=>"000000101",
  7291=>"111111111",
  7292=>"100100100",
  7293=>"000000000",
  7294=>"111111111",
  7295=>"000110110",
  7296=>"000000101",
  7297=>"111111111",
  7298=>"000000000",
  7299=>"001101111",
  7300=>"111111111",
  7301=>"111111111",
  7302=>"000000000",
  7303=>"111111001",
  7304=>"111111101",
  7305=>"000011011",
  7306=>"000000000",
  7307=>"111011000",
  7308=>"001011111",
  7309=>"111111111",
  7310=>"101001000",
  7311=>"011000000",
  7312=>"000000000",
  7313=>"111000000",
  7314=>"000000000",
  7315=>"110111111",
  7316=>"111111110",
  7317=>"111111111",
  7318=>"000000000",
  7319=>"000000000",
  7320=>"111111111",
  7321=>"011111000",
  7322=>"000000000",
  7323=>"011111001",
  7324=>"111110110",
  7325=>"000000111",
  7326=>"111111111",
  7327=>"011111011",
  7328=>"001101000",
  7329=>"001100000",
  7330=>"011110110",
  7331=>"000000000",
  7332=>"011111111",
  7333=>"101000011",
  7334=>"000000010",
  7335=>"000000000",
  7336=>"000111111",
  7337=>"111000000",
  7338=>"111111111",
  7339=>"101101111",
  7340=>"111111111",
  7341=>"111101011",
  7342=>"101001001",
  7343=>"000000000",
  7344=>"000110000",
  7345=>"111110110",
  7346=>"010111111",
  7347=>"111111111",
  7348=>"000000001",
  7349=>"011111110",
  7350=>"111111111",
  7351=>"110010110",
  7352=>"111111111",
  7353=>"100111111",
  7354=>"111111110",
  7355=>"111111111",
  7356=>"110111010",
  7357=>"101100000",
  7358=>"111111111",
  7359=>"111000000",
  7360=>"111111111",
  7361=>"000000000",
  7362=>"111110110",
  7363=>"111111111",
  7364=>"000001001",
  7365=>"000000000",
  7366=>"000000000",
  7367=>"001000000",
  7368=>"111111111",
  7369=>"000000000",
  7370=>"111111101",
  7371=>"000000000",
  7372=>"111110100",
  7373=>"111111111",
  7374=>"011011111",
  7375=>"111110100",
  7376=>"000011111",
  7377=>"000111111",
  7378=>"111011111",
  7379=>"000000000",
  7380=>"111101001",
  7381=>"100000000",
  7382=>"110111111",
  7383=>"100110111",
  7384=>"111111111",
  7385=>"110111001",
  7386=>"000101111",
  7387=>"101111110",
  7388=>"110111111",
  7389=>"111111111",
  7390=>"000000000",
  7391=>"111001000",
  7392=>"000110111",
  7393=>"010011111",
  7394=>"111111110",
  7395=>"000000010",
  7396=>"111111111",
  7397=>"010110000",
  7398=>"000101110",
  7399=>"000001111",
  7400=>"000000000",
  7401=>"000000000",
  7402=>"111111111",
  7403=>"000001111",
  7404=>"000000000",
  7405=>"110000111",
  7406=>"000000100",
  7407=>"111000000",
  7408=>"111101100",
  7409=>"111111111",
  7410=>"111111111",
  7411=>"010111111",
  7412=>"111111111",
  7413=>"111000000",
  7414=>"111111111",
  7415=>"111111111",
  7416=>"100000100",
  7417=>"010000000",
  7418=>"110111111",
  7419=>"000011111",
  7420=>"001000001",
  7421=>"111111111",
  7422=>"010000000",
  7423=>"111111111",
  7424=>"101111111",
  7425=>"010010010",
  7426=>"010111111",
  7427=>"000000000",
  7428=>"000000000",
  7429=>"111111111",
  7430=>"000000100",
  7431=>"000000000",
  7432=>"111111011",
  7433=>"000000010",
  7434=>"000000000",
  7435=>"001011111",
  7436=>"000000000",
  7437=>"000111000",
  7438=>"101101100",
  7439=>"111111111",
  7440=>"001111100",
  7441=>"000000011",
  7442=>"111111111",
  7443=>"101111111",
  7444=>"000011011",
  7445=>"010111111",
  7446=>"000000000",
  7447=>"111111111",
  7448=>"000000000",
  7449=>"000010011",
  7450=>"001000000",
  7451=>"111010011",
  7452=>"000000110",
  7453=>"001000000",
  7454=>"111111111",
  7455=>"001000000",
  7456=>"110110111",
  7457=>"101110100",
  7458=>"111111111",
  7459=>"000000000",
  7460=>"000000000",
  7461=>"000100000",
  7462=>"110110111",
  7463=>"000000000",
  7464=>"100000000",
  7465=>"011111111",
  7466=>"000011111",
  7467=>"000000000",
  7468=>"111111111",
  7469=>"000000000",
  7470=>"111111111",
  7471=>"010010000",
  7472=>"111111111",
  7473=>"000000000",
  7474=>"000000000",
  7475=>"000000011",
  7476=>"111111111",
  7477=>"001111110",
  7478=>"111111100",
  7479=>"111111111",
  7480=>"111110000",
  7481=>"111000111",
  7482=>"110111111",
  7483=>"000000100",
  7484=>"001001111",
  7485=>"101100000",
  7486=>"111111101",
  7487=>"110111110",
  7488=>"111111000",
  7489=>"010100110",
  7490=>"111111111",
  7491=>"111111111",
  7492=>"000110111",
  7493=>"100111111",
  7494=>"111111100",
  7495=>"111110100",
  7496=>"111111110",
  7497=>"011000000",
  7498=>"111111111",
  7499=>"000000000",
  7500=>"010000001",
  7501=>"111111111",
  7502=>"101000000",
  7503=>"111111111",
  7504=>"110100111",
  7505=>"100100100",
  7506=>"000111011",
  7507=>"001000000",
  7508=>"000100000",
  7509=>"011001001",
  7510=>"100000000",
  7511=>"001000000",
  7512=>"111111111",
  7513=>"000001111",
  7514=>"111111001",
  7515=>"110111111",
  7516=>"111111111",
  7517=>"100000000",
  7518=>"000100000",
  7519=>"000100010",
  7520=>"111111111",
  7521=>"000000000",
  7522=>"001011011",
  7523=>"111111111",
  7524=>"000110110",
  7525=>"111101111",
  7526=>"000000000",
  7527=>"100001000",
  7528=>"000011001",
  7529=>"111111111",
  7530=>"101100100",
  7531=>"100111111",
  7532=>"110110100",
  7533=>"001111100",
  7534=>"000000000",
  7535=>"000001000",
  7536=>"000000000",
  7537=>"010010000",
  7538=>"000000000",
  7539=>"000000000",
  7540=>"011010011",
  7541=>"111010000",
  7542=>"100000111",
  7543=>"111111010",
  7544=>"111111111",
  7545=>"111111111",
  7546=>"110111111",
  7547=>"000001000",
  7548=>"111110100",
  7549=>"111111101",
  7550=>"111101000",
  7551=>"000000000",
  7552=>"000100110",
  7553=>"100100100",
  7554=>"100110111",
  7555=>"000000000",
  7556=>"000000001",
  7557=>"111111111",
  7558=>"001111000",
  7559=>"111111111",
  7560=>"111111111",
  7561=>"000110110",
  7562=>"101111101",
  7563=>"111111110",
  7564=>"111111111",
  7565=>"111111111",
  7566=>"000000000",
  7567=>"111111111",
  7568=>"000000000",
  7569=>"111110111",
  7570=>"111101101",
  7571=>"100100111",
  7572=>"000000111",
  7573=>"010010010",
  7574=>"101101100",
  7575=>"000100000",
  7576=>"111111111",
  7577=>"000000000",
  7578=>"111111011",
  7579=>"101111111",
  7580=>"111111000",
  7581=>"111111100",
  7582=>"111111111",
  7583=>"111111011",
  7584=>"000010011",
  7585=>"011011011",
  7586=>"000100111",
  7587=>"111111111",
  7588=>"000000000",
  7589=>"000110111",
  7590=>"111111111",
  7591=>"111111111",
  7592=>"000000000",
  7593=>"000001111",
  7594=>"100110110",
  7595=>"000000110",
  7596=>"000000111",
  7597=>"111101000",
  7598=>"000111111",
  7599=>"000000000",
  7600=>"010111111",
  7601=>"000111100",
  7602=>"100100000",
  7603=>"000000000",
  7604=>"111101111",
  7605=>"111111111",
  7606=>"100100000",
  7607=>"000000010",
  7608=>"000000001",
  7609=>"000000000",
  7610=>"000000110",
  7611=>"000000010",
  7612=>"111111111",
  7613=>"011111100",
  7614=>"001000000",
  7615=>"111111110",
  7616=>"000000000",
  7617=>"000000000",
  7618=>"000000000",
  7619=>"000000000",
  7620=>"011001111",
  7621=>"111111100",
  7622=>"100100000",
  7623=>"000111111",
  7624=>"100110110",
  7625=>"111111000",
  7626=>"000111011",
  7627=>"111111110",
  7628=>"110110000",
  7629=>"000000111",
  7630=>"111100101",
  7631=>"100000000",
  7632=>"000000000",
  7633=>"011011011",
  7634=>"000101111",
  7635=>"000000000",
  7636=>"000000000",
  7637=>"111111111",
  7638=>"111101101",
  7639=>"100100110",
  7640=>"000001111",
  7641=>"111111101",
  7642=>"000000000",
  7643=>"111011111",
  7644=>"000000000",
  7645=>"000000100",
  7646=>"111111111",
  7647=>"011001011",
  7648=>"100111111",
  7649=>"010010000",
  7650=>"111111010",
  7651=>"100110000",
  7652=>"000000000",
  7653=>"111011001",
  7654=>"001111111",
  7655=>"010011010",
  7656=>"111111111",
  7657=>"001000100",
  7658=>"010111011",
  7659=>"100111111",
  7660=>"110110111",
  7661=>"000100110",
  7662=>"111111111",
  7663=>"000000000",
  7664=>"111011011",
  7665=>"111111111",
  7666=>"000001100",
  7667=>"000010111",
  7668=>"000000000",
  7669=>"110000000",
  7670=>"100000000",
  7671=>"101101101",
  7672=>"000000000",
  7673=>"000000001",
  7674=>"110110110",
  7675=>"111111001",
  7676=>"111111100",
  7677=>"111001000",
  7678=>"101111111",
  7679=>"110100100",
  7680=>"010010111",
  7681=>"011000000",
  7682=>"000000100",
  7683=>"111111111",
  7684=>"111111111",
  7685=>"011110110",
  7686=>"000000000",
  7687=>"100111111",
  7688=>"010010011",
  7689=>"000111111",
  7690=>"111111111",
  7691=>"011000000",
  7692=>"000111110",
  7693=>"111111111",
  7694=>"100100001",
  7695=>"000000000",
  7696=>"110110110",
  7697=>"000111111",
  7698=>"111111111",
  7699=>"000100000",
  7700=>"000000000",
  7701=>"111111111",
  7702=>"110111110",
  7703=>"100110100",
  7704=>"111111111",
  7705=>"000011110",
  7706=>"000000000",
  7707=>"111110000",
  7708=>"000001001",
  7709=>"000100000",
  7710=>"000000000",
  7711=>"000000010",
  7712=>"101000000",
  7713=>"000000000",
  7714=>"001011111",
  7715=>"011111111",
  7716=>"011000000",
  7717=>"001001011",
  7718=>"000100100",
  7719=>"011000000",
  7720=>"000000000",
  7721=>"000111111",
  7722=>"111111111",
  7723=>"111111111",
  7724=>"111111110",
  7725=>"111111000",
  7726=>"111111110",
  7727=>"000000000",
  7728=>"000000000",
  7729=>"000000000",
  7730=>"000000100",
  7731=>"111111111",
  7732=>"001101001",
  7733=>"011011011",
  7734=>"111101000",
  7735=>"001001011",
  7736=>"000000010",
  7737=>"111011110",
  7738=>"110111111",
  7739=>"000000101",
  7740=>"000000000",
  7741=>"110111111",
  7742=>"000001001",
  7743=>"111100000",
  7744=>"000000001",
  7745=>"100100000",
  7746=>"111111000",
  7747=>"011000000",
  7748=>"111111111",
  7749=>"110110111",
  7750=>"000000000",
  7751=>"000000000",
  7752=>"111111111",
  7753=>"111111111",
  7754=>"111111111",
  7755=>"000111000",
  7756=>"000000000",
  7757=>"011011011",
  7758=>"000000101",
  7759=>"111111111",
  7760=>"000000001",
  7761=>"111111111",
  7762=>"111111110",
  7763=>"111001001",
  7764=>"001111111",
  7765=>"111110110",
  7766=>"010111111",
  7767=>"101101001",
  7768=>"110000000",
  7769=>"000000000",
  7770=>"000010111",
  7771=>"001011011",
  7772=>"111111111",
  7773=>"000111001",
  7774=>"011001111",
  7775=>"111001001",
  7776=>"000000000",
  7777=>"000000111",
  7778=>"111111111",
  7779=>"101001000",
  7780=>"111110110",
  7781=>"000000001",
  7782=>"000101101",
  7783=>"000100101",
  7784=>"000000000",
  7785=>"001001000",
  7786=>"010000000",
  7787=>"000000000",
  7788=>"110100100",
  7789=>"111111111",
  7790=>"000000000",
  7791=>"110111111",
  7792=>"111111110",
  7793=>"001000000",
  7794=>"100100111",
  7795=>"111100100",
  7796=>"110110011",
  7797=>"000110110",
  7798=>"111111110",
  7799=>"000111111",
  7800=>"001000001",
  7801=>"111111111",
  7802=>"000000000",
  7803=>"110000000",
  7804=>"111111111",
  7805=>"000000000",
  7806=>"100000000",
  7807=>"111111111",
  7808=>"000010000",
  7809=>"011000001",
  7810=>"000000000",
  7811=>"000001000",
  7812=>"000111111",
  7813=>"000100111",
  7814=>"111111111",
  7815=>"000001001",
  7816=>"000000000",
  7817=>"000000000",
  7818=>"111111110",
  7819=>"000000000",
  7820=>"100100110",
  7821=>"000000000",
  7822=>"000000110",
  7823=>"000000000",
  7824=>"101111111",
  7825=>"000100000",
  7826=>"000010000",
  7827=>"000000000",
  7828=>"110000000",
  7829=>"111111111",
  7830=>"111111111",
  7831=>"111000000",
  7832=>"000000000",
  7833=>"111111111",
  7834=>"111101101",
  7835=>"000000000",
  7836=>"111011111",
  7837=>"011000111",
  7838=>"111111111",
  7839=>"000101100",
  7840=>"001111000",
  7841=>"000000000",
  7842=>"000111111",
  7843=>"111111111",
  7844=>"000011111",
  7845=>"001111100",
  7846=>"101101001",
  7847=>"110110110",
  7848=>"111011010",
  7849=>"000000001",
  7850=>"111111111",
  7851=>"000011000",
  7852=>"111111010",
  7853=>"000000000",
  7854=>"000000000",
  7855=>"000000000",
  7856=>"011111110",
  7857=>"000000011",
  7858=>"011111111",
  7859=>"101000100",
  7860=>"000000000",
  7861=>"100111111",
  7862=>"001101000",
  7863=>"001001111",
  7864=>"001001000",
  7865=>"000000000",
  7866=>"000110110",
  7867=>"011011000",
  7868=>"111111111",
  7869=>"000000000",
  7870=>"110110110",
  7871=>"000000100",
  7872=>"111111111",
  7873=>"110110111",
  7874=>"111110111",
  7875=>"110110000",
  7876=>"111111111",
  7877=>"011001000",
  7878=>"000001011",
  7879=>"000000000",
  7880=>"000010011",
  7881=>"101101111",
  7882=>"000000000",
  7883=>"000001000",
  7884=>"001111100",
  7885=>"100110110",
  7886=>"000000000",
  7887=>"000000000",
  7888=>"000000110",
  7889=>"100100000",
  7890=>"111111101",
  7891=>"000000001",
  7892=>"101111101",
  7893=>"111100111",
  7894=>"111111000",
  7895=>"111000000",
  7896=>"111010011",
  7897=>"000000000",
  7898=>"111111111",
  7899=>"111111111",
  7900=>"001111111",
  7901=>"000100100",
  7902=>"000101110",
  7903=>"001011000",
  7904=>"000000000",
  7905=>"110110110",
  7906=>"111110000",
  7907=>"111111111",
  7908=>"001000000",
  7909=>"000111110",
  7910=>"111111111",
  7911=>"000000000",
  7912=>"111111111",
  7913=>"001111111",
  7914=>"000000110",
  7915=>"000000000",
  7916=>"000000000",
  7917=>"000000000",
  7918=>"000100101",
  7919=>"000000000",
  7920=>"111111000",
  7921=>"001000000",
  7922=>"111111111",
  7923=>"101101001",
  7924=>"111011010",
  7925=>"111000000",
  7926=>"010000000",
  7927=>"111001000",
  7928=>"000000000",
  7929=>"011111111",
  7930=>"111111111",
  7931=>"100000100",
  7932=>"001001011",
  7933=>"000000001",
  7934=>"000111000",
  7935=>"010000000",
  7936=>"000001001",
  7937=>"000000001",
  7938=>"001001000",
  7939=>"000110111",
  7940=>"000000000",
  7941=>"111100111",
  7942=>"000000000",
  7943=>"111111111",
  7944=>"000001011",
  7945=>"000000000",
  7946=>"000001000",
  7947=>"110000000",
  7948=>"000000000",
  7949=>"111000000",
  7950=>"111111001",
  7951=>"000101111",
  7952=>"011111001",
  7953=>"000011111",
  7954=>"111101101",
  7955=>"000111111",
  7956=>"110000000",
  7957=>"011011111",
  7958=>"000001001",
  7959=>"000000000",
  7960=>"000000000",
  7961=>"111000000",
  7962=>"111111111",
  7963=>"000000000",
  7964=>"110111111",
  7965=>"000011000",
  7966=>"000000000",
  7967=>"011101101",
  7968=>"110111010",
  7969=>"001101100",
  7970=>"111110000",
  7971=>"100000001",
  7972=>"110000000",
  7973=>"111111111",
  7974=>"111111111",
  7975=>"111100000",
  7976=>"000000111",
  7977=>"101101111",
  7978=>"111100100",
  7979=>"111000000",
  7980=>"001001000",
  7981=>"001001001",
  7982=>"000000000",
  7983=>"000000000",
  7984=>"111111111",
  7985=>"110100100",
  7986=>"000011001",
  7987=>"110110111",
  7988=>"000000100",
  7989=>"000001011",
  7990=>"000111000",
  7991=>"000000000",
  7992=>"000000000",
  7993=>"001000111",
  7994=>"000010000",
  7995=>"000000000",
  7996=>"000001000",
  7997=>"000010000",
  7998=>"000000000",
  7999=>"000110111",
  8000=>"111111111",
  8001=>"111111110",
  8002=>"111111111",
  8003=>"010011000",
  8004=>"100000000",
  8005=>"000000000",
  8006=>"011011011",
  8007=>"010110100",
  8008=>"000000000",
  8009=>"000000000",
  8010=>"001001001",
  8011=>"111011011",
  8012=>"000001011",
  8013=>"111111000",
  8014=>"000101000",
  8015=>"001011111",
  8016=>"000010010",
  8017=>"110110110",
  8018=>"001001111",
  8019=>"011010010",
  8020=>"000111111",
  8021=>"011011011",
  8022=>"001000111",
  8023=>"110110000",
  8024=>"000000001",
  8025=>"010111111",
  8026=>"000000000",
  8027=>"000001001",
  8028=>"011111111",
  8029=>"111001101",
  8030=>"001001001",
  8031=>"001011111",
  8032=>"000000011",
  8033=>"111111111",
  8034=>"000001001",
  8035=>"111001111",
  8036=>"111110000",
  8037=>"111111111",
  8038=>"000000000",
  8039=>"100000000",
  8040=>"111111111",
  8041=>"000000111",
  8042=>"000000000",
  8043=>"011000000",
  8044=>"100110111",
  8045=>"001000000",
  8046=>"000111111",
  8047=>"000000000",
  8048=>"000000000",
  8049=>"110000000",
  8050=>"000000101",
  8051=>"000010000",
  8052=>"011011000",
  8053=>"110110000",
  8054=>"000111111",
  8055=>"000000011",
  8056=>"011111111",
  8057=>"000000000",
  8058=>"111000001",
  8059=>"011111000",
  8060=>"111111101",
  8061=>"111101111",
  8062=>"000000111",
  8063=>"000000000",
  8064=>"000000000",
  8065=>"111111111",
  8066=>"001001001",
  8067=>"111111111",
  8068=>"000001001",
  8069=>"111111111",
  8070=>"000000000",
  8071=>"000000100",
  8072=>"111111111",
  8073=>"111110100",
  8074=>"000000000",
  8075=>"001000000",
  8076=>"000111111",
  8077=>"000011011",
  8078=>"000010010",
  8079=>"000000000",
  8080=>"000000000",
  8081=>"111111111",
  8082=>"101000000",
  8083=>"000000000",
  8084=>"000001111",
  8085=>"000001000",
  8086=>"111111111",
  8087=>"011011011",
  8088=>"111111111",
  8089=>"100000000",
  8090=>"111111111",
  8091=>"111111111",
  8092=>"000001000",
  8093=>"101000010",
  8094=>"000000000",
  8095=>"010010000",
  8096=>"000000000",
  8097=>"110000000",
  8098=>"001101101",
  8099=>"111111111",
  8100=>"101101000",
  8101=>"110111110",
  8102=>"101001111",
  8103=>"111111000",
  8104=>"000000100",
  8105=>"011001000",
  8106=>"011111111",
  8107=>"111111111",
  8108=>"011000111",
  8109=>"111011111",
  8110=>"111001000",
  8111=>"001111011",
  8112=>"111110110",
  8113=>"111110110",
  8114=>"000000100",
  8115=>"000110111",
  8116=>"000111011",
  8117=>"101111000",
  8118=>"111110000",
  8119=>"000000000",
  8120=>"000000000",
  8121=>"111111011",
  8122=>"000000100",
  8123=>"111100101",
  8124=>"000000000",
  8125=>"101000001",
  8126=>"011000100",
  8127=>"011011011",
  8128=>"000000000",
  8129=>"110111111",
  8130=>"000011111",
  8131=>"000111111",
  8132=>"000111111",
  8133=>"010111110",
  8134=>"111111111",
  8135=>"100111110",
  8136=>"000101000",
  8137=>"001011111",
  8138=>"111111000",
  8139=>"000000000",
  8140=>"000000000",
  8141=>"000000000",
  8142=>"111111111",
  8143=>"111111111",
  8144=>"000000000",
  8145=>"001001101",
  8146=>"110110111",
  8147=>"111111000",
  8148=>"010011001",
  8149=>"011001000",
  8150=>"000001000",
  8151=>"010111111",
  8152=>"001000000",
  8153=>"001001011",
  8154=>"111000000",
  8155=>"111111111",
  8156=>"000000000",
  8157=>"111111001",
  8158=>"000000110",
  8159=>"011011001",
  8160=>"100000000",
  8161=>"000000000",
  8162=>"000000000",
  8163=>"000000111",
  8164=>"111111111",
  8165=>"111111111",
  8166=>"101001111",
  8167=>"000000011",
  8168=>"101100101",
  8169=>"000000000",
  8170=>"111111110",
  8171=>"000000000",
  8172=>"111110111",
  8173=>"100100100",
  8174=>"111101001",
  8175=>"001000000",
  8176=>"000000000",
  8177=>"000001001",
  8178=>"000000100",
  8179=>"000000000",
  8180=>"111111111",
  8181=>"011011011",
  8182=>"110011000",
  8183=>"110110000",
  8184=>"111111111",
  8185=>"110010000",
  8186=>"111111000",
  8187=>"111001100",
  8188=>"000100110",
  8189=>"000111111",
  8190=>"001001000",
  8191=>"000000000",
  8192=>"111110111",
  8193=>"111110000",
  8194=>"111111000",
  8195=>"111000000",
  8196=>"000000000",
  8197=>"000100110",
  8198=>"111000000",
  8199=>"000000000",
  8200=>"111111011",
  8201=>"000000110",
  8202=>"100000000",
  8203=>"111111001",
  8204=>"111010111",
  8205=>"111000000",
  8206=>"000000011",
  8207=>"111100111",
  8208=>"001001111",
  8209=>"111111100",
  8210=>"111000000",
  8211=>"011000000",
  8212=>"000000111",
  8213=>"010000000",
  8214=>"001000000",
  8215=>"101111111",
  8216=>"110000001",
  8217=>"111111000",
  8218=>"111000000",
  8219=>"000000011",
  8220=>"000111111",
  8221=>"000000111",
  8222=>"100000000",
  8223=>"111000000",
  8224=>"000000000",
  8225=>"111111111",
  8226=>"000001111",
  8227=>"111011001",
  8228=>"000000000",
  8229=>"111111110",
  8230=>"111110000",
  8231=>"100111011",
  8232=>"101101011",
  8233=>"111111000",
  8234=>"000000111",
  8235=>"001000111",
  8236=>"001101111",
  8237=>"010111111",
  8238=>"000000000",
  8239=>"111111111",
  8240=>"000000000",
  8241=>"111101001",
  8242=>"100001111",
  8243=>"111101111",
  8244=>"000110000",
  8245=>"110000001",
  8246=>"001011111",
  8247=>"111000000",
  8248=>"010110111",
  8249=>"111110000",
  8250=>"000000101",
  8251=>"111010111",
  8252=>"000111010",
  8253=>"000000100",
  8254=>"111111110",
  8255=>"000000000",
  8256=>"100100011",
  8257=>"000111111",
  8258=>"111111111",
  8259=>"111111001",
  8260=>"000001101",
  8261=>"110000000",
  8262=>"000000101",
  8263=>"000000111",
  8264=>"011110100",
  8265=>"000001111",
  8266=>"000000001",
  8267=>"100100000",
  8268=>"110000010",
  8269=>"111100100",
  8270=>"000001111",
  8271=>"001000000",
  8272=>"101111111",
  8273=>"100100100",
  8274=>"000111111",
  8275=>"111100100",
  8276=>"000000110",
  8277=>"000100111",
  8278=>"110000111",
  8279=>"111111111",
  8280=>"000100000",
  8281=>"000101101",
  8282=>"000000010",
  8283=>"111001001",
  8284=>"100010000",
  8285=>"000110111",
  8286=>"000000000",
  8287=>"111111001",
  8288=>"000110000",
  8289=>"101111111",
  8290=>"000110110",
  8291=>"111000000",
  8292=>"001001001",
  8293=>"111111000",
  8294=>"111111111",
  8295=>"100110000",
  8296=>"111001111",
  8297=>"110110000",
  8298=>"010000000",
  8299=>"000000111",
  8300=>"010000000",
  8301=>"000000111",
  8302=>"000000111",
  8303=>"000110111",
  8304=>"111111111",
  8305=>"000000111",
  8306=>"000100111",
  8307=>"111111000",
  8308=>"000000000",
  8309=>"000111011",
  8310=>"111000001",
  8311=>"001000111",
  8312=>"111111100",
  8313=>"111101101",
  8314=>"000000000",
  8315=>"001010111",
  8316=>"000011110",
  8317=>"000100000",
  8318=>"000000000",
  8319=>"000000000",
  8320=>"111001000",
  8321=>"111101100",
  8322=>"000111111",
  8323=>"111111010",
  8324=>"110111111",
  8325=>"000000101",
  8326=>"000110111",
  8327=>"010111111",
  8328=>"111101000",
  8329=>"011000101",
  8330=>"001000010",
  8331=>"111110000",
  8332=>"000111111",
  8333=>"110110110",
  8334=>"111111000",
  8335=>"110110111",
  8336=>"000000000",
  8337=>"111111000",
  8338=>"111111111",
  8339=>"000000111",
  8340=>"111111111",
  8341=>"000000000",
  8342=>"111100000",
  8343=>"000000000",
  8344=>"000000101",
  8345=>"111111010",
  8346=>"000000101",
  8347=>"010110010",
  8348=>"011000000",
  8349=>"111100100",
  8350=>"000000001",
  8351=>"001111010",
  8352=>"111110000",
  8353=>"111100111",
  8354=>"000000000",
  8355=>"000000111",
  8356=>"011110110",
  8357=>"111000000",
  8358=>"110000000",
  8359=>"000100100",
  8360=>"000000111",
  8361=>"111011000",
  8362=>"000111111",
  8363=>"000111111",
  8364=>"111100000",
  8365=>"111111001",
  8366=>"111111111",
  8367=>"111111100",
  8368=>"000000111",
  8369=>"111011000",
  8370=>"010010011",
  8371=>"111000000",
  8372=>"111000000",
  8373=>"101100000",
  8374=>"111000000",
  8375=>"111100000",
  8376=>"111001111",
  8377=>"000111111",
  8378=>"111001001",
  8379=>"111111001",
  8380=>"101011011",
  8381=>"111000000",
  8382=>"000111111",
  8383=>"000110111",
  8384=>"010001000",
  8385=>"100000100",
  8386=>"111000000",
  8387=>"111111000",
  8388=>"110011111",
  8389=>"111111000",
  8390=>"111001001",
  8391=>"110110001",
  8392=>"010111000",
  8393=>"111111111",
  8394=>"000101111",
  8395=>"001000000",
  8396=>"001111110",
  8397=>"000000000",
  8398=>"000000111",
  8399=>"000101111",
  8400=>"000000000",
  8401=>"100100111",
  8402=>"111100111",
  8403=>"000000111",
  8404=>"111111111",
  8405=>"011001011",
  8406=>"000111111",
  8407=>"110111111",
  8408=>"111111000",
  8409=>"110111111",
  8410=>"000000111",
  8411=>"100111111",
  8412=>"111111010",
  8413=>"000000111",
  8414=>"000000011",
  8415=>"100100111",
  8416=>"000101111",
  8417=>"000100010",
  8418=>"111111110",
  8419=>"111101000",
  8420=>"000000000",
  8421=>"001001011",
  8422=>"000011001",
  8423=>"111111000",
  8424=>"111111011",
  8425=>"100000001",
  8426=>"000100100",
  8427=>"111111110",
  8428=>"000011000",
  8429=>"001111111",
  8430=>"111011111",
  8431=>"001000000",
  8432=>"000111111",
  8433=>"111111111",
  8434=>"111111111",
  8435=>"111000001",
  8436=>"111111111",
  8437=>"011111111",
  8438=>"011000000",
  8439=>"111100100",
  8440=>"001011111",
  8441=>"111111110",
  8442=>"000000111",
  8443=>"100110111",
  8444=>"000110010",
  8445=>"111111111",
  8446=>"111000000",
  8447=>"100100111",
  8448=>"101011111",
  8449=>"000001011",
  8450=>"000001111",
  8451=>"000000111",
  8452=>"111101111",
  8453=>"000000110",
  8454=>"111000111",
  8455=>"000100100",
  8456=>"111010000",
  8457=>"111111110",
  8458=>"001000111",
  8459=>"111101000",
  8460=>"100110111",
  8461=>"100000000",
  8462=>"111111100",
  8463=>"110000000",
  8464=>"000111111",
  8465=>"001101111",
  8466=>"000000101",
  8467=>"000110111",
  8468=>"111111111",
  8469=>"111001111",
  8470=>"111000000",
  8471=>"111111111",
  8472=>"000000000",
  8473=>"111111110",
  8474=>"000000000",
  8475=>"111001000",
  8476=>"111110111",
  8477=>"111000000",
  8478=>"111111011",
  8479=>"011100100",
  8480=>"111011000",
  8481=>"111010000",
  8482=>"000000111",
  8483=>"111101000",
  8484=>"100111011",
  8485=>"001000000",
  8486=>"100100111",
  8487=>"111100000",
  8488=>"100110110",
  8489=>"000000001",
  8490=>"001000101",
  8491=>"111111000",
  8492=>"111000000",
  8493=>"111111001",
  8494=>"000000111",
  8495=>"000110110",
  8496=>"000000110",
  8497=>"000000000",
  8498=>"111111111",
  8499=>"000000001",
  8500=>"100110110",
  8501=>"000000000",
  8502=>"111010000",
  8503=>"101000100",
  8504=>"111111000",
  8505=>"000100000",
  8506=>"111111111",
  8507=>"000011000",
  8508=>"010111111",
  8509=>"100100111",
  8510=>"111111011",
  8511=>"111000111",
  8512=>"011011011",
  8513=>"100110111",
  8514=>"000000000",
  8515=>"000000000",
  8516=>"010000110",
  8517=>"000000111",
  8518=>"000111111",
  8519=>"000000111",
  8520=>"000001000",
  8521=>"000000000",
  8522=>"000000111",
  8523=>"100000110",
  8524=>"000000000",
  8525=>"000000000",
  8526=>"000100110",
  8527=>"111110100",
  8528=>"111111111",
  8529=>"000101100",
  8530=>"100100001",
  8531=>"000111011",
  8532=>"000001101",
  8533=>"011000000",
  8534=>"111110100",
  8535=>"000000101",
  8536=>"111111110",
  8537=>"001011111",
  8538=>"111100000",
  8539=>"000000100",
  8540=>"000000000",
  8541=>"111111111",
  8542=>"000000111",
  8543=>"100100111",
  8544=>"011010000",
  8545=>"000000000",
  8546=>"111010000",
  8547=>"000111110",
  8548=>"111011000",
  8549=>"101000001",
  8550=>"000111101",
  8551=>"000000111",
  8552=>"100110010",
  8553=>"000000111",
  8554=>"101000000",
  8555=>"000000000",
  8556=>"111000000",
  8557=>"001000100",
  8558=>"111010000",
  8559=>"111000000",
  8560=>"000000011",
  8561=>"001000001",
  8562=>"011100100",
  8563=>"111110110",
  8564=>"011000000",
  8565=>"000000001",
  8566=>"000000001",
  8567=>"001111111",
  8568=>"000011011",
  8569=>"000001000",
  8570=>"000000001",
  8571=>"000111000",
  8572=>"000000011",
  8573=>"000010111",
  8574=>"000000000",
  8575=>"111100110",
  8576=>"000000000",
  8577=>"111110101",
  8578=>"111001001",
  8579=>"000000000",
  8580=>"110111111",
  8581=>"110100000",
  8582=>"000000000",
  8583=>"000000000",
  8584=>"000111111",
  8585=>"110000000",
  8586=>"101000101",
  8587=>"000110111",
  8588=>"100000101",
  8589=>"111111010",
  8590=>"011111111",
  8591=>"111111111",
  8592=>"111000000",
  8593=>"111111111",
  8594=>"010100111",
  8595=>"111111111",
  8596=>"000000000",
  8597=>"110000000",
  8598=>"100100111",
  8599=>"000000001",
  8600=>"111111111",
  8601=>"000000001",
  8602=>"000000111",
  8603=>"000000111",
  8604=>"000111000",
  8605=>"010010011",
  8606=>"000111111",
  8607=>"000000001",
  8608=>"001000000",
  8609=>"111111011",
  8610=>"111000100",
  8611=>"000000111",
  8612=>"000100111",
  8613=>"111111111",
  8614=>"000100111",
  8615=>"111000000",
  8616=>"000111111",
  8617=>"111100100",
  8618=>"111001001",
  8619=>"111111111",
  8620=>"111011001",
  8621=>"111111000",
  8622=>"111111100",
  8623=>"010111111",
  8624=>"111110111",
  8625=>"111000011",
  8626=>"000000001",
  8627=>"111011000",
  8628=>"111101000",
  8629=>"111111011",
  8630=>"000000000",
  8631=>"000000000",
  8632=>"000000111",
  8633=>"111111011",
  8634=>"000000000",
  8635=>"001000000",
  8636=>"111111111",
  8637=>"100111111",
  8638=>"000000000",
  8639=>"001001001",
  8640=>"000100111",
  8641=>"000111011",
  8642=>"111111111",
  8643=>"110110111",
  8644=>"111001111",
  8645=>"011001001",
  8646=>"111110000",
  8647=>"111000000",
  8648=>"001000111",
  8649=>"111111100",
  8650=>"111000111",
  8651=>"000111111",
  8652=>"100000000",
  8653=>"111111110",
  8654=>"100000000",
  8655=>"110111111",
  8656=>"000101111",
  8657=>"000110111",
  8658=>"001111010",
  8659=>"000000000",
  8660=>"101110010",
  8661=>"111111110",
  8662=>"111110110",
  8663=>"001110111",
  8664=>"000001011",
  8665=>"111100000",
  8666=>"100100111",
  8667=>"111100100",
  8668=>"111011011",
  8669=>"111111100",
  8670=>"010011111",
  8671=>"111111000",
  8672=>"000001001",
  8673=>"100000000",
  8674=>"110011000",
  8675=>"101101000",
  8676=>"000000000",
  8677=>"000000110",
  8678=>"111111111",
  8679=>"111101111",
  8680=>"000100001",
  8681=>"111001000",
  8682=>"000111111",
  8683=>"111111111",
  8684=>"111111000",
  8685=>"100000100",
  8686=>"101111011",
  8687=>"000111111",
  8688=>"001110111",
  8689=>"111111111",
  8690=>"000000100",
  8691=>"000110111",
  8692=>"000001111",
  8693=>"000111111",
  8694=>"001111011",
  8695=>"011111101",
  8696=>"000101111",
  8697=>"001011011",
  8698=>"100000111",
  8699=>"111011000",
  8700=>"000000111",
  8701=>"111111111",
  8702=>"111011000",
  8703=>"001001001",
  8704=>"101111111",
  8705=>"100000001",
  8706=>"111111111",
  8707=>"000000111",
  8708=>"011111111",
  8709=>"100101111",
  8710=>"100100100",
  8711=>"010111111",
  8712=>"111001111",
  8713=>"101001111",
  8714=>"111101000",
  8715=>"000000001",
  8716=>"000011001",
  8717=>"100111111",
  8718=>"110111011",
  8719=>"000000110",
  8720=>"111000000",
  8721=>"000101101",
  8722=>"000100111",
  8723=>"111111111",
  8724=>"111111111",
  8725=>"111011111",
  8726=>"000000000",
  8727=>"110100100",
  8728=>"011011011",
  8729=>"001111110",
  8730=>"000000000",
  8731=>"100000100",
  8732=>"111111111",
  8733=>"000110011",
  8734=>"000000000",
  8735=>"111001101",
  8736=>"111111000",
  8737=>"000000000",
  8738=>"100000000",
  8739=>"111111000",
  8740=>"111111111",
  8741=>"111110110",
  8742=>"111101111",
  8743=>"111111111",
  8744=>"000000000",
  8745=>"000101100",
  8746=>"111111111",
  8747=>"110111111",
  8748=>"100101111",
  8749=>"000000000",
  8750=>"111010000",
  8751=>"001100110",
  8752=>"111111111",
  8753=>"111111111",
  8754=>"000000000",
  8755=>"111010110",
  8756=>"000000000",
  8757=>"110111000",
  8758=>"101000000",
  8759=>"111110101",
  8760=>"100111111",
  8761=>"111111110",
  8762=>"111111111",
  8763=>"111110110",
  8764=>"100000000",
  8765=>"111100100",
  8766=>"000000010",
  8767=>"100000000",
  8768=>"001001000",
  8769=>"000100000",
  8770=>"010000001",
  8771=>"111101111",
  8772=>"011000111",
  8773=>"111111111",
  8774=>"111111111",
  8775=>"100111111",
  8776=>"000000010",
  8777=>"000011111",
  8778=>"000000011",
  8779=>"000000010",
  8780=>"100000000",
  8781=>"011001111",
  8782=>"000111110",
  8783=>"000000000",
  8784=>"000000001",
  8785=>"000011111",
  8786=>"111111111",
  8787=>"010000000",
  8788=>"000100000",
  8789=>"000000000",
  8790=>"101000000",
  8791=>"010111010",
  8792=>"111111111",
  8793=>"000000000",
  8794=>"000000000",
  8795=>"110111111",
  8796=>"010000000",
  8797=>"111011111",
  8798=>"111000000",
  8799=>"000000110",
  8800=>"000000100",
  8801=>"000000000",
  8802=>"100100000",
  8803=>"000110000",
  8804=>"001011111",
  8805=>"000000000",
  8806=>"111101111",
  8807=>"001101101",
  8808=>"111111111",
  8809=>"000000000",
  8810=>"111111111",
  8811=>"000001101",
  8812=>"110111001",
  8813=>"100111110",
  8814=>"000000000",
  8815=>"001001111",
  8816=>"110111111",
  8817=>"111000000",
  8818=>"111111000",
  8819=>"111001000",
  8820=>"111111101",
  8821=>"011001001",
  8822=>"111010000",
  8823=>"110100000",
  8824=>"000000000",
  8825=>"010000111",
  8826=>"000000001",
  8827=>"111111111",
  8828=>"000000100",
  8829=>"000000001",
  8830=>"111101000",
  8831=>"000010000",
  8832=>"111111111",
  8833=>"111111000",
  8834=>"100111110",
  8835=>"110110000",
  8836=>"100100111",
  8837=>"000000100",
  8838=>"101000000",
  8839=>"111111111",
  8840=>"101111111",
  8841=>"001011011",
  8842=>"111111101",
  8843=>"100100110",
  8844=>"100000000",
  8845=>"111110111",
  8846=>"100111111",
  8847=>"101111111",
  8848=>"000000000",
  8849=>"100111111",
  8850=>"111101000",
  8851=>"011111111",
  8852=>"111111110",
  8853=>"010111111",
  8854=>"111111111",
  8855=>"101000001",
  8856=>"001001111",
  8857=>"110000000",
  8858=>"001001001",
  8859=>"000000111",
  8860=>"111110110",
  8861=>"011111111",
  8862=>"000000000",
  8863=>"100101111",
  8864=>"101001000",
  8865=>"000000000",
  8866=>"000000000",
  8867=>"011111101",
  8868=>"000000001",
  8869=>"000011111",
  8870=>"110111010",
  8871=>"000000000",
  8872=>"110110111",
  8873=>"001111011",
  8874=>"111111101",
  8875=>"111111111",
  8876=>"000000000",
  8877=>"000000011",
  8878=>"000000000",
  8879=>"110100111",
  8880=>"000010000",
  8881=>"111111111",
  8882=>"000000000",
  8883=>"000111111",
  8884=>"011111101",
  8885=>"111111111",
  8886=>"100000001",
  8887=>"000000101",
  8888=>"000000000",
  8889=>"000000000",
  8890=>"000000000",
  8891=>"000000001",
  8892=>"011000100",
  8893=>"111001000",
  8894=>"111111111",
  8895=>"001111111",
  8896=>"000000110",
  8897=>"111001000",
  8898=>"111111111",
  8899=>"111111110",
  8900=>"011001111",
  8901=>"001010011",
  8902=>"000000111",
  8903=>"000011011",
  8904=>"000001001",
  8905=>"111110110",
  8906=>"001001011",
  8907=>"101111111",
  8908=>"111110010",
  8909=>"000111111",
  8910=>"111110111",
  8911=>"000110100",
  8912=>"111111111",
  8913=>"100101101",
  8914=>"011001111",
  8915=>"001000000",
  8916=>"111111111",
  8917=>"000011001",
  8918=>"000000111",
  8919=>"111111010",
  8920=>"000000000",
  8921=>"111000000",
  8922=>"000000000",
  8923=>"111001011",
  8924=>"101000001",
  8925=>"110110110",
  8926=>"000001111",
  8927=>"110000000",
  8928=>"111111111",
  8929=>"111111111",
  8930=>"011001101",
  8931=>"111111111",
  8932=>"001001001",
  8933=>"111000100",
  8934=>"011001000",
  8935=>"000000000",
  8936=>"101100110",
  8937=>"100110111",
  8938=>"100110111",
  8939=>"001100110",
  8940=>"011000000",
  8941=>"111101111",
  8942=>"100101111",
  8943=>"001001010",
  8944=>"000000000",
  8945=>"000000100",
  8946=>"111111111",
  8947=>"111111111",
  8948=>"000001000",
  8949=>"000001001",
  8950=>"100000000",
  8951=>"111111111",
  8952=>"110111111",
  8953=>"111111101",
  8954=>"111001011",
  8955=>"110111110",
  8956=>"000000000",
  8957=>"111000001",
  8958=>"101101111",
  8959=>"000111000",
  8960=>"001001001",
  8961=>"011000000",
  8962=>"001111111",
  8963=>"000000000",
  8964=>"110100110",
  8965=>"111111101",
  8966=>"110000000",
  8967=>"111111000",
  8968=>"111100011",
  8969=>"001101101",
  8970=>"111001101",
  8971=>"111111010",
  8972=>"000000000",
  8973=>"100000000",
  8974=>"000010100",
  8975=>"000000000",
  8976=>"000001111",
  8977=>"111000111",
  8978=>"110111001",
  8979=>"010000000",
  8980=>"101111111",
  8981=>"101101101",
  8982=>"000000001",
  8983=>"111111111",
  8984=>"000000111",
  8985=>"111111111",
  8986=>"000000000",
  8987=>"101000001",
  8988=>"000000000",
  8989=>"001101111",
  8990=>"000000101",
  8991=>"111111000",
  8992=>"110000000",
  8993=>"000000100",
  8994=>"111000001",
  8995=>"000000010",
  8996=>"000000000",
  8997=>"110110000",
  8998=>"000000000",
  8999=>"111111111",
  9000=>"000000000",
  9001=>"000000001",
  9002=>"000000000",
  9003=>"111111111",
  9004=>"111111111",
  9005=>"010011011",
  9006=>"000000111",
  9007=>"000000000",
  9008=>"011011111",
  9009=>"111111001",
  9010=>"000011000",
  9011=>"000111111",
  9012=>"110110110",
  9013=>"011011011",
  9014=>"010011011",
  9015=>"111001001",
  9016=>"000000010",
  9017=>"000000000",
  9018=>"001000000",
  9019=>"000000001",
  9020=>"011001000",
  9021=>"110000100",
  9022=>"011000101",
  9023=>"101001001",
  9024=>"011111000",
  9025=>"111111000",
  9026=>"111111110",
  9027=>"000010000",
  9028=>"000010010",
  9029=>"111111111",
  9030=>"111111111",
  9031=>"000000000",
  9032=>"110000000",
  9033=>"111101111",
  9034=>"000000000",
  9035=>"100100000",
  9036=>"011001111",
  9037=>"101111111",
  9038=>"001000000",
  9039=>"100110100",
  9040=>"000110110",
  9041=>"000000000",
  9042=>"111000010",
  9043=>"000000000",
  9044=>"111111111",
  9045=>"111111101",
  9046=>"111000000",
  9047=>"111100100",
  9048=>"000111111",
  9049=>"000000000",
  9050=>"111111000",
  9051=>"100100111",
  9052=>"111111111",
  9053=>"111111111",
  9054=>"111101101",
  9055=>"000000011",
  9056=>"000000000",
  9057=>"000100111",
  9058=>"000000000",
  9059=>"000000000",
  9060=>"000000110",
  9061=>"010111001",
  9062=>"111111111",
  9063=>"001000000",
  9064=>"011011001",
  9065=>"000000000",
  9066=>"000111111",
  9067=>"100110111",
  9068=>"001001001",
  9069=>"001111111",
  9070=>"000001101",
  9071=>"001000000",
  9072=>"111111111",
  9073=>"111111010",
  9074=>"000000100",
  9075=>"010000000",
  9076=>"111111111",
  9077=>"000100000",
  9078=>"111111111",
  9079=>"111110111",
  9080=>"000000000",
  9081=>"111111111",
  9082=>"000000111",
  9083=>"010111000",
  9084=>"000000000",
  9085=>"010010000",
  9086=>"111111100",
  9087=>"000011111",
  9088=>"011001000",
  9089=>"111000000",
  9090=>"111111111",
  9091=>"111111111",
  9092=>"000100111",
  9093=>"000000000",
  9094=>"000000000",
  9095=>"110110110",
  9096=>"000000011",
  9097=>"111011110",
  9098=>"111111111",
  9099=>"000000000",
  9100=>"111111111",
  9101=>"000000000",
  9102=>"100100100",
  9103=>"000000110",
  9104=>"000111111",
  9105=>"111111001",
  9106=>"001000001",
  9107=>"100110000",
  9108=>"111111111",
  9109=>"000111111",
  9110=>"001111001",
  9111=>"000001000",
  9112=>"111111111",
  9113=>"000000000",
  9114=>"000011011",
  9115=>"000000110",
  9116=>"111111111",
  9117=>"010011000",
  9118=>"111111011",
  9119=>"000000000",
  9120=>"111111111",
  9121=>"111011001",
  9122=>"000000000",
  9123=>"111000000",
  9124=>"000000000",
  9125=>"111111111",
  9126=>"110111110",
  9127=>"011001111",
  9128=>"111001111",
  9129=>"000000010",
  9130=>"000111110",
  9131=>"110100111",
  9132=>"111111111",
  9133=>"101111111",
  9134=>"111011001",
  9135=>"111111111",
  9136=>"111111111",
  9137=>"111001011",
  9138=>"111111111",
  9139=>"111111100",
  9140=>"110100111",
  9141=>"100110100",
  9142=>"111000000",
  9143=>"100000101",
  9144=>"111111111",
  9145=>"000111111",
  9146=>"001001000",
  9147=>"010110110",
  9148=>"111000100",
  9149=>"111111111",
  9150=>"011011000",
  9151=>"010010000",
  9152=>"111110111",
  9153=>"111111100",
  9154=>"000000000",
  9155=>"110000111",
  9156=>"111110111",
  9157=>"111110000",
  9158=>"111111111",
  9159=>"011111111",
  9160=>"111110110",
  9161=>"100100000",
  9162=>"000001011",
  9163=>"111111111",
  9164=>"111111111",
  9165=>"000100100",
  9166=>"000011000",
  9167=>"000011111",
  9168=>"110111110",
  9169=>"000000000",
  9170=>"001111111",
  9171=>"100101001",
  9172=>"000000000",
  9173=>"100100000",
  9174=>"001000000",
  9175=>"100100100",
  9176=>"111001001",
  9177=>"101111110",
  9178=>"111111111",
  9179=>"111100000",
  9180=>"000001001",
  9181=>"111000111",
  9182=>"111110111",
  9183=>"011011001",
  9184=>"001000010",
  9185=>"000000000",
  9186=>"000000000",
  9187=>"110111111",
  9188=>"111110111",
  9189=>"000100100",
  9190=>"000000011",
  9191=>"111111111",
  9192=>"010110110",
  9193=>"000000000",
  9194=>"010000000",
  9195=>"111111000",
  9196=>"101111111",
  9197=>"100100110",
  9198=>"110100111",
  9199=>"111000000",
  9200=>"010000000",
  9201=>"111111111",
  9202=>"000000000",
  9203=>"101111010",
  9204=>"101011111",
  9205=>"111111111",
  9206=>"000011000",
  9207=>"000000010",
  9208=>"000010010",
  9209=>"000000100",
  9210=>"111111111",
  9211=>"000000000",
  9212=>"100111111",
  9213=>"011011111",
  9214=>"101010000",
  9215=>"000000010",
  9216=>"000010111",
  9217=>"111111110",
  9218=>"000000001",
  9219=>"111111111",
  9220=>"011100100",
  9221=>"110011111",
  9222=>"100111111",
  9223=>"111111111",
  9224=>"111111101",
  9225=>"111000000",
  9226=>"000100111",
  9227=>"111110000",
  9228=>"000111110",
  9229=>"111111011",
  9230=>"111110110",
  9231=>"111110111",
  9232=>"000000011",
  9233=>"000000000",
  9234=>"000000000",
  9235=>"111111111",
  9236=>"111101000",
  9237=>"111111110",
  9238=>"111111000",
  9239=>"110111000",
  9240=>"100010111",
  9241=>"111001000",
  9242=>"111111001",
  9243=>"100100111",
  9244=>"000000000",
  9245=>"000000111",
  9246=>"011111001",
  9247=>"000100101",
  9248=>"111000000",
  9249=>"111111000",
  9250=>"100100000",
  9251=>"011111111",
  9252=>"000000111",
  9253=>"111111111",
  9254=>"001111111",
  9255=>"001001100",
  9256=>"001001000",
  9257=>"110110000",
  9258=>"000000000",
  9259=>"110000000",
  9260=>"111001001",
  9261=>"100110000",
  9262=>"000000111",
  9263=>"111100000",
  9264=>"011111111",
  9265=>"000000101",
  9266=>"000000000",
  9267=>"110100100",
  9268=>"010000000",
  9269=>"000000100",
  9270=>"000000000",
  9271=>"110110110",
  9272=>"000000111",
  9273=>"001000111",
  9274=>"111111111",
  9275=>"000000000",
  9276=>"000100100",
  9277=>"001111111",
  9278=>"000100111",
  9279=>"111111110",
  9280=>"000000001",
  9281=>"111000100",
  9282=>"000000000",
  9283=>"111011111",
  9284=>"001001100",
  9285=>"111111111",
  9286=>"111000000",
  9287=>"111111111",
  9288=>"100000000",
  9289=>"001101111",
  9290=>"010011111",
  9291=>"111000000",
  9292=>"000010000",
  9293=>"001101101",
  9294=>"111000000",
  9295=>"000000000",
  9296=>"000000000",
  9297=>"000000000",
  9298=>"000011000",
  9299=>"111101110",
  9300=>"000000000",
  9301=>"100000000",
  9302=>"001111101",
  9303=>"111011111",
  9304=>"110110111",
  9305=>"101111111",
  9306=>"101111111",
  9307=>"001000101",
  9308=>"111111111",
  9309=>"001001111",
  9310=>"110110000",
  9311=>"000000000",
  9312=>"000000000",
  9313=>"100110110",
  9314=>"111000110",
  9315=>"001111111",
  9316=>"111111000",
  9317=>"001000000",
  9318=>"001000000",
  9319=>"000000000",
  9320=>"000000111",
  9321=>"000011111",
  9322=>"101001011",
  9323=>"111111111",
  9324=>"110111101",
  9325=>"100000100",
  9326=>"000000010",
  9327=>"000000011",
  9328=>"111011011",
  9329=>"000001000",
  9330=>"001000000",
  9331=>"111000100",
  9332=>"100100000",
  9333=>"011101101",
  9334=>"111111000",
  9335=>"100111111",
  9336=>"111111110",
  9337=>"111111111",
  9338=>"001001101",
  9339=>"000000000",
  9340=>"110100000",
  9341=>"111111111",
  9342=>"001001101",
  9343=>"111111011",
  9344=>"000000000",
  9345=>"000011111",
  9346=>"000000001",
  9347=>"101100100",
  9348=>"100000000",
  9349=>"001000000",
  9350=>"000110111",
  9351=>"000011000",
  9352=>"111111011",
  9353=>"110111111",
  9354=>"000000000",
  9355=>"111101101",
  9356=>"001000000",
  9357=>"111111111",
  9358=>"110110000",
  9359=>"111101101",
  9360=>"110111111",
  9361=>"000000100",
  9362=>"010111111",
  9363=>"111111011",
  9364=>"000000100",
  9365=>"000000110",
  9366=>"011010000",
  9367=>"000111111",
  9368=>"000001000",
  9369=>"111111111",
  9370=>"000011111",
  9371=>"110000000",
  9372=>"111111110",
  9373=>"000000001",
  9374=>"001001000",
  9375=>"000000000",
  9376=>"110100111",
  9377=>"111011010",
  9378=>"000001100",
  9379=>"111111011",
  9380=>"000001000",
  9381=>"101111111",
  9382=>"111111111",
  9383=>"000000011",
  9384=>"001100000",
  9385=>"000000000",
  9386=>"000000000",
  9387=>"000000100",
  9388=>"101000100",
  9389=>"000000000",
  9390=>"111111111",
  9391=>"001001000",
  9392=>"111111111",
  9393=>"100111111",
  9394=>"111111111",
  9395=>"000000000",
  9396=>"111101101",
  9397=>"111111101",
  9398=>"000001001",
  9399=>"111011000",
  9400=>"101110111",
  9401=>"000000000",
  9402=>"000000101",
  9403=>"101001100",
  9404=>"111110111",
  9405=>"110111111",
  9406=>"000000000",
  9407=>"111011011",
  9408=>"000000000",
  9409=>"110110110",
  9410=>"111111011",
  9411=>"001000000",
  9412=>"000000011",
  9413=>"010011011",
  9414=>"001000001",
  9415=>"000000110",
  9416=>"000000000",
  9417=>"111111111",
  9418=>"000000010",
  9419=>"101001111",
  9420=>"000001100",
  9421=>"001000111",
  9422=>"101001000",
  9423=>"000000000",
  9424=>"000000100",
  9425=>"011011111",
  9426=>"000000000",
  9427=>"100100000",
  9428=>"110111011",
  9429=>"111111010",
  9430=>"111111111",
  9431=>"000000111",
  9432=>"010010010",
  9433=>"111111101",
  9434=>"000000111",
  9435=>"000000000",
  9436=>"000100101",
  9437=>"000000000",
  9438=>"000000000",
  9439=>"111111011",
  9440=>"000000000",
  9441=>"010000000",
  9442=>"001011000",
  9443=>"011011000",
  9444=>"000000000",
  9445=>"000000111",
  9446=>"000110111",
  9447=>"110111111",
  9448=>"000001000",
  9449=>"100000001",
  9450=>"111000000",
  9451=>"111111000",
  9452=>"000000000",
  9453=>"000010000",
  9454=>"001100000",
  9455=>"000000000",
  9456=>"001000000",
  9457=>"110111111",
  9458=>"011110111",
  9459=>"111111101",
  9460=>"111111111",
  9461=>"000000000",
  9462=>"100110110",
  9463=>"000000000",
  9464=>"000000001",
  9465=>"111111111",
  9466=>"000000000",
  9467=>"101101111",
  9468=>"100100000",
  9469=>"111011100",
  9470=>"000001111",
  9471=>"100100101",
  9472=>"011111001",
  9473=>"110110110",
  9474=>"111110000",
  9475=>"111000110",
  9476=>"111111111",
  9477=>"000000000",
  9478=>"000000000",
  9479=>"000110110",
  9480=>"000000110",
  9481=>"000000000",
  9482=>"001011100",
  9483=>"111111001",
  9484=>"000000000",
  9485=>"000000010",
  9486=>"111111001",
  9487=>"101100100",
  9488=>"000010011",
  9489=>"000000000",
  9490=>"001001000",
  9491=>"111010001",
  9492=>"000000011",
  9493=>"000010111",
  9494=>"111110100",
  9495=>"100110111",
  9496=>"001000000",
  9497=>"000000001",
  9498=>"111111011",
  9499=>"000111111",
  9500=>"000000000",
  9501=>"000000000",
  9502=>"111000001",
  9503=>"111111111",
  9504=>"111101111",
  9505=>"111110110",
  9506=>"111111111",
  9507=>"011010010",
  9508=>"111111011",
  9509=>"111101100",
  9510=>"111111111",
  9511=>"011011111",
  9512=>"000110010",
  9513=>"111111111",
  9514=>"111010000",
  9515=>"000000001",
  9516=>"000100101",
  9517=>"011000110",
  9518=>"000000000",
  9519=>"001001111",
  9520=>"000010011",
  9521=>"000000011",
  9522=>"000000000",
  9523=>"111110000",
  9524=>"000000000",
  9525=>"110111111",
  9526=>"000000011",
  9527=>"011001000",
  9528=>"000000000",
  9529=>"101000000",
  9530=>"000000000",
  9531=>"001000000",
  9532=>"110111111",
  9533=>"000000000",
  9534=>"000000000",
  9535=>"111111000",
  9536=>"010000000",
  9537=>"111111001",
  9538=>"100110100",
  9539=>"010000000",
  9540=>"000000000",
  9541=>"111000000",
  9542=>"001000110",
  9543=>"100100000",
  9544=>"111111100",
  9545=>"111110110",
  9546=>"111000000",
  9547=>"111001011",
  9548=>"000000000",
  9549=>"111110111",
  9550=>"000100000",
  9551=>"001001001",
  9552=>"000100100",
  9553=>"111101101",
  9554=>"000000111",
  9555=>"111111111",
  9556=>"001000111",
  9557=>"000110110",
  9558=>"111111111",
  9559=>"001111110",
  9560=>"000000011",
  9561=>"001000000",
  9562=>"110000100",
  9563=>"111101111",
  9564=>"110000000",
  9565=>"000000111",
  9566=>"000000000",
  9567=>"000000000",
  9568=>"111111111",
  9569=>"000110110",
  9570=>"010110011",
  9571=>"000100111",
  9572=>"111111111",
  9573=>"111011000",
  9574=>"000110111",
  9575=>"001000000",
  9576=>"010011011",
  9577=>"001011000",
  9578=>"111111111",
  9579=>"111010010",
  9580=>"001011000",
  9581=>"101111010",
  9582=>"000000000",
  9583=>"000000000",
  9584=>"000000000",
  9585=>"111111000",
  9586=>"111111111",
  9587=>"111101100",
  9588=>"100101101",
  9589=>"100000000",
  9590=>"001011000",
  9591=>"000000000",
  9592=>"000000000",
  9593=>"111011000",
  9594=>"111111111",
  9595=>"111111011",
  9596=>"000100111",
  9597=>"111110111",
  9598=>"011111110",
  9599=>"000000000",
  9600=>"011000110",
  9601=>"000000000",
  9602=>"111111111",
  9603=>"100000000",
  9604=>"101001101",
  9605=>"000000101",
  9606=>"000000000",
  9607=>"000011110",
  9608=>"000000000",
  9609=>"001011111",
  9610=>"000000000",
  9611=>"111101101",
  9612=>"000100111",
  9613=>"111000000",
  9614=>"000000000",
  9615=>"111011011",
  9616=>"111111111",
  9617=>"000011011",
  9618=>"000000000",
  9619=>"000110110",
  9620=>"101111111",
  9621=>"000111111",
  9622=>"111101111",
  9623=>"111111111",
  9624=>"000000000",
  9625=>"000000110",
  9626=>"111111100",
  9627=>"011111111",
  9628=>"111111111",
  9629=>"010000000",
  9630=>"011111111",
  9631=>"110110000",
  9632=>"111111111",
  9633=>"000100100",
  9634=>"011000100",
  9635=>"000000111",
  9636=>"011000100",
  9637=>"101101111",
  9638=>"001000000",
  9639=>"111011010",
  9640=>"000010111",
  9641=>"111111100",
  9642=>"001111111",
  9643=>"011001000",
  9644=>"110000000",
  9645=>"000011000",
  9646=>"001100111",
  9647=>"000000011",
  9648=>"000000111",
  9649=>"110110110",
  9650=>"001001000",
  9651=>"000011111",
  9652=>"111000011",
  9653=>"011001101",
  9654=>"111010001",
  9655=>"101101111",
  9656=>"101111111",
  9657=>"111110110",
  9658=>"000110110",
  9659=>"010000000",
  9660=>"001000000",
  9661=>"001000100",
  9662=>"001000001",
  9663=>"001001001",
  9664=>"111001000",
  9665=>"010010000",
  9666=>"000000000",
  9667=>"111111010",
  9668=>"111111111",
  9669=>"000010001",
  9670=>"010000000",
  9671=>"101101111",
  9672=>"001000000",
  9673=>"000000011",
  9674=>"000000000",
  9675=>"010111111",
  9676=>"100100000",
  9677=>"111111010",
  9678=>"110010010",
  9679=>"111100000",
  9680=>"111000000",
  9681=>"011111000",
  9682=>"010010111",
  9683=>"000100100",
  9684=>"110110111",
  9685=>"100111110",
  9686=>"000101111",
  9687=>"111111111",
  9688=>"111111000",
  9689=>"110001011",
  9690=>"110010000",
  9691=>"011011111",
  9692=>"010000000",
  9693=>"000000111",
  9694=>"110110100",
  9695=>"001000100",
  9696=>"111111111",
  9697=>"000000110",
  9698=>"000001001",
  9699=>"111111010",
  9700=>"010000000",
  9701=>"010000000",
  9702=>"000000001",
  9703=>"110110010",
  9704=>"001001001",
  9705=>"111111111",
  9706=>"000000000",
  9707=>"001000000",
  9708=>"001000000",
  9709=>"000000110",
  9710=>"011011111",
  9711=>"000000111",
  9712=>"000000000",
  9713=>"000111111",
  9714=>"001100001",
  9715=>"111111111",
  9716=>"001001000",
  9717=>"111111110",
  9718=>"110111111",
  9719=>"100010000",
  9720=>"001101111",
  9721=>"000000000",
  9722=>"111111111",
  9723=>"111111110",
  9724=>"001000100",
  9725=>"000000000",
  9726=>"011000011",
  9727=>"111000000",
  9728=>"000000000",
  9729=>"111111011",
  9730=>"011000000",
  9731=>"000010001",
  9732=>"100001001",
  9733=>"000000000",
  9734=>"000001011",
  9735=>"111111111",
  9736=>"000000000",
  9737=>"011111000",
  9738=>"111000000",
  9739=>"011001101",
  9740=>"000000001",
  9741=>"000111111",
  9742=>"100110111",
  9743=>"001001111",
  9744=>"001111111",
  9745=>"000010111",
  9746=>"111111111",
  9747=>"000000000",
  9748=>"001001111",
  9749=>"000000000",
  9750=>"000000000",
  9751=>"111111001",
  9752=>"100000100",
  9753=>"111100100",
  9754=>"000000100",
  9755=>"100100100",
  9756=>"111100000",
  9757=>"001001111",
  9758=>"110111111",
  9759=>"101000000",
  9760=>"111111111",
  9761=>"000000000",
  9762=>"111111111",
  9763=>"111001011",
  9764=>"111111011",
  9765=>"000000100",
  9766=>"011111111",
  9767=>"111111111",
  9768=>"000000100",
  9769=>"001000000",
  9770=>"000000001",
  9771=>"100000111",
  9772=>"111111111",
  9773=>"110110000",
  9774=>"111111111",
  9775=>"000010000",
  9776=>"000000100",
  9777=>"101001001",
  9778=>"001000000",
  9779=>"111101111",
  9780=>"110111111",
  9781=>"001110000",
  9782=>"111001001",
  9783=>"000110100",
  9784=>"000000001",
  9785=>"100001111",
  9786=>"000000000",
  9787=>"111111111",
  9788=>"111111111",
  9789=>"000000000",
  9790=>"000000100",
  9791=>"000001111",
  9792=>"000000001",
  9793=>"011001011",
  9794=>"111111101",
  9795=>"111111111",
  9796=>"010111111",
  9797=>"000000001",
  9798=>"000000000",
  9799=>"000010010",
  9800=>"001001011",
  9801=>"110000110",
  9802=>"011011111",
  9803=>"011111111",
  9804=>"000000110",
  9805=>"000000000",
  9806=>"000001101",
  9807=>"111111111",
  9808=>"111001000",
  9809=>"111001111",
  9810=>"111111111",
  9811=>"010010000",
  9812=>"000001000",
  9813=>"000000000",
  9814=>"000000000",
  9815=>"101111111",
  9816=>"000000000",
  9817=>"100000000",
  9818=>"000000000",
  9819=>"011011001",
  9820=>"010000000",
  9821=>"000000000",
  9822=>"111100000",
  9823=>"111000000",
  9824=>"000000000",
  9825=>"000000111",
  9826=>"110110110",
  9827=>"000000000",
  9828=>"111111000",
  9829=>"001000000",
  9830=>"111111110",
  9831=>"110111001",
  9832=>"000000000",
  9833=>"000000000",
  9834=>"111111000",
  9835=>"111111100",
  9836=>"111001100",
  9837=>"111111011",
  9838=>"101101000",
  9839=>"111111111",
  9840=>"000000000",
  9841=>"111100111",
  9842=>"000000000",
  9843=>"111111111",
  9844=>"110100000",
  9845=>"110111011",
  9846=>"111110110",
  9847=>"000000000",
  9848=>"111111111",
  9849=>"101001111",
  9850=>"111111000",
  9851=>"000000000",
  9852=>"010011111",
  9853=>"111111001",
  9854=>"000011111",
  9855=>"000000000",
  9856=>"000000000",
  9857=>"111111111",
  9858=>"010010000",
  9859=>"111111011",
  9860=>"000010110",
  9861=>"111111111",
  9862=>"000000000",
  9863=>"111011001",
  9864=>"111111111",
  9865=>"000000111",
  9866=>"000000000",
  9867=>"111101101",
  9868=>"111111001",
  9869=>"111111111",
  9870=>"100111111",
  9871=>"100000000",
  9872=>"000010111",
  9873=>"000000000",
  9874=>"110000000",
  9875=>"111111111",
  9876=>"100000000",
  9877=>"001001011",
  9878=>"000000100",
  9879=>"000000000",
  9880=>"000000111",
  9881=>"100111111",
  9882=>"000000001",
  9883=>"011000111",
  9884=>"111111100",
  9885=>"110100100",
  9886=>"111111011",
  9887=>"111111111",
  9888=>"000000000",
  9889=>"000001101",
  9890=>"111110000",
  9891=>"000000000",
  9892=>"000000001",
  9893=>"000010011",
  9894=>"111111111",
  9895=>"111111000",
  9896=>"111111111",
  9897=>"000100111",
  9898=>"000000000",
  9899=>"100000100",
  9900=>"001101000",
  9901=>"111011011",
  9902=>"111101111",
  9903=>"111111101",
  9904=>"000000000",
  9905=>"011011011",
  9906=>"000000000",
  9907=>"111111111",
  9908=>"001001000",
  9909=>"000000000",
  9910=>"000000000",
  9911=>"000000110",
  9912=>"111111111",
  9913=>"110111111",
  9914=>"010001000",
  9915=>"011001111",
  9916=>"100000000",
  9917=>"100111111",
  9918=>"111111111",
  9919=>"000000000",
  9920=>"000001101",
  9921=>"111000000",
  9922=>"111111000",
  9923=>"111111111",
  9924=>"110111111",
  9925=>"111011000",
  9926=>"111111111",
  9927=>"000000000",
  9928=>"000110110",
  9929=>"111111111",
  9930=>"110101000",
  9931=>"011011000",
  9932=>"000100000",
  9933=>"000000000",
  9934=>"000011111",
  9935=>"111111111",
  9936=>"010000100",
  9937=>"000000000",
  9938=>"111000000",
  9939=>"101000000",
  9940=>"100000100",
  9941=>"111111111",
  9942=>"000000010",
  9943=>"000000000",
  9944=>"111111100",
  9945=>"100110000",
  9946=>"100100100",
  9947=>"100000000",
  9948=>"001000000",
  9949=>"000000000",
  9950=>"111111111",
  9951=>"100101100",
  9952=>"000000111",
  9953=>"000001001",
  9954=>"111110000",
  9955=>"000000000",
  9956=>"000000000",
  9957=>"111111111",
  9958=>"111111111",
  9959=>"100100110",
  9960=>"000000001",
  9961=>"001000000",
  9962=>"111111111",
  9963=>"111111111",
  9964=>"011111111",
  9965=>"000100111",
  9966=>"000111111",
  9967=>"011111111",
  9968=>"001101000",
  9969=>"010000000",
  9970=>"111111111",
  9971=>"001001000",
  9972=>"000111111",
  9973=>"110100000",
  9974=>"111100000",
  9975=>"000000000",
  9976=>"111111111",
  9977=>"000000000",
  9978=>"000000000",
  9979=>"001011111",
  9980=>"000000000",
  9981=>"000000110",
  9982=>"111011000",
  9983=>"111111111",
  9984=>"111111101",
  9985=>"000000011",
  9986=>"000000000",
  9987=>"001111111",
  9988=>"111100100",
  9989=>"000000000",
  9990=>"000000000",
  9991=>"000000111",
  9992=>"100001111",
  9993=>"010000111",
  9994=>"111111111",
  9995=>"000000110",
  9996=>"000000000",
  9997=>"111111111",
  9998=>"000000000",
  9999=>"000000000",
  10000=>"001001001",
  10001=>"000000000",
  10002=>"100000000",
  10003=>"110110111",
  10004=>"111101111",
  10005=>"000000000",
  10006=>"111111000",
  10007=>"110010000",
  10008=>"100100101",
  10009=>"111111111",
  10010=>"000000001",
  10011=>"100000000",
  10012=>"010010000",
  10013=>"000000000",
  10014=>"000000000",
  10015=>"111011001",
  10016=>"000110011",
  10017=>"010011000",
  10018=>"111111111",
  10019=>"001111111",
  10020=>"110000011",
  10021=>"000000000",
  10022=>"000000000",
  10023=>"001001000",
  10024=>"000000000",
  10025=>"000000000",
  10026=>"111111111",
  10027=>"111111000",
  10028=>"011111000",
  10029=>"000000000",
  10030=>"111110111",
  10031=>"101001001",
  10032=>"111111110",
  10033=>"000010011",
  10034=>"111111111",
  10035=>"111111010",
  10036=>"000000110",
  10037=>"111111110",
  10038=>"111111111",
  10039=>"111001001",
  10040=>"000000000",
  10041=>"110111111",
  10042=>"000010010",
  10043=>"000000000",
  10044=>"111101101",
  10045=>"001000000",
  10046=>"000000000",
  10047=>"000000100",
  10048=>"001000110",
  10049=>"000000010",
  10050=>"000000011",
  10051=>"111111111",
  10052=>"000111111",
  10053=>"101111111",
  10054=>"101111111",
  10055=>"000000000",
  10056=>"001011011",
  10057=>"000000000",
  10058=>"111110100",
  10059=>"110100110",
  10060=>"000000000",
  10061=>"000000000",
  10062=>"000000100",
  10063=>"011001000",
  10064=>"011001000",
  10065=>"111111110",
  10066=>"111111111",
  10067=>"111111000",
  10068=>"000000000",
  10069=>"011011011",
  10070=>"000000000",
  10071=>"101000000",
  10072=>"000000000",
  10073=>"011010000",
  10074=>"001001001",
  10075=>"101111111",
  10076=>"000000000",
  10077=>"000000000",
  10078=>"111111000",
  10079=>"111111011",
  10080=>"000001111",
  10081=>"000000000",
  10082=>"000101110",
  10083=>"000101111",
  10084=>"111011001",
  10085=>"101000000",
  10086=>"000000000",
  10087=>"110110000",
  10088=>"111111011",
  10089=>"111111111",
  10090=>"101001111",
  10091=>"000000100",
  10092=>"011111111",
  10093=>"111111111",
  10094=>"100100000",
  10095=>"000000000",
  10096=>"000000000",
  10097=>"110010000",
  10098=>"000000000",
  10099=>"110111110",
  10100=>"001001001",
  10101=>"100000000",
  10102=>"011000001",
  10103=>"111111111",
  10104=>"111111111",
  10105=>"000110111",
  10106=>"000000000",
  10107=>"000000000",
  10108=>"010010000",
  10109=>"000000000",
  10110=>"000000000",
  10111=>"111111111",
  10112=>"101000000",
  10113=>"001001101",
  10114=>"000000000",
  10115=>"001011110",
  10116=>"001111111",
  10117=>"000100100",
  10118=>"100110110",
  10119=>"111111100",
  10120=>"111111111",
  10121=>"001000111",
  10122=>"111111111",
  10123=>"000000000",
  10124=>"101011111",
  10125=>"100100100",
  10126=>"111111011",
  10127=>"000000000",
  10128=>"011111111",
  10129=>"111111111",
  10130=>"010000000",
  10131=>"111111111",
  10132=>"111000000",
  10133=>"011111011",
  10134=>"111110111",
  10135=>"000011011",
  10136=>"111111010",
  10137=>"101001001",
  10138=>"110110111",
  10139=>"111111111",
  10140=>"001101100",
  10141=>"000000000",
  10142=>"000000000",
  10143=>"100000110",
  10144=>"000000000",
  10145=>"000000000",
  10146=>"000000000",
  10147=>"011111111",
  10148=>"100101111",
  10149=>"000000000",
  10150=>"000000111",
  10151=>"100000000",
  10152=>"111001000",
  10153=>"000010001",
  10154=>"111111111",
  10155=>"010111000",
  10156=>"000000000",
  10157=>"011011111",
  10158=>"000111111",
  10159=>"000000000",
  10160=>"111111111",
  10161=>"001000001",
  10162=>"010111111",
  10163=>"000000000",
  10164=>"000000111",
  10165=>"100000000",
  10166=>"111111111",
  10167=>"110000000",
  10168=>"000111111",
  10169=>"010010000",
  10170=>"000000000",
  10171=>"000000000",
  10172=>"111111111",
  10173=>"110000101",
  10174=>"111101111",
  10175=>"111111111",
  10176=>"001111111",
  10177=>"100100111",
  10178=>"110111111",
  10179=>"000000000",
  10180=>"000000000",
  10181=>"111111100",
  10182=>"000000000",
  10183=>"000000000",
  10184=>"101111111",
  10185=>"100101000",
  10186=>"001001001",
  10187=>"111111111",
  10188=>"101000000",
  10189=>"000000001",
  10190=>"001111111",
  10191=>"000001110",
  10192=>"000111111",
  10193=>"100000000",
  10194=>"000000000",
  10195=>"111111111",
  10196=>"110110000",
  10197=>"111000000",
  10198=>"001001100",
  10199=>"110100111",
  10200=>"110110111",
  10201=>"000000000",
  10202=>"111111011",
  10203=>"111111000",
  10204=>"111000000",
  10205=>"011011001",
  10206=>"000000000",
  10207=>"101000000",
  10208=>"111111110",
  10209=>"110100000",
  10210=>"000000000",
  10211=>"000100101",
  10212=>"000000011",
  10213=>"011111011",
  10214=>"000000000",
  10215=>"000010000",
  10216=>"000000000",
  10217=>"111111111",
  10218=>"000110000",
  10219=>"000101111",
  10220=>"000000110",
  10221=>"000000100",
  10222=>"000001111",
  10223=>"101101111",
  10224=>"111111111",
  10225=>"000000011",
  10226=>"111111111",
  10227=>"111111111",
  10228=>"011011111",
  10229=>"000000111",
  10230=>"111000000",
  10231=>"000000000",
  10232=>"001000000",
  10233=>"111101101",
  10234=>"111111111",
  10235=>"000000000",
  10236=>"000000000",
  10237=>"100111100",
  10238=>"001001001",
  10239=>"000000000",
  10240=>"101111001",
  10241=>"000000000",
  10242=>"000000100",
  10243=>"000000000",
  10244=>"000000110",
  10245=>"100000100",
  10246=>"001101001",
  10247=>"111101101",
  10248=>"100111111",
  10249=>"110110100",
  10250=>"111111110",
  10251=>"111111111",
  10252=>"111110110",
  10253=>"111111111",
  10254=>"111101111",
  10255=>"111111011",
  10256=>"000000100",
  10257=>"000011111",
  10258=>"100000000",
  10259=>"111111111",
  10260=>"111111111",
  10261=>"000000000",
  10262=>"111111111",
  10263=>"110110110",
  10264=>"101101000",
  10265=>"100000000",
  10266=>"111111111",
  10267=>"000000001",
  10268=>"111111111",
  10269=>"011001001",
  10270=>"000100100",
  10271=>"000000000",
  10272=>"011110111",
  10273=>"000110100",
  10274=>"000000100",
  10275=>"111111011",
  10276=>"111111011",
  10277=>"000000000",
  10278=>"000000000",
  10279=>"000000000",
  10280=>"111111111",
  10281=>"000001001",
  10282=>"000110110",
  10283=>"111110100",
  10284=>"000000000",
  10285=>"000000101",
  10286=>"000000000",
  10287=>"111010000",
  10288=>"000000000",
  10289=>"000000000",
  10290=>"010010000",
  10291=>"000010010",
  10292=>"000000001",
  10293=>"001101111",
  10294=>"100000000",
  10295=>"101101011",
  10296=>"000000000",
  10297=>"010000000",
  10298=>"101100000",
  10299=>"010110000",
  10300=>"000000000",
  10301=>"010111111",
  10302=>"111111111",
  10303=>"000000000",
  10304=>"010000010",
  10305=>"001001001",
  10306=>"000000000",
  10307=>"000000110",
  10308=>"001001001",
  10309=>"111111000",
  10310=>"000000000",
  10311=>"111111111",
  10312=>"111111011",
  10313=>"111111000",
  10314=>"000000000",
  10315=>"111111101",
  10316=>"101111110",
  10317=>"000000000",
  10318=>"000100110",
  10319=>"111111001",
  10320=>"000000000",
  10321=>"111111111",
  10322=>"000000000",
  10323=>"111011111",
  10324=>"101000000",
  10325=>"000000000",
  10326=>"000101100",
  10327=>"000001111",
  10328=>"111111110",
  10329=>"111111111",
  10330=>"111111111",
  10331=>"100100100",
  10332=>"000000000",
  10333=>"010011011",
  10334=>"001000110",
  10335=>"111000110",
  10336=>"111111000",
  10337=>"000000100",
  10338=>"000000000",
  10339=>"000000111",
  10340=>"111111110",
  10341=>"111111111",
  10342=>"000000000",
  10343=>"110010000",
  10344=>"000001001",
  10345=>"100100111",
  10346=>"001011011",
  10347=>"111110100",
  10348=>"111111110",
  10349=>"111011000",
  10350=>"111001111",
  10351=>"111111111",
  10352=>"000000111",
  10353=>"000000011",
  10354=>"101100101",
  10355=>"000000000",
  10356=>"000000000",
  10357=>"000000111",
  10358=>"100111000",
  10359=>"111111111",
  10360=>"111010000",
  10361=>"111111111",
  10362=>"000000000",
  10363=>"111111111",
  10364=>"111111110",
  10365=>"000000000",
  10366=>"111111011",
  10367=>"000000000",
  10368=>"110111111",
  10369=>"111111111",
  10370=>"001000000",
  10371=>"000000100",
  10372=>"000000100",
  10373=>"111000000",
  10374=>"100111000",
  10375=>"000000110",
  10376=>"111111111",
  10377=>"000000000",
  10378=>"110111011",
  10379=>"111111111",
  10380=>"000000000",
  10381=>"000000000",
  10382=>"111011100",
  10383=>"000000000",
  10384=>"110010111",
  10385=>"000000000",
  10386=>"000111001",
  10387=>"000000000",
  10388=>"010011111",
  10389=>"000000001",
  10390=>"000000000",
  10391=>"001000000",
  10392=>"111011011",
  10393=>"000000000",
  10394=>"111111111",
  10395=>"000000000",
  10396=>"111111111",
  10397=>"100100100",
  10398=>"111111111",
  10399=>"011011011",
  10400=>"111111111",
  10401=>"000001000",
  10402=>"000000110",
  10403=>"110000000",
  10404=>"111101110",
  10405=>"111111111",
  10406=>"100000000",
  10407=>"110110000",
  10408=>"000000000",
  10409=>"000100111",
  10410=>"111000100",
  10411=>"110101000",
  10412=>"001111110",
  10413=>"100110110",
  10414=>"010000111",
  10415=>"111111111",
  10416=>"110111000",
  10417=>"111111111",
  10418=>"110100110",
  10419=>"111100001",
  10420=>"100000001",
  10421=>"111010000",
  10422=>"000100000",
  10423=>"000000000",
  10424=>"111111111",
  10425=>"111010111",
  10426=>"000000000",
  10427=>"100000101",
  10428=>"110000000",
  10429=>"000111111",
  10430=>"111111000",
  10431=>"000000010",
  10432=>"000000000",
  10433=>"110110110",
  10434=>"111111111",
  10435=>"111111111",
  10436=>"111010000",
  10437=>"000000000",
  10438=>"011001001",
  10439=>"000000000",
  10440=>"010010010",
  10441=>"100100100",
  10442=>"100100100",
  10443=>"010000000",
  10444=>"100000110",
  10445=>"100110111",
  10446=>"111011011",
  10447=>"000000000",
  10448=>"110111011",
  10449=>"000001111",
  10450=>"111111111",
  10451=>"000000110",
  10452=>"000000000",
  10453=>"111001001",
  10454=>"000000000",
  10455=>"000000000",
  10456=>"000000000",
  10457=>"111111111",
  10458=>"111111111",
  10459=>"000000000",
  10460=>"111111111",
  10461=>"000111111",
  10462=>"010000000",
  10463=>"100100110",
  10464=>"111111111",
  10465=>"000000000",
  10466=>"011001000",
  10467=>"110111111",
  10468=>"111111111",
  10469=>"100000000",
  10470=>"000110110",
  10471=>"000100111",
  10472=>"000001111",
  10473=>"111111111",
  10474=>"111111111",
  10475=>"000000000",
  10476=>"111111111",
  10477=>"111111011",
  10478=>"000000000",
  10479=>"010000000",
  10480=>"110110110",
  10481=>"000000000",
  10482=>"101000000",
  10483=>"000000001",
  10484=>"000000001",
  10485=>"000000000",
  10486=>"000000000",
  10487=>"111111111",
  10488=>"000000000",
  10489=>"000000000",
  10490=>"000110010",
  10491=>"000000000",
  10492=>"001001001",
  10493=>"111110111",
  10494=>"000110100",
  10495=>"111011001",
  10496=>"111111111",
  10497=>"010010100",
  10498=>"000000110",
  10499=>"110110110",
  10500=>"111111111",
  10501=>"000000000",
  10502=>"111111110",
  10503=>"000000000",
  10504=>"010000000",
  10505=>"000100100",
  10506=>"111111011",
  10507=>"011001111",
  10508=>"000000100",
  10509=>"111111111",
  10510=>"100010010",
  10511=>"011000000",
  10512=>"111111111",
  10513=>"111001111",
  10514=>"111111111",
  10515=>"001011111",
  10516=>"111111111",
  10517=>"000000011",
  10518=>"111111111",
  10519=>"111111111",
  10520=>"000000010",
  10521=>"111111111",
  10522=>"000000000",
  10523=>"000010011",
  10524=>"100100111",
  10525=>"000000000",
  10526=>"111111111",
  10527=>"110101011",
  10528=>"111111110",
  10529=>"111111011",
  10530=>"111111111",
  10531=>"000000111",
  10532=>"001010010",
  10533=>"110110110",
  10534=>"111111111",
  10535=>"111111110",
  10536=>"111111011",
  10537=>"111111111",
  10538=>"100100110",
  10539=>"111111111",
  10540=>"011111111",
  10541=>"000000001",
  10542=>"101101111",
  10543=>"000000000",
  10544=>"000100100",
  10545=>"100111111",
  10546=>"111111111",
  10547=>"111111111",
  10548=>"100100000",
  10549=>"000000000",
  10550=>"010111110",
  10551=>"111000000",
  10552=>"011001000",
  10553=>"011010111",
  10554=>"111111000",
  10555=>"001111111",
  10556=>"001111111",
  10557=>"100111110",
  10558=>"111111111",
  10559=>"000000001",
  10560=>"000000100",
  10561=>"000000000",
  10562=>"100000000",
  10563=>"111111111",
  10564=>"010010011",
  10565=>"000000000",
  10566=>"111111111",
  10567=>"000000000",
  10568=>"111111111",
  10569=>"110000000",
  10570=>"111101000",
  10571=>"010010010",
  10572=>"011010011",
  10573=>"111111111",
  10574=>"111111111",
  10575=>"000000000",
  10576=>"100000000",
  10577=>"000000000",
  10578=>"010000000",
  10579=>"000000000",
  10580=>"000000000",
  10581=>"011011011",
  10582=>"111111011",
  10583=>"000001000",
  10584=>"000101111",
  10585=>"110111111",
  10586=>"000010111",
  10587=>"111011011",
  10588=>"000000000",
  10589=>"000000000",
  10590=>"100001001",
  10591=>"010111110",
  10592=>"110111111",
  10593=>"100000111",
  10594=>"001001101",
  10595=>"000000000",
  10596=>"111101111",
  10597=>"000000000",
  10598=>"001111111",
  10599=>"110110110",
  10600=>"100100100",
  10601=>"000000000",
  10602=>"000001111",
  10603=>"111001001",
  10604=>"000100100",
  10605=>"001100100",
  10606=>"111111111",
  10607=>"001011111",
  10608=>"000000011",
  10609=>"111011011",
  10610=>"111000001",
  10611=>"000000000",
  10612=>"111001000",
  10613=>"000000000",
  10614=>"000000110",
  10615=>"000000000",
  10616=>"111001000",
  10617=>"000111111",
  10618=>"000000000",
  10619=>"111111111",
  10620=>"011011000",
  10621=>"000000000",
  10622=>"111111000",
  10623=>"001000000",
  10624=>"101001100",
  10625=>"000000100",
  10626=>"100100000",
  10627=>"000000000",
  10628=>"000000010",
  10629=>"000000000",
  10630=>"110111111",
  10631=>"111111001",
  10632=>"000000001",
  10633=>"000000000",
  10634=>"000000100",
  10635=>"001001000",
  10636=>"101101101",
  10637=>"001000000",
  10638=>"000000000",
  10639=>"000000000",
  10640=>"111111001",
  10641=>"100000000",
  10642=>"000000000",
  10643=>"000000100",
  10644=>"111111111",
  10645=>"000111111",
  10646=>"000000110",
  10647=>"001001000",
  10648=>"111011000",
  10649=>"111110110",
  10650=>"000000111",
  10651=>"011011110",
  10652=>"000000000",
  10653=>"000000000",
  10654=>"000011011",
  10655=>"000000100",
  10656=>"111111011",
  10657=>"111111110",
  10658=>"000000000",
  10659=>"111111111",
  10660=>"111111111",
  10661=>"000001111",
  10662=>"111111111",
  10663=>"000000000",
  10664=>"110000011",
  10665=>"000100000",
  10666=>"100000100",
  10667=>"101001000",
  10668=>"000000101",
  10669=>"000000001",
  10670=>"000000000",
  10671=>"111000000",
  10672=>"111111111",
  10673=>"000000000",
  10674=>"000000000",
  10675=>"000111111",
  10676=>"111111110",
  10677=>"000000000",
  10678=>"000000000",
  10679=>"111111111",
  10680=>"000000000",
  10681=>"000000000",
  10682=>"000000001",
  10683=>"111111110",
  10684=>"111111111",
  10685=>"100111100",
  10686=>"011001101",
  10687=>"101111100",
  10688=>"110110111",
  10689=>"000000000",
  10690=>"000100111",
  10691=>"111111100",
  10692=>"000110111",
  10693=>"101101001",
  10694=>"110000000",
  10695=>"111111111",
  10696=>"011111001",
  10697=>"111111111",
  10698=>"011001011",
  10699=>"011111011",
  10700=>"001000000",
  10701=>"110100111",
  10702=>"110111111",
  10703=>"100010000",
  10704=>"110000000",
  10705=>"000000010",
  10706=>"101000000",
  10707=>"000001001",
  10708=>"111110000",
  10709=>"001011000",
  10710=>"000111110",
  10711=>"000011001",
  10712=>"000000000",
  10713=>"000000000",
  10714=>"000000000",
  10715=>"011100110",
  10716=>"000000000",
  10717=>"111110110",
  10718=>"010000000",
  10719=>"000000000",
  10720=>"000000111",
  10721=>"010010000",
  10722=>"000000000",
  10723=>"111111101",
  10724=>"111111111",
  10725=>"001011001",
  10726=>"001011110",
  10727=>"000000000",
  10728=>"110111111",
  10729=>"101111111",
  10730=>"111011100",
  10731=>"000110111",
  10732=>"111111111",
  10733=>"000001001",
  10734=>"111111111",
  10735=>"000000000",
  10736=>"000000000",
  10737=>"000000000",
  10738=>"111111111",
  10739=>"000001011",
  10740=>"000000011",
  10741=>"011001001",
  10742=>"000000000",
  10743=>"101101101",
  10744=>"000000000",
  10745=>"100100000",
  10746=>"111111111",
  10747=>"111111111",
  10748=>"100101000",
  10749=>"100110100",
  10750=>"001000000",
  10751=>"111111111",
  10752=>"000000000",
  10753=>"000000000",
  10754=>"110101000",
  10755=>"011010111",
  10756=>"001111111",
  10757=>"111101100",
  10758=>"111110100",
  10759=>"000000000",
  10760=>"000000000",
  10761=>"111111101",
  10762=>"000100111",
  10763=>"111110110",
  10764=>"001011001",
  10765=>"011011011",
  10766=>"000000111",
  10767=>"000000000",
  10768=>"111111100",
  10769=>"111111111",
  10770=>"001011011",
  10771=>"111111111",
  10772=>"000000101",
  10773=>"111111111",
  10774=>"111111111",
  10775=>"110110110",
  10776=>"111111001",
  10777=>"000000000",
  10778=>"100000000",
  10779=>"001000000",
  10780=>"000000000",
  10781=>"000100001",
  10782=>"011111110",
  10783=>"000000000",
  10784=>"110000011",
  10785=>"000000000",
  10786=>"111110110",
  10787=>"011111111",
  10788=>"101111111",
  10789=>"001001011",
  10790=>"111111111",
  10791=>"000000000",
  10792=>"001000011",
  10793=>"111111111",
  10794=>"000000000",
  10795=>"101000000",
  10796=>"101111000",
  10797=>"111111110",
  10798=>"100000000",
  10799=>"110000000",
  10800=>"000000110",
  10801=>"111111101",
  10802=>"110110110",
  10803=>"111110110",
  10804=>"000000000",
  10805=>"111100110",
  10806=>"000010000",
  10807=>"010010110",
  10808=>"100101100",
  10809=>"000011111",
  10810=>"000001111",
  10811=>"100000111",
  10812=>"000000000",
  10813=>"000000100",
  10814=>"001001001",
  10815=>"000000000",
  10816=>"101011000",
  10817=>"101111111",
  10818=>"000100000",
  10819=>"110110000",
  10820=>"011000000",
  10821=>"011000000",
  10822=>"111011011",
  10823=>"000110111",
  10824=>"101000000",
  10825=>"111111111",
  10826=>"111111111",
  10827=>"100000000",
  10828=>"001100101",
  10829=>"000000111",
  10830=>"111000000",
  10831=>"111111111",
  10832=>"011001001",
  10833=>"000000100",
  10834=>"000000111",
  10835=>"110110010",
  10836=>"000000000",
  10837=>"111110110",
  10838=>"000000100",
  10839=>"011000000",
  10840=>"111111000",
  10841=>"111100100",
  10842=>"110110000",
  10843=>"000000000",
  10844=>"100111111",
  10845=>"011011011",
  10846=>"111101101",
  10847=>"000100011",
  10848=>"000000000",
  10849=>"111111111",
  10850=>"111111111",
  10851=>"000000111",
  10852=>"001000001",
  10853=>"111111111",
  10854=>"011000000",
  10855=>"100100000",
  10856=>"100110111",
  10857=>"000000101",
  10858=>"111111110",
  10859=>"000000000",
  10860=>"110110011",
  10861=>"111111111",
  10862=>"000000000",
  10863=>"000111111",
  10864=>"111111001",
  10865=>"010100100",
  10866=>"100001011",
  10867=>"000000010",
  10868=>"111010000",
  10869=>"000000000",
  10870=>"111100111",
  10871=>"100000000",
  10872=>"100100001",
  10873=>"110110111",
  10874=>"100000000",
  10875=>"111111111",
  10876=>"110110000",
  10877=>"011011011",
  10878=>"110000010",
  10879=>"100000000",
  10880=>"100000000",
  10881=>"110110000",
  10882=>"000000000",
  10883=>"011111111",
  10884=>"110111000",
  10885=>"000000000",
  10886=>"010010110",
  10887=>"010010000",
  10888=>"111110110",
  10889=>"110110111",
  10890=>"100111111",
  10891=>"000000000",
  10892=>"111111111",
  10893=>"111111111",
  10894=>"110110110",
  10895=>"111011001",
  10896=>"011010000",
  10897=>"000000000",
  10898=>"101101111",
  10899=>"000000000",
  10900=>"110111000",
  10901=>"010010000",
  10902=>"100000000",
  10903=>"111111111",
  10904=>"111111111",
  10905=>"000000000",
  10906=>"111111111",
  10907=>"111111101",
  10908=>"011011000",
  10909=>"000100011",
  10910=>"000100100",
  10911=>"000000101",
  10912=>"011001001",
  10913=>"011111111",
  10914=>"001000100",
  10915=>"111111011",
  10916=>"011011011",
  10917=>"011111000",
  10918=>"100000100",
  10919=>"001011110",
  10920=>"000000100",
  10921=>"011011001",
  10922=>"111111111",
  10923=>"000000100",
  10924=>"100000111",
  10925=>"000010110",
  10926=>"110010110",
  10927=>"000000011",
  10928=>"000000110",
  10929=>"011010111",
  10930=>"000000000",
  10931=>"010100000",
  10932=>"111000000",
  10933=>"111000100",
  10934=>"000011011",
  10935=>"000000001",
  10936=>"000011011",
  10937=>"101100110",
  10938=>"011000001",
  10939=>"110010000",
  10940=>"011001001",
  10941=>"011001000",
  10942=>"000000000",
  10943=>"100000000",
  10944=>"001111111",
  10945=>"000010110",
  10946=>"100000000",
  10947=>"000000000",
  10948=>"111111111",
  10949=>"111010000",
  10950=>"000000010",
  10951=>"100000100",
  10952=>"000000000",
  10953=>"111111100",
  10954=>"111101100",
  10955=>"111101100",
  10956=>"000001011",
  10957=>"111100000",
  10958=>"111000000",
  10959=>"001000000",
  10960=>"100000011",
  10961=>"111110111",
  10962=>"011011010",
  10963=>"000000000",
  10964=>"001011011",
  10965=>"111100100",
  10966=>"111111111",
  10967=>"000000000",
  10968=>"000111111",
  10969=>"011111111",
  10970=>"000000111",
  10971=>"001011011",
  10972=>"110000000",
  10973=>"000000110",
  10974=>"000000011",
  10975=>"000000011",
  10976=>"000000110",
  10977=>"111111111",
  10978=>"110110110",
  10979=>"001001001",
  10980=>"000000000",
  10981=>"000000110",
  10982=>"000000000",
  10983=>"111111111",
  10984=>"111111111",
  10985=>"100000000",
  10986=>"000000000",
  10987=>"000000000",
  10988=>"000000001",
  10989=>"000000011",
  10990=>"011000000",
  10991=>"010111111",
  10992=>"010000000",
  10993=>"110110111",
  10994=>"111111111",
  10995=>"010100101",
  10996=>"111110111",
  10997=>"000000000",
  10998=>"011011010",
  10999=>"000110111",
  11000=>"101100111",
  11001=>"111111111",
  11002=>"001111111",
  11003=>"000000000",
  11004=>"000000001",
  11005=>"011001001",
  11006=>"001111111",
  11007=>"100100111",
  11008=>"111011111",
  11009=>"001010010",
  11010=>"111111111",
  11011=>"111110110",
  11012=>"111111111",
  11013=>"100110010",
  11014=>"100100101",
  11015=>"111111101",
  11016=>"000011111",
  11017=>"110110110",
  11018=>"000010000",
  11019=>"000001001",
  11020=>"000000000",
  11021=>"000001001",
  11022=>"011011000",
  11023=>"111111111",
  11024=>"001011111",
  11025=>"001000000",
  11026=>"100000000",
  11027=>"100000000",
  11028=>"111111111",
  11029=>"000001001",
  11030=>"010000001",
  11031=>"010111000",
  11032=>"011011011",
  11033=>"000000000",
  11034=>"111111111",
  11035=>"011011000",
  11036=>"000010010",
  11037=>"001011011",
  11038=>"110111111",
  11039=>"111111001",
  11040=>"110111111",
  11041=>"111111111",
  11042=>"101101111",
  11043=>"011011101",
  11044=>"011011011",
  11045=>"110110110",
  11046=>"111010000",
  11047=>"111011111",
  11048=>"011010010",
  11049=>"000000000",
  11050=>"000011000",
  11051=>"101100100",
  11052=>"000000000",
  11053=>"001001111",
  11054=>"000000000",
  11055=>"110110111",
  11056=>"110110100",
  11057=>"000000001",
  11058=>"000000000",
  11059=>"111110111",
  11060=>"000000000",
  11061=>"000000000",
  11062=>"011011000",
  11063=>"111110001",
  11064=>"100000000",
  11065=>"110100100",
  11066=>"111111110",
  11067=>"100100111",
  11068=>"000000000",
  11069=>"110000000",
  11070=>"011011011",
  11071=>"110100110",
  11072=>"111101111",
  11073=>"000000000",
  11074=>"001111111",
  11075=>"111010110",
  11076=>"010000001",
  11077=>"011000110",
  11078=>"010110000",
  11079=>"000000100",
  11080=>"111110010",
  11081=>"000000000",
  11082=>"111111010",
  11083=>"100001000",
  11084=>"000000010",
  11085=>"011000000",
  11086=>"001011111",
  11087=>"101111111",
  11088=>"111110010",
  11089=>"111111100",
  11090=>"001000000",
  11091=>"000000000",
  11092=>"100100110",
  11093=>"111011011",
  11094=>"111111001",
  11095=>"011100000",
  11096=>"111000000",
  11097=>"111111110",
  11098=>"111011011",
  11099=>"000000000",
  11100=>"000000101",
  11101=>"011011011",
  11102=>"011010000",
  11103=>"111110110",
  11104=>"110111100",
  11105=>"111111111",
  11106=>"010001101",
  11107=>"111111111",
  11108=>"111110100",
  11109=>"011000000",
  11110=>"111111111",
  11111=>"000000000",
  11112=>"011011000",
  11113=>"010010010",
  11114=>"111111111",
  11115=>"111001001",
  11116=>"001000000",
  11117=>"010110101",
  11118=>"100000000",
  11119=>"011011000",
  11120=>"111011011",
  11121=>"110111001",
  11122=>"011000000",
  11123=>"001000000",
  11124=>"000100111",
  11125=>"100000000",
  11126=>"000001001",
  11127=>"111111111",
  11128=>"111000000",
  11129=>"111111111",
  11130=>"000110111",
  11131=>"000011000",
  11132=>"111000000",
  11133=>"100110010",
  11134=>"011000001",
  11135=>"000000000",
  11136=>"010110100",
  11137=>"000010010",
  11138=>"000000000",
  11139=>"001000011",
  11140=>"000000000",
  11141=>"111111110",
  11142=>"110000010",
  11143=>"011000000",
  11144=>"111010110",
  11145=>"111111011",
  11146=>"111111111",
  11147=>"100110111",
  11148=>"010000000",
  11149=>"000011011",
  11150=>"000000000",
  11151=>"000000000",
  11152=>"111000001",
  11153=>"000001001",
  11154=>"101000000",
  11155=>"000000000",
  11156=>"000000000",
  11157=>"101000000",
  11158=>"111000000",
  11159=>"110111111",
  11160=>"100000000",
  11161=>"100011011",
  11162=>"011110100",
  11163=>"110010000",
  11164=>"000000010",
  11165=>"111111111",
  11166=>"011011000",
  11167=>"110111111",
  11168=>"111111000",
  11169=>"111000110",
  11170=>"111100100",
  11171=>"111111111",
  11172=>"000001000",
  11173=>"111111111",
  11174=>"000000000",
  11175=>"111011000",
  11176=>"000000001",
  11177=>"111111111",
  11178=>"111110011",
  11179=>"110110110",
  11180=>"111111111",
  11181=>"101101100",
  11182=>"100000000",
  11183=>"000000111",
  11184=>"000000000",
  11185=>"100100000",
  11186=>"000001001",
  11187=>"000000010",
  11188=>"000111111",
  11189=>"000111111",
  11190=>"111111111",
  11191=>"111111111",
  11192=>"111101001",
  11193=>"111111110",
  11194=>"011001011",
  11195=>"011111011",
  11196=>"111111111",
  11197=>"000000110",
  11198=>"100100000",
  11199=>"010010001",
  11200=>"000001001",
  11201=>"111111111",
  11202=>"100000000",
  11203=>"000000000",
  11204=>"000001101",
  11205=>"000001101",
  11206=>"111110100",
  11207=>"110000000",
  11208=>"111101111",
  11209=>"000000111",
  11210=>"110111111",
  11211=>"111011000",
  11212=>"000000000",
  11213=>"000000000",
  11214=>"111011111",
  11215=>"100100110",
  11216=>"001100110",
  11217=>"000111111",
  11218=>"111111111",
  11219=>"111000000",
  11220=>"000110110",
  11221=>"000000011",
  11222=>"111111111",
  11223=>"100010000",
  11224=>"001111111",
  11225=>"000000100",
  11226=>"111111111",
  11227=>"011001011",
  11228=>"011011111",
  11229=>"010100100",
  11230=>"111111011",
  11231=>"011011011",
  11232=>"100100100",
  11233=>"001000000",
  11234=>"111111000",
  11235=>"111011010",
  11236=>"011011111",
  11237=>"101000011",
  11238=>"110011010",
  11239=>"100011011",
  11240=>"111111111",
  11241=>"110100100",
  11242=>"100111111",
  11243=>"000000000",
  11244=>"111111011",
  11245=>"111111111",
  11246=>"111101101",
  11247=>"111111011",
  11248=>"010000011",
  11249=>"111111111",
  11250=>"000001001",
  11251=>"101101111",
  11252=>"000000000",
  11253=>"000000010",
  11254=>"111110110",
  11255=>"001000011",
  11256=>"000000000",
  11257=>"110010110",
  11258=>"111111111",
  11259=>"111111111",
  11260=>"111111111",
  11261=>"111111110",
  11262=>"111111111",
  11263=>"000000000",
  11264=>"000111111",
  11265=>"000000000",
  11266=>"000000000",
  11267=>"000000000",
  11268=>"000011011",
  11269=>"111100000",
  11270=>"000000001",
  11271=>"111111111",
  11272=>"111111011",
  11273=>"000000111",
  11274=>"000000000",
  11275=>"111111111",
  11276=>"100110010",
  11277=>"111011001",
  11278=>"111111110",
  11279=>"111101111",
  11280=>"111011111",
  11281=>"111111101",
  11282=>"000000000",
  11283=>"000000000",
  11284=>"011010000",
  11285=>"000000000",
  11286=>"001000111",
  11287=>"001001000",
  11288=>"111111111",
  11289=>"111111011",
  11290=>"100111111",
  11291=>"100110100",
  11292=>"100110111",
  11293=>"101111011",
  11294=>"011100110",
  11295=>"000001000",
  11296=>"001000000",
  11297=>"000000111",
  11298=>"110100111",
  11299=>"111101111",
  11300=>"111111011",
  11301=>"111000000",
  11302=>"000000001",
  11303=>"000000000",
  11304=>"111111111",
  11305=>"000000000",
  11306=>"110100000",
  11307=>"000010111",
  11308=>"111111111",
  11309=>"111000000",
  11310=>"000000000",
  11311=>"000000000",
  11312=>"001000101",
  11313=>"111001000",
  11314=>"111001001",
  11315=>"010000001",
  11316=>"001010000",
  11317=>"000000001",
  11318=>"111001101",
  11319=>"111100100",
  11320=>"111110000",
  11321=>"110010000",
  11322=>"011001111",
  11323=>"110000000",
  11324=>"000000000",
  11325=>"111111111",
  11326=>"010010000",
  11327=>"111101100",
  11328=>"001000011",
  11329=>"111000000",
  11330=>"000000000",
  11331=>"111111010",
  11332=>"111111111",
  11333=>"000000000",
  11334=>"111000000",
  11335=>"000001001",
  11336=>"011111001",
  11337=>"000000111",
  11338=>"111111111",
  11339=>"000000000",
  11340=>"111111001",
  11341=>"000011001",
  11342=>"111110100",
  11343=>"110111111",
  11344=>"110000000",
  11345=>"110000000",
  11346=>"000111111",
  11347=>"100011001",
  11348=>"110111111",
  11349=>"000110111",
  11350=>"111111111",
  11351=>"000000000",
  11352=>"000000000",
  11353=>"100000000",
  11354=>"000001000",
  11355=>"111001001",
  11356=>"000000000",
  11357=>"111111111",
  11358=>"011011111",
  11359=>"011011011",
  11360=>"000111111",
  11361=>"010110100",
  11362=>"101101111",
  11363=>"000000101",
  11364=>"111111111",
  11365=>"100100111",
  11366=>"011001101",
  11367=>"000000000",
  11368=>"011001100",
  11369=>"111111011",
  11370=>"111100000",
  11371=>"001000000",
  11372=>"001011111",
  11373=>"000011100",
  11374=>"001000000",
  11375=>"111000000",
  11376=>"111111111",
  11377=>"001001110",
  11378=>"001011111",
  11379=>"001001000",
  11380=>"111010000",
  11381=>"000000000",
  11382=>"001001000",
  11383=>"010111111",
  11384=>"000000000",
  11385=>"000000011",
  11386=>"000001001",
  11387=>"000000000",
  11388=>"000111111",
  11389=>"000011001",
  11390=>"010111011",
  11391=>"000000000",
  11392=>"111111110",
  11393=>"000001000",
  11394=>"011001111",
  11395=>"001000110",
  11396=>"000000101",
  11397=>"000000000",
  11398=>"111111101",
  11399=>"000000000",
  11400=>"000000000",
  11401=>"001000000",
  11402=>"011000001",
  11403=>"000000000",
  11404=>"111111011",
  11405=>"111001111",
  11406=>"011011111",
  11407=>"011011011",
  11408=>"111110100",
  11409=>"000110000",
  11410=>"100111111",
  11411=>"000110011",
  11412=>"111111110",
  11413=>"111111111",
  11414=>"111111110",
  11415=>"000000000",
  11416=>"011000000",
  11417=>"110110111",
  11418=>"000010010",
  11419=>"111111111",
  11420=>"000000100",
  11421=>"111111111",
  11422=>"100000000",
  11423=>"111111010",
  11424=>"000000110",
  11425=>"110100100",
  11426=>"111101001",
  11427=>"111111111",
  11428=>"111111011",
  11429=>"010000011",
  11430=>"111111111",
  11431=>"001101111",
  11432=>"111000000",
  11433=>"111111101",
  11434=>"111111111",
  11435=>"111111111",
  11436=>"111111111",
  11437=>"111111111",
  11438=>"111110111",
  11439=>"001001001",
  11440=>"111010000",
  11441=>"011001100",
  11442=>"000111000",
  11443=>"111111111",
  11444=>"000000000",
  11445=>"100100100",
  11446=>"111000111",
  11447=>"111100100",
  11448=>"000000100",
  11449=>"111100000",
  11450=>"100001111",
  11451=>"111111111",
  11452=>"000000000",
  11453=>"000000000",
  11454=>"000000000",
  11455=>"000001001",
  11456=>"111111111",
  11457=>"110111001",
  11458=>"111111111",
  11459=>"000000111",
  11460=>"111111111",
  11461=>"000000000",
  11462=>"101000000",
  11463=>"000011011",
  11464=>"001000011",
  11465=>"111111111",
  11466=>"111111101",
  11467=>"000000000",
  11468=>"111111111",
  11469=>"111111110",
  11470=>"111111111",
  11471=>"100000000",
  11472=>"000000000",
  11473=>"011111111",
  11474=>"111111111",
  11475=>"111111000",
  11476=>"111111111",
  11477=>"110110000",
  11478=>"100010000",
  11479=>"111111111",
  11480=>"000000000",
  11481=>"111111111",
  11482=>"000000000",
  11483=>"000100111",
  11484=>"000000001",
  11485=>"000000111",
  11486=>"000000000",
  11487=>"111001000",
  11488=>"000000000",
  11489=>"111111111",
  11490=>"111111111",
  11491=>"100000011",
  11492=>"111111111",
  11493=>"110100000",
  11494=>"111111111",
  11495=>"000000001",
  11496=>"100001001",
  11497=>"111111111",
  11498=>"111001000",
  11499=>"111000000",
  11500=>"111111111",
  11501=>"000000000",
  11502=>"011101111",
  11503=>"110100111",
  11504=>"000000111",
  11505=>"000000000",
  11506=>"000010111",
  11507=>"110110111",
  11508=>"101101101",
  11509=>"111110000",
  11510=>"111111111",
  11511=>"001000000",
  11512=>"111111111",
  11513=>"111111111",
  11514=>"100000111",
  11515=>"111111000",
  11516=>"111111110",
  11517=>"111111111",
  11518=>"111111111",
  11519=>"011000000",
  11520=>"010000000",
  11521=>"111111011",
  11522=>"000000011",
  11523=>"000000000",
  11524=>"000000000",
  11525=>"111100100",
  11526=>"000000001",
  11527=>"111111000",
  11528=>"111111111",
  11529=>"111111000",
  11530=>"111111111",
  11531=>"111101111",
  11532=>"000000100",
  11533=>"111111111",
  11534=>"110100111",
  11535=>"001000000",
  11536=>"111000000",
  11537=>"111001000",
  11538=>"100000000",
  11539=>"000000000",
  11540=>"111011000",
  11541=>"001001111",
  11542=>"110111111",
  11543=>"000000000",
  11544=>"111111111",
  11545=>"000011000",
  11546=>"000000001",
  11547=>"000000000",
  11548=>"000000000",
  11549=>"000011001",
  11550=>"111111111",
  11551=>"111111000",
  11552=>"111111111",
  11553=>"111111111",
  11554=>"000000010",
  11555=>"110111111",
  11556=>"001001111",
  11557=>"000000100",
  11558=>"000111111",
  11559=>"111001000",
  11560=>"000000000",
  11561=>"110000101",
  11562=>"000000000",
  11563=>"010110010",
  11564=>"000000000",
  11565=>"100100100",
  11566=>"111111111",
  11567=>"111001000",
  11568=>"001001011",
  11569=>"101101111",
  11570=>"100110110",
  11571=>"110111010",
  11572=>"111110110",
  11573=>"000000011",
  11574=>"001001011",
  11575=>"111111100",
  11576=>"000000011",
  11577=>"111101111",
  11578=>"111011001",
  11579=>"100110110",
  11580=>"110000000",
  11581=>"000001001",
  11582=>"111111111",
  11583=>"110111111",
  11584=>"000000000",
  11585=>"000011000",
  11586=>"110010001",
  11587=>"000000000",
  11588=>"111001111",
  11589=>"101100000",
  11590=>"000000000",
  11591=>"000000000",
  11592=>"111111111",
  11593=>"000111101",
  11594=>"110000100",
  11595=>"001001101",
  11596=>"000000000",
  11597=>"111111011",
  11598=>"111000111",
  11599=>"111100110",
  11600=>"000000001",
  11601=>"000000000",
  11602=>"000000000",
  11603=>"111111110",
  11604=>"001001000",
  11605=>"111011011",
  11606=>"111111011",
  11607=>"001001000",
  11608=>"000100010",
  11609=>"000111111",
  11610=>"000001000",
  11611=>"000000000",
  11612=>"000000101",
  11613=>"111111111",
  11614=>"000001101",
  11615=>"011111111",
  11616=>"000000000",
  11617=>"111111111",
  11618=>"000001011",
  11619=>"111011011",
  11620=>"111001011",
  11621=>"111111011",
  11622=>"000010011",
  11623=>"000000111",
  11624=>"000000110",
  11625=>"000000000",
  11626=>"111111011",
  11627=>"111111000",
  11628=>"101101001",
  11629=>"111011011",
  11630=>"111111111",
  11631=>"011000000",
  11632=>"001000001",
  11633=>"111111110",
  11634=>"000110111",
  11635=>"000000001",
  11636=>"111111111",
  11637=>"100000000",
  11638=>"110111101",
  11639=>"001011000",
  11640=>"111000000",
  11641=>"111111010",
  11642=>"100000000",
  11643=>"111001001",
  11644=>"000000101",
  11645=>"000011111",
  11646=>"100000111",
  11647=>"111111011",
  11648=>"101110111",
  11649=>"000000000",
  11650=>"000000000",
  11651=>"101000100",
  11652=>"111111111",
  11653=>"000000000",
  11654=>"100000000",
  11655=>"110111111",
  11656=>"000000101",
  11657=>"001001011",
  11658=>"000001001",
  11659=>"000001000",
  11660=>"011001101",
  11661=>"011000000",
  11662=>"111111111",
  11663=>"000000000",
  11664=>"111111111",
  11665=>"000000100",
  11666=>"111111111",
  11667=>"000000000",
  11668=>"001001000",
  11669=>"011100000",
  11670=>"111111111",
  11671=>"100111111",
  11672=>"110111111",
  11673=>"101001011",
  11674=>"000000011",
  11675=>"110011001",
  11676=>"000000001",
  11677=>"000000000",
  11678=>"000000000",
  11679=>"000010010",
  11680=>"111111111",
  11681=>"111111111",
  11682=>"110000000",
  11683=>"111000000",
  11684=>"111011111",
  11685=>"011111111",
  11686=>"000111111",
  11687=>"110110110",
  11688=>"110000000",
  11689=>"000000000",
  11690=>"100100000",
  11691=>"000000100",
  11692=>"000000000",
  11693=>"101100111",
  11694=>"111111111",
  11695=>"001111011",
  11696=>"000111111",
  11697=>"000010000",
  11698=>"011111101",
  11699=>"101001000",
  11700=>"100100100",
  11701=>"111111111",
  11702=>"010000010",
  11703=>"001000000",
  11704=>"000011111",
  11705=>"110110111",
  11706=>"001001001",
  11707=>"100000111",
  11708=>"111111111",
  11709=>"111111111",
  11710=>"000010001",
  11711=>"000000001",
  11712=>"000000000",
  11713=>"111111111",
  11714=>"111111111",
  11715=>"111011011",
  11716=>"111000111",
  11717=>"111001111",
  11718=>"000000101",
  11719=>"000000011",
  11720=>"000000000",
  11721=>"000000001",
  11722=>"111111001",
  11723=>"111111111",
  11724=>"111100111",
  11725=>"010110010",
  11726=>"000000000",
  11727=>"000000000",
  11728=>"111000100",
  11729=>"011000011",
  11730=>"011000000",
  11731=>"000010000",
  11732=>"111110111",
  11733=>"111111111",
  11734=>"011011011",
  11735=>"000000000",
  11736=>"000000000",
  11737=>"111110111",
  11738=>"111111111",
  11739=>"111111111",
  11740=>"000011011",
  11741=>"000000101",
  11742=>"111111111",
  11743=>"000000000",
  11744=>"001000100",
  11745=>"111111000",
  11746=>"111110111",
  11747=>"101000110",
  11748=>"000000000",
  11749=>"010000010",
  11750=>"001001000",
  11751=>"000000000",
  11752=>"000000001",
  11753=>"000101111",
  11754=>"000000000",
  11755=>"111111111",
  11756=>"111001000",
  11757=>"011111111",
  11758=>"000000000",
  11759=>"000000000",
  11760=>"100000000",
  11761=>"111111111",
  11762=>"111111011",
  11763=>"000000000",
  11764=>"110000000",
  11765=>"000000000",
  11766=>"111111111",
  11767=>"001000001",
  11768=>"000000111",
  11769=>"101001000",
  11770=>"110111111",
  11771=>"111111111",
  11772=>"001000100",
  11773=>"000100110",
  11774=>"100000111",
  11775=>"100000000",
  11776=>"000000001",
  11777=>"000000111",
  11778=>"000111111",
  11779=>"111011001",
  11780=>"111111111",
  11781=>"000000000",
  11782=>"011111111",
  11783=>"111000000",
  11784=>"000111111",
  11785=>"111111111",
  11786=>"111011011",
  11787=>"011011001",
  11788=>"101011010",
  11789=>"100000000",
  11790=>"110000000",
  11791=>"100001011",
  11792=>"110111111",
  11793=>"010100000",
  11794=>"000000000",
  11795=>"000000000",
  11796=>"000000101",
  11797=>"111000000",
  11798=>"000000000",
  11799=>"111010000",
  11800=>"000000110",
  11801=>"000111111",
  11802=>"111101101",
  11803=>"011011011",
  11804=>"111101111",
  11805=>"111111111",
  11806=>"000001001",
  11807=>"000001000",
  11808=>"001000001",
  11809=>"000110111",
  11810=>"100111111",
  11811=>"111111111",
  11812=>"001001011",
  11813=>"111111111",
  11814=>"110000111",
  11815=>"000000000",
  11816=>"101111001",
  11817=>"011011000",
  11818=>"100100100",
  11819=>"000111100",
  11820=>"000111101",
  11821=>"000000000",
  11822=>"011001000",
  11823=>"000000000",
  11824=>"000000001",
  11825=>"000111001",
  11826=>"000111111",
  11827=>"000000110",
  11828=>"111001111",
  11829=>"110110110",
  11830=>"000000000",
  11831=>"000000001",
  11832=>"111111111",
  11833=>"000001001",
  11834=>"000000000",
  11835=>"111000000",
  11836=>"000000001",
  11837=>"110111101",
  11838=>"000000000",
  11839=>"001000101",
  11840=>"100001011",
  11841=>"011000000",
  11842=>"000000000",
  11843=>"000000000",
  11844=>"100111111",
  11845=>"000000000",
  11846=>"000000100",
  11847=>"111111111",
  11848=>"110111111",
  11849=>"001000100",
  11850=>"111111111",
  11851=>"100000110",
  11852=>"001000000",
  11853=>"111110000",
  11854=>"000000000",
  11855=>"111111111",
  11856=>"001000000",
  11857=>"111111111",
  11858=>"000100100",
  11859=>"000111111",
  11860=>"000000000",
  11861=>"100111101",
  11862=>"110111000",
  11863=>"101111111",
  11864=>"001000000",
  11865=>"111111111",
  11866=>"000000000",
  11867=>"100100000",
  11868=>"000111111",
  11869=>"110110000",
  11870=>"000111100",
  11871=>"000011110",
  11872=>"111110111",
  11873=>"000000000",
  11874=>"000000010",
  11875=>"100101111",
  11876=>"011111111",
  11877=>"000000000",
  11878=>"111111111",
  11879=>"000000000",
  11880=>"100111111",
  11881=>"110110111",
  11882=>"000111111",
  11883=>"111111110",
  11884=>"110110011",
  11885=>"111111110",
  11886=>"111111111",
  11887=>"110110110",
  11888=>"000000001",
  11889=>"111011000",
  11890=>"001000001",
  11891=>"100011011",
  11892=>"011011111",
  11893=>"000000000",
  11894=>"111111111",
  11895=>"010111011",
  11896=>"000000000",
  11897=>"101101000",
  11898=>"000000000",
  11899=>"000000000",
  11900=>"000000000",
  11901=>"000000000",
  11902=>"000000000",
  11903=>"000000011",
  11904=>"000000000",
  11905=>"000100000",
  11906=>"100000101",
  11907=>"000000000",
  11908=>"111111110",
  11909=>"111000000",
  11910=>"001011111",
  11911=>"101000000",
  11912=>"000000000",
  11913=>"000000000",
  11914=>"100100111",
  11915=>"000000000",
  11916=>"111111111",
  11917=>"000000000",
  11918=>"000111101",
  11919=>"111101110",
  11920=>"111111111",
  11921=>"101001000",
  11922=>"111101111",
  11923=>"110111110",
  11924=>"000000110",
  11925=>"000000010",
  11926=>"101111111",
  11927=>"111111000",
  11928=>"111001001",
  11929=>"110110101",
  11930=>"011011000",
  11931=>"000100100",
  11932=>"000110111",
  11933=>"000000000",
  11934=>"111000000",
  11935=>"111111111",
  11936=>"111111111",
  11937=>"111111111",
  11938=>"111111111",
  11939=>"111011000",
  11940=>"111001000",
  11941=>"000000111",
  11942=>"101000001",
  11943=>"000000000",
  11944=>"000000100",
  11945=>"000000000",
  11946=>"000000000",
  11947=>"111111011",
  11948=>"001001110",
  11949=>"001011011",
  11950=>"111110100",
  11951=>"111111110",
  11952=>"000000000",
  11953=>"000000000",
  11954=>"110110110",
  11955=>"000000111",
  11956=>"000000000",
  11957=>"111111111",
  11958=>"000000010",
  11959=>"111011000",
  11960=>"000100010",
  11961=>"111101100",
  11962=>"111001111",
  11963=>"100000000",
  11964=>"110100100",
  11965=>"000011000",
  11966=>"000000000",
  11967=>"111000000",
  11968=>"100000000",
  11969=>"000100110",
  11970=>"111000000",
  11971=>"000000000",
  11972=>"111000000",
  11973=>"111101111",
  11974=>"000001001",
  11975=>"000000000",
  11976=>"000111111",
  11977=>"011111000",
  11978=>"000000010",
  11979=>"111111111",
  11980=>"111111100",
  11981=>"100000000",
  11982=>"110100100",
  11983=>"000001011",
  11984=>"111000000",
  11985=>"000000000",
  11986=>"100000000",
  11987=>"111111111",
  11988=>"110011001",
  11989=>"111110110",
  11990=>"111111111",
  11991=>"000110110",
  11992=>"000100110",
  11993=>"000001101",
  11994=>"111101111",
  11995=>"000000000",
  11996=>"110111101",
  11997=>"000000000",
  11998=>"110000111",
  11999=>"011111111",
  12000=>"010111101",
  12001=>"011111100",
  12002=>"111011111",
  12003=>"110111101",
  12004=>"111111011",
  12005=>"001001011",
  12006=>"001100100",
  12007=>"111111000",
  12008=>"000000000",
  12009=>"000000011",
  12010=>"000010111",
  12011=>"100100000",
  12012=>"000001111",
  12013=>"111101100",
  12014=>"111000110",
  12015=>"111000101",
  12016=>"110000010",
  12017=>"111111111",
  12018=>"111100000",
  12019=>"101001000",
  12020=>"000001111",
  12021=>"001000000",
  12022=>"111111100",
  12023=>"111010000",
  12024=>"000000000",
  12025=>"000000111",
  12026=>"000000000",
  12027=>"101000000",
  12028=>"000011000",
  12029=>"001011010",
  12030=>"111111000",
  12031=>"000111111",
  12032=>"111111111",
  12033=>"011011011",
  12034=>"111111111",
  12035=>"011111100",
  12036=>"110110110",
  12037=>"110011111",
  12038=>"000000000",
  12039=>"000011111",
  12040=>"111111100",
  12041=>"000100110",
  12042=>"111111111",
  12043=>"111111110",
  12044=>"110110110",
  12045=>"000001001",
  12046=>"111111111",
  12047=>"111100000",
  12048=>"001001111",
  12049=>"101001111",
  12050=>"111111001",
  12051=>"111111111",
  12052=>"000001011",
  12053=>"000000111",
  12054=>"001001001",
  12055=>"111111100",
  12056=>"010000011",
  12057=>"111111111",
  12058=>"000000000",
  12059=>"000000110",
  12060=>"111011011",
  12061=>"111111110",
  12062=>"111111111",
  12063=>"110000101",
  12064=>"110111000",
  12065=>"011110111",
  12066=>"000000000",
  12067=>"000011001",
  12068=>"001001001",
  12069=>"101111111",
  12070=>"111111111",
  12071=>"111111101",
  12072=>"000000000",
  12073=>"000000000",
  12074=>"101001111",
  12075=>"100100111",
  12076=>"100110100",
  12077=>"000000000",
  12078=>"000101111",
  12079=>"110111111",
  12080=>"110000000",
  12081=>"000000000",
  12082=>"110111111",
  12083=>"001000011",
  12084=>"111110110",
  12085=>"000000000",
  12086=>"000110000",
  12087=>"000000111",
  12088=>"000000000",
  12089=>"000000000",
  12090=>"011011111",
  12091=>"000000000",
  12092=>"111111110",
  12093=>"000001111",
  12094=>"101101101",
  12095=>"000001111",
  12096=>"000001000",
  12097=>"110000000",
  12098=>"000000000",
  12099=>"111110000",
  12100=>"111111110",
  12101=>"000000000",
  12102=>"000000111",
  12103=>"111111011",
  12104=>"000000000",
  12105=>"111000001",
  12106=>"000000010",
  12107=>"000000000",
  12108=>"001000000",
  12109=>"101111111",
  12110=>"110010111",
  12111=>"111111111",
  12112=>"000000001",
  12113=>"011010110",
  12114=>"000010010",
  12115=>"111111111",
  12116=>"000100100",
  12117=>"011011001",
  12118=>"111110011",
  12119=>"000000000",
  12120=>"000100110",
  12121=>"001000111",
  12122=>"000111111",
  12123=>"111111111",
  12124=>"000010000",
  12125=>"111111111",
  12126=>"000011111",
  12127=>"011111111",
  12128=>"111111111",
  12129=>"000001000",
  12130=>"000000000",
  12131=>"101000101",
  12132=>"000010010",
  12133=>"000000000",
  12134=>"111111111",
  12135=>"011001111",
  12136=>"000000000",
  12137=>"000111111",
  12138=>"110110110",
  12139=>"110011001",
  12140=>"000000000",
  12141=>"111000001",
  12142=>"001000100",
  12143=>"100101111",
  12144=>"001001010",
  12145=>"000101001",
  12146=>"111111110",
  12147=>"111111111",
  12148=>"011111111",
  12149=>"000000000",
  12150=>"000000000",
  12151=>"000011001",
  12152=>"111000000",
  12153=>"110111000",
  12154=>"000000000",
  12155=>"111111111",
  12156=>"111111111",
  12157=>"111111111",
  12158=>"110110110",
  12159=>"000000000",
  12160=>"110010000",
  12161=>"111111110",
  12162=>"010000000",
  12163=>"000000111",
  12164=>"101101111",
  12165=>"100111001",
  12166=>"101101111",
  12167=>"010011000",
  12168=>"001000101",
  12169=>"111010010",
  12170=>"111001000",
  12171=>"001000000",
  12172=>"101100111",
  12173=>"000000000",
  12174=>"110001100",
  12175=>"000000000",
  12176=>"000000000",
  12177=>"000100100",
  12178=>"111111111",
  12179=>"110000000",
  12180=>"011111111",
  12181=>"000000001",
  12182=>"000011010",
  12183=>"011001001",
  12184=>"111000111",
  12185=>"111001000",
  12186=>"110110100",
  12187=>"000000000",
  12188=>"000000000",
  12189=>"000100111",
  12190=>"111111111",
  12191=>"000000000",
  12192=>"000000000",
  12193=>"000000000",
  12194=>"000111001",
  12195=>"111111111",
  12196=>"100111011",
  12197=>"000000000",
  12198=>"100111111",
  12199=>"000010000",
  12200=>"100001011",
  12201=>"011111111",
  12202=>"101100000",
  12203=>"111111111",
  12204=>"000000000",
  12205=>"011000000",
  12206=>"000111000",
  12207=>"000000000",
  12208=>"111111111",
  12209=>"111111111",
  12210=>"111111111",
  12211=>"000100000",
  12212=>"111110111",
  12213=>"111111111",
  12214=>"001111110",
  12215=>"000010000",
  12216=>"100111111",
  12217=>"000100001",
  12218=>"110110000",
  12219=>"110000000",
  12220=>"111011000",
  12221=>"110111110",
  12222=>"111111111",
  12223=>"111011010",
  12224=>"011111111",
  12225=>"000001011",
  12226=>"000000000",
  12227=>"000000000",
  12228=>"000011111",
  12229=>"000101111",
  12230=>"000000000",
  12231=>"000111001",
  12232=>"011001100",
  12233=>"000000000",
  12234=>"110111111",
  12235=>"100111111",
  12236=>"000000111",
  12237=>"000100111",
  12238=>"110111111",
  12239=>"000110111",
  12240=>"000111111",
  12241=>"110001001",
  12242=>"110000000",
  12243=>"111111111",
  12244=>"000110100",
  12245=>"100101000",
  12246=>"111111001",
  12247=>"111100000",
  12248=>"001001000",
  12249=>"000011001",
  12250=>"000000000",
  12251=>"000000000",
  12252=>"111111111",
  12253=>"110111111",
  12254=>"000000100",
  12255=>"000000011",
  12256=>"111111111",
  12257=>"000000010",
  12258=>"000000100",
  12259=>"110111111",
  12260=>"111111011",
  12261=>"110110100",
  12262=>"001000100",
  12263=>"000000100",
  12264=>"000000010",
  12265=>"000001011",
  12266=>"001000000",
  12267=>"001001001",
  12268=>"101000001",
  12269=>"110010010",
  12270=>"111111111",
  12271=>"000100111",
  12272=>"111111111",
  12273=>"000000000",
  12274=>"010011011",
  12275=>"111001111",
  12276=>"100001111",
  12277=>"011000000",
  12278=>"000110111",
  12279=>"100101111",
  12280=>"011010000",
  12281=>"100000000",
  12282=>"000111011",
  12283=>"111111111",
  12284=>"000000000",
  12285=>"000000000",
  12286=>"111110000",
  12287=>"110110110",
  12288=>"010010110",
  12289=>"011011011",
  12290=>"011011010",
  12291=>"111011001",
  12292=>"111000100",
  12293=>"111101001",
  12294=>"111111111",
  12295=>"111111101",
  12296=>"011111111",
  12297=>"111111111",
  12298=>"111001111",
  12299=>"001001010",
  12300=>"000000000",
  12301=>"111101101",
  12302=>"111101101",
  12303=>"111101101",
  12304=>"010000000",
  12305=>"111001001",
  12306=>"010010011",
  12307=>"000111111",
  12308=>"010010110",
  12309=>"010000000",
  12310=>"110010111",
  12311=>"011001000",
  12312=>"001001001",
  12313=>"000001000",
  12314=>"101000000",
  12315=>"011111111",
  12316=>"111111000",
  12317=>"110000110",
  12318=>"111100100",
  12319=>"101000000",
  12320=>"000010001",
  12321=>"000000111",
  12322=>"100100101",
  12323=>"110010010",
  12324=>"110111111",
  12325=>"010010111",
  12326=>"000000000",
  12327=>"001001111",
  12328=>"110110111",
  12329=>"010010010",
  12330=>"011111111",
  12331=>"111111100",
  12332=>"000111111",
  12333=>"001101000",
  12334=>"111011011",
  12335=>"010011111",
  12336=>"100000000",
  12337=>"011010110",
  12338=>"101001000",
  12339=>"101000000",
  12340=>"000000000",
  12341=>"101001001",
  12342=>"111100100",
  12343=>"000010010",
  12344=>"011011111",
  12345=>"101101101",
  12346=>"001001001",
  12347=>"000100100",
  12348=>"101000111",
  12349=>"101001101",
  12350=>"001001011",
  12351=>"001111101",
  12352=>"000001100",
  12353=>"000010010",
  12354=>"011001111",
  12355=>"011001010",
  12356=>"001001010",
  12357=>"011111110",
  12358=>"011011111",
  12359=>"111111111",
  12360=>"001001001",
  12361=>"000000000",
  12362=>"000000111",
  12363=>"111010011",
  12364=>"100100111",
  12365=>"110110010",
  12366=>"000100101",
  12367=>"001111111",
  12368=>"101000000",
  12369=>"101010110",
  12370=>"000000101",
  12371=>"000001001",
  12372=>"001001001",
  12373=>"001111111",
  12374=>"101011001",
  12375=>"100000000",
  12376=>"111000100",
  12377=>"000000100",
  12378=>"110111111",
  12379=>"111001000",
  12380=>"011000100",
  12381=>"100101111",
  12382=>"011111110",
  12383=>"000001001",
  12384=>"000000000",
  12385=>"000000101",
  12386=>"111001101",
  12387=>"000000000",
  12388=>"000000001",
  12389=>"100001101",
  12390=>"111111111",
  12391=>"000101111",
  12392=>"111000000",
  12393=>"000100100",
  12394=>"000011010",
  12395=>"110010000",
  12396=>"000000000",
  12397=>"100100111",
  12398=>"111111111",
  12399=>"011011011",
  12400=>"000001101",
  12401=>"110010010",
  12402=>"101101100",
  12403=>"111000011",
  12404=>"111101100",
  12405=>"111110110",
  12406=>"010010010",
  12407=>"001011010",
  12408=>"000000000",
  12409=>"101000100",
  12410=>"110110110",
  12411=>"000000001",
  12412=>"001001001",
  12413=>"000000000",
  12414=>"111010000",
  12415=>"011011011",
  12416=>"000000001",
  12417=>"001000000",
  12418=>"010111011",
  12419=>"000001000",
  12420=>"100100111",
  12421=>"000000000",
  12422=>"100000000",
  12423=>"001011111",
  12424=>"111111001",
  12425=>"000001001",
  12426=>"111111111",
  12427=>"011001001",
  12428=>"011011111",
  12429=>"000000000",
  12430=>"111001001",
  12431=>"111111111",
  12432=>"001101101",
  12433=>"001001101",
  12434=>"101101000",
  12435=>"111100110",
  12436=>"000001000",
  12437=>"101001101",
  12438=>"011011111",
  12439=>"000000011",
  12440=>"110010010",
  12441=>"010110110",
  12442=>"111010010",
  12443=>"001011111",
  12444=>"110000111",
  12445=>"000000010",
  12446=>"100000000",
  12447=>"111001101",
  12448=>"111110000",
  12449=>"000000111",
  12450=>"011011011",
  12451=>"100100100",
  12452=>"110010110",
  12453=>"011111111",
  12454=>"011111111",
  12455=>"100100100",
  12456=>"101111010",
  12457=>"111111100",
  12458=>"011011001",
  12459=>"000000111",
  12460=>"100000000",
  12461=>"101101101",
  12462=>"000000011",
  12463=>"001101101",
  12464=>"000000110",
  12465=>"001101101",
  12466=>"000101101",
  12467=>"000000001",
  12468=>"011010010",
  12469=>"110010011",
  12470=>"101001101",
  12471=>"111101100",
  12472=>"100111110",
  12473=>"000011001",
  12474=>"000000110",
  12475=>"001001111",
  12476=>"000000111",
  12477=>"001000000",
  12478=>"000000000",
  12479=>"000011011",
  12480=>"100100000",
  12481=>"001000010",
  12482=>"111011011",
  12483=>"101101111",
  12484=>"111111000",
  12485=>"010010111",
  12486=>"000000000",
  12487=>"001000100",
  12488=>"001000001",
  12489=>"101100000",
  12490=>"100101111",
  12491=>"111001001",
  12492=>"101101100",
  12493=>"011011011",
  12494=>"010000000",
  12495=>"111001000",
  12496=>"100000111",
  12497=>"001001101",
  12498=>"001001111",
  12499=>"101000000",
  12500=>"101101000",
  12501=>"101110111",
  12502=>"010010010",
  12503=>"111110110",
  12504=>"111101101",
  12505=>"111011001",
  12506=>"010010011",
  12507=>"001101111",
  12508=>"101000001",
  12509=>"001001001",
  12510=>"101111100",
  12511=>"111000100",
  12512=>"000010010",
  12513=>"010011011",
  12514=>"010100000",
  12515=>"111111110",
  12516=>"111000000",
  12517=>"100110010",
  12518=>"011001000",
  12519=>"100000000",
  12520=>"111111110",
  12521=>"111110110",
  12522=>"010000110",
  12523=>"111000000",
  12524=>"101100100",
  12525=>"000111011",
  12526=>"111001111",
  12527=>"011010000",
  12528=>"110111000",
  12529=>"010000101",
  12530=>"010110110",
  12531=>"000011011",
  12532=>"111111111",
  12533=>"000100100",
  12534=>"111111001",
  12535=>"011010111",
  12536=>"100111111",
  12537=>"100100101",
  12538=>"000010010",
  12539=>"000000010",
  12540=>"111111000",
  12541=>"011100000",
  12542=>"101001000",
  12543=>"111110111",
  12544=>"101000010",
  12545=>"101101101",
  12546=>"000101000",
  12547=>"101101100",
  12548=>"111000100",
  12549=>"000000111",
  12550=>"011111000",
  12551=>"111110110",
  12552=>"001001111",
  12553=>"000000000",
  12554=>"111011110",
  12555=>"011001111",
  12556=>"000000000",
  12557=>"000000000",
  12558=>"000010111",
  12559=>"111110110",
  12560=>"111101101",
  12561=>"000000001",
  12562=>"010111111",
  12563=>"001000000",
  12564=>"000100110",
  12565=>"100000001",
  12566=>"100100100",
  12567=>"001001111",
  12568=>"001001001",
  12569=>"010011011",
  12570=>"111011000",
  12571=>"111011010",
  12572=>"100101111",
  12573=>"010011011",
  12574=>"011111111",
  12575=>"111001101",
  12576=>"110011001",
  12577=>"001000000",
  12578=>"010010000",
  12579=>"000111111",
  12580=>"000111111",
  12581=>"101101100",
  12582=>"100100100",
  12583=>"010111111",
  12584=>"101001101",
  12585=>"111111101",
  12586=>"000011011",
  12587=>"000000010",
  12588=>"111111000",
  12589=>"000100000",
  12590=>"011001111",
  12591=>"100000100",
  12592=>"011011000",
  12593=>"111110110",
  12594=>"100001111",
  12595=>"010011011",
  12596=>"000000000",
  12597=>"101111111",
  12598=>"100100110",
  12599=>"110110110",
  12600=>"000010000",
  12601=>"000000011",
  12602=>"001001111",
  12603=>"110010000",
  12604=>"110110111",
  12605=>"001001100",
  12606=>"101101101",
  12607=>"111000001",
  12608=>"000000000",
  12609=>"000001101",
  12610=>"000000000",
  12611=>"000000000",
  12612=>"001101100",
  12613=>"011000000",
  12614=>"011111000",
  12615=>"110000111",
  12616=>"111100000",
  12617=>"000000111",
  12618=>"011010111",
  12619=>"001001001",
  12620=>"110011110",
  12621=>"000011011",
  12622=>"011010011",
  12623=>"001011011",
  12624=>"001001001",
  12625=>"111011000",
  12626=>"101111111",
  12627=>"000000101",
  12628=>"100100100",
  12629=>"001011001",
  12630=>"000000010",
  12631=>"111111100",
  12632=>"111111111",
  12633=>"000000101",
  12634=>"100000101",
  12635=>"011011011",
  12636=>"010010010",
  12637=>"000110111",
  12638=>"000000111",
  12639=>"101100110",
  12640=>"010010010",
  12641=>"001001111",
  12642=>"000011001",
  12643=>"100000000",
  12644=>"101101101",
  12645=>"001011111",
  12646=>"011111011",
  12647=>"001001110",
  12648=>"101100100",
  12649=>"111111101",
  12650=>"111001001",
  12651=>"011011001",
  12652=>"001011001",
  12653=>"111000000",
  12654=>"111101101",
  12655=>"111101001",
  12656=>"111001111",
  12657=>"111100111",
  12658=>"011011111",
  12659=>"111111100",
  12660=>"011010010",
  12661=>"111001111",
  12662=>"101000000",
  12663=>"101101001",
  12664=>"101101111",
  12665=>"011111001",
  12666=>"111101111",
  12667=>"101101101",
  12668=>"011110111",
  12669=>"111111110",
  12670=>"110010010",
  12671=>"111111111",
  12672=>"110110110",
  12673=>"000000000",
  12674=>"110010001",
  12675=>"010010011",
  12676=>"001000000",
  12677=>"000000000",
  12678=>"110110111",
  12679=>"010010010",
  12680=>"111110111",
  12681=>"011000001",
  12682=>"011011011",
  12683=>"010010010",
  12684=>"111111111",
  12685=>"100100101",
  12686=>"101101101",
  12687=>"101100101",
  12688=>"111101000",
  12689=>"000101101",
  12690=>"101111110",
  12691=>"111111010",
  12692=>"000111111",
  12693=>"000000000",
  12694=>"101101100",
  12695=>"010000000",
  12696=>"100000111",
  12697=>"111101100",
  12698=>"011111110",
  12699=>"101001001",
  12700=>"001001000",
  12701=>"110110100",
  12702=>"000010000",
  12703=>"000000111",
  12704=>"011000000",
  12705=>"101101100",
  12706=>"001000110",
  12707=>"011111010",
  12708=>"000000000",
  12709=>"000101000",
  12710=>"010000111",
  12711=>"000000101",
  12712=>"010000000",
  12713=>"011111111",
  12714=>"110111100",
  12715=>"000011101",
  12716=>"111101101",
  12717=>"111001011",
  12718=>"111101101",
  12719=>"001100111",
  12720=>"000000000",
  12721=>"111111101",
  12722=>"111111111",
  12723=>"011111111",
  12724=>"100111111",
  12725=>"100111111",
  12726=>"000000101",
  12727=>"111111000",
  12728=>"000110010",
  12729=>"101101111",
  12730=>"101101101",
  12731=>"000000000",
  12732=>"000100010",
  12733=>"001010010",
  12734=>"000000000",
  12735=>"100100101",
  12736=>"111111101",
  12737=>"101101001",
  12738=>"001101100",
  12739=>"111111111",
  12740=>"100010010",
  12741=>"001000001",
  12742=>"100101100",
  12743=>"010010010",
  12744=>"111011010",
  12745=>"100100000",
  12746=>"011111010",
  12747=>"000000111",
  12748=>"000000000",
  12749=>"111111000",
  12750=>"101101101",
  12751=>"111111101",
  12752=>"101001101",
  12753=>"000001000",
  12754=>"111101111",
  12755=>"101101101",
  12756=>"000000000",
  12757=>"111010000",
  12758=>"000001000",
  12759=>"001100100",
  12760=>"000101101",
  12761=>"011001101",
  12762=>"001001111",
  12763=>"011000101",
  12764=>"011010111",
  12765=>"111110100",
  12766=>"111101111",
  12767=>"100100100",
  12768=>"000000000",
  12769=>"101001101",
  12770=>"000011111",
  12771=>"111111111",
  12772=>"100111110",
  12773=>"111111111",
  12774=>"100000000",
  12775=>"011111000",
  12776=>"001000000",
  12777=>"111101110",
  12778=>"000101101",
  12779=>"101101101",
  12780=>"011000111",
  12781=>"001000000",
  12782=>"000000100",
  12783=>"011011011",
  12784=>"111111111",
  12785=>"001000111",
  12786=>"111111111",
  12787=>"010000000",
  12788=>"100110110",
  12789=>"000000001",
  12790=>"111111111",
  12791=>"111111100",
  12792=>"011000000",
  12793=>"001001000",
  12794=>"000000111",
  12795=>"000111000",
  12796=>"011111001",
  12797=>"001001000",
  12798=>"000000000",
  12799=>"000001001",
  12800=>"000000000",
  12801=>"000111011",
  12802=>"000000000",
  12803=>"000111111",
  12804=>"111000100",
  12805=>"011000011",
  12806=>"111111111",
  12807=>"111111111",
  12808=>"001111111",
  12809=>"000000000",
  12810=>"111110110",
  12811=>"010111100",
  12812=>"000000100",
  12813=>"111111010",
  12814=>"001001111",
  12815=>"110110111",
  12816=>"011000000",
  12817=>"111101101",
  12818=>"100100000",
  12819=>"000000000",
  12820=>"011101101",
  12821=>"100000100",
  12822=>"010000000",
  12823=>"000100100",
  12824=>"001001100",
  12825=>"011111111",
  12826=>"000000000",
  12827=>"001001000",
  12828=>"111111111",
  12829=>"000000000",
  12830=>"111001100",
  12831=>"111000111",
  12832=>"000000000",
  12833=>"001000000",
  12834=>"000010111",
  12835=>"000000000",
  12836=>"000000000",
  12837=>"100000111",
  12838=>"011011000",
  12839=>"101100101",
  12840=>"001000110",
  12841=>"111111111",
  12842=>"111111101",
  12843=>"000000000",
  12844=>"111111110",
  12845=>"111111111",
  12846=>"111111111",
  12847=>"011011011",
  12848=>"110110110",
  12849=>"111111111",
  12850=>"000011011",
  12851=>"001111111",
  12852=>"100100100",
  12853=>"000000000",
  12854=>"000000111",
  12855=>"001000100",
  12856=>"111111111",
  12857=>"111100000",
  12858=>"010000111",
  12859=>"000111011",
  12860=>"001000000",
  12861=>"000100100",
  12862=>"111111101",
  12863=>"000000100",
  12864=>"000000100",
  12865=>"100000000",
  12866=>"000000011",
  12867=>"001000001",
  12868=>"100111101",
  12869=>"111111111",
  12870=>"110100110",
  12871=>"111100100",
  12872=>"111010111",
  12873=>"111111111",
  12874=>"100000000",
  12875=>"000000000",
  12876=>"111001011",
  12877=>"110101101",
  12878=>"110010000",
  12879=>"111101001",
  12880=>"111111111",
  12881=>"001000000",
  12882=>"000000000",
  12883=>"111011111",
  12884=>"000000000",
  12885=>"011111111",
  12886=>"111111011",
  12887=>"100111110",
  12888=>"111111100",
  12889=>"111111111",
  12890=>"000000000",
  12891=>"000110101",
  12892=>"111111111",
  12893=>"011111011",
  12894=>"111111001",
  12895=>"010110110",
  12896=>"111111000",
  12897=>"010010010",
  12898=>"011000000",
  12899=>"000000000",
  12900=>"111111011",
  12901=>"000011111",
  12902=>"001000000",
  12903=>"000000000",
  12904=>"000000001",
  12905=>"111000000",
  12906=>"010100000",
  12907=>"111111111",
  12908=>"000011110",
  12909=>"111100100",
  12910=>"110000000",
  12911=>"011110110",
  12912=>"010111111",
  12913=>"110111111",
  12914=>"110111110",
  12915=>"111111110",
  12916=>"011101100",
  12917=>"110110100",
  12918=>"000000111",
  12919=>"000000000",
  12920=>"100000000",
  12921=>"000100110",
  12922=>"111111111",
  12923=>"000010110",
  12924=>"111000001",
  12925=>"111000100",
  12926=>"111111111",
  12927=>"000000000",
  12928=>"111110110",
  12929=>"001000110",
  12930=>"011001011",
  12931=>"011011000",
  12932=>"111100001",
  12933=>"111111111",
  12934=>"110110000",
  12935=>"110100000",
  12936=>"111111000",
  12937=>"000000000",
  12938=>"001101000",
  12939=>"100100111",
  12940=>"000110010",
  12941=>"000011011",
  12942=>"011001000",
  12943=>"100101111",
  12944=>"011000011",
  12945=>"111111111",
  12946=>"011111111",
  12947=>"000010010",
  12948=>"011111111",
  12949=>"110000000",
  12950=>"111111111",
  12951=>"010000000",
  12952=>"010111110",
  12953=>"101111011",
  12954=>"111111111",
  12955=>"010110000",
  12956=>"110100110",
  12957=>"001001000",
  12958=>"000000111",
  12959=>"111010011",
  12960=>"111111111",
  12961=>"111011010",
  12962=>"011011011",
  12963=>"111000000",
  12964=>"100000001",
  12965=>"011111111",
  12966=>"000000000",
  12967=>"111111100",
  12968=>"000000110",
  12969=>"100110111",
  12970=>"011000001",
  12971=>"000000000",
  12972=>"010000000",
  12973=>"000011011",
  12974=>"001000001",
  12975=>"000010000",
  12976=>"000000111",
  12977=>"111100000",
  12978=>"110110110",
  12979=>"000000000",
  12980=>"011011011",
  12981=>"010110100",
  12982=>"111100100",
  12983=>"011011111",
  12984=>"000000100",
  12985=>"110000000",
  12986=>"110100111",
  12987=>"001100000",
  12988=>"000100111",
  12989=>"011011111",
  12990=>"010111111",
  12991=>"000000100",
  12992=>"000000000",
  12993=>"111010010",
  12994=>"110111110",
  12995=>"111111111",
  12996=>"111110111",
  12997=>"111111000",
  12998=>"111000111",
  12999=>"000000111",
  13000=>"110111111",
  13001=>"001111111",
  13002=>"111011011",
  13003=>"000000000",
  13004=>"011001000",
  13005=>"111000000",
  13006=>"111000000",
  13007=>"000111111",
  13008=>"000011111",
  13009=>"011111011",
  13010=>"000010010",
  13011=>"111111111",
  13012=>"001101101",
  13013=>"000000001",
  13014=>"111111111",
  13015=>"001011001",
  13016=>"010000100",
  13017=>"000101000",
  13018=>"000000000",
  13019=>"001001111",
  13020=>"111111111",
  13021=>"001001111",
  13022=>"011011011",
  13023=>"000110100",
  13024=>"000110111",
  13025=>"110111111",
  13026=>"111111111",
  13027=>"011111111",
  13028=>"100000000",
  13029=>"011111110",
  13030=>"001000000",
  13031=>"001000000",
  13032=>"000001000",
  13033=>"111110100",
  13034=>"100100100",
  13035=>"111110111",
  13036=>"110111111",
  13037=>"110010000",
  13038=>"001000000",
  13039=>"000011000",
  13040=>"000000000",
  13041=>"111111100",
  13042=>"011011001",
  13043=>"011011111",
  13044=>"100000000",
  13045=>"000010000",
  13046=>"000111111",
  13047=>"010011111",
  13048=>"111001011",
  13049=>"000000000",
  13050=>"011111111",
  13051=>"000000001",
  13052=>"100011001",
  13053=>"000000000",
  13054=>"011111011",
  13055=>"000000000",
  13056=>"001111111",
  13057=>"100111101",
  13058=>"111111110",
  13059=>"111111000",
  13060=>"010010000",
  13061=>"000110000",
  13062=>"100100001",
  13063=>"110000111",
  13064=>"011111111",
  13065=>"000000000",
  13066=>"000010110",
  13067=>"000000000",
  13068=>"110110100",
  13069=>"111111011",
  13070=>"111111110",
  13071=>"000001000",
  13072=>"111111100",
  13073=>"000110110",
  13074=>"000000000",
  13075=>"011111111",
  13076=>"110111111",
  13077=>"000110010",
  13078=>"100111111",
  13079=>"000100100",
  13080=>"011111011",
  13081=>"000101001",
  13082=>"011111111",
  13083=>"000110110",
  13084=>"011111111",
  13085=>"000000000",
  13086=>"111111111",
  13087=>"000000011",
  13088=>"111001011",
  13089=>"000000010",
  13090=>"000111100",
  13091=>"111110011",
  13092=>"000000100",
  13093=>"000000100",
  13094=>"000000000",
  13095=>"111111111",
  13096=>"110000000",
  13097=>"111111111",
  13098=>"111111111",
  13099=>"111111111",
  13100=>"111111110",
  13101=>"101100100",
  13102=>"000000000",
  13103=>"000100000",
  13104=>"111111110",
  13105=>"110000110",
  13106=>"010000000",
  13107=>"011000000",
  13108=>"000000000",
  13109=>"111011110",
  13110=>"111111101",
  13111=>"000111111",
  13112=>"000000000",
  13113=>"000101111",
  13114=>"100111111",
  13115=>"000000000",
  13116=>"111111111",
  13117=>"011011111",
  13118=>"000100000",
  13119=>"011000000",
  13120=>"101111111",
  13121=>"011011001",
  13122=>"000110000",
  13123=>"111111000",
  13124=>"000111111",
  13125=>"000000001",
  13126=>"111000101",
  13127=>"111111000",
  13128=>"000000000",
  13129=>"011111111",
  13130=>"010010010",
  13131=>"011111110",
  13132=>"011100100",
  13133=>"000000000",
  13134=>"011111110",
  13135=>"001110100",
  13136=>"111111111",
  13137=>"111110000",
  13138=>"000000111",
  13139=>"110111100",
  13140=>"111000000",
  13141=>"111001111",
  13142=>"011000011",
  13143=>"111000001",
  13144=>"000000000",
  13145=>"110111111",
  13146=>"000000011",
  13147=>"011111000",
  13148=>"000000010",
  13149=>"111100100",
  13150=>"000000011",
  13151=>"110111011",
  13152=>"000000000",
  13153=>"000000000",
  13154=>"111111011",
  13155=>"111111111",
  13156=>"000011111",
  13157=>"111111111",
  13158=>"000001001",
  13159=>"000000111",
  13160=>"101111111",
  13161=>"111111111",
  13162=>"000000111",
  13163=>"001001011",
  13164=>"111000000",
  13165=>"110011111",
  13166=>"100111111",
  13167=>"111101111",
  13168=>"110111111",
  13169=>"001000100",
  13170=>"000000011",
  13171=>"000001000",
  13172=>"110110011",
  13173=>"111111111",
  13174=>"001001100",
  13175=>"111111011",
  13176=>"111001000",
  13177=>"011100100",
  13178=>"111100101",
  13179=>"010000100",
  13180=>"000000000",
  13181=>"111100000",
  13182=>"001001011",
  13183=>"001000000",
  13184=>"110011111",
  13185=>"111111110",
  13186=>"110110000",
  13187=>"000110001",
  13188=>"111111111",
  13189=>"010010000",
  13190=>"000000000",
  13191=>"000010000",
  13192=>"111111110",
  13193=>"000110110",
  13194=>"001001011",
  13195=>"111111111",
  13196=>"111111111",
  13197=>"000001000",
  13198=>"000110110",
  13199=>"011000000",
  13200=>"000000000",
  13201=>"001001001",
  13202=>"000011011",
  13203=>"001001000",
  13204=>"000000000",
  13205=>"111100000",
  13206=>"111011111",
  13207=>"011011001",
  13208=>"100110110",
  13209=>"111111111",
  13210=>"000000000",
  13211=>"000100111",
  13212=>"111111011",
  13213=>"101111111",
  13214=>"110000000",
  13215=>"101111000",
  13216=>"111111000",
  13217=>"010011011",
  13218=>"001111111",
  13219=>"011000111",
  13220=>"000000000",
  13221=>"000000000",
  13222=>"000000000",
  13223=>"110110110",
  13224=>"011111110",
  13225=>"000000111",
  13226=>"001011111",
  13227=>"111111000",
  13228=>"010000110",
  13229=>"000111111",
  13230=>"001000110",
  13231=>"111000000",
  13232=>"011000000",
  13233=>"000000110",
  13234=>"110111001",
  13235=>"000011111",
  13236=>"111111111",
  13237=>"000110110",
  13238=>"001000000",
  13239=>"011011000",
  13240=>"011111111",
  13241=>"101001000",
  13242=>"000100111",
  13243=>"001000000",
  13244=>"111111111",
  13245=>"111001001",
  13246=>"100110111",
  13247=>"101101100",
  13248=>"000000000",
  13249=>"001000000",
  13250=>"000000000",
  13251=>"111111111",
  13252=>"001001011",
  13253=>"111111111",
  13254=>"000111111",
  13255=>"111111111",
  13256=>"000000110",
  13257=>"111111111",
  13258=>"011110110",
  13259=>"111101101",
  13260=>"111111010",
  13261=>"011111111",
  13262=>"000111111",
  13263=>"000000000",
  13264=>"001010111",
  13265=>"110000110",
  13266=>"001000000",
  13267=>"010000000",
  13268=>"000000000",
  13269=>"000100111",
  13270=>"111001001",
  13271=>"111101011",
  13272=>"001001001",
  13273=>"111001000",
  13274=>"110001011",
  13275=>"111111110",
  13276=>"000111110",
  13277=>"011111110",
  13278=>"111000000",
  13279=>"100110110",
  13280=>"110100000",
  13281=>"110100100",
  13282=>"111111111",
  13283=>"000000000",
  13284=>"011011011",
  13285=>"111101001",
  13286=>"111111000",
  13287=>"000000111",
  13288=>"111011110",
  13289=>"000000000",
  13290=>"011111111",
  13291=>"010000100",
  13292=>"010011111",
  13293=>"111111101",
  13294=>"110111110",
  13295=>"110011111",
  13296=>"111100100",
  13297=>"001001101",
  13298=>"011011111",
  13299=>"111110110",
  13300=>"011000000",
  13301=>"011011001",
  13302=>"111110000",
  13303=>"011111110",
  13304=>"111111111",
  13305=>"111110110",
  13306=>"110111111",
  13307=>"110111000",
  13308=>"000000000",
  13309=>"100100111",
  13310=>"011111111",
  13311=>"000001001",
  13312=>"001000000",
  13313=>"111111001",
  13314=>"000101101",
  13315=>"111111111",
  13316=>"010110110",
  13317=>"111110110",
  13318=>"111001000",
  13319=>"111000101",
  13320=>"000111000",
  13321=>"100111111",
  13322=>"011000000",
  13323=>"000000000",
  13324=>"000110000",
  13325=>"101111111",
  13326=>"111010011",
  13327=>"000111000",
  13328=>"000000110",
  13329=>"000001010",
  13330=>"010000111",
  13331=>"000111111",
  13332=>"010000000",
  13333=>"111111000",
  13334=>"000000111",
  13335=>"000000001",
  13336=>"001000000",
  13337=>"001101101",
  13338=>"101001111",
  13339=>"001000010",
  13340=>"000011011",
  13341=>"111000000",
  13342=>"000001001",
  13343=>"000111000",
  13344=>"000000000",
  13345=>"111110110",
  13346=>"111011110",
  13347=>"111001001",
  13348=>"110011110",
  13349=>"000100000",
  13350=>"001001000",
  13351=>"101001001",
  13352=>"000001000",
  13353=>"111000000",
  13354=>"111111111",
  13355=>"111100100",
  13356=>"111010111",
  13357=>"000000111",
  13358=>"001100101",
  13359=>"000000011",
  13360=>"101100001",
  13361=>"111000001",
  13362=>"001000001",
  13363=>"000000010",
  13364=>"000000111",
  13365=>"000001001",
  13366=>"101101000",
  13367=>"110110000",
  13368=>"001001000",
  13369=>"000111111",
  13370=>"000000000",
  13371=>"111111111",
  13372=>"000000001",
  13373=>"111100110",
  13374=>"011111111",
  13375=>"111000000",
  13376=>"100000000",
  13377=>"111111111",
  13378=>"000111111",
  13379=>"000110111",
  13380=>"000000000",
  13381=>"100111110",
  13382=>"101000000",
  13383=>"111111000",
  13384=>"111111111",
  13385=>"011000111",
  13386=>"111001111",
  13387=>"101001011",
  13388=>"000000000",
  13389=>"111111000",
  13390=>"000001011",
  13391=>"000000010",
  13392=>"001000001",
  13393=>"000111011",
  13394=>"100000000",
  13395=>"000001011",
  13396=>"011111010",
  13397=>"111000000",
  13398=>"001001101",
  13399=>"111100110",
  13400=>"000000001",
  13401=>"001000100",
  13402=>"000000000",
  13403=>"000000000",
  13404=>"111000000",
  13405=>"000111111",
  13406=>"000000000",
  13407=>"111111111",
  13408=>"000111111",
  13409=>"010000000",
  13410=>"111111101",
  13411=>"000101111",
  13412=>"001000000",
  13413=>"000111010",
  13414=>"000000000",
  13415=>"000010000",
  13416=>"111111111",
  13417=>"000011110",
  13418=>"000001011",
  13419=>"000001011",
  13420=>"011011011",
  13421=>"111111000",
  13422=>"111110000",
  13423=>"000000011",
  13424=>"111111000",
  13425=>"001001000",
  13426=>"111111111",
  13427=>"000000001",
  13428=>"011011011",
  13429=>"000010000",
  13430=>"000111010",
  13431=>"011000000",
  13432=>"110000000",
  13433=>"111111111",
  13434=>"001000000",
  13435=>"111110110",
  13436=>"000001001",
  13437=>"110100110",
  13438=>"000000000",
  13439=>"110010001",
  13440=>"000000000",
  13441=>"000000111",
  13442=>"111000000",
  13443=>"110100111",
  13444=>"111000000",
  13445=>"111000110",
  13446=>"111111111",
  13447=>"001000000",
  13448=>"001001001",
  13449=>"111111111",
  13450=>"000000000",
  13451=>"000000111",
  13452=>"111011001",
  13453=>"100000111",
  13454=>"111000000",
  13455=>"000000000",
  13456=>"000000111",
  13457=>"000000111",
  13458=>"010000000",
  13459=>"000000100",
  13460=>"000000000",
  13461=>"000111111",
  13462=>"111000000",
  13463=>"111001000",
  13464=>"001000000",
  13465=>"111100101",
  13466=>"000000000",
  13467=>"000000000",
  13468=>"111001000",
  13469=>"111100000",
  13470=>"000000000",
  13471=>"110111010",
  13472=>"000000000",
  13473=>"000000000",
  13474=>"111111000",
  13475=>"010000000",
  13476=>"000000000",
  13477=>"111111101",
  13478=>"001111111",
  13479=>"000110100",
  13480=>"110000100",
  13481=>"000000110",
  13482=>"000000000",
  13483=>"000100100",
  13484=>"000011111",
  13485=>"000100111",
  13486=>"111101111",
  13487=>"111101000",
  13488=>"011000111",
  13489=>"100110111",
  13490=>"010111010",
  13491=>"000000111",
  13492=>"000000101",
  13493=>"101000000",
  13494=>"001000000",
  13495=>"111101100",
  13496=>"111111101",
  13497=>"111111000",
  13498=>"000001111",
  13499=>"001111100",
  13500=>"111111011",
  13501=>"111000000",
  13502=>"111001000",
  13503=>"110111111",
  13504=>"111000000",
  13505=>"011100101",
  13506=>"111000001",
  13507=>"001001000",
  13508=>"000000110",
  13509=>"100100000",
  13510=>"110000010",
  13511=>"000000111",
  13512=>"111111000",
  13513=>"111011000",
  13514=>"000000000",
  13515=>"000000000",
  13516=>"100101000",
  13517=>"000001110",
  13518=>"111000000",
  13519=>"111010001",
  13520=>"000100000",
  13521=>"110100111",
  13522=>"011010000",
  13523=>"000000111",
  13524=>"000000000",
  13525=>"000111111",
  13526=>"101111111",
  13527=>"110110111",
  13528=>"000000011",
  13529=>"001001111",
  13530=>"100000000",
  13531=>"000000000",
  13532=>"000111111",
  13533=>"000000111",
  13534=>"001011011",
  13535=>"000000000",
  13536=>"000011011",
  13537=>"000000110",
  13538=>"101101000",
  13539=>"111111111",
  13540=>"111000110",
  13541=>"110111000",
  13542=>"000000000",
  13543=>"001111111",
  13544=>"111011000",
  13545=>"111111000",
  13546=>"101001111",
  13547=>"111000001",
  13548=>"111010011",
  13549=>"000000000",
  13550=>"011111110",
  13551=>"111111111",
  13552=>"111111111",
  13553=>"000001000",
  13554=>"001111101",
  13555=>"000001111",
  13556=>"111110000",
  13557=>"111111100",
  13558=>"000111111",
  13559=>"111000000",
  13560=>"011000000",
  13561=>"000001000",
  13562=>"111001000",
  13563=>"000000110",
  13564=>"000100111",
  13565=>"111011111",
  13566=>"001111101",
  13567=>"111111111",
  13568=>"111111101",
  13569=>"100001001",
  13570=>"000000000",
  13571=>"000111010",
  13572=>"111111111",
  13573=>"111011001",
  13574=>"111111111",
  13575=>"000000000",
  13576=>"000000111",
  13577=>"011000000",
  13578=>"111111000",
  13579=>"000100100",
  13580=>"000000100",
  13581=>"000000000",
  13582=>"000000011",
  13583=>"000000010",
  13584=>"000111111",
  13585=>"111111001",
  13586=>"111000001",
  13587=>"111001000",
  13588=>"000100111",
  13589=>"111011000",
  13590=>"011001101",
  13591=>"000000000",
  13592=>"001011111",
  13593=>"111000101",
  13594=>"111010000",
  13595=>"000000000",
  13596=>"000000110",
  13597=>"000000000",
  13598=>"000001111",
  13599=>"000110111",
  13600=>"100100000",
  13601=>"000110111",
  13602=>"000010000",
  13603=>"101000000",
  13604=>"111100110",
  13605=>"001001111",
  13606=>"111111000",
  13607=>"100000110",
  13608=>"000111111",
  13609=>"000000000",
  13610=>"000000001",
  13611=>"000100111",
  13612=>"001000000",
  13613=>"010011110",
  13614=>"000000011",
  13615=>"001111111",
  13616=>"000111111",
  13617=>"110000000",
  13618=>"000111111",
  13619=>"000000000",
  13620=>"011000001",
  13621=>"111100000",
  13622=>"000111111",
  13623=>"001000000",
  13624=>"000010000",
  13625=>"111111000",
  13626=>"011111000",
  13627=>"000101101",
  13628=>"111111111",
  13629=>"111111100",
  13630=>"111110110",
  13631=>"111111000",
  13632=>"111110000",
  13633=>"100100101",
  13634=>"100000111",
  13635=>"000100100",
  13636=>"101111111",
  13637=>"001000000",
  13638=>"111111011",
  13639=>"111001101",
  13640=>"110111111",
  13641=>"010000111",
  13642=>"000100001",
  13643=>"000100110",
  13644=>"111111000",
  13645=>"111111000",
  13646=>"111000000",
  13647=>"101001111",
  13648=>"100111001",
  13649=>"111000001",
  13650=>"000001111",
  13651=>"000000011",
  13652=>"000000110",
  13653=>"010000001",
  13654=>"000111000",
  13655=>"000111111",
  13656=>"101111000",
  13657=>"001000111",
  13658=>"010000001",
  13659=>"111111111",
  13660=>"111111000",
  13661=>"111000000",
  13662=>"111001001",
  13663=>"111000000",
  13664=>"000000010",
  13665=>"000100000",
  13666=>"100000100",
  13667=>"111100100",
  13668=>"000011111",
  13669=>"001001001",
  13670=>"000000000",
  13671=>"000000100",
  13672=>"000011111",
  13673=>"111001001",
  13674=>"000011000",
  13675=>"111001001",
  13676=>"011011011",
  13677=>"000110001",
  13678=>"000000110",
  13679=>"111111000",
  13680=>"000000011",
  13681=>"000000000",
  13682=>"001011000",
  13683=>"000000100",
  13684=>"111111111",
  13685=>"101100111",
  13686=>"000000000",
  13687=>"111000001",
  13688=>"100000101",
  13689=>"000000000",
  13690=>"111010000",
  13691=>"000001001",
  13692=>"111111000",
  13693=>"111111111",
  13694=>"000011111",
  13695=>"000001011",
  13696=>"111001001",
  13697=>"001000000",
  13698=>"100111011",
  13699=>"111000000",
  13700=>"001111111",
  13701=>"001000001",
  13702=>"100000000",
  13703=>"110000000",
  13704=>"111111000",
  13705=>"111111101",
  13706=>"101000000",
  13707=>"111111111",
  13708=>"111111111",
  13709=>"000011110",
  13710=>"111001000",
  13711=>"000000000",
  13712=>"000111111",
  13713=>"001000000",
  13714=>"010110010",
  13715=>"100100100",
  13716=>"000000000",
  13717=>"000000000",
  13718=>"111111101",
  13719=>"000101001",
  13720=>"111111110",
  13721=>"000000111",
  13722=>"111111110",
  13723=>"000000111",
  13724=>"111011111",
  13725=>"011111111",
  13726=>"000000001",
  13727=>"111000000",
  13728=>"000011000",
  13729=>"110100000",
  13730=>"001000000",
  13731=>"000111111",
  13732=>"111100100",
  13733=>"000000100",
  13734=>"111000000",
  13735=>"000111111",
  13736=>"111111111",
  13737=>"001111111",
  13738=>"111111111",
  13739=>"000000001",
  13740=>"000110111",
  13741=>"001111111",
  13742=>"000000111",
  13743=>"000001001",
  13744=>"000000100",
  13745=>"000000000",
  13746=>"000000000",
  13747=>"011111011",
  13748=>"111000000",
  13749=>"101001010",
  13750=>"111100100",
  13751=>"111101000",
  13752=>"111111000",
  13753=>"111001000",
  13754=>"101101001",
  13755=>"111000000",
  13756=>"111111110",
  13757=>"101000000",
  13758=>"000110001",
  13759=>"001101101",
  13760=>"110111000",
  13761=>"111011000",
  13762=>"111111111",
  13763=>"111111111",
  13764=>"111111101",
  13765=>"000111111",
  13766=>"000111110",
  13767=>"100110110",
  13768=>"000100111",
  13769=>"111001000",
  13770=>"000000111",
  13771=>"111000000",
  13772=>"111111000",
  13773=>"111111100",
  13774=>"001111111",
  13775=>"011000000",
  13776=>"100000000",
  13777=>"000100000",
  13778=>"100001111",
  13779=>"111111111",
  13780=>"000100100",
  13781=>"111111111",
  13782=>"110111111",
  13783=>"000000111",
  13784=>"111000000",
  13785=>"000001001",
  13786=>"000000000",
  13787=>"000101101",
  13788=>"001001000",
  13789=>"001011010",
  13790=>"111000001",
  13791=>"001011100",
  13792=>"111000000",
  13793=>"000010000",
  13794=>"100000000",
  13795=>"111011010",
  13796=>"000000000",
  13797=>"111111111",
  13798=>"111001000",
  13799=>"000000111",
  13800=>"001111111",
  13801=>"111111111",
  13802=>"011000000",
  13803=>"000000111",
  13804=>"110100111",
  13805=>"000001010",
  13806=>"111111000",
  13807=>"111111111",
  13808=>"011111111",
  13809=>"001001000",
  13810=>"111111111",
  13811=>"000000011",
  13812=>"000110111",
  13813=>"011000000",
  13814=>"000000111",
  13815=>"011001000",
  13816=>"000000000",
  13817=>"110000111",
  13818=>"111011001",
  13819=>"111111000",
  13820=>"001111111",
  13821=>"000001011",
  13822=>"111101111",
  13823=>"101000000",
  13824=>"001001001",
  13825=>"000000100",
  13826=>"111100111",
  13827=>"000000000",
  13828=>"111111000",
  13829=>"000000111",
  13830=>"000001011",
  13831=>"111000111",
  13832=>"001000111",
  13833=>"111000000",
  13834=>"000000000",
  13835=>"000110000",
  13836=>"000111110",
  13837=>"000100111",
  13838=>"110001000",
  13839=>"111111100",
  13840=>"111111000",
  13841=>"111111111",
  13842=>"000101111",
  13843=>"101011001",
  13844=>"000000111",
  13845=>"100100111",
  13846=>"111111000",
  13847=>"111111001",
  13848=>"101111110",
  13849=>"011111110",
  13850=>"000000111",
  13851=>"111110100",
  13852=>"100111001",
  13853=>"111111000",
  13854=>"110001111",
  13855=>"010111010",
  13856=>"000100111",
  13857=>"111111111",
  13858=>"000000000",
  13859=>"111111110",
  13860=>"110111111",
  13861=>"111111000",
  13862=>"111110111",
  13863=>"111110000",
  13864=>"110111111",
  13865=>"100000111",
  13866=>"100101001",
  13867=>"101000000",
  13868=>"011111011",
  13869=>"111111010",
  13870=>"000001001",
  13871=>"000010110",
  13872=>"101101000",
  13873=>"000000111",
  13874=>"110000000",
  13875=>"111111111",
  13876=>"011111111",
  13877=>"010010000",
  13878=>"001000001",
  13879=>"011111001",
  13880=>"111111110",
  13881=>"111110100",
  13882=>"110111111",
  13883=>"111111111",
  13884=>"000000001",
  13885=>"111111111",
  13886=>"000111111",
  13887=>"111011111",
  13888=>"000111110",
  13889=>"110000111",
  13890=>"000000000",
  13891=>"110000000",
  13892=>"111011000",
  13893=>"110110110",
  13894=>"000001101",
  13895=>"000000000",
  13896=>"111111001",
  13897=>"100000111",
  13898=>"001000000",
  13899=>"111111111",
  13900=>"000000000",
  13901=>"000000000",
  13902=>"101111011",
  13903=>"111111001",
  13904=>"001100111",
  13905=>"111101000",
  13906=>"111111000",
  13907=>"111111110",
  13908=>"000000000",
  13909=>"110100100",
  13910=>"000000001",
  13911=>"000000101",
  13912=>"101111111",
  13913=>"101001111",
  13914=>"000000111",
  13915=>"000000111",
  13916=>"111111111",
  13917=>"111000100",
  13918=>"111111111",
  13919=>"110110000",
  13920=>"100111111",
  13921=>"110111000",
  13922=>"100000000",
  13923=>"000000010",
  13924=>"111110000",
  13925=>"111100000",
  13926=>"011000000",
  13927=>"100000000",
  13928=>"001111111",
  13929=>"000001001",
  13930=>"111111111",
  13931=>"000000000",
  13932=>"011000011",
  13933=>"000110000",
  13934=>"111001001",
  13935=>"001111111",
  13936=>"010000000",
  13937=>"001000111",
  13938=>"000000001",
  13939=>"001111111",
  13940=>"011111011",
  13941=>"000100000",
  13942=>"111011001",
  13943=>"000001000",
  13944=>"000000000",
  13945=>"111111110",
  13946=>"100000000",
  13947=>"101001111",
  13948=>"110100000",
  13949=>"000000000",
  13950=>"000000000",
  13951=>"101110000",
  13952=>"001000000",
  13953=>"111111111",
  13954=>"111000000",
  13955=>"111111111",
  13956=>"000000000",
  13957=>"001000000",
  13958=>"001000000",
  13959=>"001101111",
  13960=>"000000111",
  13961=>"100101101",
  13962=>"101111111",
  13963=>"111111000",
  13964=>"100111111",
  13965=>"000001000",
  13966=>"011000000",
  13967=>"000111110",
  13968=>"000000000",
  13969=>"000000100",
  13970=>"111111111",
  13971=>"010000000",
  13972=>"000000000",
  13973=>"000100000",
  13974=>"100101100",
  13975=>"000000100",
  13976=>"001000000",
  13977=>"000000011",
  13978=>"000000001",
  13979=>"011001011",
  13980=>"101000000",
  13981=>"001000000",
  13982=>"111111000",
  13983=>"110111111",
  13984=>"000110111",
  13985=>"000000001",
  13986=>"111111000",
  13987=>"001000000",
  13988=>"001001001",
  13989=>"110111111",
  13990=>"101101101",
  13991=>"001001001",
  13992=>"110000110",
  13993=>"001000000",
  13994=>"000000001",
  13995=>"111111000",
  13996=>"100000000",
  13997=>"110110111",
  13998=>"111111111",
  13999=>"001111000",
  14000=>"111111111",
  14001=>"100111001",
  14002=>"111111010",
  14003=>"111111001",
  14004=>"110000110",
  14005=>"000100000",
  14006=>"010111111",
  14007=>"000000111",
  14008=>"111111111",
  14009=>"111111000",
  14010=>"101001101",
  14011=>"011010001",
  14012=>"100000001",
  14013=>"111111000",
  14014=>"110110000",
  14015=>"000011111",
  14016=>"000100111",
  14017=>"001000001",
  14018=>"000111010",
  14019=>"001000000",
  14020=>"111000100",
  14021=>"000111000",
  14022=>"101000011",
  14023=>"000011100",
  14024=>"111011000",
  14025=>"111011111",
  14026=>"001000010",
  14027=>"000011111",
  14028=>"011111000",
  14029=>"000110010",
  14030=>"110100100",
  14031=>"000111111",
  14032=>"111000000",
  14033=>"110100000",
  14034=>"000000000",
  14035=>"100000111",
  14036=>"011100100",
  14037=>"111111111",
  14038=>"000000000",
  14039=>"000000001",
  14040=>"010000111",
  14041=>"000110011",
  14042=>"111111111",
  14043=>"111111111",
  14044=>"111111000",
  14045=>"101101111",
  14046=>"111111101",
  14047=>"000000001",
  14048=>"011111000",
  14049=>"001001011",
  14050=>"010000000",
  14051=>"000000111",
  14052=>"000001011",
  14053=>"000000100",
  14054=>"000111000",
  14055=>"010010111",
  14056=>"111111000",
  14057=>"111001100",
  14058=>"000000111",
  14059=>"110111111",
  14060=>"011001000",
  14061=>"000000111",
  14062=>"011000111",
  14063=>"000000000",
  14064=>"000011011",
  14065=>"111000000",
  14066=>"000100000",
  14067=>"000000000",
  14068=>"111111111",
  14069=>"001001001",
  14070=>"011110000",
  14071=>"101111111",
  14072=>"110110000",
  14073=>"111111000",
  14074=>"011000000",
  14075=>"000100000",
  14076=>"001011011",
  14077=>"001001000",
  14078=>"000000110",
  14079=>"000111111",
  14080=>"111111010",
  14081=>"101001000",
  14082=>"111110111",
  14083=>"111000111",
  14084=>"111111110",
  14085=>"101111001",
  14086=>"111000101",
  14087=>"001000111",
  14088=>"001000000",
  14089=>"110100000",
  14090=>"000000101",
  14091=>"111111111",
  14092=>"000000000",
  14093=>"000000001",
  14094=>"000000001",
  14095=>"001000000",
  14096=>"000000000",
  14097=>"001000000",
  14098=>"111111111",
  14099=>"001011111",
  14100=>"001000000",
  14101=>"000000000",
  14102=>"001101101",
  14103=>"000000111",
  14104=>"111111110",
  14105=>"111111100",
  14106=>"111101000",
  14107=>"000111111",
  14108=>"001111111",
  14109=>"111111111",
  14110=>"000000100",
  14111=>"111111100",
  14112=>"110111000",
  14113=>"001001000",
  14114=>"000000001",
  14115=>"111111000",
  14116=>"111101001",
  14117=>"000000000",
  14118=>"111111111",
  14119=>"000000000",
  14120=>"000000000",
  14121=>"000001001",
  14122=>"111111000",
  14123=>"000111111",
  14124=>"110100101",
  14125=>"111101000",
  14126=>"111111111",
  14127=>"000001111",
  14128=>"001111110",
  14129=>"110111001",
  14130=>"111111111",
  14131=>"111111010",
  14132=>"000000000",
  14133=>"000000111",
  14134=>"000000000",
  14135=>"001000000",
  14136=>"111110000",
  14137=>"100000111",
  14138=>"000000000",
  14139=>"111111100",
  14140=>"000000111",
  14141=>"010010000",
  14142=>"111100001",
  14143=>"111011001",
  14144=>"111011000",
  14145=>"000000111",
  14146=>"111111010",
  14147=>"110111111",
  14148=>"111011111",
  14149=>"010100000",
  14150=>"000110110",
  14151=>"001000111",
  14152=>"101001001",
  14153=>"000000000",
  14154=>"111111000",
  14155=>"100001001",
  14156=>"000000100",
  14157=>"111110000",
  14158=>"111111000",
  14159=>"000111000",
  14160=>"110010011",
  14161=>"000100100",
  14162=>"110110111",
  14163=>"111111111",
  14164=>"101111010",
  14165=>"011011111",
  14166=>"111111110",
  14167=>"001000001",
  14168=>"100000000",
  14169=>"111111001",
  14170=>"001000000",
  14171=>"000000000",
  14172=>"000010000",
  14173=>"011111111",
  14174=>"001000000",
  14175=>"000000000",
  14176=>"000000000",
  14177=>"111111000",
  14178=>"001011011",
  14179=>"111101111",
  14180=>"000011001",
  14181=>"001001000",
  14182=>"000000000",
  14183=>"111111111",
  14184=>"001001001",
  14185=>"001000000",
  14186=>"001000000",
  14187=>"101101001",
  14188=>"000000111",
  14189=>"101001101",
  14190=>"010010010",
  14191=>"111000000",
  14192=>"000101111",
  14193=>"111111001",
  14194=>"001011111",
  14195=>"111111100",
  14196=>"100000101",
  14197=>"000000101",
  14198=>"111111011",
  14199=>"100110100",
  14200=>"000000000",
  14201=>"000000111",
  14202=>"000000001",
  14203=>"000000110",
  14204=>"111101000",
  14205=>"000100000",
  14206=>"111100000",
  14207=>"000001001",
  14208=>"001000000",
  14209=>"000110111",
  14210=>"000000111",
  14211=>"101001011",
  14212=>"000011111",
  14213=>"100100000",
  14214=>"000010000",
  14215=>"111100000",
  14216=>"111111111",
  14217=>"111111001",
  14218=>"001011111",
  14219=>"000001111",
  14220=>"001000000",
  14221=>"000000000",
  14222=>"111111000",
  14223=>"000000000",
  14224=>"000000000",
  14225=>"000110110",
  14226=>"001111001",
  14227=>"000000001",
  14228=>"001000000",
  14229=>"000000010",
  14230=>"000000011",
  14231=>"001001000",
  14232=>"000000001",
  14233=>"111111000",
  14234=>"111111111",
  14235=>"001001111",
  14236=>"000000100",
  14237=>"011111111",
  14238=>"001000000",
  14239=>"110111111",
  14240=>"110111111",
  14241=>"111111000",
  14242=>"111111111",
  14243=>"000000010",
  14244=>"111011111",
  14245=>"111111000",
  14246=>"111101000",
  14247=>"010010000",
  14248=>"001001101",
  14249=>"000000001",
  14250=>"111111000",
  14251=>"111111000",
  14252=>"000000000",
  14253=>"000000000",
  14254=>"011001111",
  14255=>"000000100",
  14256=>"100000111",
  14257=>"111101000",
  14258=>"111111110",
  14259=>"111001000",
  14260=>"000000001",
  14261=>"000000001",
  14262=>"000000001",
  14263=>"000111000",
  14264=>"011110000",
  14265=>"111001000",
  14266=>"000000000",
  14267=>"111000000",
  14268=>"100111110",
  14269=>"000111111",
  14270=>"111111111",
  14271=>"001000001",
  14272=>"000000101",
  14273=>"111111111",
  14274=>"000000000",
  14275=>"111001111",
  14276=>"001001111",
  14277=>"111000100",
  14278=>"001000111",
  14279=>"000000000",
  14280=>"000000111",
  14281=>"110111010",
  14282=>"001001101",
  14283=>"000000101",
  14284=>"000000000",
  14285=>"000000000",
  14286=>"110100000",
  14287=>"111111110",
  14288=>"111111000",
  14289=>"111111011",
  14290=>"000000100",
  14291=>"000000000",
  14292=>"111101101",
  14293=>"111111111",
  14294=>"000000100",
  14295=>"111110100",
  14296=>"011011001",
  14297=>"111111110",
  14298=>"000000000",
  14299=>"111010011",
  14300=>"000000000",
  14301=>"001000001",
  14302=>"101000001",
  14303=>"000100011",
  14304=>"000100000",
  14305=>"000000000",
  14306=>"001001000",
  14307=>"101000000",
  14308=>"101000111",
  14309=>"000000000",
  14310=>"111111111",
  14311=>"000000000",
  14312=>"000000000",
  14313=>"000000000",
  14314=>"100100110",
  14315=>"010000000",
  14316=>"010000000",
  14317=>"001011001",
  14318=>"101001111",
  14319=>"000000001",
  14320=>"000000000",
  14321=>"000001101",
  14322=>"111111000",
  14323=>"111011001",
  14324=>"111111111",
  14325=>"000000000",
  14326=>"000000000",
  14327=>"111111100",
  14328=>"000000000",
  14329=>"000000010",
  14330=>"001000001",
  14331=>"000000101",
  14332=>"111011010",
  14333=>"000100111",
  14334=>"000000000",
  14335=>"100100110",
  14336=>"111111111",
  14337=>"111111111",
  14338=>"000100000",
  14339=>"111100000",
  14340=>"000000000",
  14341=>"010000000",
  14342=>"000000100",
  14343=>"111111111",
  14344=>"000000000",
  14345=>"000000000",
  14346=>"110111111",
  14347=>"000001000",
  14348=>"100110101",
  14349=>"111111010",
  14350=>"111101001",
  14351=>"001001001",
  14352=>"001111010",
  14353=>"111011011",
  14354=>"100100111",
  14355=>"010010000",
  14356=>"111111111",
  14357=>"100000000",
  14358=>"001101111",
  14359=>"000011011",
  14360=>"001101000",
  14361=>"000100001",
  14362=>"111101001",
  14363=>"000000000",
  14364=>"110111000",
  14365=>"000111111",
  14366=>"000000000",
  14367=>"011010010",
  14368=>"100100111",
  14369=>"111111111",
  14370=>"000100000",
  14371=>"000000000",
  14372=>"001000000",
  14373=>"111000000",
  14374=>"100000000",
  14375=>"000000000",
  14376=>"111111111",
  14377=>"000000000",
  14378=>"111001000",
  14379=>"000000000",
  14380=>"000000100",
  14381=>"111111111",
  14382=>"000100110",
  14383=>"111110010",
  14384=>"000000011",
  14385=>"000000111",
  14386=>"000100101",
  14387=>"111011011",
  14388=>"110110111",
  14389=>"000000001",
  14390=>"000010000",
  14391=>"000000000",
  14392=>"000001111",
  14393=>"111000111",
  14394=>"000001001",
  14395=>"111001000",
  14396=>"000010111",
  14397=>"000000000",
  14398=>"010111110",
  14399=>"110111111",
  14400=>"000000000",
  14401=>"000000000",
  14402=>"100110111",
  14403=>"000000000",
  14404=>"000000000",
  14405=>"110110100",
  14406=>"111111111",
  14407=>"111111111",
  14408=>"001000000",
  14409=>"000000000",
  14410=>"000000000",
  14411=>"001001000",
  14412=>"000000000",
  14413=>"000000000",
  14414=>"000000000",
  14415=>"000000000",
  14416=>"000000000",
  14417=>"011111111",
  14418=>"000100111",
  14419=>"111111000",
  14420=>"000000000",
  14421=>"001000110",
  14422=>"000100000",
  14423=>"110110111",
  14424=>"111111111",
  14425=>"111101111",
  14426=>"000000001",
  14427=>"001001001",
  14428=>"110110000",
  14429=>"000000000",
  14430=>"000010110",
  14431=>"000000000",
  14432=>"100100000",
  14433=>"011111000",
  14434=>"111111000",
  14435=>"110111111",
  14436=>"000000000",
  14437=>"000000000",
  14438=>"111000000",
  14439=>"000001001",
  14440=>"000000000",
  14441=>"000001101",
  14442=>"111111011",
  14443=>"111110100",
  14444=>"010111111",
  14445=>"111111011",
  14446=>"111111111",
  14447=>"000000000",
  14448=>"001000000",
  14449=>"111111000",
  14450=>"111111110",
  14451=>"111111111",
  14452=>"000000000",
  14453=>"000000001",
  14454=>"110110010",
  14455=>"001000000",
  14456=>"111100000",
  14457=>"000000000",
  14458=>"111100101",
  14459=>"000011001",
  14460=>"000111011",
  14461=>"110110111",
  14462=>"111111111",
  14463=>"000000000",
  14464=>"001000000",
  14465=>"000000000",
  14466=>"000010111",
  14467=>"100011011",
  14468=>"000000000",
  14469=>"000000000",
  14470=>"000000000",
  14471=>"000000000",
  14472=>"001000000",
  14473=>"100100000",
  14474=>"000000000",
  14475=>"111011000",
  14476=>"111111101",
  14477=>"111111111",
  14478=>"111111111",
  14479=>"111111111",
  14480=>"111111111",
  14481=>"000000000",
  14482=>"000001001",
  14483=>"111111111",
  14484=>"110000100",
  14485=>"000000000",
  14486=>"000000000",
  14487=>"111011011",
  14488=>"111111111",
  14489=>"111111111",
  14490=>"111111111",
  14491=>"000000000",
  14492=>"100111011",
  14493=>"001001000",
  14494=>"000000000",
  14495=>"000000110",
  14496=>"011000000",
  14497=>"111111000",
  14498=>"111111111",
  14499=>"000000000",
  14500=>"001001001",
  14501=>"000000110",
  14502=>"000100101",
  14503=>"000000100",
  14504=>"000001000",
  14505=>"011011001",
  14506=>"000000000",
  14507=>"111111110",
  14508=>"111111111",
  14509=>"000000000",
  14510=>"110111111",
  14511=>"000000000",
  14512=>"111111111",
  14513=>"000011111",
  14514=>"111111111",
  14515=>"000000000",
  14516=>"001001010",
  14517=>"011011111",
  14518=>"000001111",
  14519=>"111110000",
  14520=>"000110111",
  14521=>"001001001",
  14522=>"001000000",
  14523=>"111110101",
  14524=>"000000000",
  14525=>"000000000",
  14526=>"111111110",
  14527=>"111111111",
  14528=>"010111111",
  14529=>"000000000",
  14530=>"111111111",
  14531=>"000000100",
  14532=>"000000000",
  14533=>"111111111",
  14534=>"111111111",
  14535=>"000010111",
  14536=>"111111111",
  14537=>"111111111",
  14538=>"111100000",
  14539=>"001011111",
  14540=>"000000010",
  14541=>"000000000",
  14542=>"000000111",
  14543=>"110101100",
  14544=>"001001000",
  14545=>"000000000",
  14546=>"110111000",
  14547=>"111111111",
  14548=>"111111111",
  14549=>"000110001",
  14550=>"111011011",
  14551=>"011000000",
  14552=>"011011001",
  14553=>"000001011",
  14554=>"011111111",
  14555=>"000001001",
  14556=>"000000000",
  14557=>"000000001",
  14558=>"000000000",
  14559=>"001001000",
  14560=>"000000000",
  14561=>"000100111",
  14562=>"010010111",
  14563=>"000001000",
  14564=>"111111111",
  14565=>"110111111",
  14566=>"000000000",
  14567=>"000000000",
  14568=>"111111101",
  14569=>"000000000",
  14570=>"111111111",
  14571=>"000000000",
  14572=>"111111111",
  14573=>"000110010",
  14574=>"111001000",
  14575=>"000111000",
  14576=>"000000000",
  14577=>"000000000",
  14578=>"000111101",
  14579=>"001000100",
  14580=>"111111111",
  14581=>"011111100",
  14582=>"111101001",
  14583=>"000000000",
  14584=>"000000000",
  14585=>"111111111",
  14586=>"000110111",
  14587=>"000111111",
  14588=>"111111101",
  14589=>"111011111",
  14590=>"110000000",
  14591=>"001011111",
  14592=>"000000000",
  14593=>"110111111",
  14594=>"111001001",
  14595=>"111111111",
  14596=>"000000011",
  14597=>"011011000",
  14598=>"101000000",
  14599=>"001111111",
  14600=>"000010001",
  14601=>"000000000",
  14602=>"000000000",
  14603=>"000000011",
  14604=>"001101101",
  14605=>"011111110",
  14606=>"000111111",
  14607=>"101111101",
  14608=>"010010000",
  14609=>"111111010",
  14610=>"000000000",
  14611=>"001001000",
  14612=>"111111001",
  14613=>"000000111",
  14614=>"111100100",
  14615=>"000000000",
  14616=>"000000000",
  14617=>"000000000",
  14618=>"000000000",
  14619=>"000001111",
  14620=>"110110100",
  14621=>"111111001",
  14622=>"100000000",
  14623=>"110100111",
  14624=>"000101111",
  14625=>"111111111",
  14626=>"010000010",
  14627=>"010001011",
  14628=>"011111011",
  14629=>"000000000",
  14630=>"100111111",
  14631=>"010000010",
  14632=>"111111100",
  14633=>"111000000",
  14634=>"001111110",
  14635=>"011011000",
  14636=>"000000000",
  14637=>"100000100",
  14638=>"111000000",
  14639=>"000000111",
  14640=>"111110000",
  14641=>"110111010",
  14642=>"001000111",
  14643=>"011110111",
  14644=>"011000111",
  14645=>"000011110",
  14646=>"111111111",
  14647=>"111011111",
  14648=>"000000000",
  14649=>"010000001",
  14650=>"100100110",
  14651=>"011001000",
  14652=>"011111110",
  14653=>"111000000",
  14654=>"110110000",
  14655=>"100111001",
  14656=>"000001111",
  14657=>"111111010",
  14658=>"000000000",
  14659=>"000000000",
  14660=>"000000000",
  14661=>"000001011",
  14662=>"001000100",
  14663=>"001100111",
  14664=>"001000100",
  14665=>"111111000",
  14666=>"000010110",
  14667=>"000000000",
  14668=>"000000000",
  14669=>"111111000",
  14670=>"000000000",
  14671=>"111001011",
  14672=>"110100100",
  14673=>"000000111",
  14674=>"110111111",
  14675=>"111111111",
  14676=>"111111111",
  14677=>"011011001",
  14678=>"111111011",
  14679=>"000110010",
  14680=>"000000000",
  14681=>"111101000",
  14682=>"111111110",
  14683=>"001000001",
  14684=>"111111011",
  14685=>"000000000",
  14686=>"000000000",
  14687=>"100111111",
  14688=>"001101111",
  14689=>"011011111",
  14690=>"000000000",
  14691=>"000000000",
  14692=>"111111111",
  14693=>"000000111",
  14694=>"111111111",
  14695=>"011111111",
  14696=>"000000000",
  14697=>"111111111",
  14698=>"000000000",
  14699=>"000111110",
  14700=>"000010010",
  14701=>"101111111",
  14702=>"111111110",
  14703=>"100110000",
  14704=>"101000000",
  14705=>"000000000",
  14706=>"111111000",
  14707=>"000110111",
  14708=>"011001001",
  14709=>"111101001",
  14710=>"111111001",
  14711=>"111111111",
  14712=>"001001000",
  14713=>"000111111",
  14714=>"000000000",
  14715=>"000110101",
  14716=>"000000011",
  14717=>"111111111",
  14718=>"111111111",
  14719=>"100000000",
  14720=>"001111011",
  14721=>"111101111",
  14722=>"001001011",
  14723=>"000000000",
  14724=>"011000000",
  14725=>"110110100",
  14726=>"000011011",
  14727=>"100110000",
  14728=>"011011000",
  14729=>"111111001",
  14730=>"011001100",
  14731=>"000000001",
  14732=>"001000000",
  14733=>"111111111",
  14734=>"111111001",
  14735=>"111000001",
  14736=>"000000000",
  14737=>"111111111",
  14738=>"000000011",
  14739=>"111111011",
  14740=>"000000000",
  14741=>"000011011",
  14742=>"111111010",
  14743=>"001000000",
  14744=>"000100110",
  14745=>"000001011",
  14746=>"000000000",
  14747=>"000010001",
  14748=>"111111000",
  14749=>"111111111",
  14750=>"001000111",
  14751=>"000100000",
  14752=>"000000000",
  14753=>"110110110",
  14754=>"100110110",
  14755=>"000001111",
  14756=>"010000000",
  14757=>"000000000",
  14758=>"000100100",
  14759=>"011111111",
  14760=>"011000000",
  14761=>"100100110",
  14762=>"111111000",
  14763=>"000010011",
  14764=>"000100010",
  14765=>"111111000",
  14766=>"000000000",
  14767=>"110000000",
  14768=>"011111000",
  14769=>"111110000",
  14770=>"000101111",
  14771=>"000011111",
  14772=>"001111111",
  14773=>"111100000",
  14774=>"000000000",
  14775=>"110110000",
  14776=>"111011010",
  14777=>"000000000",
  14778=>"110111111",
  14779=>"000111111",
  14780=>"000000000",
  14781=>"111011011",
  14782=>"000000001",
  14783=>"000000000",
  14784=>"000000000",
  14785=>"111111111",
  14786=>"111111000",
  14787=>"111111110",
  14788=>"111111001",
  14789=>"111111111",
  14790=>"000000111",
  14791=>"111111111",
  14792=>"100111111",
  14793=>"001000000",
  14794=>"011000000",
  14795=>"000000000",
  14796=>"000110000",
  14797=>"111111111",
  14798=>"111111111",
  14799=>"000000100",
  14800=>"011001001",
  14801=>"111111010",
  14802=>"111011011",
  14803=>"111111111",
  14804=>"110110100",
  14805=>"000111111",
  14806=>"111011111",
  14807=>"000000000",
  14808=>"111111111",
  14809=>"000010000",
  14810=>"111111100",
  14811=>"000000100",
  14812=>"100110110",
  14813=>"111111101",
  14814=>"111011000",
  14815=>"000001101",
  14816=>"111111111",
  14817=>"001011011",
  14818=>"010010110",
  14819=>"111111111",
  14820=>"111011000",
  14821=>"111111111",
  14822=>"111011000",
  14823=>"111000000",
  14824=>"000110110",
  14825=>"000011110",
  14826=>"000000110",
  14827=>"000111111",
  14828=>"001101000",
  14829=>"000000000",
  14830=>"111111111",
  14831=>"000000000",
  14832=>"111111111",
  14833=>"110111111",
  14834=>"000000101",
  14835=>"111000100",
  14836=>"111111111",
  14837=>"110110000",
  14838=>"100000000",
  14839=>"001000000",
  14840=>"000100111",
  14841=>"111111011",
  14842=>"111111111",
  14843=>"000000000",
  14844=>"111111111",
  14845=>"110110100",
  14846=>"111111111",
  14847=>"000000000",
  14848=>"111110101",
  14849=>"000000001",
  14850=>"000000101",
  14851=>"000000011",
  14852=>"100100101",
  14853=>"111111011",
  14854=>"000000100",
  14855=>"111111111",
  14856=>"111111111",
  14857=>"110110000",
  14858=>"111111111",
  14859=>"111111110",
  14860=>"000000100",
  14861=>"001011111",
  14862=>"000111111",
  14863=>"000000000",
  14864=>"100100110",
  14865=>"111111011",
  14866=>"111111000",
  14867=>"011000000",
  14868=>"010000000",
  14869=>"000000111",
  14870=>"111111111",
  14871=>"010110110",
  14872=>"000001111",
  14873=>"110111110",
  14874=>"001001001",
  14875=>"111101101",
  14876=>"000000000",
  14877=>"100011011",
  14878=>"000100110",
  14879=>"010000110",
  14880=>"011110110",
  14881=>"000001111",
  14882=>"001000000",
  14883=>"000000100",
  14884=>"111111111",
  14885=>"000011011",
  14886=>"011000000",
  14887=>"111111111",
  14888=>"000000111",
  14889=>"000111111",
  14890=>"011111111",
  14891=>"011011111",
  14892=>"111111111",
  14893=>"011111111",
  14894=>"000000000",
  14895=>"101000000",
  14896=>"111111111",
  14897=>"100100100",
  14898=>"100111111",
  14899=>"001000110",
  14900=>"010111111",
  14901=>"100100100",
  14902=>"111000000",
  14903=>"000001001",
  14904=>"010000111",
  14905=>"111111111",
  14906=>"001001001",
  14907=>"101000000",
  14908=>"111111111",
  14909=>"111011111",
  14910=>"111111111",
  14911=>"111111111",
  14912=>"001001000",
  14913=>"111111111",
  14914=>"001000000",
  14915=>"111000111",
  14916=>"101000000",
  14917=>"111111111",
  14918=>"000000000",
  14919=>"111111111",
  14920=>"101111110",
  14921=>"111000111",
  14922=>"010010000",
  14923=>"011011100",
  14924=>"011111000",
  14925=>"100100111",
  14926=>"001000001",
  14927=>"111111111",
  14928=>"000000000",
  14929=>"011111111",
  14930=>"000000000",
  14931=>"100110000",
  14932=>"100100000",
  14933=>"011111111",
  14934=>"111111111",
  14935=>"111111111",
  14936=>"111111110",
  14937=>"000000000",
  14938=>"111000001",
  14939=>"111111001",
  14940=>"000000000",
  14941=>"011000000",
  14942=>"111111000",
  14943=>"111111011",
  14944=>"011011000",
  14945=>"100100010",
  14946=>"110111111",
  14947=>"111111111",
  14948=>"000000000",
  14949=>"000000001",
  14950=>"000010001",
  14951=>"000000000",
  14952=>"000000101",
  14953=>"111111000",
  14954=>"011011011",
  14955=>"111111111",
  14956=>"111111111",
  14957=>"111111101",
  14958=>"000000000",
  14959=>"111111000",
  14960=>"000000111",
  14961=>"010110110",
  14962=>"011111111",
  14963=>"100110110",
  14964=>"111000100",
  14965=>"111111010",
  14966=>"111111111",
  14967=>"100100000",
  14968=>"000000000",
  14969=>"100100111",
  14970=>"000000000",
  14971=>"000000000",
  14972=>"110110110",
  14973=>"001011000",
  14974=>"100000000",
  14975=>"111111111",
  14976=>"111111000",
  14977=>"111111111",
  14978=>"111111111",
  14979=>"001011011",
  14980=>"000000100",
  14981=>"111111111",
  14982=>"111111111",
  14983=>"011011111",
  14984=>"111111111",
  14985=>"111111110",
  14986=>"111111100",
  14987=>"001101111",
  14988=>"000100110",
  14989=>"111111000",
  14990=>"110111111",
  14991=>"111111111",
  14992=>"000000000",
  14993=>"111111111",
  14994=>"100000000",
  14995=>"001001111",
  14996=>"111111110",
  14997=>"110110000",
  14998=>"001000101",
  14999=>"000000000",
  15000=>"011000111",
  15001=>"100110100",
  15002=>"111111111",
  15003=>"011011000",
  15004=>"111011111",
  15005=>"000000011",
  15006=>"111111111",
  15007=>"101101101",
  15008=>"111111111",
  15009=>"001001001",
  15010=>"011011011",
  15011=>"000100000",
  15012=>"100100000",
  15013=>"100111000",
  15014=>"111111111",
  15015=>"111111111",
  15016=>"011000111",
  15017=>"000000000",
  15018=>"000000000",
  15019=>"100000011",
  15020=>"000000000",
  15021=>"001011111",
  15022=>"111000000",
  15023=>"111111111",
  15024=>"111010000",
  15025=>"111111111",
  15026=>"001001111",
  15027=>"011111111",
  15028=>"000000000",
  15029=>"110111110",
  15030=>"000000000",
  15031=>"011111111",
  15032=>"101000000",
  15033=>"000000000",
  15034=>"000000000",
  15035=>"111111111",
  15036=>"111111111",
  15037=>"000000000",
  15038=>"111111111",
  15039=>"000000000",
  15040=>"111000000",
  15041=>"111111110",
  15042=>"001001000",
  15043=>"000000011",
  15044=>"000000000",
  15045=>"000000000",
  15046=>"000000000",
  15047=>"111000110",
  15048=>"000000000",
  15049=>"001000000",
  15050=>"111101100",
  15051=>"000000000",
  15052=>"000000000",
  15053=>"111111111",
  15054=>"000001011",
  15055=>"000000000",
  15056=>"110101000",
  15057=>"000001000",
  15058=>"000000000",
  15059=>"100100100",
  15060=>"010000110",
  15061=>"000000000",
  15062=>"111111000",
  15063=>"001001000",
  15064=>"001011111",
  15065=>"110110111",
  15066=>"111111000",
  15067=>"111100000",
  15068=>"000000000",
  15069=>"101101001",
  15070=>"000000000",
  15071=>"100101101",
  15072=>"011001011",
  15073=>"000000011",
  15074=>"111111111",
  15075=>"111111110",
  15076=>"000010000",
  15077=>"100100000",
  15078=>"011111111",
  15079=>"110110100",
  15080=>"111111111",
  15081=>"000010000",
  15082=>"111011000",
  15083=>"111111011",
  15084=>"010011011",
  15085=>"111111111",
  15086=>"001110100",
  15087=>"011000000",
  15088=>"000000000",
  15089=>"000000101",
  15090=>"111111111",
  15091=>"010010111",
  15092=>"001000000",
  15093=>"111111111",
  15094=>"011111111",
  15095=>"111111111",
  15096=>"001000100",
  15097=>"111111111",
  15098=>"110000011",
  15099=>"001000000",
  15100=>"100000010",
  15101=>"011011011",
  15102=>"110000011",
  15103=>"110010000",
  15104=>"010100000",
  15105=>"001001011",
  15106=>"000000000",
  15107=>"000001111",
  15108=>"101100101",
  15109=>"011011000",
  15110=>"110110100",
  15111=>"001000000",
  15112=>"000000000",
  15113=>"000001001",
  15114=>"111111111",
  15115=>"010000000",
  15116=>"111111111",
  15117=>"111011000",
  15118=>"111101111",
  15119=>"001111000",
  15120=>"110100000",
  15121=>"011111111",
  15122=>"111111000",
  15123=>"000111011",
  15124=>"111111100",
  15125=>"000011111",
  15126=>"110010000",
  15127=>"011111111",
  15128=>"111111110",
  15129=>"111111000",
  15130=>"111001111",
  15131=>"111001000",
  15132=>"011111111",
  15133=>"001001001",
  15134=>"011111011",
  15135=>"110001111",
  15136=>"001011000",
  15137=>"000000000",
  15138=>"100000000",
  15139=>"111111111",
  15140=>"000111111",
  15141=>"111000100",
  15142=>"000000000",
  15143=>"111111100",
  15144=>"100111111",
  15145=>"111111111",
  15146=>"100011111",
  15147=>"001000000",
  15148=>"100100011",
  15149=>"101101101",
  15150=>"111111111",
  15151=>"000000000",
  15152=>"000000110",
  15153=>"111111111",
  15154=>"111111111",
  15155=>"000110110",
  15156=>"000001001",
  15157=>"111011011",
  15158=>"000001001",
  15159=>"000000011",
  15160=>"000000000",
  15161=>"001000100",
  15162=>"110100100",
  15163=>"111101111",
  15164=>"111111110",
  15165=>"001111010",
  15166=>"000000110",
  15167=>"111110100",
  15168=>"100100000",
  15169=>"111011000",
  15170=>"110100100",
  15171=>"111111111",
  15172=>"000000000",
  15173=>"001011000",
  15174=>"000000000",
  15175=>"101001001",
  15176=>"000000000",
  15177=>"000111111",
  15178=>"000011011",
  15179=>"111100000",
  15180=>"011111000",
  15181=>"111110000",
  15182=>"000000000",
  15183=>"000000100",
  15184=>"110110100",
  15185=>"010000110",
  15186=>"010110000",
  15187=>"100111000",
  15188=>"110111110",
  15189=>"011111111",
  15190=>"001011111",
  15191=>"000000000",
  15192=>"111111111",
  15193=>"001000000",
  15194=>"011100000",
  15195=>"000000000",
  15196=>"111111100",
  15197=>"000010111",
  15198=>"000000011",
  15199=>"011011001",
  15200=>"000000000",
  15201=>"111000000",
  15202=>"000000011",
  15203=>"000000000",
  15204=>"000000000",
  15205=>"000000000",
  15206=>"000100111",
  15207=>"011111111",
  15208=>"000011001",
  15209=>"111111111",
  15210=>"010111000",
  15211=>"111111111",
  15212=>"100000001",
  15213=>"000000000",
  15214=>"000000001",
  15215=>"000000000",
  15216=>"001000000",
  15217=>"111111111",
  15218=>"110100000",
  15219=>"111111111",
  15220=>"111101101",
  15221=>"111111111",
  15222=>"011001000",
  15223=>"001011111",
  15224=>"000000000",
  15225=>"111111111",
  15226=>"111111111",
  15227=>"001000110",
  15228=>"100100100",
  15229=>"000111111",
  15230=>"111111000",
  15231=>"111111111",
  15232=>"000011110",
  15233=>"000000000",
  15234=>"111111111",
  15235=>"000000000",
  15236=>"001111101",
  15237=>"000000000",
  15238=>"111011011",
  15239=>"000010000",
  15240=>"000000000",
  15241=>"100100110",
  15242=>"000000000",
  15243=>"111000001",
  15244=>"111111111",
  15245=>"000101101",
  15246=>"111111000",
  15247=>"000000000",
  15248=>"011111111",
  15249=>"001111111",
  15250=>"111111111",
  15251=>"111111111",
  15252=>"111000000",
  15253=>"000000000",
  15254=>"100100000",
  15255=>"100100110",
  15256=>"111111111",
  15257=>"000100100",
  15258=>"000000000",
  15259=>"000111111",
  15260=>"100000100",
  15261=>"001001011",
  15262=>"000000000",
  15263=>"000000000",
  15264=>"111001111",
  15265=>"001001000",
  15266=>"111100100",
  15267=>"111110111",
  15268=>"011011111",
  15269=>"111111111",
  15270=>"000000000",
  15271=>"111111011",
  15272=>"100111001",
  15273=>"000001001",
  15274=>"111111110",
  15275=>"010011010",
  15276=>"000111001",
  15277=>"111111111",
  15278=>"000000001",
  15279=>"100100100",
  15280=>"000000011",
  15281=>"000111111",
  15282=>"011011001",
  15283=>"111111111",
  15284=>"000000000",
  15285=>"111000001",
  15286=>"000000000",
  15287=>"111000000",
  15288=>"111111110",
  15289=>"111111110",
  15290=>"111111111",
  15291=>"000000011",
  15292=>"011001000",
  15293=>"000000000",
  15294=>"000000000",
  15295=>"001001001",
  15296=>"000110011",
  15297=>"010010010",
  15298=>"000000011",
  15299=>"000000000",
  15300=>"011101000",
  15301=>"010110100",
  15302=>"011001001",
  15303=>"000000000",
  15304=>"010000000",
  15305=>"000000100",
  15306=>"000000011",
  15307=>"000001111",
  15308=>"011010111",
  15309=>"000000001",
  15310=>"111111111",
  15311=>"100000010",
  15312=>"000010010",
  15313=>"001001001",
  15314=>"000111111",
  15315=>"000000000",
  15316=>"110111111",
  15317=>"100000011",
  15318=>"000000111",
  15319=>"000000110",
  15320=>"001000000",
  15321=>"111111111",
  15322=>"111111110",
  15323=>"111111111",
  15324=>"111111111",
  15325=>"000001101",
  15326=>"000000111",
  15327=>"000101001",
  15328=>"000000011",
  15329=>"001001101",
  15330=>"000000000",
  15331=>"000000001",
  15332=>"111111000",
  15333=>"000000000",
  15334=>"000000110",
  15335=>"111101111",
  15336=>"011011011",
  15337=>"111111111",
  15338=>"001000000",
  15339=>"000111001",
  15340=>"111011000",
  15341=>"101100110",
  15342=>"000000000",
  15343=>"111001011",
  15344=>"000000000",
  15345=>"000011111",
  15346=>"111111001",
  15347=>"000000001",
  15348=>"010010010",
  15349=>"111111111",
  15350=>"111011000",
  15351=>"000110100",
  15352=>"000000000",
  15353=>"011001000",
  15354=>"111110000",
  15355=>"111011000",
  15356=>"011111001",
  15357=>"110011011",
  15358=>"110000010",
  15359=>"000000000",
  15360=>"101000100",
  15361=>"000011000",
  15362=>"110110000",
  15363=>"111001000",
  15364=>"100111111",
  15365=>"000001011",
  15366=>"000000000",
  15367=>"000010111",
  15368=>"011101000",
  15369=>"111111011",
  15370=>"111111110",
  15371=>"111111111",
  15372=>"000010000",
  15373=>"100000111",
  15374=>"000000000",
  15375=>"111111111",
  15376=>"110111111",
  15377=>"110111000",
  15378=>"101000000",
  15379=>"001111101",
  15380=>"111111000",
  15381=>"000000111",
  15382=>"111110111",
  15383=>"111111001",
  15384=>"010110000",
  15385=>"101111111",
  15386=>"110000000",
  15387=>"110110010",
  15388=>"000000000",
  15389=>"001000111",
  15390=>"101100000",
  15391=>"000001011",
  15392=>"000000000",
  15393=>"000000000",
  15394=>"111011001",
  15395=>"111111011",
  15396=>"111111111",
  15397=>"111111001",
  15398=>"111111111",
  15399=>"111111101",
  15400=>"111111000",
  15401=>"000000111",
  15402=>"100000000",
  15403=>"000000000",
  15404=>"100000000",
  15405=>"111111111",
  15406=>"001011011",
  15407=>"111111111",
  15408=>"000000000",
  15409=>"100000000",
  15410=>"111111111",
  15411=>"111111000",
  15412=>"011001011",
  15413=>"001000001",
  15414=>"111111011",
  15415=>"000000101",
  15416=>"110111110",
  15417=>"100100100",
  15418=>"111101111",
  15419=>"010000000",
  15420=>"011010111",
  15421=>"001001001",
  15422=>"100001000",
  15423=>"111111011",
  15424=>"111011111",
  15425=>"011011111",
  15426=>"000000000",
  15427=>"000111000",
  15428=>"111111000",
  15429=>"111111111",
  15430=>"100111111",
  15431=>"111111111",
  15432=>"011111111",
  15433=>"000000111",
  15434=>"000011000",
  15435=>"111111000",
  15436=>"001011000",
  15437=>"111111001",
  15438=>"111111100",
  15439=>"001111100",
  15440=>"101101110",
  15441=>"001111111",
  15442=>"000010000",
  15443=>"111001001",
  15444=>"101101111",
  15445=>"110100111",
  15446=>"000110000",
  15447=>"111111111",
  15448=>"111111100",
  15449=>"000000000",
  15450=>"011011010",
  15451=>"000110000",
  15452=>"000100000",
  15453=>"111010000",
  15454=>"000000011",
  15455=>"011111111",
  15456=>"011000000",
  15457=>"111111000",
  15458=>"000000010",
  15459=>"000010000",
  15460=>"111111011",
  15461=>"000011000",
  15462=>"100110110",
  15463=>"111000111",
  15464=>"111000110",
  15465=>"000000000",
  15466=>"000000111",
  15467=>"111000110",
  15468=>"000110110",
  15469=>"000000000",
  15470=>"000000010",
  15471=>"100110001",
  15472=>"000111110",
  15473=>"000010000",
  15474=>"001101101",
  15475=>"111100000",
  15476=>"100110111",
  15477=>"000111111",
  15478=>"010110111",
  15479=>"000000000",
  15480=>"010000100",
  15481=>"111100000",
  15482=>"100100100",
  15483=>"110100100",
  15484=>"001001010",
  15485=>"111111111",
  15486=>"111110111",
  15487=>"001001001",
  15488=>"111111110",
  15489=>"000111111",
  15490=>"111110000",
  15491=>"101000000",
  15492=>"110000000",
  15493=>"111111000",
  15494=>"000001111",
  15495=>"000000000",
  15496=>"000000000",
  15497=>"001001101",
  15498=>"000000000",
  15499=>"000100100",
  15500=>"000000000",
  15501=>"011001001",
  15502=>"011111000",
  15503=>"111111000",
  15504=>"000000001",
  15505=>"111111111",
  15506=>"000000110",
  15507=>"000000000",
  15508=>"111111000",
  15509=>"110000110",
  15510=>"110111110",
  15511=>"111111011",
  15512=>"011111101",
  15513=>"111011111",
  15514=>"100000110",
  15515=>"000000000",
  15516=>"111111011",
  15517=>"001011111",
  15518=>"001100110",
  15519=>"000000000",
  15520=>"110111111",
  15521=>"001010000",
  15522=>"000000000",
  15523=>"001000000",
  15524=>"000101100",
  15525=>"000010011",
  15526=>"000000000",
  15527=>"111001011",
  15528=>"000000000",
  15529=>"111110100",
  15530=>"111111111",
  15531=>"001000110",
  15532=>"100000111",
  15533=>"000000000",
  15534=>"001111111",
  15535=>"111011000",
  15536=>"000000000",
  15537=>"111111100",
  15538=>"000000000",
  15539=>"000000000",
  15540=>"111111111",
  15541=>"000000000",
  15542=>"101000000",
  15543=>"111111000",
  15544=>"011011000",
  15545=>"000000011",
  15546=>"100000101",
  15547=>"000000000",
  15548=>"110111000",
  15549=>"111110100",
  15550=>"110111010",
  15551=>"100110000",
  15552=>"111000000",
  15553=>"000000110",
  15554=>"000000000",
  15555=>"000000000",
  15556=>"001100111",
  15557=>"111111110",
  15558=>"000000000",
  15559=>"100100111",
  15560=>"010000100",
  15561=>"000000100",
  15562=>"101000000",
  15563=>"111111111",
  15564=>"011111110",
  15565=>"111001111",
  15566=>"010111000",
  15567=>"000000000",
  15568=>"000110111",
  15569=>"100111000",
  15570=>"000000000",
  15571=>"111111101",
  15572=>"000000011",
  15573=>"001111010",
  15574=>"010010000",
  15575=>"111111110",
  15576=>"000110100",
  15577=>"010000001",
  15578=>"100000111",
  15579=>"000000000",
  15580=>"000100110",
  15581=>"000111000",
  15582=>"011000000",
  15583=>"100100101",
  15584=>"001010001",
  15585=>"010111111",
  15586=>"000110111",
  15587=>"001000000",
  15588=>"111111111",
  15589=>"001001001",
  15590=>"011010000",
  15591=>"111111011",
  15592=>"000111111",
  15593=>"111001001",
  15594=>"111111011",
  15595=>"100000111",
  15596=>"111111111",
  15597=>"000000000",
  15598=>"000000110",
  15599=>"000000000",
  15600=>"111101001",
  15601=>"000000001",
  15602=>"111111111",
  15603=>"101100000",
  15604=>"110111000",
  15605=>"111000000",
  15606=>"000000101",
  15607=>"110111000",
  15608=>"100000000",
  15609=>"000000000",
  15610=>"000000001",
  15611=>"011111111",
  15612=>"000000111",
  15613=>"110010110",
  15614=>"001111110",
  15615=>"111011001",
  15616=>"011011000",
  15617=>"011111110",
  15618=>"100000000",
  15619=>"110111111",
  15620=>"011111110",
  15621=>"111111000",
  15622=>"010111011",
  15623=>"000000000",
  15624=>"000111001",
  15625=>"111101000",
  15626=>"111100001",
  15627=>"010101101",
  15628=>"000000000",
  15629=>"000000000",
  15630=>"100100011",
  15631=>"111111111",
  15632=>"111111000",
  15633=>"010111000",
  15634=>"110000111",
  15635=>"000001000",
  15636=>"111001000",
  15637=>"111111010",
  15638=>"000000000",
  15639=>"100101001",
  15640=>"111111111",
  15641=>"000000011",
  15642=>"000000101",
  15643=>"010111111",
  15644=>"111011001",
  15645=>"111111011",
  15646=>"110100000",
  15647=>"111111010",
  15648=>"111111011",
  15649=>"011111110",
  15650=>"110000011",
  15651=>"111111101",
  15652=>"000111000",
  15653=>"000000000",
  15654=>"111110110",
  15655=>"111011001",
  15656=>"101100000",
  15657=>"000000100",
  15658=>"001110110",
  15659=>"000001000",
  15660=>"111111111",
  15661=>"111111111",
  15662=>"000000000",
  15663=>"000000111",
  15664=>"001111001",
  15665=>"111000111",
  15666=>"011111111",
  15667=>"000000000",
  15668=>"000000000",
  15669=>"001001000",
  15670=>"001110111",
  15671=>"000100000",
  15672=>"000000111",
  15673=>"010010110",
  15674=>"000000100",
  15675=>"111001001",
  15676=>"000011111",
  15677=>"011111111",
  15678=>"111111001",
  15679=>"000000100",
  15680=>"000000000",
  15681=>"000000100",
  15682=>"010100000",
  15683=>"000000111",
  15684=>"011001011",
  15685=>"000000000",
  15686=>"100110111",
  15687=>"111110111",
  15688=>"000000111",
  15689=>"000110000",
  15690=>"111000000",
  15691=>"110110111",
  15692=>"101000100",
  15693=>"111111111",
  15694=>"000100000",
  15695=>"111111111",
  15696=>"101101111",
  15697=>"000000000",
  15698=>"001000000",
  15699=>"111111000",
  15700=>"011111111",
  15701=>"111101111",
  15702=>"011111100",
  15703=>"111101111",
  15704=>"000000100",
  15705=>"000000000",
  15706=>"011111011",
  15707=>"101101111",
  15708=>"010011000",
  15709=>"111111111",
  15710=>"000011000",
  15711=>"111100111",
  15712=>"111011000",
  15713=>"111100101",
  15714=>"011111111",
  15715=>"000010011",
  15716=>"001000001",
  15717=>"111111000",
  15718=>"111111000",
  15719=>"000001001",
  15720=>"001001011",
  15721=>"000011000",
  15722=>"000000100",
  15723=>"000001001",
  15724=>"111110111",
  15725=>"000000000",
  15726=>"111111000",
  15727=>"001011000",
  15728=>"011111011",
  15729=>"000011000",
  15730=>"111111000",
  15731=>"001000001",
  15732=>"000000000",
  15733=>"110010010",
  15734=>"000010000",
  15735=>"011101111",
  15736=>"000000110",
  15737=>"010110000",
  15738=>"111111000",
  15739=>"100111111",
  15740=>"001111001",
  15741=>"111111110",
  15742=>"110110000",
  15743=>"101000000",
  15744=>"110000000",
  15745=>"110100100",
  15746=>"111100100",
  15747=>"100100100",
  15748=>"111111001",
  15749=>"000000111",
  15750=>"111111110",
  15751=>"000000000",
  15752=>"010000000",
  15753=>"111111111",
  15754=>"000110111",
  15755=>"000000000",
  15756=>"000000000",
  15757=>"110111010",
  15758=>"001111011",
  15759=>"111111111",
  15760=>"110100111",
  15761=>"000000111",
  15762=>"111011001",
  15763=>"111111001",
  15764=>"111000111",
  15765=>"111111111",
  15766=>"111111111",
  15767=>"000001000",
  15768=>"011111011",
  15769=>"000100100",
  15770=>"111111001",
  15771=>"000000010",
  15772=>"000000110",
  15773=>"000111000",
  15774=>"111110111",
  15775=>"000000000",
  15776=>"111101000",
  15777=>"111101110",
  15778=>"001011000",
  15779=>"111111111",
  15780=>"000000100",
  15781=>"011001011",
  15782=>"110000000",
  15783=>"111111001",
  15784=>"111111110",
  15785=>"110110111",
  15786=>"000110000",
  15787=>"010110111",
  15788=>"110111111",
  15789=>"000010100",
  15790=>"111111111",
  15791=>"100000001",
  15792=>"000000000",
  15793=>"010000000",
  15794=>"000000001",
  15795=>"110100000",
  15796=>"000000000",
  15797=>"001000101",
  15798=>"000010000",
  15799=>"111110110",
  15800=>"000000000",
  15801=>"100111010",
  15802=>"001101111",
  15803=>"010111111",
  15804=>"011011111",
  15805=>"111111011",
  15806=>"011000011",
  15807=>"000010000",
  15808=>"111110111",
  15809=>"010110100",
  15810=>"000110111",
  15811=>"000000000",
  15812=>"000010111",
  15813=>"100111011",
  15814=>"111111111",
  15815=>"001111011",
  15816=>"000000000",
  15817=>"100100110",
  15818=>"011011001",
  15819=>"000000111",
  15820=>"001001000",
  15821=>"011111111",
  15822=>"100110011",
  15823=>"111100110",
  15824=>"111111001",
  15825=>"000100000",
  15826=>"110111111",
  15827=>"110111000",
  15828=>"000110011",
  15829=>"110100110",
  15830=>"000100110",
  15831=>"111111111",
  15832=>"001011011",
  15833=>"101101111",
  15834=>"001111000",
  15835=>"001000111",
  15836=>"101011111",
  15837=>"000000000",
  15838=>"110111000",
  15839=>"000001101",
  15840=>"110000111",
  15841=>"000000110",
  15842=>"111111000",
  15843=>"111000000",
  15844=>"100100110",
  15845=>"111111000",
  15846=>"011110011",
  15847=>"101111000",
  15848=>"101111111",
  15849=>"111111101",
  15850=>"010111011",
  15851=>"111101111",
  15852=>"000000000",
  15853=>"111111111",
  15854=>"001111111",
  15855=>"111110100",
  15856=>"100110111",
  15857=>"000111101",
  15858=>"000011000",
  15859=>"010111111",
  15860=>"100101001",
  15861=>"111011111",
  15862=>"111111111",
  15863=>"111111000",
  15864=>"000000000",
  15865=>"111111101",
  15866=>"000010110",
  15867=>"000000111",
  15868=>"010000110",
  15869=>"001100100",
  15870=>"110111111",
  15871=>"000001111",
  15872=>"011111111",
  15873=>"111011111",
  15874=>"000001111",
  15875=>"000000000",
  15876=>"100100000",
  15877=>"000000001",
  15878=>"001001111",
  15879=>"111111111",
  15880=>"000000111",
  15881=>"000000000",
  15882=>"111111111",
  15883=>"000000000",
  15884=>"000100111",
  15885=>"000000000",
  15886=>"000000001",
  15887=>"000000101",
  15888=>"100100111",
  15889=>"000001111",
  15890=>"000000001",
  15891=>"000000000",
  15892=>"011111001",
  15893=>"000000000",
  15894=>"000000000",
  15895=>"000011111",
  15896=>"111111111",
  15897=>"111110000",
  15898=>"001001111",
  15899=>"000101100",
  15900=>"000000001",
  15901=>"111111111",
  15902=>"101111000",
  15903=>"001000000",
  15904=>"001111111",
  15905=>"000000100",
  15906=>"111111000",
  15907=>"001001001",
  15908=>"000000111",
  15909=>"000000101",
  15910=>"000000001",
  15911=>"100000000",
  15912=>"000011001",
  15913=>"111000000",
  15914=>"000000111",
  15915=>"000011111",
  15916=>"000000000",
  15917=>"100101000",
  15918=>"000000000",
  15919=>"111011111",
  15920=>"110100101",
  15921=>"000000000",
  15922=>"011100000",
  15923=>"000000000",
  15924=>"100100111",
  15925=>"011000000",
  15926=>"000000111",
  15927=>"111011011",
  15928=>"111111011",
  15929=>"001000100",
  15930=>"011011000",
  15931=>"000000000",
  15932=>"100000000",
  15933=>"101001001",
  15934=>"000000111",
  15935=>"010011010",
  15936=>"001001001",
  15937=>"000000000",
  15938=>"000000111",
  15939=>"000000111",
  15940=>"000110111",
  15941=>"000001000",
  15942=>"011000111",
  15943=>"111100100",
  15944=>"111111001",
  15945=>"111000001",
  15946=>"000000000",
  15947=>"000000000",
  15948=>"111111010",
  15949=>"001001001",
  15950=>"000111111",
  15951=>"000000000",
  15952=>"011001000",
  15953=>"100000000",
  15954=>"000000001",
  15955=>"001000000",
  15956=>"000100110",
  15957=>"111111111",
  15958=>"000000101",
  15959=>"001111101",
  15960=>"000000000",
  15961=>"000000000",
  15962=>"111111111",
  15963=>"100100001",
  15964=>"001000000",
  15965=>"110000000",
  15966=>"000011111",
  15967=>"000001000",
  15968=>"000111111",
  15969=>"111111011",
  15970=>"111111001",
  15971=>"111000111",
  15972=>"001001000",
  15973=>"000100111",
  15974=>"100000111",
  15975=>"000000000",
  15976=>"001000000",
  15977=>"111111000",
  15978=>"000000010",
  15979=>"000111111",
  15980=>"000000000",
  15981=>"111111000",
  15982=>"000001001",
  15983=>"111111111",
  15984=>"100000000",
  15985=>"000000000",
  15986=>"110000000",
  15987=>"111111111",
  15988=>"111111111",
  15989=>"000111111",
  15990=>"111111000",
  15991=>"111001100",
  15992=>"111111110",
  15993=>"001000001",
  15994=>"001001100",
  15995=>"001001011",
  15996=>"000000101",
  15997=>"111111010",
  15998=>"000000000",
  15999=>"000000000",
  16000=>"001000000",
  16001=>"111111000",
  16002=>"001000000",
  16003=>"110000000",
  16004=>"000000101",
  16005=>"111000000",
  16006=>"000000111",
  16007=>"000001001",
  16008=>"001111111",
  16009=>"000000000",
  16010=>"101111011",
  16011=>"111111111",
  16012=>"111110100",
  16013=>"010011000",
  16014=>"111111111",
  16015=>"000000000",
  16016=>"011110000",
  16017=>"000000000",
  16018=>"110010001",
  16019=>"100000001",
  16020=>"000000101",
  16021=>"111000000",
  16022=>"000000001",
  16023=>"110110000",
  16024=>"111010111",
  16025=>"001100100",
  16026=>"000000000",
  16027=>"011000000",
  16028=>"111011111",
  16029=>"001000100",
  16030=>"111111111",
  16031=>"101111111",
  16032=>"011111111",
  16033=>"110111111",
  16034=>"111111010",
  16035=>"111111110",
  16036=>"011001001",
  16037=>"111110010",
  16038=>"000000111",
  16039=>"110111111",
  16040=>"000000001",
  16041=>"001000111",
  16042=>"011001011",
  16043=>"111111000",
  16044=>"111110010",
  16045=>"111111100",
  16046=>"100100111",
  16047=>"000000100",
  16048=>"111000000",
  16049=>"111111111",
  16050=>"111111111",
  16051=>"010000111",
  16052=>"011011000",
  16053=>"111100111",
  16054=>"011111110",
  16055=>"111111111",
  16056=>"111111111",
  16057=>"001001111",
  16058=>"000111011",
  16059=>"100100110",
  16060=>"000000101",
  16061=>"000000001",
  16062=>"000000111",
  16063=>"111100000",
  16064=>"000100111",
  16065=>"000000000",
  16066=>"000000000",
  16067=>"101101111",
  16068=>"000000000",
  16069=>"000000101",
  16070=>"111001001",
  16071=>"001000001",
  16072=>"111111100",
  16073=>"111101001",
  16074=>"000000001",
  16075=>"000000000",
  16076=>"000000111",
  16077=>"111111111",
  16078=>"000000000",
  16079=>"101101000",
  16080=>"101000000",
  16081=>"011011000",
  16082=>"111101000",
  16083=>"000000000",
  16084=>"111111110",
  16085=>"001111111",
  16086=>"000000000",
  16087=>"000000111",
  16088=>"111100000",
  16089=>"111111011",
  16090=>"111111111",
  16091=>"100000110",
  16092=>"001000001",
  16093=>"001011010",
  16094=>"111111000",
  16095=>"111001001",
  16096=>"000000000",
  16097=>"111011011",
  16098=>"111110000",
  16099=>"111111011",
  16100=>"111111101",
  16101=>"000001001",
  16102=>"111111111",
  16103=>"110011111",
  16104=>"000000111",
  16105=>"000000111",
  16106=>"000000111",
  16107=>"000000000",
  16108=>"111111111",
  16109=>"000000111",
  16110=>"111010000",
  16111=>"000101111",
  16112=>"001000000",
  16113=>"111111001",
  16114=>"000000000",
  16115=>"100000000",
  16116=>"000000001",
  16117=>"101101001",
  16118=>"001100100",
  16119=>"000000000",
  16120=>"000000101",
  16121=>"111000100",
  16122=>"000000001",
  16123=>"101000000",
  16124=>"000000100",
  16125=>"011111111",
  16126=>"011011000",
  16127=>"010111111",
  16128=>"000000111",
  16129=>"100001001",
  16130=>"111111111",
  16131=>"111111010",
  16132=>"011111001",
  16133=>"001111110",
  16134=>"111111000",
  16135=>"000000000",
  16136=>"100000000",
  16137=>"000000000",
  16138=>"001001000",
  16139=>"000100101",
  16140=>"101001111",
  16141=>"111111111",
  16142=>"111111100",
  16143=>"110110000",
  16144=>"111111101",
  16145=>"000000000",
  16146=>"111011011",
  16147=>"011111111",
  16148=>"011001110",
  16149=>"000000000",
  16150=>"001001011",
  16151=>"100100101",
  16152=>"110100100",
  16153=>"111011000",
  16154=>"000000000",
  16155=>"111101001",
  16156=>"110110100",
  16157=>"001001111",
  16158=>"011111111",
  16159=>"000000000",
  16160=>"110111001",
  16161=>"011111100",
  16162=>"111011111",
  16163=>"000000101",
  16164=>"011011011",
  16165=>"000000001",
  16166=>"100000000",
  16167=>"001111111",
  16168=>"011111111",
  16169=>"000000000",
  16170=>"111111001",
  16171=>"111000000",
  16172=>"101011111",
  16173=>"100000000",
  16174=>"001000000",
  16175=>"111001101",
  16176=>"001001111",
  16177=>"111111111",
  16178=>"000000000",
  16179=>"111111100",
  16180=>"000000000",
  16181=>"001000100",
  16182=>"111100100",
  16183=>"111000100",
  16184=>"111001000",
  16185=>"000000001",
  16186=>"111111111",
  16187=>"111000000",
  16188=>"100000000",
  16189=>"000110110",
  16190=>"000000000",
  16191=>"101110110",
  16192=>"000000000",
  16193=>"101111011",
  16194=>"100011111",
  16195=>"111111110",
  16196=>"000000100",
  16197=>"010000000",
  16198=>"000000000",
  16199=>"100101111",
  16200=>"000000001",
  16201=>"001001000",
  16202=>"101000000",
  16203=>"000000100",
  16204=>"011001001",
  16205=>"011001011",
  16206=>"000000001",
  16207=>"111000000",
  16208=>"000000000",
  16209=>"111111100",
  16210=>"111100000",
  16211=>"100000001",
  16212=>"101000000",
  16213=>"000010011",
  16214=>"000101111",
  16215=>"000000001",
  16216=>"001001001",
  16217=>"111110010",
  16218=>"110000100",
  16219=>"111111000",
  16220=>"111111111",
  16221=>"110111011",
  16222=>"000100100",
  16223=>"000000000",
  16224=>"111111111",
  16225=>"000000110",
  16226=>"111110100",
  16227=>"000000000",
  16228=>"110110111",
  16229=>"111001001",
  16230=>"100000000",
  16231=>"010000101",
  16232=>"100000100",
  16233=>"110100100",
  16234=>"100100000",
  16235=>"000000000",
  16236=>"000000001",
  16237=>"000110001",
  16238=>"000011111",
  16239=>"111100001",
  16240=>"101111011",
  16241=>"000000111",
  16242=>"111011001",
  16243=>"110110000",
  16244=>"001001011",
  16245=>"001111111",
  16246=>"011000000",
  16247=>"111111111",
  16248=>"000000011",
  16249=>"000111000",
  16250=>"000000000",
  16251=>"001000111",
  16252=>"000001000",
  16253=>"111111111",
  16254=>"100000000",
  16255=>"000000001",
  16256=>"110110010",
  16257=>"011100100",
  16258=>"011011001",
  16259=>"000000000",
  16260=>"000000000",
  16261=>"000100100",
  16262=>"000100000",
  16263=>"000000000",
  16264=>"000000011",
  16265=>"111111101",
  16266=>"110110111",
  16267=>"000000111",
  16268=>"111111100",
  16269=>"101111111",
  16270=>"000101101",
  16271=>"000000011",
  16272=>"101111111",
  16273=>"111111000",
  16274=>"000000001",
  16275=>"011011011",
  16276=>"111111001",
  16277=>"000011011",
  16278=>"111001111",
  16279=>"011001000",
  16280=>"100000011",
  16281=>"111001000",
  16282=>"001000111",
  16283=>"000000000",
  16284=>"100100101",
  16285=>"000000000",
  16286=>"100100111",
  16287=>"101111000",
  16288=>"011111111",
  16289=>"111111110",
  16290=>"111111111",
  16291=>"011111011",
  16292=>"000011111",
  16293=>"100101111",
  16294=>"001000110",
  16295=>"111111111",
  16296=>"001001000",
  16297=>"111101101",
  16298=>"111110111",
  16299=>"000000000",
  16300=>"000000111",
  16301=>"111111011",
  16302=>"011000100",
  16303=>"001111000",
  16304=>"111111111",
  16305=>"000000000",
  16306=>"111111111",
  16307=>"111011001",
  16308=>"001111100",
  16309=>"001101101",
  16310=>"011111101",
  16311=>"000000000",
  16312=>"101111010",
  16313=>"111111111",
  16314=>"011000000",
  16315=>"000000000",
  16316=>"000000011",
  16317=>"111011011",
  16318=>"101001111",
  16319=>"101101111",
  16320=>"111111111",
  16321=>"001000000",
  16322=>"001101111",
  16323=>"111111011",
  16324=>"110111111",
  16325=>"111110111",
  16326=>"100000001",
  16327=>"111111111",
  16328=>"101100111",
  16329=>"000000000",
  16330=>"000000001",
  16331=>"000000000",
  16332=>"100000000",
  16333=>"000000000",
  16334=>"111111000",
  16335=>"011000100",
  16336=>"000111110",
  16337=>"011111100",
  16338=>"000001000",
  16339=>"000000000",
  16340=>"001000000",
  16341=>"111111111",
  16342=>"000000001",
  16343=>"100000000",
  16344=>"000000000",
  16345=>"000000000",
  16346=>"000000000",
  16347=>"011011111",
  16348=>"000000001",
  16349=>"101111111",
  16350=>"111111000",
  16351=>"110111111",
  16352=>"110110111",
  16353=>"110000000",
  16354=>"000001111",
  16355=>"001001011",
  16356=>"111111000",
  16357=>"011011000",
  16358=>"111011000",
  16359=>"011111001",
  16360=>"000000000",
  16361=>"011000000",
  16362=>"000000000",
  16363=>"000000000",
  16364=>"000000100",
  16365=>"100100001",
  16366=>"000000000",
  16367=>"111111000",
  16368=>"000100111",
  16369=>"011101000",
  16370=>"000111000",
  16371=>"100001000",
  16372=>"001001000",
  16373=>"111110111",
  16374=>"101101101",
  16375=>"010000000",
  16376=>"000000100",
  16377=>"001000100",
  16378=>"111111111",
  16379=>"111111111",
  16380=>"100101000",
  16381=>"111110000",
  16382=>"111001000",
  16383=>"111111001",
  16384=>"110110110",
  16385=>"000011000",
  16386=>"111000000",
  16387=>"000010010",
  16388=>"000110111",
  16389=>"000000000",
  16390=>"110110111",
  16391=>"001001001",
  16392=>"111111111",
  16393=>"000010111",
  16394=>"111111111",
  16395=>"100000100",
  16396=>"100110111",
  16397=>"011111111",
  16398=>"000001111",
  16399=>"011011111",
  16400=>"100100101",
  16401=>"111111111",
  16402=>"000000000",
  16403=>"110111111",
  16404=>"011001000",
  16405=>"000111111",
  16406=>"111100000",
  16407=>"110100100",
  16408=>"000000000",
  16409=>"000000011",
  16410=>"111101001",
  16411=>"010010000",
  16412=>"000000000",
  16413=>"111011011",
  16414=>"011011011",
  16415=>"000000100",
  16416=>"000010111",
  16417=>"111111001",
  16418=>"000000000",
  16419=>"110111111",
  16420=>"011111111",
  16421=>"010000000",
  16422=>"110100000",
  16423=>"000000111",
  16424=>"111001000",
  16425=>"001001011",
  16426=>"011101000",
  16427=>"000000100",
  16428=>"101111111",
  16429=>"110110000",
  16430=>"000111111",
  16431=>"111110100",
  16432=>"001000000",
  16433=>"000000110",
  16434=>"000000000",
  16435=>"111000000",
  16436=>"010110111",
  16437=>"111111110",
  16438=>"111001001",
  16439=>"000011011",
  16440=>"000000111",
  16441=>"011101000",
  16442=>"000000000",
  16443=>"111111111",
  16444=>"000000000",
  16445=>"111000000",
  16446=>"000000000",
  16447=>"001001000",
  16448=>"000011001",
  16449=>"000000001",
  16450=>"100111111",
  16451=>"110100111",
  16452=>"000111100",
  16453=>"001000101",
  16454=>"001001100",
  16455=>"111111111",
  16456=>"000011011",
  16457=>"000000000",
  16458=>"000000000",
  16459=>"111101111",
  16460=>"100100110",
  16461=>"001000101",
  16462=>"011000000",
  16463=>"111111111",
  16464=>"111111111",
  16465=>"111111111",
  16466=>"000000010",
  16467=>"111111110",
  16468=>"000000000",
  16469=>"000000111",
  16470=>"001100111",
  16471=>"000000111",
  16472=>"000000000",
  16473=>"000000000",
  16474=>"111111111",
  16475=>"100000100",
  16476=>"000000000",
  16477=>"001001000",
  16478=>"100100100",
  16479=>"001000000",
  16480=>"100000000",
  16481=>"111111001",
  16482=>"000110110",
  16483=>"111111111",
  16484=>"101111111",
  16485=>"111111111",
  16486=>"011110000",
  16487=>"000000000",
  16488=>"000000000",
  16489=>"111111111",
  16490=>"000001111",
  16491=>"000000000",
  16492=>"000000000",
  16493=>"000000000",
  16494=>"000000100",
  16495=>"111111111",
  16496=>"111111111",
  16497=>"010110010",
  16498=>"011011011",
  16499=>"011000000",
  16500=>"000010010",
  16501=>"000000000",
  16502=>"000101111",
  16503=>"000000100",
  16504=>"000000000",
  16505=>"111110000",
  16506=>"100101111",
  16507=>"111111111",
  16508=>"011111111",
  16509=>"100100100",
  16510=>"100100100",
  16511=>"111011000",
  16512=>"000000001",
  16513=>"111111111",
  16514=>"000000001",
  16515=>"001100000",
  16516=>"111111111",
  16517=>"001000010",
  16518=>"000000000",
  16519=>"011011111",
  16520=>"111111111",
  16521=>"000000000",
  16522=>"000000000",
  16523=>"111111111",
  16524=>"111111101",
  16525=>"011111110",
  16526=>"111111111",
  16527=>"000000000",
  16528=>"111111111",
  16529=>"110111110",
  16530=>"011111111",
  16531=>"101001001",
  16532=>"000000000",
  16533=>"111100000",
  16534=>"000111111",
  16535=>"000000000",
  16536=>"100000000",
  16537=>"111111111",
  16538=>"111000000",
  16539=>"001000000",
  16540=>"000001011",
  16541=>"000000000",
  16542=>"110101111",
  16543=>"111111111",
  16544=>"111110110",
  16545=>"000010110",
  16546=>"111111100",
  16547=>"111111111",
  16548=>"100110111",
  16549=>"110111000",
  16550=>"110111111",
  16551=>"111111111",
  16552=>"000000111",
  16553=>"011111110",
  16554=>"000000000",
  16555=>"001111001",
  16556=>"000000000",
  16557=>"000000000",
  16558=>"000000001",
  16559=>"000000000",
  16560=>"100111000",
  16561=>"001000000",
  16562=>"111111111",
  16563=>"000000100",
  16564=>"000000000",
  16565=>"101100000",
  16566=>"000000000",
  16567=>"111111111",
  16568=>"000000000",
  16569=>"011000000",
  16570=>"100000000",
  16571=>"111111111",
  16572=>"000000000",
  16573=>"000000111",
  16574=>"110110100",
  16575=>"111101111",
  16576=>"011011111",
  16577=>"011000000",
  16578=>"000100101",
  16579=>"000000000",
  16580=>"000000000",
  16581=>"000000000",
  16582=>"100111110",
  16583=>"100100000",
  16584=>"000000000",
  16585=>"000000000",
  16586=>"011111100",
  16587=>"110100100",
  16588=>"111111000",
  16589=>"101001000",
  16590=>"000000101",
  16591=>"100111111",
  16592=>"000000000",
  16593=>"000000000",
  16594=>"111111000",
  16595=>"000000000",
  16596=>"011001011",
  16597=>"100001001",
  16598=>"100000000",
  16599=>"000000000",
  16600=>"111111010",
  16601=>"110000000",
  16602=>"011000000",
  16603=>"011011110",
  16604=>"111111111",
  16605=>"101100101",
  16606=>"111111000",
  16607=>"000000000",
  16608=>"000000000",
  16609=>"110111111",
  16610=>"000000000",
  16611=>"111111111",
  16612=>"100000100",
  16613=>"110111111",
  16614=>"111111111",
  16615=>"000000000",
  16616=>"000100100",
  16617=>"000011111",
  16618=>"100100110",
  16619=>"000000000",
  16620=>"000000000",
  16621=>"111011111",
  16622=>"111111000",
  16623=>"111000110",
  16624=>"111000000",
  16625=>"111111111",
  16626=>"111111111",
  16627=>"011011111",
  16628=>"111110110",
  16629=>"000000000",
  16630=>"100110110",
  16631=>"000111000",
  16632=>"100000000",
  16633=>"000010000",
  16634=>"011111111",
  16635=>"000000000",
  16636=>"100100110",
  16637=>"000000100",
  16638=>"111111111",
  16639=>"000000111",
  16640=>"011110000",
  16641=>"001001001",
  16642=>"101101111",
  16643=>"111111111",
  16644=>"000000000",
  16645=>"000000000",
  16646=>"000000000",
  16647=>"111011001",
  16648=>"000000000",
  16649=>"111000100",
  16650=>"111111000",
  16651=>"001011111",
  16652=>"000000000",
  16653=>"000000000",
  16654=>"111111011",
  16655=>"000000000",
  16656=>"111000111",
  16657=>"111111111",
  16658=>"000000000",
  16659=>"101100111",
  16660=>"111111000",
  16661=>"000000000",
  16662=>"011111111",
  16663=>"000000111",
  16664=>"011011111",
  16665=>"000000000",
  16666=>"011011111",
  16667=>"111000000",
  16668=>"000000110",
  16669=>"000011111",
  16670=>"111111111",
  16671=>"011000000",
  16672=>"100001000",
  16673=>"000000000",
  16674=>"000000001",
  16675=>"111111111",
  16676=>"000000000",
  16677=>"110110110",
  16678=>"001100100",
  16679=>"000000111",
  16680=>"111101000",
  16681=>"111110111",
  16682=>"110000000",
  16683=>"011001111",
  16684=>"000000101",
  16685=>"111111111",
  16686=>"111101000",
  16687=>"000000000",
  16688=>"000100000",
  16689=>"110000000",
  16690=>"111111000",
  16691=>"111110111",
  16692=>"111111111",
  16693=>"000000000",
  16694=>"001000000",
  16695=>"111111011",
  16696=>"000000000",
  16697=>"000000000",
  16698=>"110100000",
  16699=>"100111111",
  16700=>"011011111",
  16701=>"000000000",
  16702=>"000100111",
  16703=>"110110110",
  16704=>"111111111",
  16705=>"000000100",
  16706=>"101100011",
  16707=>"000000000",
  16708=>"001001100",
  16709=>"001111111",
  16710=>"000000000",
  16711=>"000100110",
  16712=>"011011111",
  16713=>"011010000",
  16714=>"010111001",
  16715=>"000000000",
  16716=>"011000000",
  16717=>"000000011",
  16718=>"000000000",
  16719=>"100100110",
  16720=>"111110110",
  16721=>"000000111",
  16722=>"111101111",
  16723=>"111100111",
  16724=>"111111011",
  16725=>"001011101",
  16726=>"111111000",
  16727=>"000000100",
  16728=>"000000111",
  16729=>"111110111",
  16730=>"000011011",
  16731=>"000010110",
  16732=>"110111111",
  16733=>"000011011",
  16734=>"010000000",
  16735=>"001111001",
  16736=>"110000000",
  16737=>"111111111",
  16738=>"100100110",
  16739=>"000000000",
  16740=>"111111011",
  16741=>"000000100",
  16742=>"010000000",
  16743=>"111110111",
  16744=>"010000000",
  16745=>"111111101",
  16746=>"000000000",
  16747=>"000000000",
  16748=>"111111111",
  16749=>"000111111",
  16750=>"000000111",
  16751=>"000000000",
  16752=>"111000000",
  16753=>"111101001",
  16754=>"010011111",
  16755=>"111101111",
  16756=>"000000000",
  16757=>"001000000",
  16758=>"001101001",
  16759=>"000000000",
  16760=>"001000000",
  16761=>"000000100",
  16762=>"100000000",
  16763=>"111111110",
  16764=>"000000100",
  16765=>"111111110",
  16766=>"111111111",
  16767=>"000000000",
  16768=>"011011000",
  16769=>"111111111",
  16770=>"111111111",
  16771=>"000100110",
  16772=>"111111111",
  16773=>"000000100",
  16774=>"011001000",
  16775=>"000000100",
  16776=>"001000000",
  16777=>"001000011",
  16778=>"001000000",
  16779=>"001001000",
  16780=>"000000000",
  16781=>"000100000",
  16782=>"000000000",
  16783=>"000000000",
  16784=>"000000000",
  16785=>"111110110",
  16786=>"110111111",
  16787=>"111111111",
  16788=>"000101111",
  16789=>"000000000",
  16790=>"111111111",
  16791=>"000000010",
  16792=>"100100111",
  16793=>"111111111",
  16794=>"000000000",
  16795=>"111111111",
  16796=>"100100011",
  16797=>"111100000",
  16798=>"111101100",
  16799=>"110110000",
  16800=>"000000000",
  16801=>"011000001",
  16802=>"100100000",
  16803=>"000001001",
  16804=>"011000000",
  16805=>"110111110",
  16806=>"000000000",
  16807=>"111111000",
  16808=>"010010001",
  16809=>"010000000",
  16810=>"111111111",
  16811=>"111000000",
  16812=>"111000000",
  16813=>"001001111",
  16814=>"111000000",
  16815=>"000000000",
  16816=>"001011000",
  16817=>"000000000",
  16818=>"111000100",
  16819=>"111111111",
  16820=>"011100100",
  16821=>"000010111",
  16822=>"111111111",
  16823=>"000100100",
  16824=>"100000000",
  16825=>"111111111",
  16826=>"111100000",
  16827=>"101100110",
  16828=>"000000100",
  16829=>"111111111",
  16830=>"000000000",
  16831=>"000000100",
  16832=>"000110111",
  16833=>"001001111",
  16834=>"001000000",
  16835=>"000000000",
  16836=>"111111110",
  16837=>"000000110",
  16838=>"010000000",
  16839=>"111111111",
  16840=>"100100000",
  16841=>"000000111",
  16842=>"000000000",
  16843=>"000000100",
  16844=>"000000111",
  16845=>"000000000",
  16846=>"001000000",
  16847=>"001111111",
  16848=>"001111001",
  16849=>"110000000",
  16850=>"000000000",
  16851=>"011111111",
  16852=>"010000000",
  16853=>"111111111",
  16854=>"111111000",
  16855=>"111111111",
  16856=>"011111111",
  16857=>"111100100",
  16858=>"000000000",
  16859=>"100100100",
  16860=>"100000101",
  16861=>"110011011",
  16862=>"010011111",
  16863=>"001001111",
  16864=>"111111111",
  16865=>"111111111",
  16866=>"111101001",
  16867=>"001000000",
  16868=>"111111101",
  16869=>"000000000",
  16870=>"010010000",
  16871=>"000000011",
  16872=>"111101111",
  16873=>"111111100",
  16874=>"000100101",
  16875=>"100111111",
  16876=>"000111011",
  16877=>"000100100",
  16878=>"111111111",
  16879=>"111111111",
  16880=>"000100110",
  16881=>"111110011",
  16882=>"110110100",
  16883=>"111100110",
  16884=>"011111110",
  16885=>"000000000",
  16886=>"111111111",
  16887=>"000000000",
  16888=>"001111111",
  16889=>"000000100",
  16890=>"011010000",
  16891=>"100000111",
  16892=>"100100100",
  16893=>"011000011",
  16894=>"000000000",
  16895=>"100100111",
  16896=>"110110110",
  16897=>"010010111",
  16898=>"111101100",
  16899=>"001000001",
  16900=>"110111101",
  16901=>"000001111",
  16902=>"101101000",
  16903=>"000000000",
  16904=>"111000101",
  16905=>"111111101",
  16906=>"001001001",
  16907=>"001001111",
  16908=>"001001001",
  16909=>"111101101",
  16910=>"100100111",
  16911=>"101000001",
  16912=>"000000001",
  16913=>"111010000",
  16914=>"110010010",
  16915=>"001001000",
  16916=>"111001001",
  16917=>"111110110",
  16918=>"001000000",
  16919=>"000000000",
  16920=>"001001001",
  16921=>"111110111",
  16922=>"000000000",
  16923=>"101100111",
  16924=>"001001001",
  16925=>"000100000",
  16926=>"110110110",
  16927=>"000000101",
  16928=>"110000000",
  16929=>"110010011",
  16930=>"001000110",
  16931=>"111111111",
  16932=>"110011000",
  16933=>"011011111",
  16934=>"010010110",
  16935=>"001101111",
  16936=>"000000000",
  16937=>"000000010",
  16938=>"001001111",
  16939=>"111001000",
  16940=>"110111111",
  16941=>"111101001",
  16942=>"001001101",
  16943=>"111101101",
  16944=>"101000000",
  16945=>"001001001",
  16946=>"111101101",
  16947=>"000000110",
  16948=>"111111001",
  16949=>"001000000",
  16950=>"000000100",
  16951=>"111111100",
  16952=>"110110110",
  16953=>"000100100",
  16954=>"101000101",
  16955=>"000001001",
  16956=>"111101000",
  16957=>"000110111",
  16958=>"110110000",
  16959=>"111111111",
  16960=>"001011011",
  16961=>"001000100",
  16962=>"001011101",
  16963=>"110111101",
  16964=>"001001011",
  16965=>"000000000",
  16966=>"001001111",
  16967=>"010111111",
  16968=>"010000100",
  16969=>"000000000",
  16970=>"110110111",
  16971=>"110111110",
  16972=>"111110110",
  16973=>"110110000",
  16974=>"000000101",
  16975=>"001101111",
  16976=>"000000001",
  16977=>"111111111",
  16978=>"000000000",
  16979=>"010110110",
  16980=>"001000000",
  16981=>"000000010",
  16982=>"000000001",
  16983=>"001001000",
  16984=>"000001110",
  16985=>"111101101",
  16986=>"010010000",
  16987=>"110100101",
  16988=>"000010110",
  16989=>"110110111",
  16990=>"000000111",
  16991=>"000000000",
  16992=>"000000000",
  16993=>"000000000",
  16994=>"100110110",
  16995=>"011111010",
  16996=>"000000000",
  16997=>"000000000",
  16998=>"011111111",
  16999=>"111111010",
  17000=>"001001001",
  17001=>"111111111",
  17002=>"010110000",
  17003=>"110000000",
  17004=>"110110111",
  17005=>"001000000",
  17006=>"001001101",
  17007=>"000000011",
  17008=>"000000111",
  17009=>"001111111",
  17010=>"000000001",
  17011=>"011001111",
  17012=>"000000000",
  17013=>"111111111",
  17014=>"111100000",
  17015=>"000000100",
  17016=>"110110110",
  17017=>"000001000",
  17018=>"001001001",
  17019=>"011001000",
  17020=>"100100100",
  17021=>"000010011",
  17022=>"101101001",
  17023=>"000001000",
  17024=>"001000101",
  17025=>"111111110",
  17026=>"010111111",
  17027=>"110010011",
  17028=>"000111111",
  17029=>"001001101",
  17030=>"100110110",
  17031=>"000000000",
  17032=>"001001001",
  17033=>"111111111",
  17034=>"111111111",
  17035=>"111001001",
  17036=>"000000000",
  17037=>"000000010",
  17038=>"010011000",
  17039=>"000000000",
  17040=>"011111111",
  17041=>"000000010",
  17042=>"000010011",
  17043=>"111001011",
  17044=>"110110110",
  17045=>"101101111",
  17046=>"110111111",
  17047=>"111010000",
  17048=>"001101001",
  17049=>"111111111",
  17050=>"111101000",
  17051=>"000000111",
  17052=>"000000000",
  17053=>"111111111",
  17054=>"111111111",
  17055=>"111101000",
  17056=>"010100000",
  17057=>"001001111",
  17058=>"000000001",
  17059=>"001101101",
  17060=>"001001001",
  17061=>"000000000",
  17062=>"110010010",
  17063=>"111111010",
  17064=>"001000000",
  17065=>"110110110",
  17066=>"111111111",
  17067=>"111001111",
  17068=>"001000001",
  17069=>"110110110",
  17070=>"111111111",
  17071=>"111010010",
  17072=>"000001001",
  17073=>"000010111",
  17074=>"111111111",
  17075=>"010000000",
  17076=>"111000000",
  17077=>"001101111",
  17078=>"001000000",
  17079=>"110110111",
  17080=>"101101101",
  17081=>"101001001",
  17082=>"001101001",
  17083=>"101100001",
  17084=>"000000000",
  17085=>"000000101",
  17086=>"010000010",
  17087=>"110110111",
  17088=>"000000000",
  17089=>"000001000",
  17090=>"000000111",
  17091=>"110110110",
  17092=>"000010011",
  17093=>"010010000",
  17094=>"000111100",
  17095=>"100100000",
  17096=>"111110110",
  17097=>"101101101",
  17098=>"001001001",
  17099=>"001001101",
  17100=>"100101111",
  17101=>"001111111",
  17102=>"110000101",
  17103=>"001000000",
  17104=>"100000111",
  17105=>"111010111",
  17106=>"000100111",
  17107=>"101101101",
  17108=>"000100111",
  17109=>"001101111",
  17110=>"001001001",
  17111=>"101101111",
  17112=>"000000010",
  17113=>"101111110",
  17114=>"000000000",
  17115=>"000000000",
  17116=>"100000100",
  17117=>"111011111",
  17118=>"010011010",
  17119=>"001111110",
  17120=>"000000000",
  17121=>"000000000",
  17122=>"111111111",
  17123=>"110100000",
  17124=>"111000000",
  17125=>"001000000",
  17126=>"011001001",
  17127=>"111111000",
  17128=>"100100100",
  17129=>"110000100",
  17130=>"111001100",
  17131=>"100100111",
  17132=>"001000000",
  17133=>"000000000",
  17134=>"111111000",
  17135=>"000110111",
  17136=>"111111110",
  17137=>"100111111",
  17138=>"101001111",
  17139=>"001001101",
  17140=>"000110000",
  17141=>"000000000",
  17142=>"011011011",
  17143=>"000000000",
  17144=>"110110110",
  17145=>"110111111",
  17146=>"000000000",
  17147=>"000101111",
  17148=>"011111001",
  17149=>"000001001",
  17150=>"011000000",
  17151=>"001001001",
  17152=>"011000100",
  17153=>"001001001",
  17154=>"000000000",
  17155=>"110011111",
  17156=>"101011111",
  17157=>"111111110",
  17158=>"000000000",
  17159=>"010010100",
  17160=>"001001101",
  17161=>"101111111",
  17162=>"101001101",
  17163=>"000000101",
  17164=>"010010000",
  17165=>"101001011",
  17166=>"111111111",
  17167=>"011011111",
  17168=>"000000100",
  17169=>"000011111",
  17170=>"101001001",
  17171=>"000001011",
  17172=>"001001000",
  17173=>"000000101",
  17174=>"100100100",
  17175=>"110111110",
  17176=>"111111110",
  17177=>"000110011",
  17178=>"010010010",
  17179=>"111000000",
  17180=>"000001011",
  17181=>"010111111",
  17182=>"111111111",
  17183=>"000000101",
  17184=>"001011110",
  17185=>"010000100",
  17186=>"000000111",
  17187=>"110111111",
  17188=>"000010111",
  17189=>"111111111",
  17190=>"101001001",
  17191=>"000000000",
  17192=>"101101111",
  17193=>"000001001",
  17194=>"101000111",
  17195=>"111111101",
  17196=>"000000110",
  17197=>"000000100",
  17198=>"000000100",
  17199=>"101100000",
  17200=>"110111110",
  17201=>"001001000",
  17202=>"111111110",
  17203=>"010110110",
  17204=>"010000010",
  17205=>"111000111",
  17206=>"000000000",
  17207=>"101111111",
  17208=>"000110110",
  17209=>"111111111",
  17210=>"001001001",
  17211=>"001101101",
  17212=>"111111111",
  17213=>"100100111",
  17214=>"010000001",
  17215=>"010110110",
  17216=>"000000010",
  17217=>"111100101",
  17218=>"111100100",
  17219=>"001001001",
  17220=>"001101000",
  17221=>"001011111",
  17222=>"000000000",
  17223=>"001001101",
  17224=>"010010000",
  17225=>"000000101",
  17226=>"000000001",
  17227=>"000000010",
  17228=>"011001001",
  17229=>"100100001",
  17230=>"111111111",
  17231=>"110110100",
  17232=>"001011000",
  17233=>"101100000",
  17234=>"110110000",
  17235=>"010010110",
  17236=>"110110110",
  17237=>"011011011",
  17238=>"111010000",
  17239=>"111111011",
  17240=>"111110110",
  17241=>"111110000",
  17242=>"110110010",
  17243=>"101000101",
  17244=>"010110111",
  17245=>"000001111",
  17246=>"101001101",
  17247=>"110110110",
  17248=>"110010010",
  17249=>"010111011",
  17250=>"011011010",
  17251=>"101101001",
  17252=>"000010110",
  17253=>"000000000",
  17254=>"000000000",
  17255=>"111111111",
  17256=>"110100100",
  17257=>"100000010",
  17258=>"111111100",
  17259=>"000101001",
  17260=>"010010110",
  17261=>"111111111",
  17262=>"111111110",
  17263=>"000000100",
  17264=>"010010111",
  17265=>"001001001",
  17266=>"111111111",
  17267=>"000000000",
  17268=>"011011100",
  17269=>"101101001",
  17270=>"000000000",
  17271=>"001000000",
  17272=>"111101101",
  17273=>"000010010",
  17274=>"011010010",
  17275=>"001001101",
  17276=>"000000000",
  17277=>"111111111",
  17278=>"001001000",
  17279=>"000000100",
  17280=>"000000111",
  17281=>"111110111",
  17282=>"000000001",
  17283=>"000000011",
  17284=>"111000000",
  17285=>"110101000",
  17286=>"011000100",
  17287=>"111000000",
  17288=>"001001000",
  17289=>"011011011",
  17290=>"101101101",
  17291=>"111101101",
  17292=>"000000000",
  17293=>"011000010",
  17294=>"000000100",
  17295=>"000000001",
  17296=>"010010000",
  17297=>"000000000",
  17298=>"111111110",
  17299=>"110110110",
  17300=>"000000000",
  17301=>"000000000",
  17302=>"000000000",
  17303=>"001001101",
  17304=>"111111111",
  17305=>"000100111",
  17306=>"000000000",
  17307=>"000001001",
  17308=>"101001001",
  17309=>"001001001",
  17310=>"001101001",
  17311=>"000000001",
  17312=>"001101111",
  17313=>"111111011",
  17314=>"111011000",
  17315=>"001000000",
  17316=>"000000100",
  17317=>"110111111",
  17318=>"000010111",
  17319=>"110110111",
  17320=>"100000110",
  17321=>"000000110",
  17322=>"000000010",
  17323=>"001001111",
  17324=>"000000000",
  17325=>"001000000",
  17326=>"010110110",
  17327=>"001111111",
  17328=>"111111111",
  17329=>"000000000",
  17330=>"111111011",
  17331=>"000001011",
  17332=>"000011111",
  17333=>"101101111",
  17334=>"111111111",
  17335=>"000000011",
  17336=>"101101000",
  17337=>"010011011",
  17338=>"000000000",
  17339=>"111000000",
  17340=>"000010111",
  17341=>"111011011",
  17342=>"000000001",
  17343=>"111110111",
  17344=>"000000000",
  17345=>"111111001",
  17346=>"001001101",
  17347=>"000000000",
  17348=>"001001000",
  17349=>"111111111",
  17350=>"110110110",
  17351=>"110001000",
  17352=>"101100100",
  17353=>"011000010",
  17354=>"000000000",
  17355=>"011111000",
  17356=>"000000000",
  17357=>"110110110",
  17358=>"001000110",
  17359=>"001001101",
  17360=>"000001111",
  17361=>"111110110",
  17362=>"110110010",
  17363=>"001011111",
  17364=>"000000000",
  17365=>"111101000",
  17366=>"000000000",
  17367=>"100100100",
  17368=>"111111111",
  17369=>"111110000",
  17370=>"000001001",
  17371=>"110110100",
  17372=>"101111011",
  17373=>"110111111",
  17374=>"110000000",
  17375=>"001001001",
  17376=>"000100100",
  17377=>"000001001",
  17378=>"101000100",
  17379=>"010100111",
  17380=>"111110110",
  17381=>"010011001",
  17382=>"010000000",
  17383=>"001000101",
  17384=>"000001111",
  17385=>"111110111",
  17386=>"001000000",
  17387=>"101001111",
  17388=>"100100111",
  17389=>"101001011",
  17390=>"111111010",
  17391=>"111111111",
  17392=>"000000001",
  17393=>"100101111",
  17394=>"111001101",
  17395=>"010000111",
  17396=>"011011110",
  17397=>"111111111",
  17398=>"110111110",
  17399=>"110110110",
  17400=>"110111111",
  17401=>"000111101",
  17402=>"100000111",
  17403=>"000000000",
  17404=>"111001111",
  17405=>"001000100",
  17406=>"111111110",
  17407=>"000001111",
  17408=>"111000100",
  17409=>"000000000",
  17410=>"000000110",
  17411=>"110111111",
  17412=>"110100110",
  17413=>"111001000",
  17414=>"110100000",
  17415=>"000000000",
  17416=>"001000011",
  17417=>"111010000",
  17418=>"110110110",
  17419=>"111111111",
  17420=>"110110110",
  17421=>"111010000",
  17422=>"100100100",
  17423=>"001101111",
  17424=>"001100111",
  17425=>"111111101",
  17426=>"110110110",
  17427=>"000000000",
  17428=>"000000111",
  17429=>"111111111",
  17430=>"100101101",
  17431=>"011001000",
  17432=>"111110110",
  17433=>"110100111",
  17434=>"111111111",
  17435=>"111100001",
  17436=>"001001000",
  17437=>"010011011",
  17438=>"100000001",
  17439=>"011001000",
  17440=>"000010111",
  17441=>"111110000",
  17442=>"000000000",
  17443=>"000000000",
  17444=>"111111111",
  17445=>"111111111",
  17446=>"110111010",
  17447=>"111110000",
  17448=>"111111010",
  17449=>"000000010",
  17450=>"111110000",
  17451=>"111000000",
  17452=>"001001111",
  17453=>"000111110",
  17454=>"001001001",
  17455=>"111011111",
  17456=>"000011111",
  17457=>"111101101",
  17458=>"111100100",
  17459=>"111011001",
  17460=>"111001100",
  17461=>"000000001",
  17462=>"111101111",
  17463=>"111111000",
  17464=>"001000000",
  17465=>"000000000",
  17466=>"000000000",
  17467=>"110110010",
  17468=>"100010000",
  17469=>"101000100",
  17470=>"101110111",
  17471=>"101101101",
  17472=>"110111111",
  17473=>"111110110",
  17474=>"101000000",
  17475=>"011010010",
  17476=>"110110110",
  17477=>"000000000",
  17478=>"010000000",
  17479=>"101101111",
  17480=>"110111000",
  17481=>"011011011",
  17482=>"111111111",
  17483=>"000000000",
  17484=>"000111111",
  17485=>"111111111",
  17486=>"000111111",
  17487=>"011110110",
  17488=>"000001100",
  17489=>"110111111",
  17490=>"110000110",
  17491=>"011001011",
  17492=>"001001001",
  17493=>"000000110",
  17494=>"111111011",
  17495=>"100000000",
  17496=>"001000001",
  17497=>"001001101",
  17498=>"111111111",
  17499=>"110110110",
  17500=>"000000000",
  17501=>"101101111",
  17502=>"010000001",
  17503=>"100111111",
  17504=>"000000011",
  17505=>"111111111",
  17506=>"000000000",
  17507=>"101001001",
  17508=>"111111011",
  17509=>"110000000",
  17510=>"111110100",
  17511=>"111111001",
  17512=>"111101111",
  17513=>"001100111",
  17514=>"001001000",
  17515=>"000000000",
  17516=>"110110110",
  17517=>"001000000",
  17518=>"000001111",
  17519=>"001111111",
  17520=>"111011011",
  17521=>"000001111",
  17522=>"101001001",
  17523=>"000000000",
  17524=>"111111110",
  17525=>"001000000",
  17526=>"110110000",
  17527=>"101100111",
  17528=>"000000000",
  17529=>"111011010",
  17530=>"001000000",
  17531=>"000000000",
  17532=>"110110110",
  17533=>"110110110",
  17534=>"000000000",
  17535=>"000000000",
  17536=>"001000000",
  17537=>"110010010",
  17538=>"111000000",
  17539=>"011011000",
  17540=>"111111111",
  17541=>"010110000",
  17542=>"000000111",
  17543=>"001000000",
  17544=>"000000010",
  17545=>"000000000",
  17546=>"101100000",
  17547=>"111111111",
  17548=>"101101111",
  17549=>"001001101",
  17550=>"001101101",
  17551=>"111000000",
  17552=>"001000100",
  17553=>"000011011",
  17554=>"111100100",
  17555=>"000000000",
  17556=>"000000000",
  17557=>"000000000",
  17558=>"000010000",
  17559=>"111111111",
  17560=>"001000100",
  17561=>"001000101",
  17562=>"001000001",
  17563=>"010000001",
  17564=>"111011001",
  17565=>"111110110",
  17566=>"111111111",
  17567=>"111100000",
  17568=>"000000111",
  17569=>"101101001",
  17570=>"111111010",
  17571=>"000000000",
  17572=>"000000110",
  17573=>"000000001",
  17574=>"000001010",
  17575=>"000000000",
  17576=>"000000100",
  17577=>"011001111",
  17578=>"001001000",
  17579=>"000000000",
  17580=>"111111001",
  17581=>"000110111",
  17582=>"000000000",
  17583=>"100100000",
  17584=>"111111101",
  17585=>"111111111",
  17586=>"110111110",
  17587=>"000000111",
  17588=>"000000000",
  17589=>"001000000",
  17590=>"111111111",
  17591=>"100111111",
  17592=>"001001000",
  17593=>"010010011",
  17594=>"001000000",
  17595=>"000000000",
  17596=>"111001001",
  17597=>"011110111",
  17598=>"000000000",
  17599=>"111110111",
  17600=>"111111111",
  17601=>"000000000",
  17602=>"110111010",
  17603=>"000110110",
  17604=>"110100111",
  17605=>"000000000",
  17606=>"000110110",
  17607=>"100100110",
  17608=>"000011001",
  17609=>"000000111",
  17610=>"000000111",
  17611=>"111100000",
  17612=>"010110100",
  17613=>"000100000",
  17614=>"100100100",
  17615=>"000000000",
  17616=>"100000000",
  17617=>"111111111",
  17618=>"000000000",
  17619=>"000000000",
  17620=>"000000001",
  17621=>"011001111",
  17622=>"001001000",
  17623=>"100101100",
  17624=>"000000111",
  17625=>"000000000",
  17626=>"110110000",
  17627=>"001000000",
  17628=>"001000000",
  17629=>"001001111",
  17630=>"001000101",
  17631=>"000000101",
  17632=>"100100111",
  17633=>"000000111",
  17634=>"010010010",
  17635=>"000000000",
  17636=>"110111000",
  17637=>"111111111",
  17638=>"111011111",
  17639=>"110110010",
  17640=>"000000000",
  17641=>"001001001",
  17642=>"111111011",
  17643=>"101100110",
  17644=>"000000000",
  17645=>"111011001",
  17646=>"000000000",
  17647=>"001000000",
  17648=>"001001100",
  17649=>"011111111",
  17650=>"111110110",
  17651=>"000010001",
  17652=>"101001101",
  17653=>"011111111",
  17654=>"011001011",
  17655=>"110111111",
  17656=>"010000010",
  17657=>"000000000",
  17658=>"001101101",
  17659=>"111111001",
  17660=>"000000000",
  17661=>"001011101",
  17662=>"000011011",
  17663=>"111000000",
  17664=>"100110000",
  17665=>"001000000",
  17666=>"001001111",
  17667=>"000000000",
  17668=>"100000110",
  17669=>"000001000",
  17670=>"000111111",
  17671=>"111111111",
  17672=>"111111000",
  17673=>"001000001",
  17674=>"000000100",
  17675=>"011001000",
  17676=>"111010110",
  17677=>"000111111",
  17678=>"001000101",
  17679=>"110110000",
  17680=>"111111111",
  17681=>"001001001",
  17682=>"000100110",
  17683=>"111101100",
  17684=>"000000000",
  17685=>"111110111",
  17686=>"111011001",
  17687=>"111111111",
  17688=>"000000111",
  17689=>"001000000",
  17690=>"110000010",
  17691=>"111111111",
  17692=>"111100000",
  17693=>"011011000",
  17694=>"000110000",
  17695=>"100101111",
  17696=>"111000001",
  17697=>"111111010",
  17698=>"000111111",
  17699=>"111001000",
  17700=>"000000000",
  17701=>"110111110",
  17702=>"111110100",
  17703=>"100100111",
  17704=>"011111111",
  17705=>"110000000",
  17706=>"001000000",
  17707=>"000000000",
  17708=>"010000000",
  17709=>"111001000",
  17710=>"110000010",
  17711=>"101100111",
  17712=>"110110110",
  17713=>"110010011",
  17714=>"111000000",
  17715=>"000001011",
  17716=>"111010010",
  17717=>"000000000",
  17718=>"011111111",
  17719=>"001011001",
  17720=>"010010010",
  17721=>"111111110",
  17722=>"000001111",
  17723=>"000000010",
  17724=>"110111111",
  17725=>"010110110",
  17726=>"110110111",
  17727=>"111111010",
  17728=>"111001000",
  17729=>"001001111",
  17730=>"010110110",
  17731=>"001001111",
  17732=>"001001001",
  17733=>"101101001",
  17734=>"110000000",
  17735=>"110111110",
  17736=>"001100111",
  17737=>"111001000",
  17738=>"001000001",
  17739=>"101101110",
  17740=>"000000000",
  17741=>"000001000",
  17742=>"000010000",
  17743=>"111110000",
  17744=>"000000000",
  17745=>"001000000",
  17746=>"111111100",
  17747=>"000000011",
  17748=>"110000000",
  17749=>"111111011",
  17750=>"000000000",
  17751=>"111111111",
  17752=>"110000011",
  17753=>"111111110",
  17754=>"000110110",
  17755=>"001000001",
  17756=>"111000000",
  17757=>"000000000",
  17758=>"110111111",
  17759=>"000100011",
  17760=>"000100000",
  17761=>"100111101",
  17762=>"001001001",
  17763=>"001000001",
  17764=>"110110111",
  17765=>"000000000",
  17766=>"110110111",
  17767=>"110110110",
  17768=>"111101111",
  17769=>"111111011",
  17770=>"001001000",
  17771=>"100001101",
  17772=>"000000100",
  17773=>"101111010",
  17774=>"000000100",
  17775=>"001101111",
  17776=>"011111010",
  17777=>"001001101",
  17778=>"000000101",
  17779=>"000000000",
  17780=>"101001101",
  17781=>"111111110",
  17782=>"111000000",
  17783=>"110110110",
  17784=>"001101111",
  17785=>"000000000",
  17786=>"110100100",
  17787=>"000000000",
  17788=>"000000000",
  17789=>"000000000",
  17790=>"111111111",
  17791=>"001101111",
  17792=>"000000000",
  17793=>"000000100",
  17794=>"100000100",
  17795=>"000000110",
  17796=>"111111111",
  17797=>"000110000",
  17798=>"100111111",
  17799=>"111001111",
  17800=>"110101000",
  17801=>"000100111",
  17802=>"111111000",
  17803=>"011011000",
  17804=>"111111111",
  17805=>"111011000",
  17806=>"110110010",
  17807=>"111000000",
  17808=>"000000000",
  17809=>"000000011",
  17810=>"100101001",
  17811=>"111111110",
  17812=>"001111111",
  17813=>"010010000",
  17814=>"001001001",
  17815=>"100100110",
  17816=>"101000000",
  17817=>"101000000",
  17818=>"000000101",
  17819=>"001001011",
  17820=>"110010000",
  17821=>"000111111",
  17822=>"011001000",
  17823=>"001000000",
  17824=>"000000100",
  17825=>"110000000",
  17826=>"111010010",
  17827=>"100110111",
  17828=>"001001001",
  17829=>"000000001",
  17830=>"111111101",
  17831=>"000100110",
  17832=>"011001000",
  17833=>"111011001",
  17834=>"001001010",
  17835=>"001001000",
  17836=>"110110000",
  17837=>"111111111",
  17838=>"000000101",
  17839=>"000000111",
  17840=>"001001000",
  17841=>"000000000",
  17842=>"001111101",
  17843=>"111111110",
  17844=>"111111111",
  17845=>"000000000",
  17846=>"000000000",
  17847=>"110010000",
  17848=>"010000110",
  17849=>"110110110",
  17850=>"000001101",
  17851=>"000000000",
  17852=>"000000100",
  17853=>"000001001",
  17854=>"000000001",
  17855=>"011011001",
  17856=>"000010000",
  17857=>"001001101",
  17858=>"000011111",
  17859=>"001001011",
  17860=>"111110110",
  17861=>"000001111",
  17862=>"101100111",
  17863=>"000000000",
  17864=>"000000000",
  17865=>"000000100",
  17866=>"111111111",
  17867=>"010000000",
  17868=>"000100100",
  17869=>"111110010",
  17870=>"000011111",
  17871=>"000001111",
  17872=>"111111011",
  17873=>"111111001",
  17874=>"000000110",
  17875=>"111111111",
  17876=>"000001001",
  17877=>"000010010",
  17878=>"000100111",
  17879=>"111111011",
  17880=>"111111111",
  17881=>"000000000",
  17882=>"001001111",
  17883=>"001000000",
  17884=>"011011000",
  17885=>"111000000",
  17886=>"001011000",
  17887=>"001001011",
  17888=>"000100111",
  17889=>"000000110",
  17890=>"000000000",
  17891=>"100100111",
  17892=>"001001000",
  17893=>"001111100",
  17894=>"000000001",
  17895=>"000001111",
  17896=>"111111111",
  17897=>"111000000",
  17898=>"001011111",
  17899=>"001000011",
  17900=>"000110111",
  17901=>"011111110",
  17902=>"000000000",
  17903=>"111111111",
  17904=>"111001100",
  17905=>"111111111",
  17906=>"111111100",
  17907=>"101101000",
  17908=>"110111111",
  17909=>"010111111",
  17910=>"111111000",
  17911=>"111111110",
  17912=>"000000010",
  17913=>"110110110",
  17914=>"111100000",
  17915=>"100000000",
  17916=>"110110111",
  17917=>"111011111",
  17918=>"000000000",
  17919=>"011000000",
  17920=>"000111111",
  17921=>"000000111",
  17922=>"000111000",
  17923=>"000000111",
  17924=>"000111111",
  17925=>"011000000",
  17926=>"110000000",
  17927=>"111111111",
  17928=>"111111000",
  17929=>"111111000",
  17930=>"000111111",
  17931=>"110111011",
  17932=>"110110000",
  17933=>"000000100",
  17934=>"111111111",
  17935=>"000000000",
  17936=>"100000111",
  17937=>"000111110",
  17938=>"000111011",
  17939=>"111110111",
  17940=>"111000010",
  17941=>"000000000",
  17942=>"000010010",
  17943=>"000111111",
  17944=>"001111111",
  17945=>"011001111",
  17946=>"000000000",
  17947=>"000111110",
  17948=>"000000100",
  17949=>"111111011",
  17950=>"111111111",
  17951=>"101111111",
  17952=>"000000001",
  17953=>"000111110",
  17954=>"001110000",
  17955=>"000000010",
  17956=>"000110010",
  17957=>"100110111",
  17958=>"011111111",
  17959=>"100000000",
  17960=>"000000000",
  17961=>"000000000",
  17962=>"000000111",
  17963=>"000000000",
  17964=>"011111111",
  17965=>"000000000",
  17966=>"111111000",
  17967=>"111000000",
  17968=>"000111101",
  17969=>"111111111",
  17970=>"000011011",
  17971=>"000000000",
  17972=>"010001001",
  17973=>"111001000",
  17974=>"100001000",
  17975=>"000000100",
  17976=>"101111111",
  17977=>"000000000",
  17978=>"111000000",
  17979=>"111000000",
  17980=>"111001000",
  17981=>"100100000",
  17982=>"000100111",
  17983=>"000000000",
  17984=>"000000000",
  17985=>"000000011",
  17986=>"000000111",
  17987=>"000000111",
  17988=>"000110000",
  17989=>"000000000",
  17990=>"111000000",
  17991=>"111111011",
  17992=>"001001001",
  17993=>"111100100",
  17994=>"111111111",
  17995=>"111000001",
  17996=>"111111111",
  17997=>"000100110",
  17998=>"000000000",
  17999=>"111100111",
  18000=>"111000101",
  18001=>"111111000",
  18002=>"111000100",
  18003=>"111000001",
  18004=>"000100000",
  18005=>"000000010",
  18006=>"101000000",
  18007=>"000000000",
  18008=>"110110011",
  18009=>"111000000",
  18010=>"001000000",
  18011=>"000000100",
  18012=>"000101000",
  18013=>"001101111",
  18014=>"111111111",
  18015=>"101011011",
  18016=>"100101011",
  18017=>"000111111",
  18018=>"110110111",
  18019=>"000000111",
  18020=>"001111000",
  18021=>"000000000",
  18022=>"111000000",
  18023=>"000000111",
  18024=>"111000000",
  18025=>"111000111",
  18026=>"111000000",
  18027=>"110111110",
  18028=>"111001001",
  18029=>"101000000",
  18030=>"111101100",
  18031=>"111110010",
  18032=>"000000000",
  18033=>"000000000",
  18034=>"111111000",
  18035=>"100111111",
  18036=>"111100111",
  18037=>"000000100",
  18038=>"000000000",
  18039=>"001000101",
  18040=>"000011000",
  18041=>"110101000",
  18042=>"010011000",
  18043=>"111111111",
  18044=>"101111111",
  18045=>"001011111",
  18046=>"000000000",
  18047=>"001011111",
  18048=>"111010000",
  18049=>"000111010",
  18050=>"010000000",
  18051=>"111110000",
  18052=>"000000000",
  18053=>"000000011",
  18054=>"000111111",
  18055=>"001111011",
  18056=>"111111000",
  18057=>"100110110",
  18058=>"111100101",
  18059=>"111111111",
  18060=>"000000011",
  18061=>"000000000",
  18062=>"111000000",
  18063=>"111111000",
  18064=>"000000000",
  18065=>"111111000",
  18066=>"111111111",
  18067=>"000110111",
  18068=>"001111110",
  18069=>"011111111",
  18070=>"110000110",
  18071=>"111111000",
  18072=>"111000000",
  18073=>"001000000",
  18074=>"111001111",
  18075=>"001000000",
  18076=>"110100111",
  18077=>"001000000",
  18078=>"111011000",
  18079=>"000000000",
  18080=>"000010010",
  18081=>"000000011",
  18082=>"111000000",
  18083=>"111100111",
  18084=>"010111000",
  18085=>"111000000",
  18086=>"111000000",
  18087=>"111100100",
  18088=>"111100110",
  18089=>"110111111",
  18090=>"111111111",
  18091=>"011111011",
  18092=>"001011000",
  18093=>"000001000",
  18094=>"111111111",
  18095=>"111111000",
  18096=>"111000000",
  18097=>"111100111",
  18098=>"110101111",
  18099=>"000000111",
  18100=>"000011111",
  18101=>"111111001",
  18102=>"111000000",
  18103=>"111100000",
  18104=>"000001001",
  18105=>"111000111",
  18106=>"000000000",
  18107=>"101000111",
  18108=>"000000000",
  18109=>"100000111",
  18110=>"111000000",
  18111=>"000110111",
  18112=>"111001000",
  18113=>"000000000",
  18114=>"000110000",
  18115=>"000000000",
  18116=>"001000000",
  18117=>"000000000",
  18118=>"000000000",
  18119=>"000111111",
  18120=>"000111111",
  18121=>"001000000",
  18122=>"000111111",
  18123=>"111011111",
  18124=>"000000001",
  18125=>"000000111",
  18126=>"110111111",
  18127=>"011111111",
  18128=>"111111111",
  18129=>"000111111",
  18130=>"000010000",
  18131=>"000000000",
  18132=>"111011110",
  18133=>"000111001",
  18134=>"111010010",
  18135=>"111111000",
  18136=>"011111111",
  18137=>"101001000",
  18138=>"111001000",
  18139=>"111000000",
  18140=>"100000000",
  18141=>"111000000",
  18142=>"111111111",
  18143=>"000000000",
  18144=>"000000001",
  18145=>"000000000",
  18146=>"010111000",
  18147=>"111111001",
  18148=>"000011111",
  18149=>"000000011",
  18150=>"111000101",
  18151=>"101111011",
  18152=>"111111111",
  18153=>"101000011",
  18154=>"111110000",
  18155=>"001111111",
  18156=>"111111000",
  18157=>"111111000",
  18158=>"100110010",
  18159=>"111110110",
  18160=>"000000111",
  18161=>"110000000",
  18162=>"100111111",
  18163=>"011111000",
  18164=>"000000000",
  18165=>"111110110",
  18166=>"000111011",
  18167=>"000000000",
  18168=>"100000001",
  18169=>"011000000",
  18170=>"111111011",
  18171=>"000011000",
  18172=>"000011001",
  18173=>"111000100",
  18174=>"111000001",
  18175=>"110100000",
  18176=>"111111000",
  18177=>"111111100",
  18178=>"000000000",
  18179=>"111110100",
  18180=>"000000000",
  18181=>"111000000",
  18182=>"011000000",
  18183=>"000000111",
  18184=>"111010000",
  18185=>"000000000",
  18186=>"111111111",
  18187=>"111000000",
  18188=>"111111101",
  18189=>"010011011",
  18190=>"000111110",
  18191=>"110110111",
  18192=>"100000000",
  18193=>"000111111",
  18194=>"111111111",
  18195=>"011111111",
  18196=>"001111000",
  18197=>"100111000",
  18198=>"000000000",
  18199=>"111111100",
  18200=>"111111111",
  18201=>"111110100",
  18202=>"111111100",
  18203=>"000000000",
  18204=>"110000000",
  18205=>"000000000",
  18206=>"000000111",
  18207=>"011011000",
  18208=>"111111011",
  18209=>"111111000",
  18210=>"000110111",
  18211=>"111111111",
  18212=>"000000100",
  18213=>"000111111",
  18214=>"110111000",
  18215=>"111111011",
  18216=>"101000000",
  18217=>"101100001",
  18218=>"111010011",
  18219=>"000000000",
  18220=>"111000111",
  18221=>"000001000",
  18222=>"111010110",
  18223=>"111001111",
  18224=>"011110111",
  18225=>"011111111",
  18226=>"000000111",
  18227=>"111000000",
  18228=>"111111111",
  18229=>"000100110",
  18230=>"000000000",
  18231=>"100100100",
  18232=>"000111000",
  18233=>"111111111",
  18234=>"000000011",
  18235=>"110100111",
  18236=>"001111111",
  18237=>"110000001",
  18238=>"000001111",
  18239=>"100000000",
  18240=>"000010111",
  18241=>"101110111",
  18242=>"111000000",
  18243=>"000111110",
  18244=>"011000000",
  18245=>"111001000",
  18246=>"000001101",
  18247=>"110000001",
  18248=>"111100000",
  18249=>"000111111",
  18250=>"000000000",
  18251=>"000111111",
  18252=>"000110110",
  18253=>"111000111",
  18254=>"111001000",
  18255=>"100000000",
  18256=>"111011001",
  18257=>"101101111",
  18258=>"000000000",
  18259=>"000000000",
  18260=>"001000000",
  18261=>"000111111",
  18262=>"000011001",
  18263=>"000000110",
  18264=>"111111111",
  18265=>"000000000",
  18266=>"111111111",
  18267=>"000000000",
  18268=>"110000000",
  18269=>"011001000",
  18270=>"111001000",
  18271=>"001101111",
  18272=>"000000111",
  18273=>"000111101",
  18274=>"101111111",
  18275=>"111111000",
  18276=>"000100001",
  18277=>"000001111",
  18278=>"000000000",
  18279=>"001000000",
  18280=>"001111100",
  18281=>"000010011",
  18282=>"000000001",
  18283=>"011000000",
  18284=>"111011000",
  18285=>"000111100",
  18286=>"111000000",
  18287=>"101001111",
  18288=>"000111010",
  18289=>"000011111",
  18290=>"110100111",
  18291=>"111101111",
  18292=>"100000111",
  18293=>"000001111",
  18294=>"111000000",
  18295=>"001000000",
  18296=>"111110111",
  18297=>"000000001",
  18298=>"000111111",
  18299=>"000000011",
  18300=>"111111111",
  18301=>"011111111",
  18302=>"111111000",
  18303=>"100100111",
  18304=>"111111111",
  18305=>"111011001",
  18306=>"001000001",
  18307=>"000000111",
  18308=>"111000001",
  18309=>"110010000",
  18310=>"000000111",
  18311=>"000000111",
  18312=>"111000000",
  18313=>"000000000",
  18314=>"110000100",
  18315=>"111111000",
  18316=>"111111011",
  18317=>"111110100",
  18318=>"111111000",
  18319=>"001000001",
  18320=>"000000010",
  18321=>"100111111",
  18322=>"111011001",
  18323=>"000111100",
  18324=>"000111111",
  18325=>"000000000",
  18326=>"001001011",
  18327=>"011111001",
  18328=>"111111111",
  18329=>"000000111",
  18330=>"111000000",
  18331=>"000000000",
  18332=>"000000111",
  18333=>"000000000",
  18334=>"001000111",
  18335=>"000001011",
  18336=>"010111111",
  18337=>"011000000",
  18338=>"101000000",
  18339=>"111000000",
  18340=>"111011000",
  18341=>"011000101",
  18342=>"110000111",
  18343=>"000110111",
  18344=>"100111111",
  18345=>"101000000",
  18346=>"111111111",
  18347=>"000000000",
  18348=>"000000000",
  18349=>"111000000",
  18350=>"100000000",
  18351=>"101111111",
  18352=>"000000000",
  18353=>"000000000",
  18354=>"000000000",
  18355=>"001000000",
  18356=>"000010110",
  18357=>"011000111",
  18358=>"000011111",
  18359=>"001000011",
  18360=>"100111111",
  18361=>"101111111",
  18362=>"110111111",
  18363=>"111011111",
  18364=>"000100010",
  18365=>"111111000",
  18366=>"111001000",
  18367=>"100100100",
  18368=>"111000100",
  18369=>"000000111",
  18370=>"111000000",
  18371=>"111111111",
  18372=>"111000000",
  18373=>"111000000",
  18374=>"000000001",
  18375=>"000111011",
  18376=>"111111000",
  18377=>"111101000",
  18378=>"101000100",
  18379=>"000000000",
  18380=>"111111100",
  18381=>"011001001",
  18382=>"010011000",
  18383=>"111110000",
  18384=>"110000000",
  18385=>"101001101",
  18386=>"110111111",
  18387=>"000000111",
  18388=>"000000000",
  18389=>"111111101",
  18390=>"111000000",
  18391=>"111111110",
  18392=>"111000000",
  18393=>"101000000",
  18394=>"101101000",
  18395=>"111111111",
  18396=>"000000110",
  18397=>"111111000",
  18398=>"100000000",
  18399=>"000000000",
  18400=>"000000000",
  18401=>"000010111",
  18402=>"111100110",
  18403=>"111000111",
  18404=>"011001000",
  18405=>"111000111",
  18406=>"111111101",
  18407=>"100000000",
  18408=>"000111111",
  18409=>"100110111",
  18410=>"010000000",
  18411=>"111111100",
  18412=>"000000000",
  18413=>"000001000",
  18414=>"111111000",
  18415=>"000000011",
  18416=>"001111111",
  18417=>"000010001",
  18418=>"111111111",
  18419=>"000000000",
  18420=>"111110000",
  18421=>"011000001",
  18422=>"000000000",
  18423=>"110110111",
  18424=>"000000111",
  18425=>"111001000",
  18426=>"000000000",
  18427=>"011000000",
  18428=>"000000000",
  18429=>"000111111",
  18430=>"100000000",
  18431=>"111001111",
  18432=>"111111111",
  18433=>"011011011",
  18434=>"110000000",
  18435=>"111000000",
  18436=>"111111001",
  18437=>"100100111",
  18438=>"111111000",
  18439=>"000000111",
  18440=>"000000000",
  18441=>"100000000",
  18442=>"111111111",
  18443=>"111100010",
  18444=>"011011011",
  18445=>"001000000",
  18446=>"100000000",
  18447=>"111111111",
  18448=>"000000000",
  18449=>"101111111",
  18450=>"111111111",
  18451=>"111110111",
  18452=>"000000000",
  18453=>"101101111",
  18454=>"000000000",
  18455=>"101101111",
  18456=>"111111111",
  18457=>"111100111",
  18458=>"000000000",
  18459=>"111111011",
  18460=>"000001111",
  18461=>"111111111",
  18462=>"000011111",
  18463=>"011111111",
  18464=>"000000101",
  18465=>"111110000",
  18466=>"001011111",
  18467=>"000000000",
  18468=>"000000000",
  18469=>"111111000",
  18470=>"001000000",
  18471=>"111001000",
  18472=>"001001111",
  18473=>"011001001",
  18474=>"101000000",
  18475=>"100000100",
  18476=>"000000000",
  18477=>"000110111",
  18478=>"100110111",
  18479=>"111110000",
  18480=>"011111000",
  18481=>"100100110",
  18482=>"000000100",
  18483=>"111000000",
  18484=>"110110000",
  18485=>"110111000",
  18486=>"011001001",
  18487=>"000010101",
  18488=>"000000000",
  18489=>"000000111",
  18490=>"101111111",
  18491=>"110110110",
  18492=>"111111000",
  18493=>"001000001",
  18494=>"000000000",
  18495=>"111001000",
  18496=>"001001111",
  18497=>"000000000",
  18498=>"000000110",
  18499=>"111111111",
  18500=>"001111111",
  18501=>"000100100",
  18502=>"111101000",
  18503=>"000000000",
  18504=>"100100101",
  18505=>"111000000",
  18506=>"111111111",
  18507=>"000000000",
  18508=>"010110010",
  18509=>"110100000",
  18510=>"010000000",
  18511=>"111001000",
  18512=>"010110000",
  18513=>"000000000",
  18514=>"000000110",
  18515=>"111111001",
  18516=>"111100100",
  18517=>"000000000",
  18518=>"000000000",
  18519=>"001000000",
  18520=>"001000000",
  18521=>"111000111",
  18522=>"100000100",
  18523=>"010000000",
  18524=>"000000000",
  18525=>"000000000",
  18526=>"111011111",
  18527=>"111111111",
  18528=>"111001011",
  18529=>"000000000",
  18530=>"111101111",
  18531=>"000000000",
  18532=>"001000000",
  18533=>"011011000",
  18534=>"100110011",
  18535=>"001100111",
  18536=>"111000000",
  18537=>"000000000",
  18538=>"111001001",
  18539=>"000110110",
  18540=>"000000000",
  18541=>"111111111",
  18542=>"011000001",
  18543=>"000000000",
  18544=>"111111111",
  18545=>"111110000",
  18546=>"110110000",
  18547=>"111001000",
  18548=>"111111111",
  18549=>"011011011",
  18550=>"100100000",
  18551=>"000000111",
  18552=>"001001001",
  18553=>"110111111",
  18554=>"000000000",
  18555=>"111100000",
  18556=>"000110110",
  18557=>"010111111",
  18558=>"000000000",
  18559=>"000101111",
  18560=>"111111111",
  18561=>"000000000",
  18562=>"110000000",
  18563=>"110111011",
  18564=>"111110100",
  18565=>"111110110",
  18566=>"111010000",
  18567=>"110000000",
  18568=>"101000000",
  18569=>"000000111",
  18570=>"101100000",
  18571=>"000000111",
  18572=>"000000000",
  18573=>"111100011",
  18574=>"000000000",
  18575=>"000000000",
  18576=>"100100111",
  18577=>"100000001",
  18578=>"111110111",
  18579=>"100110111",
  18580=>"000000100",
  18581=>"000000111",
  18582=>"000000111",
  18583=>"111000000",
  18584=>"011100100",
  18585=>"111110111",
  18586=>"011110111",
  18587=>"010000001",
  18588=>"111001111",
  18589=>"001000001",
  18590=>"111111000",
  18591=>"000110111",
  18592=>"000000000",
  18593=>"010010010",
  18594=>"111111111",
  18595=>"001011111",
  18596=>"000000000",
  18597=>"011001000",
  18598=>"111000000",
  18599=>"010010000",
  18600=>"000000010",
  18601=>"111111111",
  18602=>"000100111",
  18603=>"111111000",
  18604=>"001100110",
  18605=>"000000000",
  18606=>"111111111",
  18607=>"111111111",
  18608=>"011111111",
  18609=>"111111111",
  18610=>"000010000",
  18611=>"110000000",
  18612=>"010110100",
  18613=>"000110000",
  18614=>"111111111",
  18615=>"000000000",
  18616=>"000000000",
  18617=>"000000000",
  18618=>"000000000",
  18619=>"011010000",
  18620=>"110100100",
  18621=>"111111111",
  18622=>"000000000",
  18623=>"111110110",
  18624=>"000000000",
  18625=>"111111101",
  18626=>"000000000",
  18627=>"000110111",
  18628=>"111111000",
  18629=>"010000000",
  18630=>"000000000",
  18631=>"011110000",
  18632=>"000000000",
  18633=>"000000100",
  18634=>"111111111",
  18635=>"110110100",
  18636=>"111011111",
  18637=>"111111111",
  18638=>"000000000",
  18639=>"110000000",
  18640=>"000010111",
  18641=>"000000011",
  18642=>"000000110",
  18643=>"000000111",
  18644=>"111111111",
  18645=>"111111111",
  18646=>"000000000",
  18647=>"111110111",
  18648=>"000000111",
  18649=>"110000001",
  18650=>"000000001",
  18651=>"001000111",
  18652=>"011000000",
  18653=>"111011111",
  18654=>"011011000",
  18655=>"001100110",
  18656=>"000000000",
  18657=>"111000000",
  18658=>"000000100",
  18659=>"111111110",
  18660=>"111111011",
  18661=>"111110110",
  18662=>"000000110",
  18663=>"011011111",
  18664=>"101000001",
  18665=>"000000000",
  18666=>"111111101",
  18667=>"000000101",
  18668=>"100011111",
  18669=>"100000000",
  18670=>"000001011",
  18671=>"111111000",
  18672=>"100000000",
  18673=>"000000000",
  18674=>"111111111",
  18675=>"000111001",
  18676=>"111000111",
  18677=>"100000001",
  18678=>"111111111",
  18679=>"001000000",
  18680=>"100101111",
  18681=>"000000000",
  18682=>"111111111",
  18683=>"011011111",
  18684=>"001111111",
  18685=>"010011011",
  18686=>"011000000",
  18687=>"001001111",
  18688=>"011011011",
  18689=>"011010010",
  18690=>"001000000",
  18691=>"111011000",
  18692=>"001100000",
  18693=>"000000000",
  18694=>"100100100",
  18695=>"000000000",
  18696=>"111110000",
  18697=>"001000000",
  18698=>"000000000",
  18699=>"000000000",
  18700=>"000000000",
  18701=>"000000000",
  18702=>"111111110",
  18703=>"111001000",
  18704=>"011111111",
  18705=>"000011110",
  18706=>"000000000",
  18707=>"000000100",
  18708=>"000000000",
  18709=>"111111111",
  18710=>"010010001",
  18711=>"000000000",
  18712=>"000000001",
  18713=>"000000000",
  18714=>"100000001",
  18715=>"011001111",
  18716=>"000000111",
  18717=>"000000000",
  18718=>"000000000",
  18719=>"100000001",
  18720=>"001001001",
  18721=>"111000000",
  18722=>"111110110",
  18723=>"111111111",
  18724=>"111011011",
  18725=>"011000000",
  18726=>"101101100",
  18727=>"000000000",
  18728=>"001011011",
  18729=>"111101111",
  18730=>"100000000",
  18731=>"111111000",
  18732=>"111111001",
  18733=>"000000010",
  18734=>"000000000",
  18735=>"111111111",
  18736=>"111111111",
  18737=>"111111111",
  18738=>"001000000",
  18739=>"000000000",
  18740=>"000000000",
  18741=>"111111111",
  18742=>"000000100",
  18743=>"001000000",
  18744=>"100000000",
  18745=>"101100100",
  18746=>"000001001",
  18747=>"000000110",
  18748=>"010000010",
  18749=>"111111011",
  18750=>"000000000",
  18751=>"111111001",
  18752=>"000000000",
  18753=>"111111011",
  18754=>"111111110",
  18755=>"111111111",
  18756=>"000001011",
  18757=>"000000110",
  18758=>"000000000",
  18759=>"000000000",
  18760=>"000000000",
  18761=>"010010000",
  18762=>"111111111",
  18763=>"100110100",
  18764=>"011011011",
  18765=>"000000110",
  18766=>"010011011",
  18767=>"000100101",
  18768=>"000100100",
  18769=>"011111111",
  18770=>"000000011",
  18771=>"000111111",
  18772=>"100000000",
  18773=>"111111111",
  18774=>"011010111",
  18775=>"000000100",
  18776=>"000000000",
  18777=>"000000000",
  18778=>"111111111",
  18779=>"000000000",
  18780=>"000000000",
  18781=>"101000011",
  18782=>"111110000",
  18783=>"111111111",
  18784=>"000000110",
  18785=>"000000111",
  18786=>"011011111",
  18787=>"000000000",
  18788=>"001111111",
  18789=>"000000001",
  18790=>"000000000",
  18791=>"000000000",
  18792=>"000010010",
  18793=>"110110110",
  18794=>"011111111",
  18795=>"111111111",
  18796=>"011011011",
  18797=>"000010111",
  18798=>"000000000",
  18799=>"000011001",
  18800=>"011011000",
  18801=>"000111111",
  18802=>"111000000",
  18803=>"111111111",
  18804=>"100100100",
  18805=>"001001000",
  18806=>"000000000",
  18807=>"000000100",
  18808=>"000000000",
  18809=>"000101011",
  18810=>"000000000",
  18811=>"000000110",
  18812=>"111011011",
  18813=>"000111111",
  18814=>"000000001",
  18815=>"111011001",
  18816=>"011011011",
  18817=>"111111111",
  18818=>"111101001",
  18819=>"100100000",
  18820=>"111111111",
  18821=>"011011111",
  18822=>"000001000",
  18823=>"001111111",
  18824=>"111000000",
  18825=>"000000000",
  18826=>"001000100",
  18827=>"100101110",
  18828=>"111011001",
  18829=>"000010010",
  18830=>"011000000",
  18831=>"011011111",
  18832=>"000000000",
  18833=>"000000000",
  18834=>"111111111",
  18835=>"100000000",
  18836=>"111101110",
  18837=>"001000100",
  18838=>"001011000",
  18839=>"000000000",
  18840=>"000000000",
  18841=>"001001011",
  18842=>"111111111",
  18843=>"000010011",
  18844=>"100000011",
  18845=>"100000001",
  18846=>"101000100",
  18847=>"000000010",
  18848=>"001100111",
  18849=>"011011110",
  18850=>"111101000",
  18851=>"100100000",
  18852=>"111001000",
  18853=>"010111110",
  18854=>"111011000",
  18855=>"111111111",
  18856=>"001000110",
  18857=>"111111111",
  18858=>"111100111",
  18859=>"100100000",
  18860=>"000001000",
  18861=>"111111111",
  18862=>"011001000",
  18863=>"000000111",
  18864=>"111111111",
  18865=>"110111111",
  18866=>"000000000",
  18867=>"111100110",
  18868=>"000000100",
  18869=>"000000000",
  18870=>"011011001",
  18871=>"000000000",
  18872=>"111111000",
  18873=>"000010111",
  18874=>"111011001",
  18875=>"111111111",
  18876=>"111111111",
  18877=>"001000001",
  18878=>"000100111",
  18879=>"000000010",
  18880=>"111111111",
  18881=>"100000111",
  18882=>"000000000",
  18883=>"000000111",
  18884=>"111111111",
  18885=>"101111111",
  18886=>"000000000",
  18887=>"011001111",
  18888=>"000000000",
  18889=>"000000100",
  18890=>"100000110",
  18891=>"000000100",
  18892=>"111111000",
  18893=>"111011000",
  18894=>"111001001",
  18895=>"010111011",
  18896=>"010110110",
  18897=>"111111111",
  18898=>"110011001",
  18899=>"000000000",
  18900=>"111110111",
  18901=>"111110111",
  18902=>"001000110",
  18903=>"100110110",
  18904=>"100000111",
  18905=>"001000000",
  18906=>"111111001",
  18907=>"111111111",
  18908=>"111111111",
  18909=>"111111110",
  18910=>"110111001",
  18911=>"001011111",
  18912=>"000111111",
  18913=>"001000000",
  18914=>"111001000",
  18915=>"000000111",
  18916=>"101100111",
  18917=>"000000100",
  18918=>"111111111",
  18919=>"110110100",
  18920=>"000000101",
  18921=>"111111111",
  18922=>"000000111",
  18923=>"000000000",
  18924=>"111001001",
  18925=>"000000000",
  18926=>"111011011",
  18927=>"111100111",
  18928=>"100110111",
  18929=>"010111111",
  18930=>"000011111",
  18931=>"000000000",
  18932=>"111111001",
  18933=>"101001010",
  18934=>"001111111",
  18935=>"111100110",
  18936=>"111111111",
  18937=>"000000110",
  18938=>"000000111",
  18939=>"111000000",
  18940=>"111100001",
  18941=>"011111001",
  18942=>"000001011",
  18943=>"000000001",
  18944=>"100100100",
  18945=>"000000000",
  18946=>"111100111",
  18947=>"101101111",
  18948=>"000000000",
  18949=>"000000101",
  18950=>"111111111",
  18951=>"101100111",
  18952=>"100000000",
  18953=>"101001001",
  18954=>"001000000",
  18955=>"111011000",
  18956=>"011010000",
  18957=>"101100100",
  18958=>"000011111",
  18959=>"010110111",
  18960=>"001001000",
  18961=>"010000000",
  18962=>"111011111",
  18963=>"011111111",
  18964=>"100000000",
  18965=>"111010000",
  18966=>"111000001",
  18967=>"000000000",
  18968=>"000000111",
  18969=>"011110100",
  18970=>"111001000",
  18971=>"111010111",
  18972=>"000000000",
  18973=>"010000000",
  18974=>"111111111",
  18975=>"111111000",
  18976=>"111111111",
  18977=>"110110110",
  18978=>"110110110",
  18979=>"000000000",
  18980=>"000000000",
  18981=>"101001001",
  18982=>"111111111",
  18983=>"111101101",
  18984=>"000000000",
  18985=>"111111100",
  18986=>"000000101",
  18987=>"000111111",
  18988=>"010111111",
  18989=>"111111111",
  18990=>"000000101",
  18991=>"111111111",
  18992=>"000000001",
  18993=>"111111111",
  18994=>"000100000",
  18995=>"000011010",
  18996=>"111111111",
  18997=>"111011111",
  18998=>"111000000",
  18999=>"110110110",
  19000=>"000100101",
  19001=>"110111111",
  19002=>"111111111",
  19003=>"111111110",
  19004=>"001001001",
  19005=>"010110010",
  19006=>"001011011",
  19007=>"000000000",
  19008=>"000000000",
  19009=>"100000000",
  19010=>"011001000",
  19011=>"100001101",
  19012=>"111010000",
  19013=>"011111111",
  19014=>"000000000",
  19015=>"111000000",
  19016=>"110110000",
  19017=>"000111111",
  19018=>"000000001",
  19019=>"001111001",
  19020=>"000000111",
  19021=>"111001001",
  19022=>"101111111",
  19023=>"000000000",
  19024=>"110110010",
  19025=>"100001111",
  19026=>"000000000",
  19027=>"110100001",
  19028=>"000000000",
  19029=>"101101111",
  19030=>"111000011",
  19031=>"111111110",
  19032=>"111111011",
  19033=>"111101111",
  19034=>"000000000",
  19035=>"000000000",
  19036=>"000011111",
  19037=>"000000000",
  19038=>"000000001",
  19039=>"111011001",
  19040=>"011111111",
  19041=>"010110010",
  19042=>"000000000",
  19043=>"100110111",
  19044=>"000000010",
  19045=>"000100100",
  19046=>"000100111",
  19047=>"101101101",
  19048=>"111111010",
  19049=>"100000001",
  19050=>"110111111",
  19051=>"110011000",
  19052=>"100010010",
  19053=>"111111111",
  19054=>"000000000",
  19055=>"000001001",
  19056=>"000100000",
  19057=>"000001001",
  19058=>"001101111",
  19059=>"000000100",
  19060=>"000000000",
  19061=>"111111111",
  19062=>"000000000",
  19063=>"011001101",
  19064=>"000001001",
  19065=>"001011011",
  19066=>"000000000",
  19067=>"000001111",
  19068=>"000000000",
  19069=>"000000000",
  19070=>"000000000",
  19071=>"000000000",
  19072=>"111111111",
  19073=>"110000000",
  19074=>"111111111",
  19075=>"011010011",
  19076=>"110000111",
  19077=>"000000001",
  19078=>"000000001",
  19079=>"111110110",
  19080=>"111111111",
  19081=>"000000000",
  19082=>"001001001",
  19083=>"000000100",
  19084=>"000000000",
  19085=>"111111111",
  19086=>"110000000",
  19087=>"111111111",
  19088=>"000000000",
  19089=>"001001001",
  19090=>"011111000",
  19091=>"001011111",
  19092=>"000000111",
  19093=>"100000000",
  19094=>"111111110",
  19095=>"111101100",
  19096=>"000000101",
  19097=>"111111111",
  19098=>"111111111",
  19099=>"000000000",
  19100=>"111100010",
  19101=>"001000111",
  19102=>"000000010",
  19103=>"110110010",
  19104=>"101000001",
  19105=>"001010000",
  19106=>"111111111",
  19107=>"100101101",
  19108=>"001001101",
  19109=>"111111111",
  19110=>"100000000",
  19111=>"000111111",
  19112=>"100101000",
  19113=>"000000101",
  19114=>"000001101",
  19115=>"000000000",
  19116=>"001100110",
  19117=>"100000000",
  19118=>"000000001",
  19119=>"000000001",
  19120=>"011111111",
  19121=>"111100001",
  19122=>"111111110",
  19123=>"111101001",
  19124=>"100000000",
  19125=>"000010000",
  19126=>"011010111",
  19127=>"000000101",
  19128=>"111111111",
  19129=>"111111111",
  19130=>"001001001",
  19131=>"111110000",
  19132=>"000000000",
  19133=>"111111010",
  19134=>"000000011",
  19135=>"000000000",
  19136=>"111101111",
  19137=>"011111111",
  19138=>"111111110",
  19139=>"000000000",
  19140=>"000000111",
  19141=>"000000011",
  19142=>"000000111",
  19143=>"100100000",
  19144=>"111111000",
  19145=>"010000000",
  19146=>"000000000",
  19147=>"101000001",
  19148=>"010110100",
  19149=>"111011110",
  19150=>"111111111",
  19151=>"000111101",
  19152=>"000001000",
  19153=>"111001011",
  19154=>"000000001",
  19155=>"000000000",
  19156=>"000000101",
  19157=>"000000000",
  19158=>"000001001",
  19159=>"000000000",
  19160=>"110100110",
  19161=>"010110010",
  19162=>"111111111",
  19163=>"111111111",
  19164=>"111111000",
  19165=>"111100101",
  19166=>"000111111",
  19167=>"110110000",
  19168=>"000001001",
  19169=>"000000000",
  19170=>"000000000",
  19171=>"111111010",
  19172=>"000000000",
  19173=>"000000000",
  19174=>"001000110",
  19175=>"000000001",
  19176=>"011011011",
  19177=>"001011010",
  19178=>"010111111",
  19179=>"000000000",
  19180=>"101001011",
  19181=>"000000111",
  19182=>"001111111",
  19183=>"111111111",
  19184=>"000000000",
  19185=>"111000000",
  19186=>"100111101",
  19187=>"101000000",
  19188=>"111111111",
  19189=>"111110000",
  19190=>"000000000",
  19191=>"111111111",
  19192=>"000011101",
  19193=>"000000000",
  19194=>"000010010",
  19195=>"001001000",
  19196=>"001000001",
  19197=>"000000000",
  19198=>"111111000",
  19199=>"111111111",
  19200=>"000000000",
  19201=>"001011011",
  19202=>"000000110",
  19203=>"000101111",
  19204=>"010010000",
  19205=>"000011111",
  19206=>"111111111",
  19207=>"110111101",
  19208=>"100001111",
  19209=>"110110000",
  19210=>"000000000",
  19211=>"111111010",
  19212=>"111111110",
  19213=>"000000110",
  19214=>"101001111",
  19215=>"111000000",
  19216=>"000000000",
  19217=>"001001000",
  19218=>"000000001",
  19219=>"000111111",
  19220=>"100000000",
  19221=>"111111101",
  19222=>"101111011",
  19223=>"111110110",
  19224=>"000100111",
  19225=>"111111111",
  19226=>"000000000",
  19227=>"010010110",
  19228=>"011011011",
  19229=>"010111111",
  19230=>"000000000",
  19231=>"011111111",
  19232=>"011111000",
  19233=>"111111010",
  19234=>"111111001",
  19235=>"101000001",
  19236=>"011001001",
  19237=>"000000010",
  19238=>"111110110",
  19239=>"001000000",
  19240=>"000100100",
  19241=>"000000111",
  19242=>"010110110",
  19243=>"000000000",
  19244=>"000000011",
  19245=>"000110110",
  19246=>"111111110",
  19247=>"000000000",
  19248=>"110110000",
  19249=>"010100110",
  19250=>"000000001",
  19251=>"000000001",
  19252=>"110110000",
  19253=>"111001000",
  19254=>"000000001",
  19255=>"000000111",
  19256=>"111111010",
  19257=>"111111101",
  19258=>"000000001",
  19259=>"111000001",
  19260=>"000001000",
  19261=>"000010101",
  19262=>"101101101",
  19263=>"111001101",
  19264=>"011111000",
  19265=>"000001000",
  19266=>"000000001",
  19267=>"101001111",
  19268=>"111011011",
  19269=>"010000000",
  19270=>"000000000",
  19271=>"000000000",
  19272=>"000000101",
  19273=>"001000000",
  19274=>"000000000",
  19275=>"010000100",
  19276=>"100000000",
  19277=>"111111111",
  19278=>"111101111",
  19279=>"111111111",
  19280=>"111111111",
  19281=>"101001111",
  19282=>"111111101",
  19283=>"001000111",
  19284=>"000000000",
  19285=>"000011011",
  19286=>"110110000",
  19287=>"100101101",
  19288=>"111111010",
  19289=>"000000000",
  19290=>"110110000",
  19291=>"000000100",
  19292=>"000000000",
  19293=>"011111111",
  19294=>"111011001",
  19295=>"000000001",
  19296=>"000000001",
  19297=>"000000000",
  19298=>"011011011",
  19299=>"111111001",
  19300=>"111110110",
  19301=>"011011011",
  19302=>"110100111",
  19303=>"000000000",
  19304=>"000000001",
  19305=>"011001000",
  19306=>"000000100",
  19307=>"001000000",
  19308=>"100110110",
  19309=>"001001000",
  19310=>"111111111",
  19311=>"000111111",
  19312=>"101000000",
  19313=>"100101111",
  19314=>"000010111",
  19315=>"011011011",
  19316=>"110110000",
  19317=>"000110100",
  19318=>"000001001",
  19319=>"000000000",
  19320=>"100100100",
  19321=>"000000000",
  19322=>"101000000",
  19323=>"001001101",
  19324=>"110100000",
  19325=>"101101101",
  19326=>"000001101",
  19327=>"101101101",
  19328=>"110000001",
  19329=>"111111001",
  19330=>"111111110",
  19331=>"000000000",
  19332=>"000100111",
  19333=>"001101111",
  19334=>"011111111",
  19335=>"001000000",
  19336=>"001111111",
  19337=>"010111111",
  19338=>"100000010",
  19339=>"111111111",
  19340=>"100000111",
  19341=>"000000001",
  19342=>"111111111",
  19343=>"111111110",
  19344=>"000000000",
  19345=>"000000000",
  19346=>"111111111",
  19347=>"000100111",
  19348=>"111111111",
  19349=>"011001000",
  19350=>"000000110",
  19351=>"110000000",
  19352=>"101000000",
  19353=>"111110000",
  19354=>"111111111",
  19355=>"110110000",
  19356=>"100000000",
  19357=>"000000111",
  19358=>"101001101",
  19359=>"110110010",
  19360=>"100110010",
  19361=>"000101111",
  19362=>"110110000",
  19363=>"111101000",
  19364=>"110111101",
  19365=>"111101001",
  19366=>"100000000",
  19367=>"111000000",
  19368=>"001000100",
  19369=>"000000001",
  19370=>"110111111",
  19371=>"111111011",
  19372=>"000000000",
  19373=>"111001111",
  19374=>"111001000",
  19375=>"100100000",
  19376=>"000000000",
  19377=>"111111110",
  19378=>"011111111",
  19379=>"110111110",
  19380=>"000000000",
  19381=>"111111101",
  19382=>"000000001",
  19383=>"000000000",
  19384=>"110110111",
  19385=>"000011111",
  19386=>"011101001",
  19387=>"111111100",
  19388=>"001001000",
  19389=>"111011100",
  19390=>"101101010",
  19391=>"000000111",
  19392=>"000000000",
  19393=>"000010110",
  19394=>"000110110",
  19395=>"000110000",
  19396=>"010110111",
  19397=>"110000000",
  19398=>"000000000",
  19399=>"000000000",
  19400=>"001011111",
  19401=>"100111111",
  19402=>"111111000",
  19403=>"000000000",
  19404=>"011011000",
  19405=>"111110010",
  19406=>"100000101",
  19407=>"111100101",
  19408=>"101101001",
  19409=>"011011011",
  19410=>"111111111",
  19411=>"000000000",
  19412=>"000001000",
  19413=>"111111111",
  19414=>"011001001",
  19415=>"110111111",
  19416=>"111001001",
  19417=>"111000000",
  19418=>"111000000",
  19419=>"000000000",
  19420=>"111111110",
  19421=>"000000001",
  19422=>"000001011",
  19423=>"000111111",
  19424=>"111001000",
  19425=>"111000000",
  19426=>"101101111",
  19427=>"010000011",
  19428=>"110000000",
  19429=>"001001101",
  19430=>"011001111",
  19431=>"110000000",
  19432=>"110110110",
  19433=>"111001000",
  19434=>"000111111",
  19435=>"001110101",
  19436=>"100000001",
  19437=>"000001001",
  19438=>"000111111",
  19439=>"000010011",
  19440=>"000001000",
  19441=>"000111111",
  19442=>"000000000",
  19443=>"010110010",
  19444=>"111111110",
  19445=>"000000000",
  19446=>"111111000",
  19447=>"001111111",
  19448=>"000000000",
  19449=>"000000000",
  19450=>"010000000",
  19451=>"000000000",
  19452=>"100100111",
  19453=>"100100100",
  19454=>"111000000",
  19455=>"101001101",
  19456=>"111000000",
  19457=>"000000111",
  19458=>"111000000",
  19459=>"111111011",
  19460=>"000000110",
  19461=>"111000000",
  19462=>"000000000",
  19463=>"000001111",
  19464=>"011111100",
  19465=>"100111111",
  19466=>"000000000",
  19467=>"111111011",
  19468=>"000101001",
  19469=>"110100101",
  19470=>"101111111",
  19471=>"000000100",
  19472=>"111111001",
  19473=>"000000110",
  19474=>"110000000",
  19475=>"000000000",
  19476=>"011111111",
  19477=>"000000111",
  19478=>"011001001",
  19479=>"111111001",
  19480=>"111111000",
  19481=>"000001111",
  19482=>"100111111",
  19483=>"000101101",
  19484=>"000000000",
  19485=>"100100111",
  19486=>"111101000",
  19487=>"000001111",
  19488=>"111110000",
  19489=>"111111111",
  19490=>"111001101",
  19491=>"111100100",
  19492=>"000010011",
  19493=>"000111111",
  19494=>"000000111",
  19495=>"000111111",
  19496=>"001000000",
  19497=>"000110000",
  19498=>"000111111",
  19499=>"111111000",
  19500=>"100000000",
  19501=>"000111111",
  19502=>"001001001",
  19503=>"111111111",
  19504=>"000001001",
  19505=>"000000111",
  19506=>"000110110",
  19507=>"001001011",
  19508=>"111111001",
  19509=>"100100110",
  19510=>"101000000",
  19511=>"000100000",
  19512=>"000000100",
  19513=>"111111001",
  19514=>"001000001",
  19515=>"000111111",
  19516=>"110111111",
  19517=>"000010000",
  19518=>"011011011",
  19519=>"000000111",
  19520=>"000111111",
  19521=>"110110110",
  19522=>"000001001",
  19523=>"000000011",
  19524=>"001000100",
  19525=>"001011111",
  19526=>"111111001",
  19527=>"111111011",
  19528=>"100000000",
  19529=>"111000000",
  19530=>"111000110",
  19531=>"111110100",
  19532=>"000000000",
  19533=>"000000000",
  19534=>"001001111",
  19535=>"011111111",
  19536=>"000000000",
  19537=>"100111111",
  19538=>"111000101",
  19539=>"011111001",
  19540=>"000000000",
  19541=>"111111111",
  19542=>"111000100",
  19543=>"001111101",
  19544=>"111111111",
  19545=>"001001101",
  19546=>"111001000",
  19547=>"000001011",
  19548=>"000111000",
  19549=>"000100111",
  19550=>"000001111",
  19551=>"011000000",
  19552=>"000000000",
  19553=>"111000000",
  19554=>"111111111",
  19555=>"110111111",
  19556=>"111100110",
  19557=>"111010010",
  19558=>"111011101",
  19559=>"000101110",
  19560=>"110010001",
  19561=>"011011111",
  19562=>"111010000",
  19563=>"000000000",
  19564=>"111110110",
  19565=>"111000000",
  19566=>"011000000",
  19567=>"000000011",
  19568=>"000000111",
  19569=>"000000000",
  19570=>"111111000",
  19571=>"000000000",
  19572=>"100100000",
  19573=>"100100000",
  19574=>"111111111",
  19575=>"110110111",
  19576=>"000000000",
  19577=>"000000000",
  19578=>"000000001",
  19579=>"000111000",
  19580=>"111111110",
  19581=>"111001000",
  19582=>"000000000",
  19583=>"111111000",
  19584=>"000000111",
  19585=>"101000000",
  19586=>"111010000",
  19587=>"111111000",
  19588=>"000000111",
  19589=>"111100011",
  19590=>"111000000",
  19591=>"100110110",
  19592=>"111100001",
  19593=>"000011111",
  19594=>"000000000",
  19595=>"001000000",
  19596=>"111111001",
  19597=>"111111011",
  19598=>"001000111",
  19599=>"110111000",
  19600=>"111111000",
  19601=>"000000000",
  19602=>"000001001",
  19603=>"001111110",
  19604=>"110000000",
  19605=>"100110000",
  19606=>"000100111",
  19607=>"111111111",
  19608=>"110111111",
  19609=>"001111001",
  19610=>"111111111",
  19611=>"000000000",
  19612=>"111111111",
  19613=>"000000001",
  19614=>"111111011",
  19615=>"111111010",
  19616=>"111110100",
  19617=>"011001000",
  19618=>"000000001",
  19619=>"000000000",
  19620=>"000000000",
  19621=>"000111111",
  19622=>"111111010",
  19623=>"101101011",
  19624=>"111110100",
  19625=>"000000100",
  19626=>"001011000",
  19627=>"111111111",
  19628=>"000000000",
  19629=>"111100111",
  19630=>"111011111",
  19631=>"000000111",
  19632=>"000011001",
  19633=>"000100110",
  19634=>"111111010",
  19635=>"011111000",
  19636=>"110111111",
  19637=>"111111001",
  19638=>"111000111",
  19639=>"111010000",
  19640=>"111111111",
  19641=>"110111111",
  19642=>"000000000",
  19643=>"000000101",
  19644=>"000000110",
  19645=>"111011000",
  19646=>"000000000",
  19647=>"010110010",
  19648=>"000111111",
  19649=>"100111111",
  19650=>"111011001",
  19651=>"000111111",
  19652=>"000011111",
  19653=>"010111111",
  19654=>"010110111",
  19655=>"110110110",
  19656=>"111111110",
  19657=>"111110110",
  19658=>"100000111",
  19659=>"000000000",
  19660=>"111111111",
  19661=>"000100111",
  19662=>"000010111",
  19663=>"111111110",
  19664=>"110111111",
  19665=>"100111000",
  19666=>"111111110",
  19667=>"111010000",
  19668=>"000000111",
  19669=>"011011010",
  19670=>"000001111",
  19671=>"100100111",
  19672=>"111110000",
  19673=>"000000001",
  19674=>"000000101",
  19675=>"000100111",
  19676=>"111000000",
  19677=>"000000101",
  19678=>"000111000",
  19679=>"111111000",
  19680=>"000000000",
  19681=>"000111111",
  19682=>"000111111",
  19683=>"000000000",
  19684=>"000011111",
  19685=>"100100110",
  19686=>"111001011",
  19687=>"111001000",
  19688=>"000000000",
  19689=>"110111111",
  19690=>"111111111",
  19691=>"011010110",
  19692=>"111011001",
  19693=>"001000001",
  19694=>"010111001",
  19695=>"011000110",
  19696=>"000000000",
  19697=>"110000000",
  19698=>"111111111",
  19699=>"000001011",
  19700=>"000000000",
  19701=>"111111000",
  19702=>"100111000",
  19703=>"111000000",
  19704=>"111001000",
  19705=>"000000000",
  19706=>"000000000",
  19707=>"000000000",
  19708=>"011011111",
  19709=>"011000000",
  19710=>"000000000",
  19711=>"111101100",
  19712=>"000000111",
  19713=>"011111111",
  19714=>"111111111",
  19715=>"000000000",
  19716=>"001001100",
  19717=>"110000000",
  19718=>"000000111",
  19719=>"111010111",
  19720=>"111111110",
  19721=>"000111111",
  19722=>"111000111",
  19723=>"111111111",
  19724=>"101001001",
  19725=>"111001000",
  19726=>"111110100",
  19727=>"111111111",
  19728=>"000000000",
  19729=>"000000001",
  19730=>"111001001",
  19731=>"100100000",
  19732=>"001001000",
  19733=>"111111000",
  19734=>"111111001",
  19735=>"111111111",
  19736=>"011011111",
  19737=>"111000000",
  19738=>"111111000",
  19739=>"111110100",
  19740=>"000001101",
  19741=>"000000000",
  19742=>"001000000",
  19743=>"000111000",
  19744=>"101101111",
  19745=>"000011011",
  19746=>"000000011",
  19747=>"000111111",
  19748=>"000000000",
  19749=>"001011111",
  19750=>"100111000",
  19751=>"111111111",
  19752=>"111111111",
  19753=>"000111111",
  19754=>"000000000",
  19755=>"000000000",
  19756=>"001000111",
  19757=>"000110111",
  19758=>"000000111",
  19759=>"110000110",
  19760=>"000000000",
  19761=>"000000000",
  19762=>"110110000",
  19763=>"000000011",
  19764=>"111101011",
  19765=>"111111000",
  19766=>"110110100",
  19767=>"111111001",
  19768=>"010001000",
  19769=>"111111101",
  19770=>"111111000",
  19771=>"010000000",
  19772=>"111111000",
  19773=>"100001101",
  19774=>"000010010",
  19775=>"000000100",
  19776=>"000000111",
  19777=>"111111010",
  19778=>"000000000",
  19779=>"111001000",
  19780=>"000000000",
  19781=>"101101111",
  19782=>"000111000",
  19783=>"001011001",
  19784=>"000000000",
  19785=>"000000000",
  19786=>"111111001",
  19787=>"000000110",
  19788=>"000000000",
  19789=>"000000000",
  19790=>"110111111",
  19791=>"100111111",
  19792=>"000000000",
  19793=>"111110000",
  19794=>"110110111",
  19795=>"000000000",
  19796=>"001000000",
  19797=>"011011011",
  19798=>"000111111",
  19799=>"111111111",
  19800=>"111101111",
  19801=>"111111111",
  19802=>"111000000",
  19803=>"000000111",
  19804=>"000111110",
  19805=>"110011001",
  19806=>"011011000",
  19807=>"100111111",
  19808=>"111111000",
  19809=>"000000000",
  19810=>"111011011",
  19811=>"001001011",
  19812=>"100101000",
  19813=>"000110000",
  19814=>"000111111",
  19815=>"111111000",
  19816=>"000001111",
  19817=>"000001000",
  19818=>"000111110",
  19819=>"001011011",
  19820=>"000111100",
  19821=>"111000000",
  19822=>"111111111",
  19823=>"000000000",
  19824=>"000000000",
  19825=>"000010000",
  19826=>"100111111",
  19827=>"100100110",
  19828=>"000000000",
  19829=>"111111111",
  19830=>"000000000",
  19831=>"110111111",
  19832=>"000000101",
  19833=>"000000010",
  19834=>"000010100",
  19835=>"111110000",
  19836=>"111111111",
  19837=>"000000111",
  19838=>"111111000",
  19839=>"000111111",
  19840=>"000011000",
  19841=>"110110111",
  19842=>"000001111",
  19843=>"000111000",
  19844=>"001111111",
  19845=>"001000011",
  19846=>"111111110",
  19847=>"111111111",
  19848=>"000000000",
  19849=>"001011011",
  19850=>"110111111",
  19851=>"111011000",
  19852=>"111100111",
  19853=>"111111001",
  19854=>"111000000",
  19855=>"000000110",
  19856=>"000000000",
  19857=>"000000111",
  19858=>"110010011",
  19859=>"111111100",
  19860=>"111111111",
  19861=>"010010011",
  19862=>"000110110",
  19863=>"001000000",
  19864=>"000000000",
  19865=>"000000111",
  19866=>"001001111",
  19867=>"111111111",
  19868=>"000111111",
  19869=>"000000000",
  19870=>"000000000",
  19871=>"000000111",
  19872=>"000110000",
  19873=>"011111101",
  19874=>"111001000",
  19875=>"111111000",
  19876=>"111001001",
  19877=>"001111011",
  19878=>"100111111",
  19879=>"111111100",
  19880=>"000000000",
  19881=>"011111000",
  19882=>"111010000",
  19883=>"001000000",
  19884=>"110010000",
  19885=>"000000111",
  19886=>"011000110",
  19887=>"000100000",
  19888=>"111000000",
  19889=>"100000111",
  19890=>"001111111",
  19891=>"000110111",
  19892=>"000001000",
  19893=>"001000001",
  19894=>"111011110",
  19895=>"111011001",
  19896=>"100000000",
  19897=>"000111111",
  19898=>"110000000",
  19899=>"111100010",
  19900=>"111011111",
  19901=>"000000001",
  19902=>"000000000",
  19903=>"111100000",
  19904=>"000000110",
  19905=>"111111000",
  19906=>"000001011",
  19907=>"110111010",
  19908=>"011000101",
  19909=>"111001000",
  19910=>"111110000",
  19911=>"110111111",
  19912=>"000101000",
  19913=>"110111110",
  19914=>"111000000",
  19915=>"000111111",
  19916=>"000000001",
  19917=>"010110010",
  19918=>"110000110",
  19919=>"111110111",
  19920=>"001000000",
  19921=>"111111111",
  19922=>"110000000",
  19923=>"000111110",
  19924=>"100000000",
  19925=>"111111000",
  19926=>"000110111",
  19927=>"111111101",
  19928=>"000000111",
  19929=>"111011000",
  19930=>"010110111",
  19931=>"000000000",
  19932=>"111011000",
  19933=>"001001001",
  19934=>"111111111",
  19935=>"111110100",
  19936=>"111111111",
  19937=>"000000111",
  19938=>"111111001",
  19939=>"000000000",
  19940=>"000000000",
  19941=>"000111111",
  19942=>"011001000",
  19943=>"111000000",
  19944=>"111111101",
  19945=>"111010000",
  19946=>"000010000",
  19947=>"001111001",
  19948=>"110011111",
  19949=>"110000000",
  19950=>"000111111",
  19951=>"000000111",
  19952=>"111101001",
  19953=>"111111000",
  19954=>"111111111",
  19955=>"000000000",
  19956=>"111111111",
  19957=>"000100111",
  19958=>"111110000",
  19959=>"110111100",
  19960=>"110000111",
  19961=>"111111000",
  19962=>"000000000",
  19963=>"111111001",
  19964=>"000111110",
  19965=>"001111111",
  19966=>"110111000",
  19967=>"111111000",
  19968=>"111111101",
  19969=>"110111101",
  19970=>"000100111",
  19971=>"000000110",
  19972=>"111111000",
  19973=>"000000010",
  19974=>"111011001",
  19975=>"000000000",
  19976=>"000000000",
  19977=>"001111001",
  19978=>"101101101",
  19979=>"000000000",
  19980=>"110110100",
  19981=>"000111111",
  19982=>"010110001",
  19983=>"111111011",
  19984=>"001001000",
  19985=>"111111111",
  19986=>"000000000",
  19987=>"111111111",
  19988=>"000000100",
  19989=>"000000000",
  19990=>"111111111",
  19991=>"001011001",
  19992=>"111111110",
  19993=>"111111111",
  19994=>"010000110",
  19995=>"000000000",
  19996=>"111111111",
  19997=>"011001000",
  19998=>"111111000",
  19999=>"000001111",
  20000=>"100100110",
  20001=>"000100111",
  20002=>"001101110",
  20003=>"111111110",
  20004=>"111001000",
  20005=>"000000001",
  20006=>"000000100",
  20007=>"011000100",
  20008=>"011000101",
  20009=>"000000000",
  20010=>"101110100",
  20011=>"111111111",
  20012=>"111111011",
  20013=>"000000000",
  20014=>"000110100",
  20015=>"110111111",
  20016=>"101000111",
  20017=>"111111111",
  20018=>"001000111",
  20019=>"000000111",
  20020=>"100110000",
  20021=>"111111111",
  20022=>"111000110",
  20023=>"100000000",
  20024=>"111111000",
  20025=>"000001111",
  20026=>"011011011",
  20027=>"111111111",
  20028=>"000001111",
  20029=>"100001011",
  20030=>"111000010",
  20031=>"000000111",
  20032=>"111111001",
  20033=>"000000000",
  20034=>"011011111",
  20035=>"000000000",
  20036=>"010111111",
  20037=>"111111111",
  20038=>"111110000",
  20039=>"111111111",
  20040=>"001001001",
  20041=>"111000110",
  20042=>"111111010",
  20043=>"101001011",
  20044=>"111100000",
  20045=>"000000100",
  20046=>"010000000",
  20047=>"000000000",
  20048=>"000000000",
  20049=>"000110011",
  20050=>"000000000",
  20051=>"110111111",
  20052=>"000000000",
  20053=>"000000000",
  20054=>"111111111",
  20055=>"100110110",
  20056=>"000000101",
  20057=>"111000101",
  20058=>"111111111",
  20059=>"000000000",
  20060=>"111111111",
  20061=>"001001111",
  20062=>"100101111",
  20063=>"000000011",
  20064=>"111111000",
  20065=>"100111011",
  20066=>"111111001",
  20067=>"000000001",
  20068=>"111111110",
  20069=>"111111111",
  20070=>"110010000",
  20071=>"111110111",
  20072=>"110111111",
  20073=>"000100100",
  20074=>"010100111",
  20075=>"000000000",
  20076=>"100100000",
  20077=>"110111000",
  20078=>"000000001",
  20079=>"111011111",
  20080=>"111000000",
  20081=>"000000111",
  20082=>"000111111",
  20083=>"100101111",
  20084=>"000000000",
  20085=>"000000000",
  20086=>"001011011",
  20087=>"111111000",
  20088=>"000000011",
  20089=>"100000000",
  20090=>"000000111",
  20091=>"000000000",
  20092=>"001000000",
  20093=>"000000000",
  20094=>"111111111",
  20095=>"000110100",
  20096=>"000000000",
  20097=>"100110100",
  20098=>"010100000",
  20099=>"011011011",
  20100=>"111111011",
  20101=>"000000111",
  20102=>"000000110",
  20103=>"111111001",
  20104=>"000001001",
  20105=>"000111111",
  20106=>"111101001",
  20107=>"010111111",
  20108=>"101111111",
  20109=>"111101111",
  20110=>"000000000",
  20111=>"010000000",
  20112=>"101000111",
  20113=>"111100100",
  20114=>"001011111",
  20115=>"011111111",
  20116=>"100100111",
  20117=>"000000110",
  20118=>"000000000",
  20119=>"111111111",
  20120=>"100100111",
  20121=>"100100110",
  20122=>"000000000",
  20123=>"101100101",
  20124=>"111111111",
  20125=>"101001000",
  20126=>"111111000",
  20127=>"111111111",
  20128=>"000000000",
  20129=>"111111111",
  20130=>"111111111",
  20131=>"111111111",
  20132=>"110111110",
  20133=>"110111111",
  20134=>"100000000",
  20135=>"111010000",
  20136=>"110000000",
  20137=>"000000000",
  20138=>"111111111",
  20139=>"110000000",
  20140=>"010111111",
  20141=>"100100001",
  20142=>"111111111",
  20143=>"000000001",
  20144=>"000000001",
  20145=>"111111100",
  20146=>"111111011",
  20147=>"111010000",
  20148=>"110101011",
  20149=>"000000110",
  20150=>"001111111",
  20151=>"110000011",
  20152=>"000000000",
  20153=>"000000000",
  20154=>"110000000",
  20155=>"100111111",
  20156=>"001001000",
  20157=>"111111111",
  20158=>"110110111",
  20159=>"100100010",
  20160=>"100111111",
  20161=>"000000000",
  20162=>"111111111",
  20163=>"001111111",
  20164=>"111111111",
  20165=>"000000101",
  20166=>"100000110",
  20167=>"111111111",
  20168=>"000000010",
  20169=>"001000001",
  20170=>"101101111",
  20171=>"100000000",
  20172=>"110110100",
  20173=>"101111001",
  20174=>"111011011",
  20175=>"111000000",
  20176=>"000000000",
  20177=>"000100110",
  20178=>"101000000",
  20179=>"001001000",
  20180=>"111111011",
  20181=>"100100100",
  20182=>"000000111",
  20183=>"101100111",
  20184=>"111000000",
  20185=>"000000101",
  20186=>"100000000",
  20187=>"000011111",
  20188=>"000000011",
  20189=>"111111101",
  20190=>"111111111",
  20191=>"100000010",
  20192=>"000110000",
  20193=>"000011111",
  20194=>"111101000",
  20195=>"111111111",
  20196=>"010111110",
  20197=>"011001001",
  20198=>"000010111",
  20199=>"000000101",
  20200=>"110111111",
  20201=>"101111000",
  20202=>"000000001",
  20203=>"110101111",
  20204=>"001000000",
  20205=>"000000000",
  20206=>"111000011",
  20207=>"111111111",
  20208=>"100110000",
  20209=>"000000000",
  20210=>"111001000",
  20211=>"000000100",
  20212=>"111111111",
  20213=>"111001000",
  20214=>"100100000",
  20215=>"110111111",
  20216=>"110111111",
  20217=>"000000000",
  20218=>"000000011",
  20219=>"111110000",
  20220=>"111110000",
  20221=>"000000000",
  20222=>"000000000",
  20223=>"000000001",
  20224=>"000000100",
  20225=>"111001001",
  20226=>"011011000",
  20227=>"000001011",
  20228=>"111101111",
  20229=>"000000000",
  20230=>"111111111",
  20231=>"100111111",
  20232=>"000000000",
  20233=>"100000110",
  20234=>"111111111",
  20235=>"111111011",
  20236=>"111111111",
  20237=>"000000000",
  20238=>"111110110",
  20239=>"000000010",
  20240=>"001011000",
  20241=>"111111111",
  20242=>"000000000",
  20243=>"000111111",
  20244=>"000000000",
  20245=>"000000000",
  20246=>"011000000",
  20247=>"000000000",
  20248=>"001111000",
  20249=>"111111000",
  20250=>"111111111",
  20251=>"000000000",
  20252=>"000000000",
  20253=>"111111111",
  20254=>"000000000",
  20255=>"110000000",
  20256=>"110111011",
  20257=>"111100000",
  20258=>"111111111",
  20259=>"000011111",
  20260=>"110110000",
  20261=>"000001111",
  20262=>"111111111",
  20263=>"000000100",
  20264=>"000000111",
  20265=>"010111010",
  20266=>"110101111",
  20267=>"111111111",
  20268=>"111111001",
  20269=>"110100000",
  20270=>"101000000",
  20271=>"010010011",
  20272=>"000000000",
  20273=>"000000000",
  20274=>"000100101",
  20275=>"000000111",
  20276=>"000000000",
  20277=>"001000000",
  20278=>"000110110",
  20279=>"000000000",
  20280=>"000000000",
  20281=>"000001100",
  20282=>"000000101",
  20283=>"000000110",
  20284=>"111110110",
  20285=>"000100111",
  20286=>"000000001",
  20287=>"001001111",
  20288=>"001000000",
  20289=>"000000000",
  20290=>"111111111",
  20291=>"000110110",
  20292=>"111111111",
  20293=>"111000000",
  20294=>"110000000",
  20295=>"001111010",
  20296=>"111001001",
  20297=>"000000100",
  20298=>"111111111",
  20299=>"110000001",
  20300=>"000000001",
  20301=>"000001000",
  20302=>"000000000",
  20303=>"110110100",
  20304=>"001001001",
  20305=>"000000110",
  20306=>"111110110",
  20307=>"110110111",
  20308=>"000111111",
  20309=>"011011001",
  20310=>"001001001",
  20311=>"001111111",
  20312=>"000100010",
  20313=>"000000000",
  20314=>"000001000",
  20315=>"010010011",
  20316=>"000000000",
  20317=>"110111111",
  20318=>"110111111",
  20319=>"000001000",
  20320=>"111111100",
  20321=>"000000000",
  20322=>"001001000",
  20323=>"000100111",
  20324=>"000000000",
  20325=>"000000000",
  20326=>"000011001",
  20327=>"001000101",
  20328=>"111111110",
  20329=>"011011111",
  20330=>"000000001",
  20331=>"111010101",
  20332=>"000001000",
  20333=>"100000000",
  20334=>"110110100",
  20335=>"111000000",
  20336=>"111111111",
  20337=>"011001001",
  20338=>"000111001",
  20339=>"111111011",
  20340=>"000000000",
  20341=>"000001111",
  20342=>"000000000",
  20343=>"000000000",
  20344=>"111101111",
  20345=>"111100000",
  20346=>"100111000",
  20347=>"111111111",
  20348=>"100000000",
  20349=>"110110100",
  20350=>"000000000",
  20351=>"000000000",
  20352=>"011001000",
  20353=>"000000000",
  20354=>"111111111",
  20355=>"000000000",
  20356=>"100100000",
  20357=>"110111111",
  20358=>"011000000",
  20359=>"000000000",
  20360=>"100000000",
  20361=>"111011011",
  20362=>"111011011",
  20363=>"110100000",
  20364=>"101100111",
  20365=>"110100100",
  20366=>"101100000",
  20367=>"000000100",
  20368=>"111011111",
  20369=>"111101110",
  20370=>"011111111",
  20371=>"111110110",
  20372=>"011111111",
  20373=>"000010000",
  20374=>"001000001",
  20375=>"000001000",
  20376=>"000000000",
  20377=>"101111000",
  20378=>"100111111",
  20379=>"101100101",
  20380=>"110111000",
  20381=>"111000000",
  20382=>"000000000",
  20383=>"111111110",
  20384=>"000011001",
  20385=>"011011010",
  20386=>"000001110",
  20387=>"000010000",
  20388=>"000110100",
  20389=>"000000010",
  20390=>"111111001",
  20391=>"000111000",
  20392=>"110000000",
  20393=>"110010000",
  20394=>"111111010",
  20395=>"100100101",
  20396=>"011011011",
  20397=>"000000001",
  20398=>"000000001",
  20399=>"000000000",
  20400=>"111111111",
  20401=>"000000000",
  20402=>"000000000",
  20403=>"000000000",
  20404=>"011101111",
  20405=>"110111111",
  20406=>"000101111",
  20407=>"011000000",
  20408=>"001111000",
  20409=>"000000111",
  20410=>"111111111",
  20411=>"001000000",
  20412=>"001110111",
  20413=>"000110111",
  20414=>"000000000",
  20415=>"000110110",
  20416=>"000011011",
  20417=>"001000000",
  20418=>"000000111",
  20419=>"000000000",
  20420=>"101111111",
  20421=>"111011011",
  20422=>"000000101",
  20423=>"000000011",
  20424=>"000000000",
  20425=>"001001000",
  20426=>"000000001",
  20427=>"111111111",
  20428=>"110000010",
  20429=>"000000110",
  20430=>"111111101",
  20431=>"111111110",
  20432=>"011010000",
  20433=>"110100011",
  20434=>"000110110",
  20435=>"000000111",
  20436=>"111111111",
  20437=>"001000000",
  20438=>"000000000",
  20439=>"011011011",
  20440=>"101101111",
  20441=>"000000000",
  20442=>"001010111",
  20443=>"111001011",
  20444=>"000000000",
  20445=>"000000101",
  20446=>"000000000",
  20447=>"111111111",
  20448=>"111000000",
  20449=>"111100000",
  20450=>"000000000",
  20451=>"001000000",
  20452=>"111100110",
  20453=>"000110000",
  20454=>"000010001",
  20455=>"111011011",
  20456=>"000000001",
  20457=>"111111111",
  20458=>"111111001",
  20459=>"000001111",
  20460=>"000000000",
  20461=>"000000000",
  20462=>"000000000",
  20463=>"100110100",
  20464=>"000000000",
  20465=>"111111111",
  20466=>"111111111",
  20467=>"000001111",
  20468=>"111111111",
  20469=>"000000000",
  20470=>"000001001",
  20471=>"111111000",
  20472=>"011011011",
  20473=>"000000001",
  20474=>"001101101",
  20475=>"000000000",
  20476=>"100000000",
  20477=>"000000000",
  20478=>"000000001",
  20479=>"101111111",
  20480=>"111001000",
  20481=>"000000011",
  20482=>"000010010",
  20483=>"011011000",
  20484=>"000111111",
  20485=>"000000000",
  20486=>"111111111",
  20487=>"111010010",
  20488=>"011000000",
  20489=>"111110110",
  20490=>"100111101",
  20491=>"100101100",
  20492=>"000000000",
  20493=>"110000000",
  20494=>"111111111",
  20495=>"000000000",
  20496=>"111111011",
  20497=>"000111011",
  20498=>"000000000",
  20499=>"111111110",
  20500=>"000000000",
  20501=>"000000000",
  20502=>"111111001",
  20503=>"100100000",
  20504=>"000001001",
  20505=>"000011110",
  20506=>"111111110",
  20507=>"010011111",
  20508=>"000000000",
  20509=>"000000000",
  20510=>"001011001",
  20511=>"111111111",
  20512=>"000000000",
  20513=>"110000000",
  20514=>"100111111",
  20515=>"111111111",
  20516=>"100000000",
  20517=>"000110101",
  20518=>"000000001",
  20519=>"000000000",
  20520=>"111111111",
  20521=>"011111011",
  20522=>"111011001",
  20523=>"001001001",
  20524=>"000000111",
  20525=>"000000000",
  20526=>"000000000",
  20527=>"110010010",
  20528=>"000000000",
  20529=>"000000000",
  20530=>"000110110",
  20531=>"000111111",
  20532=>"000101111",
  20533=>"111111111",
  20534=>"111111111",
  20535=>"000001000",
  20536=>"111011000",
  20537=>"001000000",
  20538=>"000000101",
  20539=>"111000011",
  20540=>"111111111",
  20541=>"011111011",
  20542=>"000000000",
  20543=>"001000000",
  20544=>"101111011",
  20545=>"000000000",
  20546=>"110111111",
  20547=>"101001111",
  20548=>"110000000",
  20549=>"011000110",
  20550=>"001000111",
  20551=>"111111001",
  20552=>"001000000",
  20553=>"101100111",
  20554=>"011111111",
  20555=>"111111110",
  20556=>"111111111",
  20557=>"000000111",
  20558=>"000000111",
  20559=>"010000001",
  20560=>"000000000",
  20561=>"100001111",
  20562=>"100111000",
  20563=>"101100100",
  20564=>"000000000",
  20565=>"011011111",
  20566=>"100110010",
  20567=>"000000000",
  20568=>"111111000",
  20569=>"000000111",
  20570=>"111000000",
  20571=>"110100000",
  20572=>"001001001",
  20573=>"111111111",
  20574=>"111111111",
  20575=>"011001100",
  20576=>"010000000",
  20577=>"111111010",
  20578=>"011111110",
  20579=>"000110110",
  20580=>"110111111",
  20581=>"000000000",
  20582=>"111101111",
  20583=>"000000000",
  20584=>"111111111",
  20585=>"111111111",
  20586=>"101010010",
  20587=>"000000000",
  20588=>"101100000",
  20589=>"000000000",
  20590=>"111110000",
  20591=>"000000101",
  20592=>"111111010",
  20593=>"111111111",
  20594=>"011011011",
  20595=>"111101001",
  20596=>"000000001",
  20597=>"111001000",
  20598=>"111111000",
  20599=>"100000000",
  20600=>"010011000",
  20601=>"111111111",
  20602=>"111111111",
  20603=>"000000000",
  20604=>"010100111",
  20605=>"000110110",
  20606=>"100111010",
  20607=>"000001000",
  20608=>"000000000",
  20609=>"111000000",
  20610=>"000000000",
  20611=>"000000000",
  20612=>"111111101",
  20613=>"101000000",
  20614=>"000000100",
  20615=>"110111111",
  20616=>"111001000",
  20617=>"111000000",
  20618=>"000000000",
  20619=>"000000000",
  20620=>"111001011",
  20621=>"111110010",
  20622=>"001111111",
  20623=>"000000000",
  20624=>"111111011",
  20625=>"000000001",
  20626=>"111110000",
  20627=>"000000000",
  20628=>"000000110",
  20629=>"111111111",
  20630=>"111111111",
  20631=>"111111000",
  20632=>"111011011",
  20633=>"000000000",
  20634=>"000000011",
  20635=>"000000010",
  20636=>"101000010",
  20637=>"110111111",
  20638=>"000000111",
  20639=>"000000000",
  20640=>"111111110",
  20641=>"110100111",
  20642=>"000000000",
  20643=>"000000000",
  20644=>"000011000",
  20645=>"110010000",
  20646=>"000000111",
  20647=>"110111111",
  20648=>"000011111",
  20649=>"101000000",
  20650=>"000000000",
  20651=>"100101101",
  20652=>"111111111",
  20653=>"111111000",
  20654=>"011011011",
  20655=>"111111111",
  20656=>"111010000",
  20657=>"110110001",
  20658=>"111110110",
  20659=>"010111111",
  20660=>"000000101",
  20661=>"111001011",
  20662=>"000000000",
  20663=>"111111011",
  20664=>"000000000",
  20665=>"000000000",
  20666=>"001001011",
  20667=>"111000000",
  20668=>"111111111",
  20669=>"111101000",
  20670=>"110000000",
  20671=>"011000000",
  20672=>"000100111",
  20673=>"110111000",
  20674=>"010000000",
  20675=>"111111111",
  20676=>"111010111",
  20677=>"011011011",
  20678=>"000000000",
  20679=>"010001000",
  20680=>"000000000",
  20681=>"000001110",
  20682=>"000000000",
  20683=>"111110010",
  20684=>"100100000",
  20685=>"110100000",
  20686=>"111110100",
  20687=>"111111110",
  20688=>"111111011",
  20689=>"000110111",
  20690=>"111111111",
  20691=>"000000010",
  20692=>"000000000",
  20693=>"111111100",
  20694=>"000000100",
  20695=>"010000000",
  20696=>"111111000",
  20697=>"111111000",
  20698=>"000000011",
  20699=>"111111111",
  20700=>"000001111",
  20701=>"111111100",
  20702=>"111111111",
  20703=>"111011111",
  20704=>"000000000",
  20705=>"000000011",
  20706=>"111111111",
  20707=>"111111111",
  20708=>"000100110",
  20709=>"100110110",
  20710=>"111111111",
  20711=>"111011000",
  20712=>"001001000",
  20713=>"111111111",
  20714=>"001000010",
  20715=>"001111111",
  20716=>"111111111",
  20717=>"111111111",
  20718=>"010110001",
  20719=>"000010100",
  20720=>"011001000",
  20721=>"110110110",
  20722=>"111000111",
  20723=>"000000001",
  20724=>"000011000",
  20725=>"110110111",
  20726=>"100100000",
  20727=>"000000000",
  20728=>"000101111",
  20729=>"011011000",
  20730=>"000000000",
  20731=>"010000111",
  20732=>"001000000",
  20733=>"000101111",
  20734=>"100000101",
  20735=>"000001000",
  20736=>"011111110",
  20737=>"000001001",
  20738=>"000111111",
  20739=>"000000000",
  20740=>"111011000",
  20741=>"111111111",
  20742=>"110111111",
  20743=>"000111111",
  20744=>"001001011",
  20745=>"000000000",
  20746=>"101111111",
  20747=>"010000000",
  20748=>"100000100",
  20749=>"000000000",
  20750=>"011101100",
  20751=>"111111111",
  20752=>"111111001",
  20753=>"000101111",
  20754=>"111110111",
  20755=>"000100100",
  20756=>"111111111",
  20757=>"111111010",
  20758=>"110000000",
  20759=>"100111111",
  20760=>"111111111",
  20761=>"000111111",
  20762=>"000011000",
  20763=>"111110110",
  20764=>"000000001",
  20765=>"000000111",
  20766=>"111110110",
  20767=>"000000100",
  20768=>"100110111",
  20769=>"000000000",
  20770=>"000000000",
  20771=>"111111111",
  20772=>"100000000",
  20773=>"000001111",
  20774=>"011001000",
  20775=>"111111111",
  20776=>"000111111",
  20777=>"000000000",
  20778=>"110001000",
  20779=>"000000101",
  20780=>"111110100",
  20781=>"001001001",
  20782=>"000111000",
  20783=>"000000000",
  20784=>"000000000",
  20785=>"000011110",
  20786=>"000000000",
  20787=>"000000001",
  20788=>"111100111",
  20789=>"111000000",
  20790=>"011011111",
  20791=>"000000000",
  20792=>"010000000",
  20793=>"000000000",
  20794=>"000000011",
  20795=>"000000011",
  20796=>"001111011",
  20797=>"000000100",
  20798=>"000011111",
  20799=>"011000000",
  20800=>"111110110",
  20801=>"000000000",
  20802=>"000000000",
  20803=>"111111010",
  20804=>"000000111",
  20805=>"000000111",
  20806=>"110111111",
  20807=>"111111110",
  20808=>"000000000",
  20809=>"010000111",
  20810=>"111000110",
  20811=>"100101111",
  20812=>"111111101",
  20813=>"100101111",
  20814=>"000000000",
  20815=>"111110100",
  20816=>"011011110",
  20817=>"101000000",
  20818=>"110000000",
  20819=>"001001101",
  20820=>"000000000",
  20821=>"111111001",
  20822=>"111111111",
  20823=>"000000111",
  20824=>"000000000",
  20825=>"000000000",
  20826=>"111000000",
  20827=>"001011111",
  20828=>"000000000",
  20829=>"110111111",
  20830=>"100100101",
  20831=>"000011111",
  20832=>"111111111",
  20833=>"111001011",
  20834=>"111110000",
  20835=>"000000000",
  20836=>"111111111",
  20837=>"001000101",
  20838=>"000000000",
  20839=>"111111001",
  20840=>"011111111",
  20841=>"111111011",
  20842=>"001111010",
  20843=>"011011101",
  20844=>"100111111",
  20845=>"111011001",
  20846=>"000000000",
  20847=>"000011111",
  20848=>"010111110",
  20849=>"010110000",
  20850=>"111000100",
  20851=>"000000111",
  20852=>"110000000",
  20853=>"000111011",
  20854=>"000010000",
  20855=>"011001001",
  20856=>"000000111",
  20857=>"000000000",
  20858=>"000011011",
  20859=>"000000001",
  20860=>"100000000",
  20861=>"111111001",
  20862=>"000000101",
  20863=>"000000000",
  20864=>"001111111",
  20865=>"111111111",
  20866=>"000011010",
  20867=>"000000000",
  20868=>"000001111",
  20869=>"111110000",
  20870=>"000000000",
  20871=>"111111001",
  20872=>"001001111",
  20873=>"111111000",
  20874=>"000100110",
  20875=>"111001111",
  20876=>"111111111",
  20877=>"110000010",
  20878=>"001001001",
  20879=>"110111110",
  20880=>"000000000",
  20881=>"000000000",
  20882=>"011110100",
  20883=>"000010010",
  20884=>"001000000",
  20885=>"010010000",
  20886=>"111111111",
  20887=>"000000101",
  20888=>"000000100",
  20889=>"111000000",
  20890=>"000000100",
  20891=>"000000000",
  20892=>"000000110",
  20893=>"001001110",
  20894=>"000001001",
  20895=>"000110110",
  20896=>"000110100",
  20897=>"111111000",
  20898=>"111001001",
  20899=>"000000000",
  20900=>"000111111",
  20901=>"110110111",
  20902=>"111000000",
  20903=>"110111111",
  20904=>"000000101",
  20905=>"111011001",
  20906=>"000111111",
  20907=>"101000000",
  20908=>"111111100",
  20909=>"111111111",
  20910=>"000010011",
  20911=>"001100000",
  20912=>"000000000",
  20913=>"111000000",
  20914=>"110011111",
  20915=>"111111111",
  20916=>"100000111",
  20917=>"111011011",
  20918=>"000110110",
  20919=>"100000000",
  20920=>"000000101",
  20921=>"111111111",
  20922=>"000000000",
  20923=>"111111001",
  20924=>"111000111",
  20925=>"001011101",
  20926=>"000000100",
  20927=>"110010000",
  20928=>"010111111",
  20929=>"000000000",
  20930=>"001001001",
  20931=>"101100111",
  20932=>"000000111",
  20933=>"000000100",
  20934=>"001001011",
  20935=>"011000000",
  20936=>"111011011",
  20937=>"111000000",
  20938=>"000000111",
  20939=>"111111101",
  20940=>"000000001",
  20941=>"111111111",
  20942=>"000000101",
  20943=>"111111110",
  20944=>"000000000",
  20945=>"111111111",
  20946=>"111111110",
  20947=>"111111110",
  20948=>"000000000",
  20949=>"000010110",
  20950=>"110111110",
  20951=>"111110011",
  20952=>"000000000",
  20953=>"000000101",
  20954=>"000000000",
  20955=>"111111000",
  20956=>"000010000",
  20957=>"000000000",
  20958=>"111011011",
  20959=>"000000000",
  20960=>"000010110",
  20961=>"001011001",
  20962=>"110111110",
  20963=>"000010111",
  20964=>"000001111",
  20965=>"101100111",
  20966=>"111111011",
  20967=>"111111111",
  20968=>"000000000",
  20969=>"111111111",
  20970=>"000000000",
  20971=>"111111111",
  20972=>"110000001",
  20973=>"111101111",
  20974=>"000001000",
  20975=>"111111111",
  20976=>"011011001",
  20977=>"111101001",
  20978=>"000011011",
  20979=>"110010111",
  20980=>"000000000",
  20981=>"000000010",
  20982=>"001011111",
  20983=>"111011110",
  20984=>"000100110",
  20985=>"011000000",
  20986=>"000110111",
  20987=>"111111000",
  20988=>"111000000",
  20989=>"100011000",
  20990=>"111011011",
  20991=>"110110110",
  20992=>"000000100",
  20993=>"100000001",
  20994=>"111111111",
  20995=>"000000101",
  20996=>"110110111",
  20997=>"000000000",
  20998=>"111111001",
  20999=>"100101111",
  21000=>"000000000",
  21001=>"000110110",
  21002=>"101001001",
  21003=>"111111111",
  21004=>"110110110",
  21005=>"111111010",
  21006=>"110100011",
  21007=>"000000000",
  21008=>"100100110",
  21009=>"010110111",
  21010=>"000000000",
  21011=>"000000110",
  21012=>"000000100",
  21013=>"111111111",
  21014=>"111111111",
  21015=>"111100100",
  21016=>"100000101",
  21017=>"110100100",
  21018=>"101100111",
  21019=>"111111111",
  21020=>"001000001",
  21021=>"111111011",
  21022=>"100000011",
  21023=>"100000000",
  21024=>"100000000",
  21025=>"000100000",
  21026=>"000000000",
  21027=>"111011001",
  21028=>"110110010",
  21029=>"110110010",
  21030=>"000000000",
  21031=>"111111111",
  21032=>"000000000",
  21033=>"100101101",
  21034=>"000000000",
  21035=>"100111101",
  21036=>"111110000",
  21037=>"000000100",
  21038=>"001001001",
  21039=>"111111111",
  21040=>"011000000",
  21041=>"000001000",
  21042=>"101100100",
  21043=>"011011011",
  21044=>"111111000",
  21045=>"000010110",
  21046=>"111111000",
  21047=>"111110011",
  21048=>"000000000",
  21049=>"000001111",
  21050=>"011001011",
  21051=>"000001111",
  21052=>"000000000",
  21053=>"000000000",
  21054=>"011001000",
  21055=>"000000101",
  21056=>"000011011",
  21057=>"010010000",
  21058=>"111110100",
  21059=>"111111111",
  21060=>"110110100",
  21061=>"011011001",
  21062=>"100000000",
  21063=>"000000000",
  21064=>"111111001",
  21065=>"111101011",
  21066=>"001001000",
  21067=>"010000001",
  21068=>"111111101",
  21069=>"000000000",
  21070=>"000000000",
  21071=>"001000000",
  21072=>"101101001",
  21073=>"111111010",
  21074=>"000000000",
  21075=>"110110110",
  21076=>"001001101",
  21077=>"101000000",
  21078=>"000001101",
  21079=>"111111111",
  21080=>"111011010",
  21081=>"100000001",
  21082=>"000000000",
  21083=>"100000000",
  21084=>"000000011",
  21085=>"000101101",
  21086=>"010111111",
  21087=>"011010000",
  21088=>"000111011",
  21089=>"001001101",
  21090=>"111101111",
  21091=>"001000100",
  21092=>"110110010",
  21093=>"100101111",
  21094=>"001001000",
  21095=>"000000000",
  21096=>"000001100",
  21097=>"001000101",
  21098=>"010010111",
  21099=>"111001001",
  21100=>"000000000",
  21101=>"000000000",
  21102=>"000000001",
  21103=>"010000000",
  21104=>"011011000",
  21105=>"010010111",
  21106=>"101001001",
  21107=>"011001000",
  21108=>"001001001",
  21109=>"100110000",
  21110=>"111100101",
  21111=>"010111000",
  21112=>"000100000",
  21113=>"000000000",
  21114=>"001001001",
  21115=>"000000000",
  21116=>"100110100",
  21117=>"111000000",
  21118=>"110000000",
  21119=>"110111010",
  21120=>"000001001",
  21121=>"110110111",
  21122=>"011000000",
  21123=>"000000000",
  21124=>"001101001",
  21125=>"001001101",
  21126=>"001001101",
  21127=>"110110111",
  21128=>"000110110",
  21129=>"000001111",
  21130=>"111111111",
  21131=>"000001001",
  21132=>"111111111",
  21133=>"000000000",
  21134=>"000000101",
  21135=>"010010011",
  21136=>"101101101",
  21137=>"000000000",
  21138=>"111111110",
  21139=>"001000000",
  21140=>"010000000",
  21141=>"101101111",
  21142=>"000111111",
  21143=>"000000111",
  21144=>"001001000",
  21145=>"100100000",
  21146=>"101011001",
  21147=>"000001110",
  21148=>"010000011",
  21149=>"001001111",
  21150=>"111111110",
  21151=>"000000101",
  21152=>"111001000",
  21153=>"110111111",
  21154=>"000000000",
  21155=>"110010010",
  21156=>"000000000",
  21157=>"011111111",
  21158=>"000000000",
  21159=>"110110111",
  21160=>"011000001",
  21161=>"000001101",
  21162=>"001000000",
  21163=>"101101111",
  21164=>"111111111",
  21165=>"001001001",
  21166=>"111101000",
  21167=>"111100111",
  21168=>"010011010",
  21169=>"011111110",
  21170=>"111111110",
  21171=>"111101101",
  21172=>"111011011",
  21173=>"001011011",
  21174=>"111111110",
  21175=>"110110110",
  21176=>"000000000",
  21177=>"011111111",
  21178=>"110111000",
  21179=>"000000000",
  21180=>"111101111",
  21181=>"111110110",
  21182=>"011111100",
  21183=>"111111111",
  21184=>"100000000",
  21185=>"000000000",
  21186=>"010110111",
  21187=>"010010000",
  21188=>"101101111",
  21189=>"000000001",
  21190=>"101000000",
  21191=>"001101101",
  21192=>"000011011",
  21193=>"100111111",
  21194=>"101000000",
  21195=>"100000000",
  21196=>"110111111",
  21197=>"111111110",
  21198=>"100000000",
  21199=>"000111101",
  21200=>"000001000",
  21201=>"000000101",
  21202=>"110000000",
  21203=>"111111011",
  21204=>"101111111",
  21205=>"001101000",
  21206=>"000000000",
  21207=>"111111111",
  21208=>"111010000",
  21209=>"111101101",
  21210=>"111111111",
  21211=>"111001000",
  21212=>"001001111",
  21213=>"111100000",
  21214=>"000000000",
  21215=>"000000001",
  21216=>"000000001",
  21217=>"011010010",
  21218=>"000000000",
  21219=>"000010000",
  21220=>"111111110",
  21221=>"011000000",
  21222=>"110100100",
  21223=>"110110110",
  21224=>"010110010",
  21225=>"000101001",
  21226=>"110000000",
  21227=>"011111001",
  21228=>"101000101",
  21229=>"101000000",
  21230=>"010010111",
  21231=>"111101111",
  21232=>"001101101",
  21233=>"000001000",
  21234=>"000001111",
  21235=>"001001000",
  21236=>"010110110",
  21237=>"110100000",
  21238=>"011011011",
  21239=>"111111010",
  21240=>"010000010",
  21241=>"111111001",
  21242=>"000001000",
  21243=>"111111000",
  21244=>"001010110",
  21245=>"000000101",
  21246=>"100100111",
  21247=>"000001001",
  21248=>"000000001",
  21249=>"001001001",
  21250=>"100111101",
  21251=>"110000010",
  21252=>"101001001",
  21253=>"000010011",
  21254=>"100111001",
  21255=>"000110010",
  21256=>"111001000",
  21257=>"000000001",
  21258=>"111101100",
  21259=>"010111011",
  21260=>"000000000",
  21261=>"101101100",
  21262=>"111111111",
  21263=>"000000100",
  21264=>"111001001",
  21265=>"111111111",
  21266=>"111111111",
  21267=>"110110111",
  21268=>"111111111",
  21269=>"000000000",
  21270=>"001001000",
  21271=>"001001111",
  21272=>"010110110",
  21273=>"000111111",
  21274=>"110000000",
  21275=>"000000000",
  21276=>"111111111",
  21277=>"111111111",
  21278=>"000001001",
  21279=>"111111111",
  21280=>"010000000",
  21281=>"000001111",
  21282=>"111010010",
  21283=>"110110111",
  21284=>"000000000",
  21285=>"000000000",
  21286=>"000000000",
  21287=>"001000000",
  21288=>"000001001",
  21289=>"111011000",
  21290=>"010010010",
  21291=>"001001000",
  21292=>"101000000",
  21293=>"011001001",
  21294=>"011000111",
  21295=>"111000000",
  21296=>"000100111",
  21297=>"110000000",
  21298=>"000001001",
  21299=>"010000000",
  21300=>"100101101",
  21301=>"011001001",
  21302=>"000111110",
  21303=>"101001101",
  21304=>"000000000",
  21305=>"000000111",
  21306=>"111111111",
  21307=>"100000100",
  21308=>"000011101",
  21309=>"111111111",
  21310=>"110110011",
  21311=>"000000000",
  21312=>"111111110",
  21313=>"100110100",
  21314=>"110110010",
  21315=>"001001001",
  21316=>"001001100",
  21317=>"100000110",
  21318=>"001101011",
  21319=>"000110111",
  21320=>"100101101",
  21321=>"111011111",
  21322=>"111111111",
  21323=>"111111100",
  21324=>"111000010",
  21325=>"110110010",
  21326=>"111111111",
  21327=>"011010110",
  21328=>"001001000",
  21329=>"000001000",
  21330=>"111000000",
  21331=>"111111111",
  21332=>"100000001",
  21333=>"011011001",
  21334=>"000000110",
  21335=>"100101101",
  21336=>"110111111",
  21337=>"111111111",
  21338=>"000000000",
  21339=>"001000000",
  21340=>"011000000",
  21341=>"001001111",
  21342=>"100100110",
  21343=>"110110111",
  21344=>"000001100",
  21345=>"000000000",
  21346=>"000111110",
  21347=>"001101101",
  21348=>"100110100",
  21349=>"000000000",
  21350=>"000111111",
  21351=>"110000000",
  21352=>"111101100",
  21353=>"110000010",
  21354=>"011000000",
  21355=>"111111110",
  21356=>"100110110",
  21357=>"110111000",
  21358=>"111110111",
  21359=>"000001001",
  21360=>"000000001",
  21361=>"110000000",
  21362=>"111101111",
  21363=>"000010000",
  21364=>"011110110",
  21365=>"000000101",
  21366=>"000100100",
  21367=>"111100000",
  21368=>"000001000",
  21369=>"000000101",
  21370=>"000000111",
  21371=>"111010000",
  21372=>"010010010",
  21373=>"111111111",
  21374=>"001001101",
  21375=>"001001001",
  21376=>"110110110",
  21377=>"000000010",
  21378=>"110100000",
  21379=>"101101001",
  21380=>"011000101",
  21381=>"011011011",
  21382=>"000001000",
  21383=>"111111111",
  21384=>"111111110",
  21385=>"111100000",
  21386=>"000000000",
  21387=>"010111111",
  21388=>"000011111",
  21389=>"000000000",
  21390=>"111011000",
  21391=>"110110110",
  21392=>"000000000",
  21393=>"001001001",
  21394=>"110110000",
  21395=>"010110000",
  21396=>"000001111",
  21397=>"010010010",
  21398=>"101000000",
  21399=>"001001001",
  21400=>"111101101",
  21401=>"101011000",
  21402=>"000001000",
  21403=>"000000000",
  21404=>"001000000",
  21405=>"110010000",
  21406=>"000001011",
  21407=>"111111110",
  21408=>"000000000",
  21409=>"101111111",
  21410=>"111000010",
  21411=>"101111111",
  21412=>"111110010",
  21413=>"010111111",
  21414=>"101001101",
  21415=>"110011000",
  21416=>"101101101",
  21417=>"100111111",
  21418=>"010000110",
  21419=>"000000000",
  21420=>"101111101",
  21421=>"111101001",
  21422=>"000110100",
  21423=>"000100100",
  21424=>"101101100",
  21425=>"000000000",
  21426=>"000001001",
  21427=>"010000000",
  21428=>"100001101",
  21429=>"000001011",
  21430=>"000000001",
  21431=>"111001000",
  21432=>"000001000",
  21433=>"000000010",
  21434=>"010010000",
  21435=>"111111000",
  21436=>"110100101",
  21437=>"111110110",
  21438=>"111110000",
  21439=>"100000100",
  21440=>"000000010",
  21441=>"000010011",
  21442=>"000000100",
  21443=>"001001001",
  21444=>"100001001",
  21445=>"110111100",
  21446=>"000001100",
  21447=>"111100000",
  21448=>"000000000",
  21449=>"000000111",
  21450=>"101101101",
  21451=>"001001011",
  21452=>"000000100",
  21453=>"001011011",
  21454=>"001001000",
  21455=>"000000101",
  21456=>"000010110",
  21457=>"111111011",
  21458=>"000011111",
  21459=>"111101001",
  21460=>"101101101",
  21461=>"111011011",
  21462=>"000000101",
  21463=>"011011011",
  21464=>"000001101",
  21465=>"000000000",
  21466=>"100100111",
  21467=>"000000101",
  21468=>"111100000",
  21469=>"000110010",
  21470=>"000000100",
  21471=>"100000000",
  21472=>"110000000",
  21473=>"101101100",
  21474=>"010010000",
  21475=>"111111000",
  21476=>"111111111",
  21477=>"111111011",
  21478=>"111000111",
  21479=>"000001001",
  21480=>"111111111",
  21481=>"111111111",
  21482=>"111110000",
  21483=>"111111011",
  21484=>"110000001",
  21485=>"000100100",
  21486=>"101100100",
  21487=>"001001000",
  21488=>"111111001",
  21489=>"011010110",
  21490=>"011011000",
  21491=>"000000000",
  21492=>"110000100",
  21493=>"011011011",
  21494=>"111111110",
  21495=>"110110110",
  21496=>"111011001",
  21497=>"000000000",
  21498=>"000001000",
  21499=>"101101101",
  21500=>"110110101",
  21501=>"111111111",
  21502=>"111001000",
  21503=>"001111111",
  21504=>"111101111",
  21505=>"111111111",
  21506=>"111011001",
  21507=>"100000111",
  21508=>"000110111",
  21509=>"111110110",
  21510=>"001000011",
  21511=>"000000000",
  21512=>"000000000",
  21513=>"110111111",
  21514=>"000000111",
  21515=>"001000000",
  21516=>"000100000",
  21517=>"000000001",
  21518=>"100000100",
  21519=>"111111000",
  21520=>"000000000",
  21521=>"000100101",
  21522=>"001111111",
  21523=>"111111111",
  21524=>"000000000",
  21525=>"001000000",
  21526=>"000000011",
  21527=>"111000000",
  21528=>"111111111",
  21529=>"111001000",
  21530=>"111110000",
  21531=>"000000010",
  21532=>"000110111",
  21533=>"111111111",
  21534=>"001000000",
  21535=>"111111000",
  21536=>"111111111",
  21537=>"001001011",
  21538=>"000100000",
  21539=>"000111111",
  21540=>"110111111",
  21541=>"011111111",
  21542=>"010010111",
  21543=>"000110010",
  21544=>"010111011",
  21545=>"011000000",
  21546=>"000101100",
  21547=>"100110110",
  21548=>"111111110",
  21549=>"111000000",
  21550=>"000111111",
  21551=>"000000100",
  21552=>"111111111",
  21553=>"111000000",
  21554=>"000000000",
  21555=>"111110110",
  21556=>"100100000",
  21557=>"111110010",
  21558=>"010000000",
  21559=>"011000000",
  21560=>"111100111",
  21561=>"000110111",
  21562=>"000000000",
  21563=>"000100111",
  21564=>"000000000",
  21565=>"011000000",
  21566=>"000000000",
  21567=>"000000111",
  21568=>"111111100",
  21569=>"011111100",
  21570=>"000111111",
  21571=>"111111111",
  21572=>"111111001",
  21573=>"100100110",
  21574=>"110100100",
  21575=>"111111011",
  21576=>"001001000",
  21577=>"100000111",
  21578=>"111111011",
  21579=>"000100111",
  21580=>"110000111",
  21581=>"011011000",
  21582=>"111111000",
  21583=>"000000000",
  21584=>"111111111",
  21585=>"000000111",
  21586=>"000000000",
  21587=>"101111101",
  21588=>"011111000",
  21589=>"000000010",
  21590=>"111111111",
  21591=>"111001000",
  21592=>"111100111",
  21593=>"000000000",
  21594=>"001001000",
  21595=>"110011011",
  21596=>"111000000",
  21597=>"100100000",
  21598=>"101011111",
  21599=>"111111111",
  21600=>"000000100",
  21601=>"000110111",
  21602=>"110111100",
  21603=>"000110100",
  21604=>"000001111",
  21605=>"110100110",
  21606=>"111100000",
  21607=>"100111110",
  21608=>"000000000",
  21609=>"111111111",
  21610=>"110111110",
  21611=>"001000000",
  21612=>"000000000",
  21613=>"111111111",
  21614=>"111110110",
  21615=>"000000010",
  21616=>"000010111",
  21617=>"000000010",
  21618=>"011000000",
  21619=>"000000000",
  21620=>"000000000",
  21621=>"000001001",
  21622=>"000000111",
  21623=>"111111000",
  21624=>"000010000",
  21625=>"111111001",
  21626=>"111000000",
  21627=>"111100110",
  21628=>"100110000",
  21629=>"011000000",
  21630=>"000000001",
  21631=>"111111001",
  21632=>"111100100",
  21633=>"001001111",
  21634=>"111111111",
  21635=>"000000111",
  21636=>"100111110",
  21637=>"000101111",
  21638=>"111110110",
  21639=>"000101111",
  21640=>"111000000",
  21641=>"000111111",
  21642=>"000000000",
  21643=>"000100110",
  21644=>"011000000",
  21645=>"011010110",
  21646=>"111110000",
  21647=>"111111000",
  21648=>"000000000",
  21649=>"101001011",
  21650=>"000000000",
  21651=>"111111111",
  21652=>"000000000",
  21653=>"111010010",
  21654=>"110000000",
  21655=>"000000000",
  21656=>"000000000",
  21657=>"000000100",
  21658=>"011001000",
  21659=>"000111001",
  21660=>"011100110",
  21661=>"111110111",
  21662=>"000000000",
  21663=>"000000100",
  21664=>"000000000",
  21665=>"111000000",
  21666=>"000100111",
  21667=>"111011111",
  21668=>"110010001",
  21669=>"000111111",
  21670=>"110100000",
  21671=>"000000000",
  21672=>"000000111",
  21673=>"000000111",
  21674=>"111111101",
  21675=>"100000111",
  21676=>"000000000",
  21677=>"111000000",
  21678=>"011000000",
  21679=>"101111111",
  21680=>"000000111",
  21681=>"111011001",
  21682=>"111111000",
  21683=>"111111111",
  21684=>"000000111",
  21685=>"111000111",
  21686=>"111010000",
  21687=>"000001101",
  21688=>"011011111",
  21689=>"000000000",
  21690=>"111011111",
  21691=>"011011011",
  21692=>"011111000",
  21693=>"000000000",
  21694=>"111100111",
  21695=>"001101000",
  21696=>"100110110",
  21697=>"110111111",
  21698=>"000000000",
  21699=>"011111000",
  21700=>"000000000",
  21701=>"000000000",
  21702=>"000001000",
  21703=>"111111010",
  21704=>"000000010",
  21705=>"111111111",
  21706=>"111111110",
  21707=>"111111111",
  21708=>"111111100",
  21709=>"000000000",
  21710=>"000111111",
  21711=>"100100111",
  21712=>"100100000",
  21713=>"100000000",
  21714=>"000111111",
  21715=>"001001000",
  21716=>"111110000",
  21717=>"001010110",
  21718=>"100000000",
  21719=>"100000111",
  21720=>"000000111",
  21721=>"000101101",
  21722=>"111111111",
  21723=>"111111111",
  21724=>"110000011",
  21725=>"101100111",
  21726=>"111111111",
  21727=>"011011000",
  21728=>"000110000",
  21729=>"111111000",
  21730=>"111110000",
  21731=>"001000110",
  21732=>"010000000",
  21733=>"111110110",
  21734=>"111111111",
  21735=>"111111100",
  21736=>"111111111",
  21737=>"101100110",
  21738=>"111100111",
  21739=>"111001000",
  21740=>"001111111",
  21741=>"000110000",
  21742=>"110100110",
  21743=>"111011011",
  21744=>"110000000",
  21745=>"111100000",
  21746=>"111111111",
  21747=>"011011111",
  21748=>"000110111",
  21749=>"101101001",
  21750=>"111111011",
  21751=>"000000000",
  21752=>"110110100",
  21753=>"010011000",
  21754=>"111100000",
  21755=>"000111001",
  21756=>"100000000",
  21757=>"000000000",
  21758=>"011000111",
  21759=>"000000000",
  21760=>"000000000",
  21761=>"000000000",
  21762=>"000001000",
  21763=>"000001111",
  21764=>"100111111",
  21765=>"111011000",
  21766=>"000000000",
  21767=>"000110111",
  21768=>"011000111",
  21769=>"100100111",
  21770=>"111111111",
  21771=>"111101111",
  21772=>"100100100",
  21773=>"101101111",
  21774=>"111111111",
  21775=>"000101111",
  21776=>"111000000",
  21777=>"101000000",
  21778=>"000000000",
  21779=>"011000000",
  21780=>"111000000",
  21781=>"111100100",
  21782=>"011011010",
  21783=>"000001000",
  21784=>"111111111",
  21785=>"111111000",
  21786=>"111111000",
  21787=>"111001011",
  21788=>"000110111",
  21789=>"111000000",
  21790=>"111111100",
  21791=>"111000001",
  21792=>"000001001",
  21793=>"100000001",
  21794=>"000000111",
  21795=>"111011000",
  21796=>"111110000",
  21797=>"111111111",
  21798=>"110111111",
  21799=>"000000000",
  21800=>"101000000",
  21801=>"000101111",
  21802=>"000000000",
  21803=>"000000000",
  21804=>"001010011",
  21805=>"000000010",
  21806=>"111100111",
  21807=>"000000000",
  21808=>"001110100",
  21809=>"001011000",
  21810=>"101000000",
  21811=>"100000000",
  21812=>"111000000",
  21813=>"111111111",
  21814=>"111000010",
  21815=>"111000000",
  21816=>"000000000",
  21817=>"000000111",
  21818=>"001011011",
  21819=>"101110100",
  21820=>"001000000",
  21821=>"001000000",
  21822=>"111111111",
  21823=>"111011001",
  21824=>"000110111",
  21825=>"000000000",
  21826=>"000000110",
  21827=>"000000100",
  21828=>"000000111",
  21829=>"111111111",
  21830=>"111110111",
  21831=>"000110111",
  21832=>"111111000",
  21833=>"010110111",
  21834=>"100111111",
  21835=>"101111111",
  21836=>"011111111",
  21837=>"111011000",
  21838=>"000010010",
  21839=>"100101100",
  21840=>"111111000",
  21841=>"111111111",
  21842=>"001011111",
  21843=>"001000000",
  21844=>"000000000",
  21845=>"000011011",
  21846=>"000111111",
  21847=>"111100111",
  21848=>"000110110",
  21849=>"000000000",
  21850=>"111000000",
  21851=>"111111111",
  21852=>"000000000",
  21853=>"000000000",
  21854=>"000011001",
  21855=>"001001000",
  21856=>"000000000",
  21857=>"111100001",
  21858=>"100000000",
  21859=>"101101111",
  21860=>"111000000",
  21861=>"000000000",
  21862=>"111111111",
  21863=>"100110110",
  21864=>"110111111",
  21865=>"000000111",
  21866=>"101001000",
  21867=>"000000000",
  21868=>"101001000",
  21869=>"000001111",
  21870=>"011111111",
  21871=>"000000000",
  21872=>"010010011",
  21873=>"111000111",
  21874=>"010000001",
  21875=>"111110100",
  21876=>"111111100",
  21877=>"000000101",
  21878=>"000100111",
  21879=>"000000000",
  21880=>"000000000",
  21881=>"111111000",
  21882=>"000001011",
  21883=>"111000000",
  21884=>"111001111",
  21885=>"000000001",
  21886=>"111110110",
  21887=>"111111111",
  21888=>"000111111",
  21889=>"000000111",
  21890=>"111111101",
  21891=>"000001011",
  21892=>"111111111",
  21893=>"110111110",
  21894=>"000111000",
  21895=>"111101000",
  21896=>"000000000",
  21897=>"011011111",
  21898=>"111000001",
  21899=>"000110111",
  21900=>"111111111",
  21901=>"000000000",
  21902=>"100000000",
  21903=>"111100110",
  21904=>"000000000",
  21905=>"111111110",
  21906=>"111101101",
  21907=>"001000000",
  21908=>"001111111",
  21909=>"111001000",
  21910=>"000000000",
  21911=>"110110111",
  21912=>"111000000",
  21913=>"000000111",
  21914=>"000000111",
  21915=>"011111111",
  21916=>"000001111",
  21917=>"000000111",
  21918=>"000000010",
  21919=>"111111111",
  21920=>"111101000",
  21921=>"001010000",
  21922=>"000000000",
  21923=>"111111111",
  21924=>"101101101",
  21925=>"110000000",
  21926=>"100100100",
  21927=>"001111111",
  21928=>"010111100",
  21929=>"100000000",
  21930=>"000000000",
  21931=>"001001010",
  21932=>"111111000",
  21933=>"111110000",
  21934=>"111111111",
  21935=>"111111111",
  21936=>"000000000",
  21937=>"101000000",
  21938=>"001011111",
  21939=>"000101000",
  21940=>"000000111",
  21941=>"111000111",
  21942=>"010110110",
  21943=>"100000000",
  21944=>"000010011",
  21945=>"000010011",
  21946=>"001000000",
  21947=>"000111111",
  21948=>"000000000",
  21949=>"100000111",
  21950=>"111000000",
  21951=>"010010010",
  21952=>"011001000",
  21953=>"000000000",
  21954=>"111111011",
  21955=>"000000000",
  21956=>"000000111",
  21957=>"000000110",
  21958=>"000111111",
  21959=>"100111110",
  21960=>"000111111",
  21961=>"000000000",
  21962=>"100000000",
  21963=>"000000000",
  21964=>"111111000",
  21965=>"000000000",
  21966=>"100000000",
  21967=>"111111111",
  21968=>"100000010",
  21969=>"000100100",
  21970=>"000001111",
  21971=>"001000011",
  21972=>"100110000",
  21973=>"111111111",
  21974=>"000000011",
  21975=>"000000000",
  21976=>"100110100",
  21977=>"000000111",
  21978=>"000011111",
  21979=>"001000000",
  21980=>"000000000",
  21981=>"001001011",
  21982=>"000001000",
  21983=>"000001011",
  21984=>"000111111",
  21985=>"100100101",
  21986=>"111111000",
  21987=>"111000000",
  21988=>"000000010",
  21989=>"111001000",
  21990=>"011000011",
  21991=>"111001000",
  21992=>"111111111",
  21993=>"011010000",
  21994=>"101111011",
  21995=>"000110110",
  21996=>"110111111",
  21997=>"001000000",
  21998=>"000000001",
  21999=>"000000010",
  22000=>"001011111",
  22001=>"111111100",
  22002=>"000000000",
  22003=>"000000000",
  22004=>"000000111",
  22005=>"000000000",
  22006=>"010000000",
  22007=>"100000111",
  22008=>"111111000",
  22009=>"101000000",
  22010=>"110110011",
  22011=>"111100100",
  22012=>"000010111",
  22013=>"000011010",
  22014=>"000001000",
  22015=>"101001100",
  22016=>"000000000",
  22017=>"000000000",
  22018=>"111111000",
  22019=>"000000000",
  22020=>"000000000",
  22021=>"111111111",
  22022=>"110111100",
  22023=>"000000000",
  22024=>"000000111",
  22025=>"000001101",
  22026=>"000000000",
  22027=>"111000011",
  22028=>"000010100",
  22029=>"000000101",
  22030=>"101111111",
  22031=>"000000100",
  22032=>"111110111",
  22033=>"110111101",
  22034=>"000000000",
  22035=>"111111111",
  22036=>"111111000",
  22037=>"000000001",
  22038=>"010010010",
  22039=>"011000111",
  22040=>"001001000",
  22041=>"010000000",
  22042=>"111111001",
  22043=>"011001111",
  22044=>"000010011",
  22045=>"000000000",
  22046=>"001111111",
  22047=>"000000000",
  22048=>"011000100",
  22049=>"111110000",
  22050=>"001111111",
  22051=>"000000000",
  22052=>"000100100",
  22053=>"111111111",
  22054=>"000000000",
  22055=>"111111110",
  22056=>"100000001",
  22057=>"111111111",
  22058=>"000000000",
  22059=>"001111111",
  22060=>"111111111",
  22061=>"000100000",
  22062=>"111111111",
  22063=>"000000000",
  22064=>"000000000",
  22065=>"111111110",
  22066=>"010011011",
  22067=>"000000000",
  22068=>"100100110",
  22069=>"000100100",
  22070=>"010000000",
  22071=>"000000100",
  22072=>"000111111",
  22073=>"000000000",
  22074=>"111111111",
  22075=>"000000000",
  22076=>"111111111",
  22077=>"000000100",
  22078=>"111111000",
  22079=>"111111111",
  22080=>"000100000",
  22081=>"000000000",
  22082=>"111111111",
  22083=>"111111111",
  22084=>"111001000",
  22085=>"111111100",
  22086=>"000000000",
  22087=>"000000111",
  22088=>"111111111",
  22089=>"100111111",
  22090=>"111000000",
  22091=>"111111111",
  22092=>"100110100",
  22093=>"111111100",
  22094=>"111111111",
  22095=>"111111000",
  22096=>"000111111",
  22097=>"011011000",
  22098=>"000000000",
  22099=>"111011000",
  22100=>"111111111",
  22101=>"000000110",
  22102=>"100000000",
  22103=>"100011101",
  22104=>"000000001",
  22105=>"000000111",
  22106=>"011111111",
  22107=>"000000000",
  22108=>"000000000",
  22109=>"111111000",
  22110=>"111111001",
  22111=>"111110110",
  22112=>"000000111",
  22113=>"111111111",
  22114=>"000000000",
  22115=>"111111111",
  22116=>"000000000",
  22117=>"000111111",
  22118=>"001000000",
  22119=>"111111111",
  22120=>"001011000",
  22121=>"110111111",
  22122=>"001000000",
  22123=>"001111110",
  22124=>"111111111",
  22125=>"000000000",
  22126=>"111111101",
  22127=>"111111111",
  22128=>"000111111",
  22129=>"001000000",
  22130=>"111111111",
  22131=>"100100111",
  22132=>"100100100",
  22133=>"000000000",
  22134=>"000011111",
  22135=>"010000000",
  22136=>"000111100",
  22137=>"000011001",
  22138=>"111110100",
  22139=>"001000000",
  22140=>"000100100",
  22141=>"101000100",
  22142=>"111010000",
  22143=>"111111010",
  22144=>"000010000",
  22145=>"000000000",
  22146=>"111111111",
  22147=>"001111101",
  22148=>"000100111",
  22149=>"111111110",
  22150=>"100100000",
  22151=>"000011000",
  22152=>"000000000",
  22153=>"000000110",
  22154=>"000000000",
  22155=>"000111111",
  22156=>"000000011",
  22157=>"000000000",
  22158=>"001110000",
  22159=>"111111111",
  22160=>"101100111",
  22161=>"111111111",
  22162=>"000000000",
  22163=>"000000110",
  22164=>"000000000",
  22165=>"111111111",
  22166=>"011011001",
  22167=>"111111110",
  22168=>"000000000",
  22169=>"111000111",
  22170=>"110110111",
  22171=>"000000000",
  22172=>"011111111",
  22173=>"100000000",
  22174=>"111101111",
  22175=>"100100000",
  22176=>"001001000",
  22177=>"111111001",
  22178=>"111111111",
  22179=>"000100110",
  22180=>"000000100",
  22181=>"111111100",
  22182=>"111111111",
  22183=>"010000000",
  22184=>"000000000",
  22185=>"010001000",
  22186=>"000000100",
  22187=>"000000000",
  22188=>"110111111",
  22189=>"000000000",
  22190=>"111111111",
  22191=>"101011000",
  22192=>"000010010",
  22193=>"110110110",
  22194=>"101111011",
  22195=>"000000000",
  22196=>"000100110",
  22197=>"010011011",
  22198=>"000000000",
  22199=>"000000000",
  22200=>"111111111",
  22201=>"000000111",
  22202=>"000100100",
  22203=>"111110111",
  22204=>"000000011",
  22205=>"111111000",
  22206=>"101000000",
  22207=>"110111011",
  22208=>"000000000",
  22209=>"000100100",
  22210=>"000100110",
  22211=>"000000000",
  22212=>"111111111",
  22213=>"000000000",
  22214=>"001001000",
  22215=>"000000001",
  22216=>"111111111",
  22217=>"000110000",
  22218=>"000011111",
  22219=>"000000000",
  22220=>"000000000",
  22221=>"000010111",
  22222=>"110100111",
  22223=>"111010000",
  22224=>"110100000",
  22225=>"111111111",
  22226=>"010000010",
  22227=>"000000000",
  22228=>"000000000",
  22229=>"000001111",
  22230=>"111011000",
  22231=>"111110101",
  22232=>"000000000",
  22233=>"111100111",
  22234=>"001000000",
  22235=>"010011000",
  22236=>"000001100",
  22237=>"111000000",
  22238=>"000011001",
  22239=>"111100000",
  22240=>"000000000",
  22241=>"000000011",
  22242=>"111000000",
  22243=>"011001111",
  22244=>"110111111",
  22245=>"111111001",
  22246=>"000111001",
  22247=>"000000000",
  22248=>"000000000",
  22249=>"111111111",
  22250=>"101111111",
  22251=>"000000001",
  22252=>"000000000",
  22253=>"000000000",
  22254=>"000101111",
  22255=>"001001111",
  22256=>"111011111",
  22257=>"001100101",
  22258=>"111111111",
  22259=>"001111111",
  22260=>"111110100",
  22261=>"111111111",
  22262=>"011011011",
  22263=>"000111111",
  22264=>"111101111",
  22265=>"001000000",
  22266=>"000000101",
  22267=>"111111110",
  22268=>"100001001",
  22269=>"101101111",
  22270=>"000000100",
  22271=>"000000100",
  22272=>"001101111",
  22273=>"000010011",
  22274=>"110110111",
  22275=>"000000000",
  22276=>"111111111",
  22277=>"001001000",
  22278=>"111111111",
  22279=>"000000000",
  22280=>"000110111",
  22281=>"111111111",
  22282=>"000000000",
  22283=>"100111111",
  22284=>"111111111",
  22285=>"100000100",
  22286=>"111111011",
  22287=>"111111110",
  22288=>"111111111",
  22289=>"100100101",
  22290=>"111111100",
  22291=>"000000000",
  22292=>"011111111",
  22293=>"111111111",
  22294=>"011001000",
  22295=>"000000000",
  22296=>"101111110",
  22297=>"000000000",
  22298=>"101111111",
  22299=>"000000000",
  22300=>"100100111",
  22301=>"000000000",
  22302=>"011000000",
  22303=>"000111100",
  22304=>"100110000",
  22305=>"001111011",
  22306=>"101001001",
  22307=>"001001011",
  22308=>"011110110",
  22309=>"000000000",
  22310=>"111111111",
  22311=>"000011110",
  22312=>"100100100",
  22313=>"000000110",
  22314=>"000000000",
  22315=>"011001111",
  22316=>"111111111",
  22317=>"000111111",
  22318=>"000100000",
  22319=>"100100000",
  22320=>"000000010",
  22321=>"000110111",
  22322=>"110111111",
  22323=>"111111011",
  22324=>"000001000",
  22325=>"000000000",
  22326=>"100110000",
  22327=>"000000000",
  22328=>"011001000",
  22329=>"111111111",
  22330=>"111111111",
  22331=>"111111111",
  22332=>"110100000",
  22333=>"111111111",
  22334=>"100110110",
  22335=>"110110111",
  22336=>"001001110",
  22337=>"100111111",
  22338=>"000000000",
  22339=>"110110111",
  22340=>"000000111",
  22341=>"001101111",
  22342=>"000000000",
  22343=>"000001111",
  22344=>"000100100",
  22345=>"000000100",
  22346=>"001000000",
  22347=>"100000000",
  22348=>"010100110",
  22349=>"000000000",
  22350=>"111111101",
  22351=>"111111111",
  22352=>"110111000",
  22353=>"111111111",
  22354=>"111111111",
  22355=>"000000100",
  22356=>"111111011",
  22357=>"011011011",
  22358=>"111111111",
  22359=>"000000000",
  22360=>"101101111",
  22361=>"000101100",
  22362=>"001100111",
  22363=>"000000000",
  22364=>"000000000",
  22365=>"000100100",
  22366=>"111111111",
  22367=>"000100001",
  22368=>"000000000",
  22369=>"000000000",
  22370=>"000000111",
  22371=>"110000000",
  22372=>"111111111",
  22373=>"000000000",
  22374=>"000000000",
  22375=>"010000110",
  22376=>"000000000",
  22377=>"111000000",
  22378=>"000000000",
  22379=>"000000000",
  22380=>"100100100",
  22381=>"000000111",
  22382=>"000000010",
  22383=>"111100111",
  22384=>"000100100",
  22385=>"000000000",
  22386=>"000000000",
  22387=>"110000000",
  22388=>"111111100",
  22389=>"000000000",
  22390=>"000000001",
  22391=>"000000000",
  22392=>"111111000",
  22393=>"000001001",
  22394=>"100100100",
  22395=>"110111111",
  22396=>"111111110",
  22397=>"111111111",
  22398=>"111111111",
  22399=>"111111111",
  22400=>"000000000",
  22401=>"000110111",
  22402=>"100100111",
  22403=>"000000000",
  22404=>"000000000",
  22405=>"000000000",
  22406=>"111111110",
  22407=>"000000100",
  22408=>"000101111",
  22409=>"000000000",
  22410=>"000000101",
  22411=>"111111010",
  22412=>"111111111",
  22413=>"000000001",
  22414=>"000011001",
  22415=>"000000000",
  22416=>"101101101",
  22417=>"000000001",
  22418=>"001011001",
  22419=>"000000001",
  22420=>"000000000",
  22421=>"000000010",
  22422=>"000000100",
  22423=>"100001000",
  22424=>"000011000",
  22425=>"111100110",
  22426=>"000000000",
  22427=>"100000000",
  22428=>"111111111",
  22429=>"011000010",
  22430=>"000000000",
  22431=>"001111111",
  22432=>"100111001",
  22433=>"010011011",
  22434=>"001100100",
  22435=>"111000111",
  22436=>"100101101",
  22437=>"000000010",
  22438=>"000100111",
  22439=>"110111011",
  22440=>"101101100",
  22441=>"111010100",
  22442=>"000000111",
  22443=>"000000000",
  22444=>"000000001",
  22445=>"100100111",
  22446=>"000000111",
  22447=>"111111111",
  22448=>"000000000",
  22449=>"000011111",
  22450=>"110000000",
  22451=>"101111111",
  22452=>"000000000",
  22453=>"000000000",
  22454=>"111111111",
  22455=>"111111000",
  22456=>"111111000",
  22457=>"111111111",
  22458=>"000001111",
  22459=>"100100100",
  22460=>"111111111",
  22461=>"100000110",
  22462=>"111101100",
  22463=>"010010000",
  22464=>"101000000",
  22465=>"011111000",
  22466=>"000000111",
  22467=>"000000000",
  22468=>"000100111",
  22469=>"001001001",
  22470=>"111111000",
  22471=>"010011011",
  22472=>"000000000",
  22473=>"001001100",
  22474=>"001111111",
  22475=>"000011000",
  22476=>"111110000",
  22477=>"000000000",
  22478=>"000000100",
  22479=>"000000001",
  22480=>"000000000",
  22481=>"000111111",
  22482=>"000000110",
  22483=>"000000000",
  22484=>"111111111",
  22485=>"001011111",
  22486=>"111001000",
  22487=>"000000111",
  22488=>"111111111",
  22489=>"111111111",
  22490=>"000000111",
  22491=>"111111111",
  22492=>"000010001",
  22493=>"001001001",
  22494=>"000000001",
  22495=>"000000000",
  22496=>"011001100",
  22497=>"000100110",
  22498=>"111111000",
  22499=>"111111110",
  22500=>"111101111",
  22501=>"001001101",
  22502=>"111111111",
  22503=>"000000000",
  22504=>"111111000",
  22505=>"011111111",
  22506=>"000000001",
  22507=>"111111111",
  22508=>"000000000",
  22509=>"111000000",
  22510=>"001000000",
  22511=>"101101101",
  22512=>"100000000",
  22513=>"111111111",
  22514=>"111100100",
  22515=>"001001000",
  22516=>"111111011",
  22517=>"000000000",
  22518=>"000110111",
  22519=>"000000000",
  22520=>"111111111",
  22521=>"001001000",
  22522=>"100000000",
  22523=>"000000000",
  22524=>"000000000",
  22525=>"000000000",
  22526=>"111000000",
  22527=>"000000000",
  22528=>"110111000",
  22529=>"000000000",
  22530=>"000000111",
  22531=>"100101000",
  22532=>"000000001",
  22533=>"000000111",
  22534=>"000000001",
  22535=>"111111111",
  22536=>"000000000",
  22537=>"111101101",
  22538=>"000000001",
  22539=>"111111110",
  22540=>"001101101",
  22541=>"100000000",
  22542=>"110111001",
  22543=>"000000011",
  22544=>"111001100",
  22545=>"000110100",
  22546=>"111111110",
  22547=>"110111110",
  22548=>"111111111",
  22549=>"001001001",
  22550=>"100111111",
  22551=>"111111001",
  22552=>"111111000",
  22553=>"011000010",
  22554=>"111001000",
  22555=>"001000110",
  22556=>"111000000",
  22557=>"111111111",
  22558=>"011001111",
  22559=>"111100000",
  22560=>"000000111",
  22561=>"111100000",
  22562=>"001000000",
  22563=>"111011111",
  22564=>"000000000",
  22565=>"000000100",
  22566=>"000100111",
  22567=>"111111110",
  22568=>"101111111",
  22569=>"011001001",
  22570=>"111111111",
  22571=>"011110111",
  22572=>"111111100",
  22573=>"111111100",
  22574=>"111111111",
  22575=>"000000000",
  22576=>"000001111",
  22577=>"000000000",
  22578=>"000000000",
  22579=>"000000011",
  22580=>"110111101",
  22581=>"011011111",
  22582=>"001001011",
  22583=>"001000001",
  22584=>"000000000",
  22585=>"001001001",
  22586=>"000000111",
  22587=>"111111110",
  22588=>"100000000",
  22589=>"000110111",
  22590=>"000000100",
  22591=>"001100101",
  22592=>"011111100",
  22593=>"000100111",
  22594=>"000000000",
  22595=>"111111000",
  22596=>"000111111",
  22597=>"111100000",
  22598=>"111111110",
  22599=>"000000001",
  22600=>"111111111",
  22601=>"110111110",
  22602=>"111101111",
  22603=>"111000111",
  22604=>"000101000",
  22605=>"111111111",
  22606=>"000000000",
  22607=>"111010111",
  22608=>"000111111",
  22609=>"000001000",
  22610=>"011111110",
  22611=>"011011111",
  22612=>"011000111",
  22613=>"100000000",
  22614=>"001001000",
  22615=>"010000101",
  22616=>"000000000",
  22617=>"111001000",
  22618=>"111111000",
  22619=>"111001001",
  22620=>"000001111",
  22621=>"111011000",
  22622=>"000100111",
  22623=>"011111110",
  22624=>"000111100",
  22625=>"110111111",
  22626=>"001011011",
  22627=>"000001000",
  22628=>"111111011",
  22629=>"000010111",
  22630=>"000000000",
  22631=>"111111111",
  22632=>"111111111",
  22633=>"100000000",
  22634=>"101001111",
  22635=>"110001001",
  22636=>"010011011",
  22637=>"111111110",
  22638=>"111111000",
  22639=>"110111000",
  22640=>"000000000",
  22641=>"000000111",
  22642=>"101111110",
  22643=>"001011011",
  22644=>"000000000",
  22645=>"000000000",
  22646=>"100000000",
  22647=>"000000000",
  22648=>"000000000",
  22649=>"111100111",
  22650=>"111111111",
  22651=>"000000000",
  22652=>"010110110",
  22653=>"000111111",
  22654=>"011000000",
  22655=>"000011111",
  22656=>"111111000",
  22657=>"000000111",
  22658=>"111111111",
  22659=>"110100011",
  22660=>"000000111",
  22661=>"000001111",
  22662=>"000111000",
  22663=>"111111000",
  22664=>"111111111",
  22665=>"000000011",
  22666=>"000000011",
  22667=>"000111111",
  22668=>"000000000",
  22669=>"001000000",
  22670=>"000100100",
  22671=>"000000000",
  22672=>"011000000",
  22673=>"000001111",
  22674=>"000000001",
  22675=>"000000010",
  22676=>"001001111",
  22677=>"111111000",
  22678=>"111111011",
  22679=>"111000000",
  22680=>"001101111",
  22681=>"000000000",
  22682=>"000101000",
  22683=>"000000000",
  22684=>"000000001",
  22685=>"000000000",
  22686=>"000110000",
  22687=>"000000010",
  22688=>"001111000",
  22689=>"111011111",
  22690=>"111000000",
  22691=>"000000000",
  22692=>"000011011",
  22693=>"111111000",
  22694=>"111000000",
  22695=>"000111001",
  22696=>"111000110",
  22697=>"000000000",
  22698=>"111111111",
  22699=>"000100000",
  22700=>"111111000",
  22701=>"000111001",
  22702=>"000111111",
  22703=>"111111011",
  22704=>"111000000",
  22705=>"100100000",
  22706=>"111111111",
  22707=>"000000101",
  22708=>"000100100",
  22709=>"000000000",
  22710=>"000000110",
  22711=>"110111111",
  22712=>"111111111",
  22713=>"111000101",
  22714=>"000000011",
  22715=>"111111000",
  22716=>"000000000",
  22717=>"111111000",
  22718=>"111000000",
  22719=>"001011111",
  22720=>"000000000",
  22721=>"000000000",
  22722=>"000001111",
  22723=>"111111000",
  22724=>"110000100",
  22725=>"000000001",
  22726=>"000000001",
  22727=>"100101111",
  22728=>"111000000",
  22729=>"111110111",
  22730=>"000100000",
  22731=>"000111111",
  22732=>"111111110",
  22733=>"111111000",
  22734=>"111000000",
  22735=>"111111111",
  22736=>"111111011",
  22737=>"000111010",
  22738=>"110000000",
  22739=>"000000000",
  22740=>"001011000",
  22741=>"111111000",
  22742=>"111111000",
  22743=>"000000000",
  22744=>"000000001",
  22745=>"101000100",
  22746=>"000111111",
  22747=>"000111000",
  22748=>"000000000",
  22749=>"111110000",
  22750=>"111111111",
  22751=>"000000111",
  22752=>"111111111",
  22753=>"111001111",
  22754=>"000000000",
  22755=>"001000000",
  22756=>"111111000",
  22757=>"111100100",
  22758=>"111111111",
  22759=>"110110111",
  22760=>"111111000",
  22761=>"010011000",
  22762=>"001110111",
  22763=>"001011111",
  22764=>"001011000",
  22765=>"111000000",
  22766=>"111111111",
  22767=>"000000111",
  22768=>"111111011",
  22769=>"001011011",
  22770=>"111111111",
  22771=>"000000111",
  22772=>"010111111",
  22773=>"000000011",
  22774=>"000000010",
  22775=>"000000100",
  22776=>"000000110",
  22777=>"000000000",
  22778=>"001001011",
  22779=>"101000000",
  22780=>"000001111",
  22781=>"111111001",
  22782=>"000001001",
  22783=>"000010111",
  22784=>"000000111",
  22785=>"111001001",
  22786=>"000000000",
  22787=>"000000000",
  22788=>"000000001",
  22789=>"000000000",
  22790=>"111011111",
  22791=>"000000001",
  22792=>"000111111",
  22793=>"111111000",
  22794=>"110111000",
  22795=>"100000010",
  22796=>"111111111",
  22797=>"000000111",
  22798=>"000000000",
  22799=>"000111111",
  22800=>"111110000",
  22801=>"111100000",
  22802=>"111111111",
  22803=>"000100110",
  22804=>"000111000",
  22805=>"000000011",
  22806=>"011000000",
  22807=>"000100110",
  22808=>"110110111",
  22809=>"000000000",
  22810=>"000001111",
  22811=>"000000000",
  22812=>"000111111",
  22813=>"011000000",
  22814=>"111111000",
  22815=>"011111111",
  22816=>"111111010",
  22817=>"000000000",
  22818=>"000000111",
  22819=>"000000000",
  22820=>"111010000",
  22821=>"000110111",
  22822=>"100101000",
  22823=>"000111111",
  22824=>"100111000",
  22825=>"000000100",
  22826=>"101100111",
  22827=>"000000111",
  22828=>"111111111",
  22829=>"100110101",
  22830=>"000000000",
  22831=>"000000000",
  22832=>"111111111",
  22833=>"000001111",
  22834=>"111111010",
  22835=>"011111111",
  22836=>"011000110",
  22837=>"101000000",
  22838=>"000000101",
  22839=>"000000110",
  22840=>"100100000",
  22841=>"100000000",
  22842=>"111011000",
  22843=>"000111000",
  22844=>"000000000",
  22845=>"111111100",
  22846=>"000010111",
  22847=>"000111111",
  22848=>"000000111",
  22849=>"001001000",
  22850=>"111111111",
  22851=>"111000000",
  22852=>"111111111",
  22853=>"111110000",
  22854=>"000000000",
  22855=>"000000110",
  22856=>"000001001",
  22857=>"101000000",
  22858=>"000111100",
  22859=>"000001111",
  22860=>"100000011",
  22861=>"100101111",
  22862=>"000101111",
  22863=>"010010011",
  22864=>"000010110",
  22865=>"000000000",
  22866=>"000110111",
  22867=>"001011111",
  22868=>"000100111",
  22869=>"011111111",
  22870=>"001011001",
  22871=>"111000000",
  22872=>"111100111",
  22873=>"000001000",
  22874=>"100000100",
  22875=>"111011010",
  22876=>"000011000",
  22877=>"111111111",
  22878=>"000001100",
  22879=>"001110100",
  22880=>"000000000",
  22881=>"111111111",
  22882=>"000000111",
  22883=>"111000000",
  22884=>"000000000",
  22885=>"000000111",
  22886=>"111111111",
  22887=>"111110110",
  22888=>"000110111",
  22889=>"010000000",
  22890=>"111101011",
  22891=>"000100110",
  22892=>"000110111",
  22893=>"000000111",
  22894=>"000110111",
  22895=>"111110000",
  22896=>"000011111",
  22897=>"000001010",
  22898=>"111110000",
  22899=>"110100100",
  22900=>"110000000",
  22901=>"000100100",
  22902=>"000000000",
  22903=>"000000111",
  22904=>"111000000",
  22905=>"000000000",
  22906=>"011000111",
  22907=>"000111111",
  22908=>"111111111",
  22909=>"001000000",
  22910=>"000000000",
  22911=>"111000000",
  22912=>"110110000",
  22913=>"111000000",
  22914=>"111001000",
  22915=>"111110000",
  22916=>"000000000",
  22917=>"000000001",
  22918=>"000000000",
  22919=>"111111011",
  22920=>"111111110",
  22921=>"000000111",
  22922=>"000000000",
  22923=>"000000111",
  22924=>"111000111",
  22925=>"010000000",
  22926=>"000000000",
  22927=>"001001001",
  22928=>"101111111",
  22929=>"111000110",
  22930=>"000011010",
  22931=>"000000000",
  22932=>"000100000",
  22933=>"000011111",
  22934=>"111000001",
  22935=>"000001111",
  22936=>"111100110",
  22937=>"000000000",
  22938=>"100000000",
  22939=>"000111111",
  22940=>"000100111",
  22941=>"011111111",
  22942=>"000000111",
  22943=>"000001001",
  22944=>"000000000",
  22945=>"000111111",
  22946=>"000000000",
  22947=>"001010010",
  22948=>"000000000",
  22949=>"100111111",
  22950=>"000000001",
  22951=>"000111111",
  22952=>"000101000",
  22953=>"101000011",
  22954=>"001011011",
  22955=>"000011000",
  22956=>"001001001",
  22957=>"011001000",
  22958=>"001111111",
  22959=>"000000000",
  22960=>"111111000",
  22961=>"110000101",
  22962=>"110111111",
  22963=>"000000111",
  22964=>"111110000",
  22965=>"101000000",
  22966=>"100100100",
  22967=>"111111111",
  22968=>"101000111",
  22969=>"000000111",
  22970=>"000000001",
  22971=>"110000000",
  22972=>"111111000",
  22973=>"111111100",
  22974=>"101111000",
  22975=>"011111011",
  22976=>"101101111",
  22977=>"111111100",
  22978=>"111111111",
  22979=>"000000001",
  22980=>"101111111",
  22981=>"111111000",
  22982=>"111111101",
  22983=>"000000000",
  22984=>"101111111",
  22985=>"111111111",
  22986=>"000000111",
  22987=>"010111000",
  22988=>"100110000",
  22989=>"000000000",
  22990=>"110000000",
  22991=>"111011111",
  22992=>"111111111",
  22993=>"111100000",
  22994=>"111111111",
  22995=>"111111111",
  22996=>"101100100",
  22997=>"111001000",
  22998=>"000100010",
  22999=>"100100011",
  23000=>"000101000",
  23001=>"000111111",
  23002=>"100011011",
  23003=>"000000000",
  23004=>"000111111",
  23005=>"111110000",
  23006=>"001111111",
  23007=>"001001000",
  23008=>"011000000",
  23009=>"000000101",
  23010=>"001000000",
  23011=>"101100000",
  23012=>"000000000",
  23013=>"111111000",
  23014=>"001001011",
  23015=>"000000111",
  23016=>"110111111",
  23017=>"111111000",
  23018=>"110110001",
  23019=>"000110111",
  23020=>"111011111",
  23021=>"000100110",
  23022=>"111111111",
  23023=>"000000000",
  23024=>"000000111",
  23025=>"000111111",
  23026=>"101111000",
  23027=>"100110110",
  23028=>"000000110",
  23029=>"110100000",
  23030=>"111111001",
  23031=>"111111111",
  23032=>"000000000",
  23033=>"100000000",
  23034=>"010110110",
  23035=>"111111111",
  23036=>"111101111",
  23037=>"011111111",
  23038=>"111000101",
  23039=>"111000000",
  23040=>"110111111",
  23041=>"000000000",
  23042=>"000110111",
  23043=>"000000010",
  23044=>"110101111",
  23045=>"101111111",
  23046=>"001001000",
  23047=>"111111111",
  23048=>"000000000",
  23049=>"000000000",
  23050=>"000001111",
  23051=>"000000111",
  23052=>"000000100",
  23053=>"111111111",
  23054=>"110100111",
  23055=>"000100011",
  23056=>"111111111",
  23057=>"000000000",
  23058=>"111111111",
  23059=>"110111111",
  23060=>"010110111",
  23061=>"011000000",
  23062=>"111110010",
  23063=>"011111111",
  23064=>"011111111",
  23065=>"100101000",
  23066=>"111111101",
  23067=>"000000100",
  23068=>"111111110",
  23069=>"111111111",
  23070=>"000000000",
  23071=>"000000101",
  23072=>"000000100",
  23073=>"000110111",
  23074=>"111100110",
  23075=>"110110111",
  23076=>"111011000",
  23077=>"111100100",
  23078=>"001000111",
  23079=>"111000101",
  23080=>"111100100",
  23081=>"011111111",
  23082=>"111111001",
  23083=>"111111000",
  23084=>"000000000",
  23085=>"011111011",
  23086=>"000001000",
  23087=>"100001111",
  23088=>"000110111",
  23089=>"111111111",
  23090=>"000000000",
  23091=>"100100000",
  23092=>"000000000",
  23093=>"111111000",
  23094=>"000000001",
  23095=>"111100000",
  23096=>"111111100",
  23097=>"100000100",
  23098=>"000100000",
  23099=>"010000000",
  23100=>"111111111",
  23101=>"000000000",
  23102=>"010010000",
  23103=>"001111001",
  23104=>"001001101",
  23105=>"000000000",
  23106=>"000000000",
  23107=>"100000101",
  23108=>"000000100",
  23109=>"011110111",
  23110=>"000000100",
  23111=>"111001000",
  23112=>"100100001",
  23113=>"000000001",
  23114=>"111111111",
  23115=>"111111000",
  23116=>"000011111",
  23117=>"001001101",
  23118=>"000000000",
  23119=>"001001000",
  23120=>"000000000",
  23121=>"111111000",
  23122=>"000100100",
  23123=>"011011100",
  23124=>"111101000",
  23125=>"000000111",
  23126=>"000000111",
  23127=>"000000001",
  23128=>"110000111",
  23129=>"010000000",
  23130=>"110000110",
  23131=>"000001011",
  23132=>"000000000",
  23133=>"000000000",
  23134=>"101001111",
  23135=>"000011111",
  23136=>"111111111",
  23137=>"001111000",
  23138=>"001001000",
  23139=>"111000000",
  23140=>"001010110",
  23141=>"101000000",
  23142=>"100000111",
  23143=>"000000110",
  23144=>"111111111",
  23145=>"111110100",
  23146=>"000000000",
  23147=>"000000111",
  23148=>"000001000",
  23149=>"000100110",
  23150=>"101100111",
  23151=>"001000101",
  23152=>"110101000",
  23153=>"111011000",
  23154=>"101011011",
  23155=>"000111111",
  23156=>"000100000",
  23157=>"111111000",
  23158=>"111111111",
  23159=>"000101111",
  23160=>"000000100",
  23161=>"111000000",
  23162=>"001000000",
  23163=>"000111111",
  23164=>"101111111",
  23165=>"010000100",
  23166=>"000000000",
  23167=>"000000000",
  23168=>"111110100",
  23169=>"101111101",
  23170=>"111111000",
  23171=>"000000001",
  23172=>"000000100",
  23173=>"111100000",
  23174=>"111000001",
  23175=>"111110000",
  23176=>"111101100",
  23177=>"001001001",
  23178=>"000001011",
  23179=>"000011011",
  23180=>"000010110",
  23181=>"000000000",
  23182=>"111100101",
  23183=>"000000000",
  23184=>"111001000",
  23185=>"000101111",
  23186=>"000011011",
  23187=>"111111111",
  23188=>"111111111",
  23189=>"001001001",
  23190=>"111111000",
  23191=>"001001111",
  23192=>"011000000",
  23193=>"000000000",
  23194=>"111000000",
  23195=>"000111011",
  23196=>"000000000",
  23197=>"111110111",
  23198=>"001111111",
  23199=>"000100000",
  23200=>"000001000",
  23201=>"111001000",
  23202=>"111000000",
  23203=>"000000000",
  23204=>"101000000",
  23205=>"111111000",
  23206=>"111111000",
  23207=>"110110100",
  23208=>"000000000",
  23209=>"000000000",
  23210=>"000000101",
  23211=>"000111111",
  23212=>"000000011",
  23213=>"000100100",
  23214=>"000001111",
  23215=>"000000000",
  23216=>"100110000",
  23217=>"100100100",
  23218=>"110111111",
  23219=>"111111100",
  23220=>"111000110",
  23221=>"000000001",
  23222=>"000000001",
  23223=>"001000000",
  23224=>"111111001",
  23225=>"111000100",
  23226=>"111000110",
  23227=>"001000010",
  23228=>"000000000",
  23229=>"011000000",
  23230=>"111000000",
  23231=>"111010000",
  23232=>"111111111",
  23233=>"111111000",
  23234=>"000001111",
  23235=>"111101001",
  23236=>"111111111",
  23237=>"000111111",
  23238=>"111101111",
  23239=>"000000000",
  23240=>"111001000",
  23241=>"111111000",
  23242=>"000000101",
  23243=>"011011000",
  23244=>"111110000",
  23245=>"101000111",
  23246=>"000000000",
  23247=>"111111001",
  23248=>"111000000",
  23249=>"111000000",
  23250=>"111001111",
  23251=>"000000000",
  23252=>"111101111",
  23253=>"100110111",
  23254=>"111111111",
  23255=>"000000001",
  23256=>"000000110",
  23257=>"000000101",
  23258=>"111111000",
  23259=>"111111000",
  23260=>"000011001",
  23261=>"100101100",
  23262=>"111111010",
  23263=>"000111001",
  23264=>"000000100",
  23265=>"010000011",
  23266=>"000000011",
  23267=>"111110000",
  23268=>"101111101",
  23269=>"000000110",
  23270=>"001001001",
  23271=>"011000000",
  23272=>"110111111",
  23273=>"111011000",
  23274=>"011111111",
  23275=>"000000000",
  23276=>"111111000",
  23277=>"000000001",
  23278=>"001000111",
  23279=>"000000000",
  23280=>"000110110",
  23281=>"000000001",
  23282=>"111000000",
  23283=>"101000111",
  23284=>"011001000",
  23285=>"000001001",
  23286=>"111111111",
  23287=>"000000000",
  23288=>"001000000",
  23289=>"111101000",
  23290=>"111011011",
  23291=>"010000111",
  23292=>"000001001",
  23293=>"000101001",
  23294=>"000000110",
  23295=>"111000000",
  23296=>"100111111",
  23297=>"111110000",
  23298=>"111111111",
  23299=>"000110110",
  23300=>"001001011",
  23301=>"001000000",
  23302=>"111111111",
  23303=>"000000011",
  23304=>"110101111",
  23305=>"011001111",
  23306=>"001111111",
  23307=>"101001000",
  23308=>"111110110",
  23309=>"000000000",
  23310=>"110011111",
  23311=>"000110000",
  23312=>"000000000",
  23313=>"100100001",
  23314=>"111100000",
  23315=>"001010111",
  23316=>"111111111",
  23317=>"111101101",
  23318=>"100000000",
  23319=>"000000000",
  23320=>"111111000",
  23321=>"000001111",
  23322=>"000000010",
  23323=>"000000110",
  23324=>"111110100",
  23325=>"000000111",
  23326=>"111111111",
  23327=>"000111111",
  23328=>"011001100",
  23329=>"010100111",
  23330=>"110110010",
  23331=>"111000001",
  23332=>"111111000",
  23333=>"100111011",
  23334=>"111111000",
  23335=>"111111000",
  23336=>"000000000",
  23337=>"111000000",
  23338=>"111111000",
  23339=>"111111101",
  23340=>"000000001",
  23341=>"110111111",
  23342=>"000111111",
  23343=>"111111000",
  23344=>"101011011",
  23345=>"000011011",
  23346=>"111111011",
  23347=>"111111000",
  23348=>"111111111",
  23349=>"111000001",
  23350=>"110111111",
  23351=>"000111111",
  23352=>"111111111",
  23353=>"101000000",
  23354=>"111111111",
  23355=>"110000000",
  23356=>"111100000",
  23357=>"000000000",
  23358=>"001000111",
  23359=>"111111111",
  23360=>"011111001",
  23361=>"110000100",
  23362=>"000000011",
  23363=>"111111000",
  23364=>"110100111",
  23365=>"111110000",
  23366=>"000001001",
  23367=>"000000000",
  23368=>"000011111",
  23369=>"001111111",
  23370=>"111000001",
  23371=>"111111001",
  23372=>"000001001",
  23373=>"111111000",
  23374=>"011011001",
  23375=>"011111100",
  23376=>"000001011",
  23377=>"111111111",
  23378=>"111000000",
  23379=>"111111000",
  23380=>"111001000",
  23381=>"011011011",
  23382=>"110000000",
  23383=>"001000000",
  23384=>"000001111",
  23385=>"111111111",
  23386=>"000000111",
  23387=>"001000001",
  23388=>"111111000",
  23389=>"111111000",
  23390=>"000001111",
  23391=>"110000000",
  23392=>"110000001",
  23393=>"111111000",
  23394=>"001000000",
  23395=>"111111111",
  23396=>"111110100",
  23397=>"000111001",
  23398=>"010000000",
  23399=>"110000000",
  23400=>"110111011",
  23401=>"111110000",
  23402=>"001001111",
  23403=>"000101101",
  23404=>"000010111",
  23405=>"000000111",
  23406=>"001000000",
  23407=>"000000111",
  23408=>"000000111",
  23409=>"000111111",
  23410=>"111101101",
  23411=>"100010111",
  23412=>"111000000",
  23413=>"001000000",
  23414=>"000000000",
  23415=>"001001111",
  23416=>"111111100",
  23417=>"000111000",
  23418=>"111001000",
  23419=>"001101000",
  23420=>"000000110",
  23421=>"111100000",
  23422=>"000000000",
  23423=>"111111001",
  23424=>"111001000",
  23425=>"001000000",
  23426=>"100100111",
  23427=>"000000111",
  23428=>"111110111",
  23429=>"111111111",
  23430=>"110011011",
  23431=>"111111111",
  23432=>"110000010",
  23433=>"000000000",
  23434=>"000111111",
  23435=>"111111111",
  23436=>"100000111",
  23437=>"111011000",
  23438=>"110000000",
  23439=>"111111111",
  23440=>"000000110",
  23441=>"111110100",
  23442=>"111000111",
  23443=>"111111111",
  23444=>"111111000",
  23445=>"011000000",
  23446=>"101100111",
  23447=>"111110000",
  23448=>"111111000",
  23449=>"111011001",
  23450=>"111000000",
  23451=>"111000000",
  23452=>"111111111",
  23453=>"000011000",
  23454=>"111111000",
  23455=>"110110111",
  23456=>"001110111",
  23457=>"000001001",
  23458=>"110000000",
  23459=>"000000111",
  23460=>"111111111",
  23461=>"111111110",
  23462=>"111111110",
  23463=>"000000111",
  23464=>"101000000",
  23465=>"011000001",
  23466=>"111111111",
  23467=>"111111111",
  23468=>"111111111",
  23469=>"001101001",
  23470=>"111111011",
  23471=>"110000000",
  23472=>"111111111",
  23473=>"000000000",
  23474=>"111001000",
  23475=>"000000000",
  23476=>"111010000",
  23477=>"000010110",
  23478=>"000111111",
  23479=>"000000000",
  23480=>"111010100",
  23481=>"000000110",
  23482=>"101101000",
  23483=>"000001000",
  23484=>"000110110",
  23485=>"100100110",
  23486=>"101000010",
  23487=>"111011011",
  23488=>"000000000",
  23489=>"111010000",
  23490=>"010000000",
  23491=>"111111111",
  23492=>"011110111",
  23493=>"011000000",
  23494=>"100000000",
  23495=>"011111111",
  23496=>"000101111",
  23497=>"000000000",
  23498=>"100000000",
  23499=>"111111111",
  23500=>"010000110",
  23501=>"001000000",
  23502=>"111111111",
  23503=>"111111111",
  23504=>"101001011",
  23505=>"111111100",
  23506=>"111010000",
  23507=>"111111111",
  23508=>"111101000",
  23509=>"000111111",
  23510=>"000111111",
  23511=>"000000000",
  23512=>"101111001",
  23513=>"101111101",
  23514=>"001101101",
  23515=>"111101111",
  23516=>"111100000",
  23517=>"000000000",
  23518=>"111110111",
  23519=>"110000000",
  23520=>"110010000",
  23521=>"000000000",
  23522=>"000011111",
  23523=>"101111111",
  23524=>"100001011",
  23525=>"111111000",
  23526=>"000000111",
  23527=>"010111111",
  23528=>"001000000",
  23529=>"001000000",
  23530=>"000000000",
  23531=>"000000000",
  23532=>"111111000",
  23533=>"110001001",
  23534=>"111110010",
  23535=>"111110000",
  23536=>"111001111",
  23537=>"000000000",
  23538=>"100110111",
  23539=>"101000000",
  23540=>"001000000",
  23541=>"000111111",
  23542=>"000000111",
  23543=>"000100100",
  23544=>"111111111",
  23545=>"000000001",
  23546=>"111111111",
  23547=>"000000111",
  23548=>"000000100",
  23549=>"110000000",
  23550=>"011000000",
  23551=>"111000000",
  23552=>"110010000",
  23553=>"101111000",
  23554=>"111000000",
  23555=>"010011111",
  23556=>"111101111",
  23557=>"111110000",
  23558=>"110111000",
  23559=>"111111111",
  23560=>"110110111",
  23561=>"111001000",
  23562=>"100110111",
  23563=>"111111111",
  23564=>"110111110",
  23565=>"000000000",
  23566=>"000100100",
  23567=>"101111111",
  23568=>"101011111",
  23569=>"001111100",
  23570=>"001101111",
  23571=>"000000000",
  23572=>"111111000",
  23573=>"001001111",
  23574=>"100000111",
  23575=>"110110111",
  23576=>"000000010",
  23577=>"001101111",
  23578=>"110000000",
  23579=>"110100000",
  23580=>"111100000",
  23581=>"001111111",
  23582=>"111001000",
  23583=>"110000000",
  23584=>"000111011",
  23585=>"100000000",
  23586=>"111111111",
  23587=>"000000000",
  23588=>"000000001",
  23589=>"111000000",
  23590=>"010000110",
  23591=>"110000000",
  23592=>"000101111",
  23593=>"111111111",
  23594=>"010001111",
  23595=>"111111111",
  23596=>"000000111",
  23597=>"001111100",
  23598=>"000000110",
  23599=>"000111111",
  23600=>"000100000",
  23601=>"011011011",
  23602=>"111111111",
  23603=>"000000000",
  23604=>"001001100",
  23605=>"000001111",
  23606=>"100000101",
  23607=>"100000000",
  23608=>"000010000",
  23609=>"110100111",
  23610=>"111111001",
  23611=>"111111111",
  23612=>"111110111",
  23613=>"111111111",
  23614=>"010111111",
  23615=>"110111111",
  23616=>"111111111",
  23617=>"001100000",
  23618=>"110110000",
  23619=>"111000000",
  23620=>"010000000",
  23621=>"001111111",
  23622=>"111011000",
  23623=>"000000000",
  23624=>"011010010",
  23625=>"111111001",
  23626=>"111111111",
  23627=>"011000000",
  23628=>"000101111",
  23629=>"111111101",
  23630=>"000010000",
  23631=>"000000000",
  23632=>"110000000",
  23633=>"111110000",
  23634=>"000000000",
  23635=>"001110000",
  23636=>"101001001",
  23637=>"000000000",
  23638=>"100000010",
  23639=>"000000000",
  23640=>"001101111",
  23641=>"111100000",
  23642=>"011000000",
  23643=>"100101000",
  23644=>"110000110",
  23645=>"111101001",
  23646=>"000000010",
  23647=>"100001111",
  23648=>"111000110",
  23649=>"000000000",
  23650=>"000110111",
  23651=>"000000100",
  23652=>"111111000",
  23653=>"111111111",
  23654=>"001000000",
  23655=>"111000000",
  23656=>"101111111",
  23657=>"000000000",
  23658=>"111011111",
  23659=>"000111111",
  23660=>"000000110",
  23661=>"000000000",
  23662=>"111001111",
  23663=>"000111011",
  23664=>"111111000",
  23665=>"000100111",
  23666=>"101111111",
  23667=>"000000111",
  23668=>"100100100",
  23669=>"110111111",
  23670=>"001111111",
  23671=>"111001111",
  23672=>"111000000",
  23673=>"111001000",
  23674=>"000000001",
  23675=>"111001011",
  23676=>"111001000",
  23677=>"000000000",
  23678=>"000000000",
  23679=>"101011100",
  23680=>"000000001",
  23681=>"111111101",
  23682=>"000010111",
  23683=>"111110000",
  23684=>"110000001",
  23685=>"111111000",
  23686=>"100100010",
  23687=>"111111001",
  23688=>"001011011",
  23689=>"100111111",
  23690=>"111111111",
  23691=>"111100000",
  23692=>"001001111",
  23693=>"101000000",
  23694=>"000000000",
  23695=>"100000000",
  23696=>"000000000",
  23697=>"001000000",
  23698=>"000000111",
  23699=>"111000000",
  23700=>"111111111",
  23701=>"111000001",
  23702=>"111111010",
  23703=>"011001000",
  23704=>"001000000",
  23705=>"001010000",
  23706=>"110111010",
  23707=>"000000000",
  23708=>"111100000",
  23709=>"110110111",
  23710=>"110110001",
  23711=>"000011011",
  23712=>"111011011",
  23713=>"000000000",
  23714=>"111111111",
  23715=>"000000000",
  23716=>"110111001",
  23717=>"111000100",
  23718=>"111000000",
  23719=>"100100100",
  23720=>"111111111",
  23721=>"001000000",
  23722=>"010000000",
  23723=>"011111111",
  23724=>"000000011",
  23725=>"000001000",
  23726=>"111111110",
  23727=>"001101111",
  23728=>"111111111",
  23729=>"111111111",
  23730=>"111111000",
  23731=>"110100000",
  23732=>"000011011",
  23733=>"000111111",
  23734=>"000000000",
  23735=>"000000000",
  23736=>"101101000",
  23737=>"000000000",
  23738=>"111000000",
  23739=>"001001001",
  23740=>"000000000",
  23741=>"111100111",
  23742=>"111111111",
  23743=>"000100101",
  23744=>"000001001",
  23745=>"111111111",
  23746=>"000000000",
  23747=>"111111111",
  23748=>"111111111",
  23749=>"100100000",
  23750=>"111011001",
  23751=>"000001001",
  23752=>"111000000",
  23753=>"000011000",
  23754=>"111111111",
  23755=>"000010011",
  23756=>"111011111",
  23757=>"100101111",
  23758=>"111111011",
  23759=>"111000000",
  23760=>"110010011",
  23761=>"000000000",
  23762=>"111000000",
  23763=>"000000000",
  23764=>"111111101",
  23765=>"111111000",
  23766=>"010010010",
  23767=>"000000000",
  23768=>"011111111",
  23769=>"101001101",
  23770=>"111111111",
  23771=>"100111000",
  23772=>"011000000",
  23773=>"101000000",
  23774=>"011111111",
  23775=>"000111010",
  23776=>"000110111",
  23777=>"000100000",
  23778=>"000000000",
  23779=>"111110100",
  23780=>"000001001",
  23781=>"011011000",
  23782=>"100000000",
  23783=>"111111110",
  23784=>"111111110",
  23785=>"111110110",
  23786=>"111000000",
  23787=>"011111111",
  23788=>"111101101",
  23789=>"000110000",
  23790=>"000000000",
  23791=>"111100010",
  23792=>"000000011",
  23793=>"111111111",
  23794=>"111110010",
  23795=>"001111111",
  23796=>"000000111",
  23797=>"111111011",
  23798=>"100100101",
  23799=>"111111000",
  23800=>"000000000",
  23801=>"101101100",
  23802=>"111001000",
  23803=>"111101111",
  23804=>"111010000",
  23805=>"110000000",
  23806=>"000001000",
  23807=>"110111110",
  23808=>"101101001",
  23809=>"101100101",
  23810=>"111011111",
  23811=>"000000000",
  23812=>"111111111",
  23813=>"101111111",
  23814=>"001111011",
  23815=>"000000000",
  23816=>"111111111",
  23817=>"000000000",
  23818=>"000000000",
  23819=>"111111110",
  23820=>"000000000",
  23821=>"101000011",
  23822=>"100000111",
  23823=>"011111111",
  23824=>"111110001",
  23825=>"011001001",
  23826=>"001000000",
  23827=>"111111111",
  23828=>"000000000",
  23829=>"100100111",
  23830=>"101111111",
  23831=>"111111000",
  23832=>"101111111",
  23833=>"111000000",
  23834=>"011000000",
  23835=>"111111111",
  23836=>"110100101",
  23837=>"110000000",
  23838=>"111111111",
  23839=>"111111111",
  23840=>"111111111",
  23841=>"111111010",
  23842=>"011111111",
  23843=>"111111111",
  23844=>"111010010",
  23845=>"110111111",
  23846=>"001111011",
  23847=>"011111110",
  23848=>"000000000",
  23849=>"100000000",
  23850=>"000010000",
  23851=>"000000110",
  23852=>"111111111",
  23853=>"110110110",
  23854=>"000000000",
  23855=>"111101101",
  23856=>"001000000",
  23857=>"100000000",
  23858=>"000010011",
  23859=>"111111111",
  23860=>"000000000",
  23861=>"011001000",
  23862=>"111111000",
  23863=>"100000001",
  23864=>"111111000",
  23865=>"111000111",
  23866=>"110000111",
  23867=>"000000000",
  23868=>"111111111",
  23869=>"011011000",
  23870=>"110110000",
  23871=>"000001000",
  23872=>"000111110",
  23873=>"000000111",
  23874=>"000000000",
  23875=>"111111010",
  23876=>"000000001",
  23877=>"111101111",
  23878=>"010000000",
  23879=>"111111000",
  23880=>"111101100",
  23881=>"111100000",
  23882=>"000000111",
  23883=>"000100100",
  23884=>"111111101",
  23885=>"100000000",
  23886=>"001000000",
  23887=>"010010011",
  23888=>"011011011",
  23889=>"011000011",
  23890=>"111111111",
  23891=>"000000000",
  23892=>"111111000",
  23893=>"111010000",
  23894=>"001011011",
  23895=>"111001011",
  23896=>"111111111",
  23897=>"000010111",
  23898=>"111111111",
  23899=>"111000000",
  23900=>"111110000",
  23901=>"111111011",
  23902=>"011111111",
  23903=>"111111111",
  23904=>"111000000",
  23905=>"111101101",
  23906=>"111100100",
  23907=>"111001000",
  23908=>"100111111",
  23909=>"101101111",
  23910=>"001000100",
  23911=>"001001000",
  23912=>"111011111",
  23913=>"011111111",
  23914=>"111101100",
  23915=>"111101111",
  23916=>"111111111",
  23917=>"001001100",
  23918=>"000000000",
  23919=>"100100000",
  23920=>"111000001",
  23921=>"111101111",
  23922=>"011001000",
  23923=>"100100100",
  23924=>"111110111",
  23925=>"100100000",
  23926=>"011011111",
  23927=>"111111111",
  23928=>"000000001",
  23929=>"101001000",
  23930=>"001001101",
  23931=>"111111000",
  23932=>"001001011",
  23933=>"111111101",
  23934=>"111111011",
  23935=>"000100111",
  23936=>"100000000",
  23937=>"001000001",
  23938=>"110110111",
  23939=>"000000000",
  23940=>"111111111",
  23941=>"000010000",
  23942=>"000011000",
  23943=>"111110011",
  23944=>"011011110",
  23945=>"011001110",
  23946=>"101000000",
  23947=>"000011000",
  23948=>"111111001",
  23949=>"100100101",
  23950=>"111101000",
  23951=>"110111100",
  23952=>"111111100",
  23953=>"000000111",
  23954=>"001101111",
  23955=>"111111110",
  23956=>"000000111",
  23957=>"101101101",
  23958=>"000000000",
  23959=>"100000000",
  23960=>"000000000",
  23961=>"111001000",
  23962=>"001000000",
  23963=>"111111111",
  23964=>"111111110",
  23965=>"000000000",
  23966=>"111111111",
  23967=>"011111111",
  23968=>"011000000",
  23969=>"111011101",
  23970=>"000000000",
  23971=>"011000000",
  23972=>"000000000",
  23973=>"011101111",
  23974=>"000000000",
  23975=>"011011011",
  23976=>"000000000",
  23977=>"111111111",
  23978=>"111100111",
  23979=>"101101001",
  23980=>"111111111",
  23981=>"111000000",
  23982=>"100000001",
  23983=>"111111111",
  23984=>"111011111",
  23985=>"011111111",
  23986=>"000000000",
  23987=>"111111111",
  23988=>"110000000",
  23989=>"011000000",
  23990=>"000110010",
  23991=>"111111010",
  23992=>"000000000",
  23993=>"111011111",
  23994=>"111000000",
  23995=>"000000000",
  23996=>"000000000",
  23997=>"100000000",
  23998=>"000000000",
  23999=>"100100001",
  24000=>"000111011",
  24001=>"111111111",
  24002=>"000000000",
  24003=>"111111110",
  24004=>"000100000",
  24005=>"111111100",
  24006=>"000000000",
  24007=>"000100000",
  24008=>"011000000",
  24009=>"110100101",
  24010=>"111000000",
  24011=>"000000111",
  24012=>"000000000",
  24013=>"111111110",
  24014=>"100000000",
  24015=>"110000000",
  24016=>"000111000",
  24017=>"011011011",
  24018=>"000000000",
  24019=>"000000111",
  24020=>"100111111",
  24021=>"111111000",
  24022=>"000000001",
  24023=>"010011011",
  24024=>"111111111",
  24025=>"110011011",
  24026=>"100100110",
  24027=>"110000000",
  24028=>"011111111",
  24029=>"001001011",
  24030=>"110111010",
  24031=>"110100111",
  24032=>"100110110",
  24033=>"111111111",
  24034=>"000000000",
  24035=>"111011010",
  24036=>"000000000",
  24037=>"111111111",
  24038=>"001001101",
  24039=>"011111111",
  24040=>"010111111",
  24041=>"111100000",
  24042=>"111111111",
  24043=>"000111111",
  24044=>"001000100",
  24045=>"000100000",
  24046=>"000001111",
  24047=>"000000111",
  24048=>"111111111",
  24049=>"110111111",
  24050=>"100000000",
  24051=>"110111111",
  24052=>"101000001",
  24053=>"111001000",
  24054=>"111111111",
  24055=>"001000000",
  24056=>"110000000",
  24057=>"011011010",
  24058=>"110111111",
  24059=>"001001001",
  24060=>"000000110",
  24061=>"101000001",
  24062=>"100111111",
  24063=>"101111111",
  24064=>"000001111",
  24065=>"001000000",
  24066=>"000000000",
  24067=>"000100000",
  24068=>"100000111",
  24069=>"000000000",
  24070=>"000000000",
  24071=>"011111110",
  24072=>"111111111",
  24073=>"101111001",
  24074=>"011001111",
  24075=>"110110001",
  24076=>"000000100",
  24077=>"001000000",
  24078=>"111111110",
  24079=>"001000101",
  24080=>"111000000",
  24081=>"001001111",
  24082=>"000001011",
  24083=>"000000000",
  24084=>"000000111",
  24085=>"000000000",
  24086=>"100110000",
  24087=>"000000101",
  24088=>"111111101",
  24089=>"001101001",
  24090=>"110000100",
  24091=>"000000001",
  24092=>"111111111",
  24093=>"100000110",
  24094=>"000000100",
  24095=>"100100111",
  24096=>"011101100",
  24097=>"000000000",
  24098=>"100000110",
  24099=>"111111000",
  24100=>"111100111",
  24101=>"000001000",
  24102=>"000000000",
  24103=>"000000000",
  24104=>"111000000",
  24105=>"001000000",
  24106=>"111110111",
  24107=>"110100000",
  24108=>"000000111",
  24109=>"000000011",
  24110=>"111011000",
  24111=>"000000000",
  24112=>"111111111",
  24113=>"111111001",
  24114=>"110111111",
  24115=>"111001000",
  24116=>"000000111",
  24117=>"111111000",
  24118=>"111110111",
  24119=>"000000110",
  24120=>"001011011",
  24121=>"000001111",
  24122=>"100110111",
  24123=>"011011100",
  24124=>"111001111",
  24125=>"101111111",
  24126=>"000000000",
  24127=>"111111111",
  24128=>"111111111",
  24129=>"000111111",
  24130=>"111111111",
  24131=>"000000111",
  24132=>"100000011",
  24133=>"001001001",
  24134=>"100111100",
  24135=>"000000011",
  24136=>"000000001",
  24137=>"111101100",
  24138=>"100111111",
  24139=>"000011111",
  24140=>"111111001",
  24141=>"111111011",
  24142=>"111100111",
  24143=>"111111111",
  24144=>"110110000",
  24145=>"111111000",
  24146=>"000111111",
  24147=>"001100110",
  24148=>"111111111",
  24149=>"001100000",
  24150=>"000100111",
  24151=>"000000000",
  24152=>"000000000",
  24153=>"011000111",
  24154=>"100000100",
  24155=>"110110111",
  24156=>"110111000",
  24157=>"111000000",
  24158=>"000000111",
  24159=>"111111011",
  24160=>"011000000",
  24161=>"011011100",
  24162=>"011000000",
  24163=>"001000000",
  24164=>"111111111",
  24165=>"000000000",
  24166=>"111111101",
  24167=>"000000001",
  24168=>"111111000",
  24169=>"000000000",
  24170=>"000000000",
  24171=>"000000000",
  24172=>"100111111",
  24173=>"101000000",
  24174=>"111001111",
  24175=>"111001111",
  24176=>"000001111",
  24177=>"111111000",
  24178=>"111111101",
  24179=>"111110110",
  24180=>"111111111",
  24181=>"000000111",
  24182=>"110100000",
  24183=>"000111111",
  24184=>"101001000",
  24185=>"111101001",
  24186=>"000000000",
  24187=>"000000001",
  24188=>"110000000",
  24189=>"111111111",
  24190=>"111010000",
  24191=>"000000000",
  24192=>"100000010",
  24193=>"111111110",
  24194=>"111111111",
  24195=>"001111111",
  24196=>"000000000",
  24197=>"111011000",
  24198=>"110111000",
  24199=>"000000110",
  24200=>"100000000",
  24201=>"011000111",
  24202=>"011111111",
  24203=>"111111111",
  24204=>"001000000",
  24205=>"101111001",
  24206=>"111111000",
  24207=>"000000011",
  24208=>"111100000",
  24209=>"011111100",
  24210=>"111111111",
  24211=>"111110000",
  24212=>"000110110",
  24213=>"111111101",
  24214=>"010011000",
  24215=>"000000000",
  24216=>"000000000",
  24217=>"111110111",
  24218=>"001000000",
  24219=>"000000001",
  24220=>"000000000",
  24221=>"111100000",
  24222=>"000100111",
  24223=>"000000111",
  24224=>"100111110",
  24225=>"111111110",
  24226=>"111011001",
  24227=>"010000000",
  24228=>"000110100",
  24229=>"100000000",
  24230=>"000000000",
  24231=>"111111000",
  24232=>"100000111",
  24233=>"001001011",
  24234=>"111111111",
  24235=>"111111111",
  24236=>"000101011",
  24237=>"111111111",
  24238=>"001001011",
  24239=>"000111111",
  24240=>"001001000",
  24241=>"111100110",
  24242=>"000000011",
  24243=>"010000000",
  24244=>"000000000",
  24245=>"111100111",
  24246=>"111101001",
  24247=>"111100000",
  24248=>"001000000",
  24249=>"010011111",
  24250=>"000000000",
  24251=>"001000000",
  24252=>"000000011",
  24253=>"111111100",
  24254=>"110111111",
  24255=>"000001001",
  24256=>"001001000",
  24257=>"010000000",
  24258=>"000000000",
  24259=>"000000000",
  24260=>"111111100",
  24261=>"100111111",
  24262=>"000000010",
  24263=>"000000000",
  24264=>"111001010",
  24265=>"000000111",
  24266=>"111001101",
  24267=>"001000000",
  24268=>"000010110",
  24269=>"010000000",
  24270=>"000000111",
  24271=>"000101111",
  24272=>"000000000",
  24273=>"000000011",
  24274=>"111111011",
  24275=>"000000000",
  24276=>"100100111",
  24277=>"000111110",
  24278=>"111100000",
  24279=>"000010000",
  24280=>"110111111",
  24281=>"100000000",
  24282=>"000000111",
  24283=>"111000000",
  24284=>"000000100",
  24285=>"001011000",
  24286=>"000100000",
  24287=>"000101001",
  24288=>"011000000",
  24289=>"010111001",
  24290=>"000111000",
  24291=>"111110111",
  24292=>"111111001",
  24293=>"111011110",
  24294=>"110111111",
  24295=>"010111010",
  24296=>"111001111",
  24297=>"100100011",
  24298=>"110000000",
  24299=>"000000111",
  24300=>"111010111",
  24301=>"000000000",
  24302=>"111111101",
  24303=>"111111000",
  24304=>"110000110",
  24305=>"000000111",
  24306=>"111111111",
  24307=>"000100000",
  24308=>"110110000",
  24309=>"000000000",
  24310=>"100000101",
  24311=>"010000000",
  24312=>"000000111",
  24313=>"111111001",
  24314=>"000100100",
  24315=>"110010000",
  24316=>"111110000",
  24317=>"101001001",
  24318=>"000100010",
  24319=>"000000000",
  24320=>"000000001",
  24321=>"000000101",
  24322=>"100110111",
  24323=>"000000000",
  24324=>"111111111",
  24325=>"111111111",
  24326=>"000000000",
  24327=>"000001111",
  24328=>"000000000",
  24329=>"000111000",
  24330=>"000000000",
  24331=>"111111111",
  24332=>"110100110",
  24333=>"111111111",
  24334=>"111111111",
  24335=>"111111011",
  24336=>"111100000",
  24337=>"000101111",
  24338=>"111100000",
  24339=>"110110011",
  24340=>"000000000",
  24341=>"100100111",
  24342=>"000000100",
  24343=>"000000000",
  24344=>"111001101",
  24345=>"110100000",
  24346=>"000100000",
  24347=>"000110111",
  24348=>"001001111",
  24349=>"000000111",
  24350=>"111000100",
  24351=>"011101101",
  24352=>"110100000",
  24353=>"000000000",
  24354=>"000011011",
  24355=>"000000100",
  24356=>"111100000",
  24357=>"000111000",
  24358=>"000000100",
  24359=>"110111110",
  24360=>"111111011",
  24361=>"000100111",
  24362=>"111100100",
  24363=>"100000000",
  24364=>"111111001",
  24365=>"000001001",
  24366=>"100000000",
  24367=>"000000000",
  24368=>"011011001",
  24369=>"000000000",
  24370=>"110000111",
  24371=>"111011000",
  24372=>"110011010",
  24373=>"000000000",
  24374=>"111111111",
  24375=>"111111001",
  24376=>"000111111",
  24377=>"111101111",
  24378=>"000001111",
  24379=>"111111011",
  24380=>"000000111",
  24381=>"000001110",
  24382=>"110000000",
  24383=>"000000000",
  24384=>"000011011",
  24385=>"000000000",
  24386=>"001101111",
  24387=>"111010000",
  24388=>"001101000",
  24389=>"111000000",
  24390=>"110000000",
  24391=>"110111111",
  24392=>"000000000",
  24393=>"000000000",
  24394=>"011011010",
  24395=>"111101100",
  24396=>"111111111",
  24397=>"000100000",
  24398=>"111111000",
  24399=>"111111000",
  24400=>"000000100",
  24401=>"100000000",
  24402=>"111111000",
  24403=>"110110000",
  24404=>"000011000",
  24405=>"101011011",
  24406=>"011101001",
  24407=>"111111001",
  24408=>"111110110",
  24409=>"001001000",
  24410=>"011000000",
  24411=>"000000011",
  24412=>"000000000",
  24413=>"111111100",
  24414=>"111111000",
  24415=>"000110100",
  24416=>"111111111",
  24417=>"111111111",
  24418=>"001001001",
  24419=>"000000011",
  24420=>"000000001",
  24421=>"000001111",
  24422=>"100101101",
  24423=>"111111001",
  24424=>"110000110",
  24425=>"111111111",
  24426=>"000010000",
  24427=>"111101000",
  24428=>"011011101",
  24429=>"000000000",
  24430=>"000011111",
  24431=>"000000001",
  24432=>"000111111",
  24433=>"000010010",
  24434=>"001101100",
  24435=>"001000001",
  24436=>"100111111",
  24437=>"101111111",
  24438=>"111000011",
  24439=>"001111111",
  24440=>"111000000",
  24441=>"111001001",
  24442=>"111111000",
  24443=>"110111000",
  24444=>"000000111",
  24445=>"000111000",
  24446=>"111111001",
  24447=>"000000111",
  24448=>"000000000",
  24449=>"000010111",
  24450=>"000000000",
  24451=>"000000111",
  24452=>"111000111",
  24453=>"000010010",
  24454=>"000000000",
  24455=>"000000000",
  24456=>"111111000",
  24457=>"001111000",
  24458=>"111101001",
  24459=>"011011010",
  24460=>"111111110",
  24461=>"000100100",
  24462=>"111000000",
  24463=>"110110000",
  24464=>"100000000",
  24465=>"000000000",
  24466=>"111111111",
  24467=>"000000110",
  24468=>"000000111",
  24469=>"111111111",
  24470=>"011100111",
  24471=>"000000001",
  24472=>"000000000",
  24473=>"000000001",
  24474=>"000000111",
  24475=>"001011111",
  24476=>"011001101",
  24477=>"100100111",
  24478=>"111000000",
  24479=>"000000111",
  24480=>"000000001",
  24481=>"111011000",
  24482=>"000111111",
  24483=>"111100111",
  24484=>"100000110",
  24485=>"010000000",
  24486=>"111110000",
  24487=>"000110000",
  24488=>"000010110",
  24489=>"001111111",
  24490=>"100100000",
  24491=>"011001100",
  24492=>"111000000",
  24493=>"111111100",
  24494=>"011111111",
  24495=>"000000111",
  24496=>"111000111",
  24497=>"011000000",
  24498=>"011111001",
  24499=>"111111111",
  24500=>"111111111",
  24501=>"111111110",
  24502=>"000000111",
  24503=>"001111000",
  24504=>"100111111",
  24505=>"001101111",
  24506=>"111101001",
  24507=>"111111000",
  24508=>"000010000",
  24509=>"000000000",
  24510=>"001000000",
  24511=>"000001111",
  24512=>"110100111",
  24513=>"111000000",
  24514=>"111111111",
  24515=>"000111111",
  24516=>"111111111",
  24517=>"000001111",
  24518=>"000000000",
  24519=>"110000000",
  24520=>"011001000",
  24521=>"111111100",
  24522=>"000001111",
  24523=>"000000000",
  24524=>"111111111",
  24525=>"000111011",
  24526=>"000010000",
  24527=>"110110110",
  24528=>"111011000",
  24529=>"001000000",
  24530=>"110111011",
  24531=>"010010111",
  24532=>"100000000",
  24533=>"111011000",
  24534=>"111111101",
  24535=>"001000110",
  24536=>"111111111",
  24537=>"111111001",
  24538=>"000000000",
  24539=>"111000000",
  24540=>"011011011",
  24541=>"110000000",
  24542=>"100111000",
  24543=>"000000111",
  24544=>"010000111",
  24545=>"011010011",
  24546=>"110111100",
  24547=>"011111111",
  24548=>"000000110",
  24549=>"111000111",
  24550=>"111111000",
  24551=>"110110100",
  24552=>"100000100",
  24553=>"111100000",
  24554=>"001110111",
  24555=>"000000000",
  24556=>"000110000",
  24557=>"111111100",
  24558=>"000000000",
  24559=>"001000000",
  24560=>"011111111",
  24561=>"001000101",
  24562=>"111001000",
  24563=>"110010000",
  24564=>"110000000",
  24565=>"110111101",
  24566=>"000000111",
  24567=>"001000110",
  24568=>"111011111",
  24569=>"000111111",
  24570=>"000000111",
  24571=>"000000100",
  24572=>"000001000",
  24573=>"111101000",
  24574=>"000000000",
  24575=>"111000000",
  24576=>"100111111",
  24577=>"000000000",
  24578=>"000000000",
  24579=>"111111111",
  24580=>"000011111",
  24581=>"001000101",
  24582=>"111000000",
  24583=>"100000000",
  24584=>"000000000",
  24585=>"000111111",
  24586=>"111111111",
  24587=>"000000110",
  24588=>"000011000",
  24589=>"111111011",
  24590=>"110001000",
  24591=>"000001011",
  24592=>"100000000",
  24593=>"111111100",
  24594=>"001011111",
  24595=>"100100100",
  24596=>"111111011",
  24597=>"000011111",
  24598=>"111100100",
  24599=>"000000100",
  24600=>"000111111",
  24601=>"111011011",
  24602=>"000000001",
  24603=>"111100110",
  24604=>"000000000",
  24605=>"001001000",
  24606=>"000000000",
  24607=>"000000111",
  24608=>"110111001",
  24609=>"000000101",
  24610=>"000000000",
  24611=>"000000000",
  24612=>"010000110",
  24613=>"000000000",
  24614=>"000000100",
  24615=>"111111011",
  24616=>"000100110",
  24617=>"111111100",
  24618=>"000001011",
  24619=>"000000000",
  24620=>"101101111",
  24621=>"000111110",
  24622=>"111111111",
  24623=>"100000000",
  24624=>"000001011",
  24625=>"000000001",
  24626=>"000000001",
  24627=>"000010000",
  24628=>"010101111",
  24629=>"101001111",
  24630=>"000000000",
  24631=>"010000000",
  24632=>"111111011",
  24633=>"000000110",
  24634=>"111111111",
  24635=>"111000000",
  24636=>"011001011",
  24637=>"000000000",
  24638=>"011000111",
  24639=>"111000000",
  24640=>"001001101",
  24641=>"000000000",
  24642=>"000000000",
  24643=>"101101111",
  24644=>"110111111",
  24645=>"001001000",
  24646=>"000000000",
  24647=>"111111111",
  24648=>"110110111",
  24649=>"100111111",
  24650=>"111111111",
  24651=>"111111111",
  24652=>"110101110",
  24653=>"110111111",
  24654=>"001011011",
  24655=>"110100111",
  24656=>"000110111",
  24657=>"001000000",
  24658=>"000000000",
  24659=>"000100000",
  24660=>"111111111",
  24661=>"000000000",
  24662=>"000000000",
  24663=>"111000000",
  24664=>"010110000",
  24665=>"000000111",
  24666=>"111101111",
  24667=>"000000100",
  24668=>"010000000",
  24669=>"011111111",
  24670=>"000001001",
  24671=>"111111000",
  24672=>"101000000",
  24673=>"000001000",
  24674=>"000000000",
  24675=>"000000000",
  24676=>"001001000",
  24677=>"111100000",
  24678=>"001111111",
  24679=>"011010111",
  24680=>"000000110",
  24681=>"111111111",
  24682=>"000000110",
  24683=>"101111011",
  24684=>"111110000",
  24685=>"111001000",
  24686=>"111000000",
  24687=>"000000000",
  24688=>"111111001",
  24689=>"101000000",
  24690=>"000000111",
  24691=>"000001011",
  24692=>"111111011",
  24693=>"000000001",
  24694=>"000000000",
  24695=>"111101111",
  24696=>"000011111",
  24697=>"000111111",
  24698=>"111111111",
  24699=>"111111111",
  24700=>"000000000",
  24701=>"001001011",
  24702=>"000000111",
  24703=>"001000000",
  24704=>"001001001",
  24705=>"111010000",
  24706=>"000000000",
  24707=>"000000000",
  24708=>"111111111",
  24709=>"111111111",
  24710=>"001001101",
  24711=>"001000001",
  24712=>"001111111",
  24713=>"000000000",
  24714=>"000000000",
  24715=>"110000000",
  24716=>"000000010",
  24717=>"000000000",
  24718=>"111111111",
  24719=>"111111011",
  24720=>"000000011",
  24721=>"111111111",
  24722=>"000001001",
  24723=>"000000000",
  24724=>"000010101",
  24725=>"011110111",
  24726=>"111011011",
  24727=>"111101001",
  24728=>"001000000",
  24729=>"111111110",
  24730=>"111000000",
  24731=>"000000000",
  24732=>"101110100",
  24733=>"000011011",
  24734=>"111111111",
  24735=>"010111111",
  24736=>"111010100",
  24737=>"110111111",
  24738=>"111110000",
  24739=>"111111111",
  24740=>"111001001",
  24741=>"100111111",
  24742=>"000000111",
  24743=>"000000111",
  24744=>"000000000",
  24745=>"000000000",
  24746=>"111001000",
  24747=>"000111111",
  24748=>"000000110",
  24749=>"111111111",
  24750=>"110100111",
  24751=>"101101000",
  24752=>"111100000",
  24753=>"000110110",
  24754=>"110111111",
  24755=>"000000000",
  24756=>"110110001",
  24757=>"100000101",
  24758=>"011111000",
  24759=>"000000000",
  24760=>"000011111",
  24761=>"111111101",
  24762=>"111000000",
  24763=>"111001001",
  24764=>"011001001",
  24765=>"000000000",
  24766=>"000000000",
  24767=>"111111011",
  24768=>"001000000",
  24769=>"010111111",
  24770=>"000011111",
  24771=>"001001000",
  24772=>"000000000",
  24773=>"000001111",
  24774=>"000000001",
  24775=>"111001100",
  24776=>"111001000",
  24777=>"000101101",
  24778=>"000000001",
  24779=>"111001111",
  24780=>"000101100",
  24781=>"000010000",
  24782=>"000000010",
  24783=>"000001001",
  24784=>"111011001",
  24785=>"000000000",
  24786=>"000000000",
  24787=>"111111000",
  24788=>"111111111",
  24789=>"000000001",
  24790=>"000000000",
  24791=>"000000111",
  24792=>"111111100",
  24793=>"100000000",
  24794=>"000111111",
  24795=>"111111111",
  24796=>"110000100",
  24797=>"101111111",
  24798=>"000000000",
  24799=>"010011001",
  24800=>"111000000",
  24801=>"111111110",
  24802=>"010000000",
  24803=>"000001001",
  24804=>"011111111",
  24805=>"001001000",
  24806=>"111111111",
  24807=>"011011111",
  24808=>"000000000",
  24809=>"111111000",
  24810=>"010000111",
  24811=>"111111111",
  24812=>"000011111",
  24813=>"001000000",
  24814=>"000000001",
  24815=>"000000000",
  24816=>"111110111",
  24817=>"100111111",
  24818=>"000000000",
  24819=>"101001000",
  24820=>"111101111",
  24821=>"010000000",
  24822=>"000000001",
  24823=>"001001001",
  24824=>"000000000",
  24825=>"000000000",
  24826=>"000111110",
  24827=>"110110010",
  24828=>"000000001",
  24829=>"111001000",
  24830=>"000001001",
  24831=>"000001001",
  24832=>"001000000",
  24833=>"011111100",
  24834=>"111111000",
  24835=>"000000000",
  24836=>"000000000",
  24837=>"110110010",
  24838=>"000000000",
  24839=>"000000010",
  24840=>"111111111",
  24841=>"110110111",
  24842=>"011001001",
  24843=>"111111101",
  24844=>"111101111",
  24845=>"111111111",
  24846=>"000000000",
  24847=>"000100111",
  24848=>"010111111",
  24849=>"000000000",
  24850=>"000000000",
  24851=>"110111111",
  24852=>"000000000",
  24853=>"000000000",
  24854=>"110111111",
  24855=>"001100000",
  24856=>"010100001",
  24857=>"111101111",
  24858=>"000010010",
  24859=>"100000000",
  24860=>"000101100",
  24861=>"101100001",
  24862=>"000000000",
  24863=>"011000000",
  24864=>"101111011",
  24865=>"111111111",
  24866=>"111001011",
  24867=>"000011111",
  24868=>"000000110",
  24869=>"111111111",
  24870=>"111111111",
  24871=>"101001000",
  24872=>"011000000",
  24873=>"111111111",
  24874=>"000011000",
  24875=>"000000000",
  24876=>"111111111",
  24877=>"000110100",
  24878=>"000001001",
  24879=>"111111111",
  24880=>"001111111",
  24881=>"011111111",
  24882=>"000000000",
  24883=>"001000000",
  24884=>"000000100",
  24885=>"111111111",
  24886=>"001000000",
  24887=>"100000000",
  24888=>"111111101",
  24889=>"001001111",
  24890=>"000000000",
  24891=>"000000101",
  24892=>"001001111",
  24893=>"100100110",
  24894=>"000000100",
  24895=>"011111010",
  24896=>"000000000",
  24897=>"001001111",
  24898=>"111111011",
  24899=>"100100110",
  24900=>"111111000",
  24901=>"011011011",
  24902=>"011111110",
  24903=>"111101101",
  24904=>"000000000",
  24905=>"110000000",
  24906=>"111111111",
  24907=>"000111110",
  24908=>"000000000",
  24909=>"000000000",
  24910=>"100101111",
  24911=>"100101111",
  24912=>"000111011",
  24913=>"101100001",
  24914=>"011011111",
  24915=>"111111111",
  24916=>"100000100",
  24917=>"001001001",
  24918=>"111111111",
  24919=>"000000000",
  24920=>"111111111",
  24921=>"010110110",
  24922=>"000000111",
  24923=>"111111111",
  24924=>"000000000",
  24925=>"111111111",
  24926=>"110110110",
  24927=>"000000111",
  24928=>"111111111",
  24929=>"000011111",
  24930=>"000100000",
  24931=>"111101011",
  24932=>"000000100",
  24933=>"011000000",
  24934=>"101101100",
  24935=>"000000101",
  24936=>"010011000",
  24937=>"011011000",
  24938=>"000000111",
  24939=>"111111000",
  24940=>"000000010",
  24941=>"111000001",
  24942=>"000000000",
  24943=>"100010000",
  24944=>"111000000",
  24945=>"000000011",
  24946=>"010010000",
  24947=>"111100111",
  24948=>"111110110",
  24949=>"000000100",
  24950=>"010011000",
  24951=>"100000000",
  24952=>"111000001",
  24953=>"000110111",
  24954=>"000000000",
  24955=>"011111111",
  24956=>"001010000",
  24957=>"110111111",
  24958=>"010000000",
  24959=>"000000001",
  24960=>"000000000",
  24961=>"111111001",
  24962=>"110000001",
  24963=>"000011111",
  24964=>"000000000",
  24965=>"111111000",
  24966=>"000011111",
  24967=>"011011011",
  24968=>"000000000",
  24969=>"111011000",
  24970=>"000100111",
  24971=>"111110110",
  24972=>"111111111",
  24973=>"000000000",
  24974=>"000000000",
  24975=>"000000000",
  24976=>"011000000",
  24977=>"000000000",
  24978=>"111010100",
  24979=>"000000000",
  24980=>"111111111",
  24981=>"000000000",
  24982=>"001100010",
  24983=>"111111111",
  24984=>"111101111",
  24985=>"000011011",
  24986=>"111000000",
  24987=>"111000000",
  24988=>"011011111",
  24989=>"000000000",
  24990=>"011111111",
  24991=>"000000000",
  24992=>"001000001",
  24993=>"000000000",
  24994=>"110111111",
  24995=>"111011111",
  24996=>"000000000",
  24997=>"111111111",
  24998=>"111111111",
  24999=>"000010111",
  25000=>"000000001",
  25001=>"000000100",
  25002=>"111000000",
  25003=>"110110111",
  25004=>"000000000",
  25005=>"110110100",
  25006=>"000110111",
  25007=>"110111111",
  25008=>"111111111",
  25009=>"000000000",
  25010=>"000000000",
  25011=>"000000000",
  25012=>"011001011",
  25013=>"111111100",
  25014=>"000000000",
  25015=>"000000011",
  25016=>"111111011",
  25017=>"111111111",
  25018=>"000000000",
  25019=>"011111111",
  25020=>"111111111",
  25021=>"000000100",
  25022=>"000000000",
  25023=>"110000100",
  25024=>"111111111",
  25025=>"111101111",
  25026=>"111111111",
  25027=>"010111111",
  25028=>"111111000",
  25029=>"000100100",
  25030=>"111100111",
  25031=>"111111111",
  25032=>"011000000",
  25033=>"111100000",
  25034=>"001101000",
  25035=>"111111011",
  25036=>"111111110",
  25037=>"100000111",
  25038=>"000000000",
  25039=>"000000100",
  25040=>"111111011",
  25041=>"000000001",
  25042=>"000000000",
  25043=>"111111111",
  25044=>"001001000",
  25045=>"000000111",
  25046=>"000000001",
  25047=>"100100000",
  25048=>"000100101",
  25049=>"111111111",
  25050=>"110101111",
  25051=>"100101111",
  25052=>"000000000",
  25053=>"111111111",
  25054=>"111111111",
  25055=>"010110100",
  25056=>"000000001",
  25057=>"011000000",
  25058=>"111000000",
  25059=>"000000100",
  25060=>"110000000",
  25061=>"000000111",
  25062=>"000000110",
  25063=>"011110000",
  25064=>"111110100",
  25065=>"000000000",
  25066=>"000000111",
  25067=>"111111111",
  25068=>"000111111",
  25069=>"111101111",
  25070=>"111000111",
  25071=>"111110000",
  25072=>"001001111",
  25073=>"011101111",
  25074=>"111111111",
  25075=>"000000111",
  25076=>"111110111",
  25077=>"011111111",
  25078=>"110110110",
  25079=>"000000000",
  25080=>"001111000",
  25081=>"000001000",
  25082=>"010111111",
  25083=>"000000000",
  25084=>"000000000",
  25085=>"011011111",
  25086=>"000110111",
  25087=>"111111111",
  25088=>"001001001",
  25089=>"111000000",
  25090=>"101111001",
  25091=>"000000111",
  25092=>"101111111",
  25093=>"000000000",
  25094=>"111001000",
  25095=>"000000001",
  25096=>"000000000",
  25097=>"000000111",
  25098=>"000000000",
  25099=>"111011111",
  25100=>"100100100",
  25101=>"011111111",
  25102=>"100110111",
  25103=>"000111111",
  25104=>"100110111",
  25105=>"000000000",
  25106=>"110010011",
  25107=>"000000101",
  25108=>"000001011",
  25109=>"010010011",
  25110=>"000000100",
  25111=>"101101100",
  25112=>"000000000",
  25113=>"110110100",
  25114=>"111111111",
  25115=>"100100001",
  25116=>"111001001",
  25117=>"011111000",
  25118=>"000000001",
  25119=>"111011000",
  25120=>"000000001",
  25121=>"111111000",
  25122=>"110100000",
  25123=>"000000000",
  25124=>"011011000",
  25125=>"110111111",
  25126=>"111001011",
  25127=>"011000000",
  25128=>"000000000",
  25129=>"111111101",
  25130=>"000000100",
  25131=>"111010000",
  25132=>"000000000",
  25133=>"000000000",
  25134=>"100010000",
  25135=>"011001000",
  25136=>"011010111",
  25137=>"000000000",
  25138=>"100100100",
  25139=>"001001001",
  25140=>"100110111",
  25141=>"100110110",
  25142=>"111111010",
  25143=>"110000101",
  25144=>"111111111",
  25145=>"101000000",
  25146=>"111111000",
  25147=>"001011111",
  25148=>"101101111",
  25149=>"000000000",
  25150=>"000110111",
  25151=>"000000000",
  25152=>"111011000",
  25153=>"111111100",
  25154=>"001111111",
  25155=>"111111111",
  25156=>"110111001",
  25157=>"111111111",
  25158=>"001000000",
  25159=>"000000000",
  25160=>"000011011",
  25161=>"001001111",
  25162=>"111111000",
  25163=>"000000001",
  25164=>"000110111",
  25165=>"110110110",
  25166=>"000000000",
  25167=>"101111111",
  25168=>"000000001",
  25169=>"011011000",
  25170=>"000000000",
  25171=>"000000000",
  25172=>"011111111",
  25173=>"000101001",
  25174=>"000000001",
  25175=>"100100100",
  25176=>"111001000",
  25177=>"001001000",
  25178=>"011011111",
  25179=>"000000000",
  25180=>"000000000",
  25181=>"110000010",
  25182=>"001000000",
  25183=>"001001000",
  25184=>"000000000",
  25185=>"001100000",
  25186=>"001000000",
  25187=>"000000111",
  25188=>"111111000",
  25189=>"111010111",
  25190=>"000100101",
  25191=>"011000100",
  25192=>"000000000",
  25193=>"111111111",
  25194=>"111111111",
  25195=>"000000000",
  25196=>"101111111",
  25197=>"111010000",
  25198=>"000000100",
  25199=>"000000000",
  25200=>"010000001",
  25201=>"010000111",
  25202=>"100000000",
  25203=>"000000000",
  25204=>"011000000",
  25205=>"000000000",
  25206=>"000100110",
  25207=>"000011011",
  25208=>"000000111",
  25209=>"000011011",
  25210=>"111101111",
  25211=>"000000000",
  25212=>"110110111",
  25213=>"111111111",
  25214=>"111111111",
  25215=>"110000000",
  25216=>"000000000",
  25217=>"111111111",
  25218=>"111111100",
  25219=>"111111000",
  25220=>"000000111",
  25221=>"111111111",
  25222=>"101001111",
  25223=>"111101101",
  25224=>"010010000",
  25225=>"101100100",
  25226=>"111111111",
  25227=>"000011000",
  25228=>"111111111",
  25229=>"000000000",
  25230=>"011110111",
  25231=>"000000000",
  25232=>"000111111",
  25233=>"100110111",
  25234=>"000010111",
  25235=>"111000000",
  25236=>"011000100",
  25237=>"000111111",
  25238=>"000000000",
  25239=>"000000000",
  25240=>"101000001",
  25241=>"111111000",
  25242=>"000000001",
  25243=>"000111111",
  25244=>"110000000",
  25245=>"000000101",
  25246=>"011001111",
  25247=>"111001001",
  25248=>"111111111",
  25249=>"101111001",
  25250=>"000110001",
  25251=>"000000000",
  25252=>"000001001",
  25253=>"011111111",
  25254=>"101000001",
  25255=>"000001111",
  25256=>"111111000",
  25257=>"111100000",
  25258=>"000000000",
  25259=>"000000100",
  25260=>"111111111",
  25261=>"100000001",
  25262=>"111111111",
  25263=>"000010111",
  25264=>"111011011",
  25265=>"000010010",
  25266=>"111111011",
  25267=>"111000000",
  25268=>"000101111",
  25269=>"100110111",
  25270=>"111111111",
  25271=>"111111110",
  25272=>"110111111",
  25273=>"111011010",
  25274=>"000001001",
  25275=>"100000111",
  25276=>"101101111",
  25277=>"111111000",
  25278=>"000111011",
  25279=>"001111111",
  25280=>"000000000",
  25281=>"001101111",
  25282=>"011111000",
  25283=>"000000000",
  25284=>"000001111",
  25285=>"101000101",
  25286=>"000000101",
  25287=>"110111000",
  25288=>"000000011",
  25289=>"111001000",
  25290=>"000000101",
  25291=>"111111111",
  25292=>"001000000",
  25293=>"010110110",
  25294=>"000000000",
  25295=>"000000000",
  25296=>"111111000",
  25297=>"000000000",
  25298=>"111110110",
  25299=>"111111011",
  25300=>"011000111",
  25301=>"011011000",
  25302=>"000000000",
  25303=>"111111111",
  25304=>"111111110",
  25305=>"110111001",
  25306=>"111101111",
  25307=>"011010011",
  25308=>"000111111",
  25309=>"000000001",
  25310=>"000000000",
  25311=>"111111101",
  25312=>"111000111",
  25313=>"011011111",
  25314=>"000011011",
  25315=>"000000000",
  25316=>"000001110",
  25317=>"101001000",
  25318=>"111111110",
  25319=>"101111011",
  25320=>"101111011",
  25321=>"000001111",
  25322=>"101110111",
  25323=>"000000000",
  25324=>"111111111",
  25325=>"111011000",
  25326=>"111111011",
  25327=>"111011011",
  25328=>"011011111",
  25329=>"111000000",
  25330=>"110111111",
  25331=>"000000000",
  25332=>"111111111",
  25333=>"111011000",
  25334=>"111111111",
  25335=>"111111111",
  25336=>"000000000",
  25337=>"000001111",
  25338=>"001001000",
  25339=>"010000000",
  25340=>"000000000",
  25341=>"000000101",
  25342=>"111001101",
  25343=>"000000111",
  25344=>"000000000",
  25345=>"111010011",
  25346=>"000000000",
  25347=>"000000000",
  25348=>"010111011",
  25349=>"110111010",
  25350=>"010111111",
  25351=>"000000000",
  25352=>"000000000",
  25353=>"000000011",
  25354=>"100000001",
  25355=>"000000000",
  25356=>"111011111",
  25357=>"000110000",
  25358=>"111111000",
  25359=>"111111111",
  25360=>"000001000",
  25361=>"111111111",
  25362=>"001000111",
  25363=>"000110111",
  25364=>"000111111",
  25365=>"000000000",
  25366=>"000000011",
  25367=>"000000000",
  25368=>"111011000",
  25369=>"011000000",
  25370=>"001001000",
  25371=>"100000000",
  25372=>"100100110",
  25373=>"000000000",
  25374=>"000000000",
  25375=>"000101000",
  25376=>"111111101",
  25377=>"000000000",
  25378=>"111111000",
  25379=>"001000000",
  25380=>"111000000",
  25381=>"111111111",
  25382=>"001000000",
  25383=>"111011100",
  25384=>"000000000",
  25385=>"000000100",
  25386=>"111100000",
  25387=>"000000000",
  25388=>"111111110",
  25389=>"000000001",
  25390=>"000000000",
  25391=>"111111000",
  25392=>"111111011",
  25393=>"111111111",
  25394=>"000000011",
  25395=>"000000000",
  25396=>"111111111",
  25397=>"000110111",
  25398=>"000000000",
  25399=>"111111011",
  25400=>"000011111",
  25401=>"001001010",
  25402=>"101111101",
  25403=>"011011000",
  25404=>"000000000",
  25405=>"011000111",
  25406=>"000000000",
  25407=>"111111111",
  25408=>"001011111",
  25409=>"111111100",
  25410=>"000001001",
  25411=>"111000000",
  25412=>"000100110",
  25413=>"110010110",
  25414=>"000000001",
  25415=>"000000111",
  25416=>"000000000",
  25417=>"000000000",
  25418=>"000000001",
  25419=>"101001000",
  25420=>"111000111",
  25421=>"111111111",
  25422=>"111111111",
  25423=>"000111111",
  25424=>"101100111",
  25425=>"000000000",
  25426=>"011001000",
  25427=>"000100111",
  25428=>"111111000",
  25429=>"011011011",
  25430=>"001000101",
  25431=>"101100100",
  25432=>"101001000",
  25433=>"111110110",
  25434=>"000000000",
  25435=>"111111010",
  25436=>"000000000",
  25437=>"111110110",
  25438=>"111111111",
  25439=>"011111111",
  25440=>"111111100",
  25441=>"000000000",
  25442=>"100110110",
  25443=>"111111011",
  25444=>"000000100",
  25445=>"110000000",
  25446=>"111111111",
  25447=>"000000000",
  25448=>"111111000",
  25449=>"111111010",
  25450=>"111111111",
  25451=>"000110110",
  25452=>"111101000",
  25453=>"000000000",
  25454=>"001001000",
  25455=>"000000000",
  25456=>"000000000",
  25457=>"100100110",
  25458=>"100000000",
  25459=>"001011000",
  25460=>"111001001",
  25461=>"000000000",
  25462=>"000000011",
  25463=>"111010000",
  25464=>"000000000",
  25465=>"111111111",
  25466=>"001001001",
  25467=>"110110000",
  25468=>"111100000",
  25469=>"000000000",
  25470=>"111111111",
  25471=>"111000000",
  25472=>"111111100",
  25473=>"000000001",
  25474=>"111111111",
  25475=>"001001001",
  25476=>"011001000",
  25477=>"000010110",
  25478=>"000001000",
  25479=>"001111111",
  25480=>"111111111",
  25481=>"000000110",
  25482=>"000111111",
  25483=>"111100000",
  25484=>"111101000",
  25485=>"110110110",
  25486=>"111111001",
  25487=>"000000000",
  25488=>"000000000",
  25489=>"111111010",
  25490=>"111111111",
  25491=>"000000000",
  25492=>"111111111",
  25493=>"000010110",
  25494=>"100100101",
  25495=>"111111000",
  25496=>"000110100",
  25497=>"000000000",
  25498=>"101000001",
  25499=>"000000000",
  25500=>"111111111",
  25501=>"000111111",
  25502=>"111000000",
  25503=>"111111111",
  25504=>"111100000",
  25505=>"000101110",
  25506=>"111101000",
  25507=>"111111110",
  25508=>"110000000",
  25509=>"000000000",
  25510=>"011000100",
  25511=>"000111011",
  25512=>"000000000",
  25513=>"000000111",
  25514=>"100000111",
  25515=>"010000000",
  25516=>"001000000",
  25517=>"000000001",
  25518=>"110011010",
  25519=>"000000000",
  25520=>"000000001",
  25521=>"000000000",
  25522=>"111101111",
  25523=>"111000000",
  25524=>"000000111",
  25525=>"011000000",
  25526=>"111111111",
  25527=>"111000000",
  25528=>"111111001",
  25529=>"000010000",
  25530=>"100000000",
  25531=>"111000111",
  25532=>"100100001",
  25533=>"111001000",
  25534=>"000011000",
  25535=>"011001001",
  25536=>"101000000",
  25537=>"110000000",
  25538=>"111111000",
  25539=>"111000000",
  25540=>"000000111",
  25541=>"001011001",
  25542=>"000000000",
  25543=>"010110010",
  25544=>"100000111",
  25545=>"110000111",
  25546=>"111000001",
  25547=>"000000000",
  25548=>"110011111",
  25549=>"111111111",
  25550=>"010000000",
  25551=>"001011111",
  25552=>"000100000",
  25553=>"111111111",
  25554=>"000000101",
  25555=>"111101110",
  25556=>"111110100",
  25557=>"110111111",
  25558=>"000000111",
  25559=>"011111011",
  25560=>"000000001",
  25561=>"000100001",
  25562=>"111111010",
  25563=>"101011111",
  25564=>"111111111",
  25565=>"111110000",
  25566=>"011111111",
  25567=>"101001011",
  25568=>"111111111",
  25569=>"111111111",
  25570=>"111111111",
  25571=>"000110111",
  25572=>"011000000",
  25573=>"111111111",
  25574=>"000000011",
  25575=>"111000000",
  25576=>"111111111",
  25577=>"000111111",
  25578=>"111000110",
  25579=>"111111011",
  25580=>"101000001",
  25581=>"111110110",
  25582=>"000000111",
  25583=>"000000101",
  25584=>"010111011",
  25585=>"110111111",
  25586=>"001101111",
  25587=>"100100000",
  25588=>"000000001",
  25589=>"111111011",
  25590=>"011011111",
  25591=>"000000001",
  25592=>"111111111",
  25593=>"000001000",
  25594=>"000000000",
  25595=>"000101101",
  25596=>"111111110",
  25597=>"111111111",
  25598=>"111111100",
  25599=>"000000000",
  25600=>"111111111",
  25601=>"111001000",
  25602=>"111000000",
  25603=>"101110000",
  25604=>"000111111",
  25605=>"001001101",
  25606=>"111111111",
  25607=>"000111111",
  25608=>"011111111",
  25609=>"111000000",
  25610=>"010111000",
  25611=>"000000110",
  25612=>"111001111",
  25613=>"111111011",
  25614=>"110000000",
  25615=>"000000000",
  25616=>"000101101",
  25617=>"111111111",
  25618=>"100001001",
  25619=>"100111111",
  25620=>"011000000",
  25621=>"111111111",
  25622=>"111010000",
  25623=>"000111111",
  25624=>"110111111",
  25625=>"111100100",
  25626=>"111000000",
  25627=>"111111111",
  25628=>"000111111",
  25629=>"111101100",
  25630=>"000001011",
  25631=>"111111111",
  25632=>"000000111",
  25633=>"111111011",
  25634=>"011011000",
  25635=>"111011000",
  25636=>"000000000",
  25637=>"111111111",
  25638=>"000000111",
  25639=>"000100100",
  25640=>"010000000",
  25641=>"000000000",
  25642=>"110110110",
  25643=>"111010101",
  25644=>"100101000",
  25645=>"111011000",
  25646=>"100100100",
  25647=>"110111111",
  25648=>"000000100",
  25649=>"111111000",
  25650=>"010010110",
  25651=>"000010111",
  25652=>"100000011",
  25653=>"111100000",
  25654=>"000000000",
  25655=>"110110111",
  25656=>"111000111",
  25657=>"011111111",
  25658=>"001000111",
  25659=>"100110111",
  25660=>"000000000",
  25661=>"011011001",
  25662=>"010110011",
  25663=>"111000100",
  25664=>"000010111",
  25665=>"101100111",
  25666=>"011000000",
  25667=>"011000010",
  25668=>"000000111",
  25669=>"111000000",
  25670=>"000000000",
  25671=>"111111111",
  25672=>"010000000",
  25673=>"000000111",
  25674=>"000110111",
  25675=>"001100000",
  25676=>"100000000",
  25677=>"111111111",
  25678=>"101000000",
  25679=>"111110000",
  25680=>"111111111",
  25681=>"001001110",
  25682=>"000100000",
  25683=>"110110100",
  25684=>"100000000",
  25685=>"000000000",
  25686=>"001110100",
  25687=>"000000011",
  25688=>"000111010",
  25689=>"000000001",
  25690=>"010000000",
  25691=>"101001111",
  25692=>"111111011",
  25693=>"000111111",
  25694=>"110111110",
  25695=>"000010000",
  25696=>"110000000",
  25697=>"111111100",
  25698=>"000000110",
  25699=>"000001001",
  25700=>"000000110",
  25701=>"110110110",
  25702=>"111000100",
  25703=>"000101111",
  25704=>"001000000",
  25705=>"000000000",
  25706=>"001000000",
  25707=>"000000001",
  25708=>"110111100",
  25709=>"000110000",
  25710=>"000000010",
  25711=>"011111111",
  25712=>"111111111",
  25713=>"111111111",
  25714=>"100100000",
  25715=>"100100000",
  25716=>"000000100",
  25717=>"111111110",
  25718=>"000001000",
  25719=>"110010011",
  25720=>"110000000",
  25721=>"000111111",
  25722=>"101000000",
  25723=>"111110000",
  25724=>"110111111",
  25725=>"111010000",
  25726=>"000000011",
  25727=>"001000101",
  25728=>"111111000",
  25729=>"010010111",
  25730=>"111011001",
  25731=>"000011110",
  25732=>"000110111",
  25733=>"000100100",
  25734=>"001111111",
  25735=>"011011111",
  25736=>"100000111",
  25737=>"111111111",
  25738=>"111000000",
  25739=>"111100110",
  25740=>"111111110",
  25741=>"000111111",
  25742=>"111111111",
  25743=>"000011000",
  25744=>"000001111",
  25745=>"111111001",
  25746=>"001111111",
  25747=>"101101111",
  25748=>"010101111",
  25749=>"110110100",
  25750=>"000000101",
  25751=>"000000001",
  25752=>"000000100",
  25753=>"111111000",
  25754=>"000011010",
  25755=>"100100111",
  25756=>"000000111",
  25757=>"110100110",
  25758=>"001111111",
  25759=>"011011111",
  25760=>"111111110",
  25761=>"111111000",
  25762=>"011111111",
  25763=>"111111110",
  25764=>"111001001",
  25765=>"110110000",
  25766=>"000111110",
  25767=>"011111011",
  25768=>"000000000",
  25769=>"000000000",
  25770=>"000011111",
  25771=>"110111000",
  25772=>"010010100",
  25773=>"100110110",
  25774=>"010010000",
  25775=>"000000001",
  25776=>"100000000",
  25777=>"110100000",
  25778=>"011011011",
  25779=>"000101000",
  25780=>"110000000",
  25781=>"111111000",
  25782=>"111110000",
  25783=>"111111111",
  25784=>"010011011",
  25785=>"001000111",
  25786=>"111000000",
  25787=>"110000011",
  25788=>"000000111",
  25789=>"111110110",
  25790=>"000111111",
  25791=>"111100100",
  25792=>"001100110",
  25793=>"011011011",
  25794=>"100101111",
  25795=>"111001111",
  25796=>"000000001",
  25797=>"000001111",
  25798=>"111110000",
  25799=>"000100111",
  25800=>"000000000",
  25801=>"000000110",
  25802=>"000000000",
  25803=>"111001001",
  25804=>"001011111",
  25805=>"110110100",
  25806=>"000000001",
  25807=>"110111111",
  25808=>"101100100",
  25809=>"110111001",
  25810=>"111110000",
  25811=>"000000000",
  25812=>"111110110",
  25813=>"111111000",
  25814=>"001111000",
  25815=>"010000010",
  25816=>"011000101",
  25817=>"011111100",
  25818=>"111111000",
  25819=>"000000000",
  25820=>"000000111",
  25821=>"001111001",
  25822=>"111111111",
  25823=>"011001001",
  25824=>"101111000",
  25825=>"001000111",
  25826=>"011000000",
  25827=>"000111011",
  25828=>"110111010",
  25829=>"110001111",
  25830=>"000111111",
  25831=>"000100000",
  25832=>"111111000",
  25833=>"100100111",
  25834=>"111111111",
  25835=>"010101111",
  25836=>"000101111",
  25837=>"001001000",
  25838=>"111001000",
  25839=>"111111000",
  25840=>"000000001",
  25841=>"000000111",
  25842=>"110110111",
  25843=>"000011111",
  25844=>"011100000",
  25845=>"000000100",
  25846=>"000110110",
  25847=>"001000100",
  25848=>"111111111",
  25849=>"111111111",
  25850=>"111111001",
  25851=>"111111111",
  25852=>"010110111",
  25853=>"100000101",
  25854=>"000111111",
  25855=>"000010000",
  25856=>"011011010",
  25857=>"011011011",
  25858=>"111101000",
  25859=>"000101111",
  25860=>"000000010",
  25861=>"111111000",
  25862=>"110001000",
  25863=>"010011111",
  25864=>"000010111",
  25865=>"000000000",
  25866=>"000100100",
  25867=>"111111111",
  25868=>"111001011",
  25869=>"000000000",
  25870=>"000111000",
  25871=>"000111111",
  25872=>"111000000",
  25873=>"111111111",
  25874=>"111111000",
  25875=>"111011111",
  25876=>"000000000",
  25877=>"100000110",
  25878=>"000011011",
  25879=>"000100100",
  25880=>"010011000",
  25881=>"110000000",
  25882=>"000111111",
  25883=>"000001001",
  25884=>"000111100",
  25885=>"000000000",
  25886=>"111111111",
  25887=>"111111101",
  25888=>"011111111",
  25889=>"000111111",
  25890=>"000000000",
  25891=>"000100110",
  25892=>"001001111",
  25893=>"000100111",
  25894=>"100011001",
  25895=>"000000110",
  25896=>"111110111",
  25897=>"111111111",
  25898=>"110011001",
  25899=>"100100000",
  25900=>"111011110",
  25901=>"000000111",
  25902=>"000100000",
  25903=>"011001001",
  25904=>"011110000",
  25905=>"010111110",
  25906=>"000000111",
  25907=>"011111110",
  25908=>"111101000",
  25909=>"001100110",
  25910=>"011111111",
  25911=>"110110001",
  25912=>"000000111",
  25913=>"101100111",
  25914=>"111000000",
  25915=>"111000110",
  25916=>"011111110",
  25917=>"110100100",
  25918=>"000000000",
  25919=>"110000000",
  25920=>"001111001",
  25921=>"000110111",
  25922=>"000000110",
  25923=>"111000000",
  25924=>"110111111",
  25925=>"010000011",
  25926=>"111000000",
  25927=>"111000000",
  25928=>"001001000",
  25929=>"111011101",
  25930=>"000000000",
  25931=>"001001011",
  25932=>"011111100",
  25933=>"000111011",
  25934=>"000011011",
  25935=>"011001000",
  25936=>"010011010",
  25937=>"100000001",
  25938=>"110111111",
  25939=>"011100100",
  25940=>"000011011",
  25941=>"110110111",
  25942=>"000000000",
  25943=>"110111111",
  25944=>"000000000",
  25945=>"000101000",
  25946=>"010000000",
  25947=>"000011111",
  25948=>"101101101",
  25949=>"111010111",
  25950=>"000000000",
  25951=>"110100101",
  25952=>"000101101",
  25953=>"000111111",
  25954=>"000010111",
  25955=>"000000111",
  25956=>"111110000",
  25957=>"100111111",
  25958=>"011000000",
  25959=>"110110110",
  25960=>"000000111",
  25961=>"111111010",
  25962=>"111100110",
  25963=>"111100000",
  25964=>"110011010",
  25965=>"110000111",
  25966=>"000000100",
  25967=>"000000000",
  25968=>"000001111",
  25969=>"111111011",
  25970=>"000000111",
  25971=>"111000000",
  25972=>"100111111",
  25973=>"000010000",
  25974=>"100111111",
  25975=>"000000000",
  25976=>"011000000",
  25977=>"111111111",
  25978=>"010000000",
  25979=>"111111111",
  25980=>"000000000",
  25981=>"000111111",
  25982=>"000000000",
  25983=>"111000000",
  25984=>"000010000",
  25985=>"000000100",
  25986=>"100100000",
  25987=>"100000000",
  25988=>"111111000",
  25989=>"000100111",
  25990=>"000111111",
  25991=>"011001111",
  25992=>"111000000",
  25993=>"000111111",
  25994=>"111111100",
  25995=>"101101000",
  25996=>"000111111",
  25997=>"010010011",
  25998=>"000011000",
  25999=>"000000100",
  26000=>"100000100",
  26001=>"010011001",
  26002=>"001011011",
  26003=>"110111111",
  26004=>"111111111",
  26005=>"110110010",
  26006=>"000001000",
  26007=>"110001111",
  26008=>"110111100",
  26009=>"000000111",
  26010=>"000000000",
  26011=>"110000000",
  26012=>"010110111",
  26013=>"011111111",
  26014=>"111000000",
  26015=>"100110101",
  26016=>"111101111",
  26017=>"000110010",
  26018=>"110011011",
  26019=>"000000000",
  26020=>"010000000",
  26021=>"111000000",
  26022=>"111011000",
  26023=>"111111111",
  26024=>"000000100",
  26025=>"000111000",
  26026=>"010111110",
  26027=>"111111000",
  26028=>"000000100",
  26029=>"011000000",
  26030=>"000111111",
  26031=>"100000000",
  26032=>"011011111",
  26033=>"100100111",
  26034=>"111111111",
  26035=>"000001101",
  26036=>"111111111",
  26037=>"000000011",
  26038=>"111111111",
  26039=>"000110010",
  26040=>"000000111",
  26041=>"011011001",
  26042=>"100100111",
  26043=>"111110000",
  26044=>"001111111",
  26045=>"110000000",
  26046=>"000001011",
  26047=>"100110010",
  26048=>"000000000",
  26049=>"111000000",
  26050=>"000000000",
  26051=>"000111111",
  26052=>"000000101",
  26053=>"110110111",
  26054=>"000000101",
  26055=>"101001000",
  26056=>"001111111",
  26057=>"001111111",
  26058=>"000111111",
  26059=>"001000000",
  26060=>"111110000",
  26061=>"000111111",
  26062=>"000010110",
  26063=>"000100001",
  26064=>"001011001",
  26065=>"111000110",
  26066=>"111011100",
  26067=>"001101101",
  26068=>"000110110",
  26069=>"000111111",
  26070=>"111111110",
  26071=>"111111001",
  26072=>"110100000",
  26073=>"001111111",
  26074=>"011111110",
  26075=>"010011000",
  26076=>"111111010",
  26077=>"111111101",
  26078=>"000110000",
  26079=>"110001001",
  26080=>"101101111",
  26081=>"111011001",
  26082=>"111101000",
  26083=>"110000000",
  26084=>"000111111",
  26085=>"000000001",
  26086=>"101001000",
  26087=>"111111111",
  26088=>"001010011",
  26089=>"001100000",
  26090=>"000000000",
  26091=>"000000000",
  26092=>"111100000",
  26093=>"001000000",
  26094=>"111111001",
  26095=>"000000000",
  26096=>"111000000",
  26097=>"111110000",
  26098=>"000000111",
  26099=>"001001011",
  26100=>"111011111",
  26101=>"111110100",
  26102=>"001111111",
  26103=>"100000001",
  26104=>"000000000",
  26105=>"011001001",
  26106=>"000000001",
  26107=>"000100000",
  26108=>"111111101",
  26109=>"010010000",
  26110=>"111011000",
  26111=>"111000000",
  26112=>"110110100",
  26113=>"000001000",
  26114=>"111110110",
  26115=>"111111001",
  26116=>"111111111",
  26117=>"100000000",
  26118=>"000000100",
  26119=>"001001001",
  26120=>"000000101",
  26121=>"111111111",
  26122=>"001001101",
  26123=>"000101111",
  26124=>"111110110",
  26125=>"001100000",
  26126=>"000000110",
  26127=>"111111111",
  26128=>"101101000",
  26129=>"000001001",
  26130=>"111111101",
  26131=>"000000000",
  26132=>"000011000",
  26133=>"110111111",
  26134=>"100000001",
  26135=>"111011001",
  26136=>"000000000",
  26137=>"000000100",
  26138=>"000001000",
  26139=>"100100100",
  26140=>"111111111",
  26141=>"110110111",
  26142=>"100110110",
  26143=>"110000000",
  26144=>"001000100",
  26145=>"000100000",
  26146=>"100100110",
  26147=>"111101101",
  26148=>"111111111",
  26149=>"000000000",
  26150=>"111111111",
  26151=>"011111111",
  26152=>"001011111",
  26153=>"000111111",
  26154=>"000000000",
  26155=>"000111000",
  26156=>"001000000",
  26157=>"111111111",
  26158=>"111110111",
  26159=>"111101100",
  26160=>"001110100",
  26161=>"111111000",
  26162=>"011011011",
  26163=>"000000000",
  26164=>"110110111",
  26165=>"010010011",
  26166=>"000000000",
  26167=>"000000001",
  26168=>"000100111",
  26169=>"011011000",
  26170=>"000000000",
  26171=>"000000111",
  26172=>"111111010",
  26173=>"000000000",
  26174=>"111010000",
  26175=>"111111100",
  26176=>"001000100",
  26177=>"001011111",
  26178=>"111111111",
  26179=>"000000000",
  26180=>"000100110",
  26181=>"000000000",
  26182=>"111011000",
  26183=>"111111100",
  26184=>"000010110",
  26185=>"001000101",
  26186=>"110000100",
  26187=>"000100100",
  26188=>"000000000",
  26189=>"111111110",
  26190=>"100010000",
  26191=>"000000111",
  26192=>"000001000",
  26193=>"000000000",
  26194=>"000000000",
  26195=>"010110110",
  26196=>"111110000",
  26197=>"011010000",
  26198=>"101111011",
  26199=>"110111111",
  26200=>"100111111",
  26201=>"101101111",
  26202=>"000100100",
  26203=>"001011011",
  26204=>"001001000",
  26205=>"111111011",
  26206=>"000001000",
  26207=>"001000000",
  26208=>"000000000",
  26209=>"111111111",
  26210=>"111111111",
  26211=>"011000111",
  26212=>"111100000",
  26213=>"000000000",
  26214=>"000000000",
  26215=>"111111000",
  26216=>"111111111",
  26217=>"000000110",
  26218=>"000000000",
  26219=>"000010110",
  26220=>"010000000",
  26221=>"111111101",
  26222=>"111111111",
  26223=>"111110000",
  26224=>"000000000",
  26225=>"000000000",
  26226=>"011011111",
  26227=>"000000101",
  26228=>"111111111",
  26229=>"000111111",
  26230=>"111111100",
  26231=>"000010111",
  26232=>"011111111",
  26233=>"111111000",
  26234=>"110111101",
  26235=>"111111111",
  26236=>"111111111",
  26237=>"110011011",
  26238=>"101101111",
  26239=>"111111111",
  26240=>"000111011",
  26241=>"110111111",
  26242=>"000000111",
  26243=>"000000000",
  26244=>"111101001",
  26245=>"111111111",
  26246=>"000101111",
  26247=>"000000000",
  26248=>"111111111",
  26249=>"111110000",
  26250=>"000000000",
  26251=>"101001101",
  26252=>"111001000",
  26253=>"000000111",
  26254=>"000000000",
  26255=>"000110100",
  26256=>"111011111",
  26257=>"111111111",
  26258=>"000000000",
  26259=>"010111000",
  26260=>"101101100",
  26261=>"000000000",
  26262=>"000000000",
  26263=>"001101101",
  26264=>"111100000",
  26265=>"100100110",
  26266=>"111111111",
  26267=>"011010000",
  26268=>"000001001",
  26269=>"000000000",
  26270=>"111011001",
  26271=>"000000000",
  26272=>"000100000",
  26273=>"110111111",
  26274=>"010111000",
  26275=>"111111111",
  26276=>"111101001",
  26277=>"100111111",
  26278=>"010110010",
  26279=>"000000011",
  26280=>"000011110",
  26281=>"111100100",
  26282=>"100110110",
  26283=>"110000000",
  26284=>"000000001",
  26285=>"100110000",
  26286=>"111111111",
  26287=>"000000000",
  26288=>"000000000",
  26289=>"001001001",
  26290=>"110110110",
  26291=>"000000000",
  26292=>"000000000",
  26293=>"111111100",
  26294=>"111001000",
  26295=>"100000001",
  26296=>"001000000",
  26297=>"010110010",
  26298=>"101001001",
  26299=>"111011111",
  26300=>"110111011",
  26301=>"000001001",
  26302=>"110100110",
  26303=>"101001000",
  26304=>"000000000",
  26305=>"000000000",
  26306=>"111011011",
  26307=>"111000000",
  26308=>"100000100",
  26309=>"101101001",
  26310=>"111111101",
  26311=>"111111000",
  26312=>"000110111",
  26313=>"101111111",
  26314=>"001101101",
  26315=>"110000000",
  26316=>"111111111",
  26317=>"000001111",
  26318=>"000000000",
  26319=>"111111100",
  26320=>"111110000",
  26321=>"100100000",
  26322=>"111111111",
  26323=>"110100000",
  26324=>"001000000",
  26325=>"000000100",
  26326=>"000010000",
  26327=>"100111011",
  26328=>"000000000",
  26329=>"010111111",
  26330=>"000110000",
  26331=>"000000111",
  26332=>"100110111",
  26333=>"111110111",
  26334=>"011111111",
  26335=>"100111111",
  26336=>"000000000",
  26337=>"010110111",
  26338=>"001000000",
  26339=>"111111001",
  26340=>"000000000",
  26341=>"000011011",
  26342=>"000100100",
  26343=>"111101000",
  26344=>"111111000",
  26345=>"011001001",
  26346=>"111011011",
  26347=>"111111111",
  26348=>"000000000",
  26349=>"010000011",
  26350=>"000000111",
  26351=>"110111110",
  26352=>"101001110",
  26353=>"001000001",
  26354=>"010000000",
  26355=>"001011010",
  26356=>"111111111",
  26357=>"100000000",
  26358=>"111111110",
  26359=>"111111111",
  26360=>"000000000",
  26361=>"100000000",
  26362=>"000001000",
  26363=>"101111111",
  26364=>"011111111",
  26365=>"000001001",
  26366=>"111111000",
  26367=>"100111100",
  26368=>"011001001",
  26369=>"111111111",
  26370=>"111111111",
  26371=>"100111111",
  26372=>"000101111",
  26373=>"111111111",
  26374=>"111111100",
  26375=>"111111110",
  26376=>"001011001",
  26377=>"000111000",
  26378=>"100000000",
  26379=>"000101001",
  26380=>"110110111",
  26381=>"101111111",
  26382=>"010000010",
  26383=>"001100100",
  26384=>"000000000",
  26385=>"000000000",
  26386=>"111111111",
  26387=>"111111111",
  26388=>"000111010",
  26389=>"001000110",
  26390=>"111100000",
  26391=>"000000000",
  26392=>"101101111",
  26393=>"111101000",
  26394=>"000000000",
  26395=>"000000100",
  26396=>"111111110",
  26397=>"000000000",
  26398=>"110100111",
  26399=>"000000000",
  26400=>"111111111",
  26401=>"000111100",
  26402=>"000000000",
  26403=>"111111111",
  26404=>"001000000",
  26405=>"111111111",
  26406=>"111111111",
  26407=>"100000000",
  26408=>"000100110",
  26409=>"110000000",
  26410=>"111011000",
  26411=>"001001000",
  26412=>"000010010",
  26413=>"111001111",
  26414=>"000000000",
  26415=>"000001111",
  26416=>"001000000",
  26417=>"001011011",
  26418=>"000000010",
  26419=>"111111000",
  26420=>"000000000",
  26421=>"100111111",
  26422=>"100111111",
  26423=>"111000001",
  26424=>"000000000",
  26425=>"101101111",
  26426=>"110111111",
  26427=>"111101111",
  26428=>"000010110",
  26429=>"111111110",
  26430=>"101101001",
  26431=>"000000000",
  26432=>"000000000",
  26433=>"101000000",
  26434=>"000000000",
  26435=>"111111111",
  26436=>"100110111",
  26437=>"000000000",
  26438=>"101111110",
  26439=>"100100000",
  26440=>"000111111",
  26441=>"000000000",
  26442=>"000000000",
  26443=>"111101000",
  26444=>"111001000",
  26445=>"010010000",
  26446=>"000000000",
  26447=>"011011011",
  26448=>"100010011",
  26449=>"000000100",
  26450=>"111111111",
  26451=>"000000000",
  26452=>"111111111",
  26453=>"011011011",
  26454=>"111111001",
  26455=>"000111111",
  26456=>"111111111",
  26457=>"111101111",
  26458=>"000000000",
  26459=>"011000000",
  26460=>"110110000",
  26461=>"000000000",
  26462=>"111111111",
  26463=>"011111001",
  26464=>"100000000",
  26465=>"111111100",
  26466=>"011011011",
  26467=>"000000000",
  26468=>"001001000",
  26469=>"010111111",
  26470=>"011000000",
  26471=>"000001111",
  26472=>"010010000",
  26473=>"000000000",
  26474=>"110001000",
  26475=>"100100101",
  26476=>"000000000",
  26477=>"101111111",
  26478=>"000111111",
  26479=>"000111111",
  26480=>"111111111",
  26481=>"001111111",
  26482=>"111011011",
  26483=>"111111111",
  26484=>"000111111",
  26485=>"111111111",
  26486=>"000000111",
  26487=>"111111111",
  26488=>"000000000",
  26489=>"000000000",
  26490=>"000111011",
  26491=>"000111111",
  26492=>"100100100",
  26493=>"111111111",
  26494=>"000000000",
  26495=>"000000000",
  26496=>"001011111",
  26497=>"111111111",
  26498=>"000000000",
  26499=>"111111111",
  26500=>"000001001",
  26501=>"100100101",
  26502=>"000000100",
  26503=>"101000101",
  26504=>"000111111",
  26505=>"000000001",
  26506=>"000000000",
  26507=>"001000001",
  26508=>"111111111",
  26509=>"111111110",
  26510=>"001001000",
  26511=>"000000011",
  26512=>"000000000",
  26513=>"000000000",
  26514=>"010010000",
  26515=>"100110000",
  26516=>"000100000",
  26517=>"000000001",
  26518=>"111111111",
  26519=>"111111111",
  26520=>"100000111",
  26521=>"011110100",
  26522=>"111111100",
  26523=>"000000000",
  26524=>"000000000",
  26525=>"000000010",
  26526=>"101101111",
  26527=>"110111000",
  26528=>"111111111",
  26529=>"111111111",
  26530=>"000110111",
  26531=>"000000000",
  26532=>"100100000",
  26533=>"000000000",
  26534=>"111111111",
  26535=>"000000011",
  26536=>"111000111",
  26537=>"111111111",
  26538=>"000000100",
  26539=>"011001001",
  26540=>"000000000",
  26541=>"111111111",
  26542=>"001001000",
  26543=>"111111111",
  26544=>"111111000",
  26545=>"111111100",
  26546=>"111111111",
  26547=>"111111111",
  26548=>"111111111",
  26549=>"100100101",
  26550=>"111111111",
  26551=>"111111000",
  26552=>"111111111",
  26553=>"111000000",
  26554=>"011001000",
  26555=>"111111111",
  26556=>"000000000",
  26557=>"000000000",
  26558=>"111000011",
  26559=>"001001001",
  26560=>"111011000",
  26561=>"010010000",
  26562=>"000001111",
  26563=>"011011011",
  26564=>"111111111",
  26565=>"001011001",
  26566=>"111111111",
  26567=>"000101111",
  26568=>"111111000",
  26569=>"111001101",
  26570=>"000111111",
  26571=>"000000000",
  26572=>"110010000",
  26573=>"000000000",
  26574=>"111111000",
  26575=>"111111111",
  26576=>"000111011",
  26577=>"000000000",
  26578=>"000000111",
  26579=>"011011011",
  26580=>"000000000",
  26581=>"111111111",
  26582=>"000000000",
  26583=>"111000111",
  26584=>"000010111",
  26585=>"000000000",
  26586=>"110000000",
  26587=>"111111001",
  26588=>"000000111",
  26589=>"000010110",
  26590=>"111011000",
  26591=>"100000000",
  26592=>"111111111",
  26593=>"001101100",
  26594=>"000011000",
  26595=>"000000000",
  26596=>"001000101",
  26597=>"000000000",
  26598=>"000000000",
  26599=>"011110000",
  26600=>"111111110",
  26601=>"000000011",
  26602=>"000001111",
  26603=>"000100100",
  26604=>"101111111",
  26605=>"110110110",
  26606=>"111111111",
  26607=>"111111111",
  26608=>"111111100",
  26609=>"110111111",
  26610=>"000000000",
  26611=>"111100000",
  26612=>"000000000",
  26613=>"111111000",
  26614=>"100000000",
  26615=>"000110100",
  26616=>"111111111",
  26617=>"000000000",
  26618=>"101000000",
  26619=>"000000000",
  26620=>"100000110",
  26621=>"111101100",
  26622=>"000000000",
  26623=>"000000000",
  26624=>"000110111",
  26625=>"111000000",
  26626=>"000100111",
  26627=>"011111111",
  26628=>"111011011",
  26629=>"000000000",
  26630=>"000000000",
  26631=>"111111111",
  26632=>"111111111",
  26633=>"111111000",
  26634=>"000000000",
  26635=>"111101111",
  26636=>"110100100",
  26637=>"000000000",
  26638=>"011000000",
  26639=>"011011001",
  26640=>"111000011",
  26641=>"000000001",
  26642=>"111000000",
  26643=>"111001101",
  26644=>"000000101",
  26645=>"111111111",
  26646=>"000011111",
  26647=>"111000111",
  26648=>"000000000",
  26649=>"100100110",
  26650=>"111111000",
  26651=>"111000110",
  26652=>"101001001",
  26653=>"100110000",
  26654=>"001001001",
  26655=>"000111000",
  26656=>"111000000",
  26657=>"111100010",
  26658=>"000000000",
  26659=>"000000000",
  26660=>"100110111",
  26661=>"111111111",
  26662=>"000111111",
  26663=>"001111001",
  26664=>"100000001",
  26665=>"000000000",
  26666=>"011001000",
  26667=>"000000000",
  26668=>"110101111",
  26669=>"011000000",
  26670=>"000000000",
  26671=>"100101111",
  26672=>"000000111",
  26673=>"001111000",
  26674=>"001000100",
  26675=>"111111111",
  26676=>"110110000",
  26677=>"011011000",
  26678=>"111111000",
  26679=>"010000000",
  26680=>"111111100",
  26681=>"000010111",
  26682=>"000000111",
  26683=>"111111000",
  26684=>"111110000",
  26685=>"011111000",
  26686=>"010011111",
  26687=>"000001111",
  26688=>"001001011",
  26689=>"000000000",
  26690=>"000000001",
  26691=>"000000001",
  26692=>"110000000",
  26693=>"101100111",
  26694=>"000000000",
  26695=>"111111111",
  26696=>"001111110",
  26697=>"100000000",
  26698=>"111011001",
  26699=>"010111000",
  26700=>"010111111",
  26701=>"000000011",
  26702=>"000000100",
  26703=>"000000000",
  26704=>"011001111",
  26705=>"000000000",
  26706=>"111000000",
  26707=>"100100000",
  26708=>"000000000",
  26709=>"111111000",
  26710=>"000010000",
  26711=>"011011000",
  26712=>"000000000",
  26713=>"000100111",
  26714=>"000100111",
  26715=>"111001101",
  26716=>"111010000",
  26717=>"111111111",
  26718=>"001111000",
  26719=>"000000111",
  26720=>"000111111",
  26721=>"000000000",
  26722=>"000000000",
  26723=>"110000000",
  26724=>"100111111",
  26725=>"100100000",
  26726=>"000000001",
  26727=>"111000000",
  26728=>"001111000",
  26729=>"111111111",
  26730=>"101111111",
  26731=>"000000000",
  26732=>"100110110",
  26733=>"111111000",
  26734=>"110000000",
  26735=>"111111011",
  26736=>"111111101",
  26737=>"111111111",
  26738=>"111100000",
  26739=>"001111000",
  26740=>"111111111",
  26741=>"000001101",
  26742=>"010000000",
  26743=>"000000000",
  26744=>"101000000",
  26745=>"000111111",
  26746=>"000000000",
  26747=>"111111011",
  26748=>"000000000",
  26749=>"000000001",
  26750=>"101101111",
  26751=>"010000000",
  26752=>"111111100",
  26753=>"111111110",
  26754=>"100000111",
  26755=>"011111001",
  26756=>"111101111",
  26757=>"000100111",
  26758=>"000000111",
  26759=>"111010110",
  26760=>"101100111",
  26761=>"111111111",
  26762=>"011111000",
  26763=>"111111100",
  26764=>"110000011",
  26765=>"010111000",
  26766=>"011011010",
  26767=>"001001000",
  26768=>"000001000",
  26769=>"111001000",
  26770=>"110111111",
  26771=>"010010000",
  26772=>"000000100",
  26773=>"000000100",
  26774=>"000000000",
  26775=>"000000000",
  26776=>"000000111",
  26777=>"111111111",
  26778=>"111000000",
  26779=>"000000010",
  26780=>"000000001",
  26781=>"001000000",
  26782=>"000000110",
  26783=>"000000000",
  26784=>"111100000",
  26785=>"000000000",
  26786=>"000000000",
  26787=>"111011111",
  26788=>"100000000",
  26789=>"000000010",
  26790=>"111111000",
  26791=>"010010000",
  26792=>"000111000",
  26793=>"000000000",
  26794=>"100110111",
  26795=>"110111111",
  26796=>"000011111",
  26797=>"000011011",
  26798=>"111111101",
  26799=>"101101100",
  26800=>"000100111",
  26801=>"011111001",
  26802=>"111110111",
  26803=>"111100000",
  26804=>"111111111",
  26805=>"010000000",
  26806=>"000000000",
  26807=>"000000011",
  26808=>"110111111",
  26809=>"111111000",
  26810=>"000010000",
  26811=>"000110111",
  26812=>"111110000",
  26813=>"111001001",
  26814=>"110000000",
  26815=>"111111111",
  26816=>"100000000",
  26817=>"100111111",
  26818=>"111111001",
  26819=>"000111111",
  26820=>"000111111",
  26821=>"100011000",
  26822=>"110011011",
  26823=>"111110110",
  26824=>"011101111",
  26825=>"111111111",
  26826=>"000101111",
  26827=>"101101010",
  26828=>"000111110",
  26829=>"000000100",
  26830=>"100111111",
  26831=>"000000000",
  26832=>"110111111",
  26833=>"001000111",
  26834=>"000101111",
  26835=>"000000111",
  26836=>"000000000",
  26837=>"111110110",
  26838=>"111101111",
  26839=>"111010000",
  26840=>"000111011",
  26841=>"001101100",
  26842=>"111101000",
  26843=>"111000000",
  26844=>"000000111",
  26845=>"001000110",
  26846=>"101000111",
  26847=>"000001000",
  26848=>"010110110",
  26849=>"110010000",
  26850=>"111110111",
  26851=>"111111000",
  26852=>"110110000",
  26853=>"111111111",
  26854=>"111011000",
  26855=>"000000000",
  26856=>"111111001",
  26857=>"011011000",
  26858=>"111101000",
  26859=>"101000111",
  26860=>"111111000",
  26861=>"100000101",
  26862=>"111111111",
  26863=>"111000000",
  26864=>"001000001",
  26865=>"011000111",
  26866=>"110000101",
  26867=>"111000000",
  26868=>"000011000",
  26869=>"010011000",
  26870=>"100110011",
  26871=>"111111111",
  26872=>"000110110",
  26873=>"111100100",
  26874=>"000000000",
  26875=>"000111111",
  26876=>"111010000",
  26877=>"110111010",
  26878=>"011011111",
  26879=>"000100111",
  26880=>"000000000",
  26881=>"111111000",
  26882=>"111110111",
  26883=>"001111111",
  26884=>"111100111",
  26885=>"111101101",
  26886=>"001000000",
  26887=>"000000000",
  26888=>"000000000",
  26889=>"100110110",
  26890=>"110000000",
  26891=>"000000000",
  26892=>"000100110",
  26893=>"000110111",
  26894=>"101101100",
  26895=>"110000000",
  26896=>"000000110",
  26897=>"111011000",
  26898=>"000000000",
  26899=>"000110110",
  26900=>"000100111",
  26901=>"000111111",
  26902=>"111011011",
  26903=>"001111000",
  26904=>"111001001",
  26905=>"000111111",
  26906=>"000000001",
  26907=>"111110111",
  26908=>"111111000",
  26909=>"011000010",
  26910=>"001000001",
  26911=>"111111111",
  26912=>"000110100",
  26913=>"111111000",
  26914=>"100000000",
  26915=>"111001000",
  26916=>"111111111",
  26917=>"111000000",
  26918=>"010000000",
  26919=>"000010000",
  26920=>"000000111",
  26921=>"001000000",
  26922=>"110110111",
  26923=>"011000000",
  26924=>"001001000",
  26925=>"001011111",
  26926=>"000111000",
  26927=>"011111000",
  26928=>"000000110",
  26929=>"111000001",
  26930=>"111001001",
  26931=>"101101111",
  26932=>"110000000",
  26933=>"000110111",
  26934=>"000011111",
  26935=>"000000110",
  26936=>"011011000",
  26937=>"111101000",
  26938=>"111011000",
  26939=>"001001000",
  26940=>"000000010",
  26941=>"000000000",
  26942=>"000001010",
  26943=>"111111111",
  26944=>"000000000",
  26945=>"111100000",
  26946=>"111111111",
  26947=>"111010000",
  26948=>"111111111",
  26949=>"111000000",
  26950=>"111111111",
  26951=>"000000111",
  26952=>"111111011",
  26953=>"110000000",
  26954=>"000000111",
  26955=>"111111111",
  26956=>"100100111",
  26957=>"000010010",
  26958=>"000111111",
  26959=>"001001000",
  26960=>"111011000",
  26961=>"000000000",
  26962=>"000000101",
  26963=>"110000000",
  26964=>"000000000",
  26965=>"000000011",
  26966=>"011111111",
  26967=>"111111111",
  26968=>"101111111",
  26969=>"001111111",
  26970=>"000111111",
  26971=>"000000111",
  26972=>"111101000",
  26973=>"110000000",
  26974=>"000000000",
  26975=>"000011011",
  26976=>"000000000",
  26977=>"000010001",
  26978=>"110110000",
  26979=>"111000000",
  26980=>"000000110",
  26981=>"000000001",
  26982=>"111101111",
  26983=>"000111111",
  26984=>"111111111",
  26985=>"111100100",
  26986=>"000000011",
  26987=>"110110010",
  26988=>"111111111",
  26989=>"000111110",
  26990=>"111011000",
  26991=>"010011000",
  26992=>"111111000",
  26993=>"000000000",
  26994=>"101110111",
  26995=>"000000000",
  26996=>"000001000",
  26997=>"001000001",
  26998=>"011111111",
  26999=>"111000000",
  27000=>"000000000",
  27001=>"111111000",
  27002=>"010000100",
  27003=>"000000000",
  27004=>"011011000",
  27005=>"000000000",
  27006=>"111111000",
  27007=>"000000000",
  27008=>"010011011",
  27009=>"111111111",
  27010=>"111111111",
  27011=>"111111111",
  27012=>"111000100",
  27013=>"000100100",
  27014=>"010000000",
  27015=>"111111111",
  27016=>"001010000",
  27017=>"111000000",
  27018=>"111110110",
  27019=>"110100111",
  27020=>"000000001",
  27021=>"001000010",
  27022=>"100110000",
  27023=>"101000000",
  27024=>"110010111",
  27025=>"111000001",
  27026=>"111100100",
  27027=>"000000000",
  27028=>"111111111",
  27029=>"001001000",
  27030=>"100111001",
  27031=>"000001001",
  27032=>"111111000",
  27033=>"000111000",
  27034=>"000000110",
  27035=>"111111111",
  27036=>"001000000",
  27037=>"111110111",
  27038=>"001011000",
  27039=>"000000000",
  27040=>"101100111",
  27041=>"111110001",
  27042=>"000000100",
  27043=>"000000000",
  27044=>"011111111",
  27045=>"000111111",
  27046=>"000000111",
  27047=>"111111111",
  27048=>"000000001",
  27049=>"011000000",
  27050=>"111000000",
  27051=>"000000000",
  27052=>"000000000",
  27053=>"100100110",
  27054=>"111011010",
  27055=>"011011101",
  27056=>"000110001",
  27057=>"000000111",
  27058=>"111101000",
  27059=>"000000000",
  27060=>"001111111",
  27061=>"000000000",
  27062=>"001000001",
  27063=>"000101111",
  27064=>"111111000",
  27065=>"111100000",
  27066=>"111000000",
  27067=>"101001111",
  27068=>"111111110",
  27069=>"111111111",
  27070=>"000000000",
  27071=>"011011011",
  27072=>"000000000",
  27073=>"111111111",
  27074=>"000110111",
  27075=>"111000000",
  27076=>"110110000",
  27077=>"011011110",
  27078=>"000000000",
  27079=>"110001000",
  27080=>"011000000",
  27081=>"000000000",
  27082=>"110000000",
  27083=>"000111010",
  27084=>"000000000",
  27085=>"111000111",
  27086=>"001000000",
  27087=>"110110110",
  27088=>"100100000",
  27089=>"111100111",
  27090=>"101001000",
  27091=>"111111111",
  27092=>"011000011",
  27093=>"110100000",
  27094=>"001011000",
  27095=>"001011001",
  27096=>"100111111",
  27097=>"111000000",
  27098=>"000000111",
  27099=>"000001111",
  27100=>"000000000",
  27101=>"000000000",
  27102=>"011000000",
  27103=>"000010011",
  27104=>"010111000",
  27105=>"111011000",
  27106=>"000000010",
  27107=>"011011111",
  27108=>"111001001",
  27109=>"000000111",
  27110=>"000000000",
  27111=>"000110111",
  27112=>"111111111",
  27113=>"000000000",
  27114=>"111100111",
  27115=>"000000000",
  27116=>"111000011",
  27117=>"011001100",
  27118=>"111001000",
  27119=>"111111001",
  27120=>"000000000",
  27121=>"000111111",
  27122=>"000000000",
  27123=>"011010000",
  27124=>"000000100",
  27125=>"111000000",
  27126=>"000000000",
  27127=>"111111101",
  27128=>"000111000",
  27129=>"100100000",
  27130=>"110111011",
  27131=>"000100000",
  27132=>"111011100",
  27133=>"111110110",
  27134=>"111000000",
  27135=>"100000000",
  27136=>"111000000",
  27137=>"111000000",
  27138=>"000000111",
  27139=>"111111111",
  27140=>"001000000",
  27141=>"111111111",
  27142=>"000001000",
  27143=>"100000000",
  27144=>"111111011",
  27145=>"000000000",
  27146=>"000100111",
  27147=>"111010010",
  27148=>"000000000",
  27149=>"000000000",
  27150=>"010010000",
  27151=>"111111111",
  27152=>"101101000",
  27153=>"000000000",
  27154=>"111000000",
  27155=>"010110111",
  27156=>"111111111",
  27157=>"111111111",
  27158=>"111011011",
  27159=>"111111111",
  27160=>"000000000",
  27161=>"000000010",
  27162=>"111111001",
  27163=>"001011111",
  27164=>"111000111",
  27165=>"011011000",
  27166=>"001001111",
  27167=>"000000001",
  27168=>"111111111",
  27169=>"000000111",
  27170=>"111101111",
  27171=>"111110111",
  27172=>"111011111",
  27173=>"000100000",
  27174=>"000000001",
  27175=>"000111111",
  27176=>"000000101",
  27177=>"111111110",
  27178=>"111111111",
  27179=>"111000100",
  27180=>"111111111",
  27181=>"111001000",
  27182=>"111111111",
  27183=>"111111101",
  27184=>"000000000",
  27185=>"111011111",
  27186=>"000000000",
  27187=>"011011011",
  27188=>"000000000",
  27189=>"110010100",
  27190=>"000000000",
  27191=>"001101111",
  27192=>"100000000",
  27193=>"000000000",
  27194=>"000011111",
  27195=>"000000000",
  27196=>"111111111",
  27197=>"000000000",
  27198=>"001011011",
  27199=>"111001111",
  27200=>"000011111",
  27201=>"000000000",
  27202=>"000000010",
  27203=>"111001000",
  27204=>"010000000",
  27205=>"111111011",
  27206=>"111000000",
  27207=>"100100100",
  27208=>"011000001",
  27209=>"000000111",
  27210=>"011011011",
  27211=>"100100001",
  27212=>"111011111",
  27213=>"000000000",
  27214=>"001000000",
  27215=>"000011000",
  27216=>"000000011",
  27217=>"001000000",
  27218=>"000000000",
  27219=>"111101000",
  27220=>"000000000",
  27221=>"111111011",
  27222=>"111000000",
  27223=>"111000001",
  27224=>"000000101",
  27225=>"111001111",
  27226=>"000000000",
  27227=>"000000000",
  27228=>"000000111",
  27229=>"000000111",
  27230=>"111111110",
  27231=>"111111100",
  27232=>"111000111",
  27233=>"010000000",
  27234=>"111111011",
  27235=>"100100111",
  27236=>"000000000",
  27237=>"111111000",
  27238=>"110111111",
  27239=>"111111111",
  27240=>"100000000",
  27241=>"111111111",
  27242=>"000000000",
  27243=>"111111111",
  27244=>"100100000",
  27245=>"100100111",
  27246=>"000000000",
  27247=>"011111111",
  27248=>"000000101",
  27249=>"001101010",
  27250=>"000010011",
  27251=>"110000110",
  27252=>"000000110",
  27253=>"000011111",
  27254=>"000010111",
  27255=>"101001111",
  27256=>"110110001",
  27257=>"111101001",
  27258=>"000000000",
  27259=>"000001111",
  27260=>"000000000",
  27261=>"000110111",
  27262=>"111111000",
  27263=>"000010110",
  27264=>"101111111",
  27265=>"111111111",
  27266=>"111100111",
  27267=>"111011001",
  27268=>"111001000",
  27269=>"111111111",
  27270=>"000000000",
  27271=>"000000000",
  27272=>"111111111",
  27273=>"001000000",
  27274=>"111111100",
  27275=>"010110010",
  27276=>"111111111",
  27277=>"010111111",
  27278=>"011001111",
  27279=>"110111010",
  27280=>"010000000",
  27281=>"111111111",
  27282=>"000000000",
  27283=>"110000000",
  27284=>"001111100",
  27285=>"001000001",
  27286=>"111111101",
  27287=>"111111101",
  27288=>"111111111",
  27289=>"000000000",
  27290=>"011111011",
  27291=>"000000110",
  27292=>"011000000",
  27293=>"010000000",
  27294=>"000000000",
  27295=>"000111111",
  27296=>"111000000",
  27297=>"000000000",
  27298=>"000000110",
  27299=>"111111001",
  27300=>"000000001",
  27301=>"111111111",
  27302=>"111101111",
  27303=>"011000000",
  27304=>"011110111",
  27305=>"000100000",
  27306=>"111111111",
  27307=>"110110111",
  27308=>"111111111",
  27309=>"110010000",
  27310=>"111111111",
  27311=>"111111111",
  27312=>"111111111",
  27313=>"110110111",
  27314=>"110111111",
  27315=>"111000000",
  27316=>"001000000",
  27317=>"001001111",
  27318=>"000111111",
  27319=>"000000000",
  27320=>"011111111",
  27321=>"000000000",
  27322=>"010110100",
  27323=>"101111111",
  27324=>"111011011",
  27325=>"001111111",
  27326=>"100000000",
  27327=>"111111111",
  27328=>"000000111",
  27329=>"000000000",
  27330=>"000000110",
  27331=>"110110110",
  27332=>"110000101",
  27333=>"111111110",
  27334=>"011001111",
  27335=>"000000000",
  27336=>"010010000",
  27337=>"111111111",
  27338=>"101111111",
  27339=>"000000111",
  27340=>"000000000",
  27341=>"000000111",
  27342=>"111111010",
  27343=>"001000000",
  27344=>"000000000",
  27345=>"000000110",
  27346=>"010110011",
  27347=>"000000111",
  27348=>"000000100",
  27349=>"000000000",
  27350=>"111000010",
  27351=>"111000000",
  27352=>"101000000",
  27353=>"111101101",
  27354=>"000000000",
  27355=>"000000000",
  27356=>"111111000",
  27357=>"000000000",
  27358=>"000000000",
  27359=>"111101111",
  27360=>"000000000",
  27361=>"001111111",
  27362=>"111111111",
  27363=>"000000000",
  27364=>"000000000",
  27365=>"111010111",
  27366=>"010000000",
  27367=>"001000000",
  27368=>"000001000",
  27369=>"111111111",
  27370=>"000000111",
  27371=>"111101100",
  27372=>"111111111",
  27373=>"011011011",
  27374=>"001000000",
  27375=>"000011111",
  27376=>"000100111",
  27377=>"011000000",
  27378=>"111111101",
  27379=>"000000101",
  27380=>"000000000",
  27381=>"000111111",
  27382=>"000000111",
  27383=>"000000000",
  27384=>"111111001",
  27385=>"111100000",
  27386=>"100111111",
  27387=>"011011011",
  27388=>"000000000",
  27389=>"010000000",
  27390=>"001100111",
  27391=>"000110110",
  27392=>"011011011",
  27393=>"110010000",
  27394=>"111111111",
  27395=>"110010011",
  27396=>"100100111",
  27397=>"001001111",
  27398=>"111101000",
  27399=>"000000000",
  27400=>"000000000",
  27401=>"000000000",
  27402=>"111111111",
  27403=>"001011111",
  27404=>"111111111",
  27405=>"000000000",
  27406=>"000001000",
  27407=>"100110100",
  27408=>"000000001",
  27409=>"011010000",
  27410=>"111111111",
  27411=>"000000000",
  27412=>"000001011",
  27413=>"000000000",
  27414=>"011011000",
  27415=>"111100000",
  27416=>"111000000",
  27417=>"110100101",
  27418=>"111011001",
  27419=>"000100100",
  27420=>"110111010",
  27421=>"000000100",
  27422=>"000000100",
  27423=>"010111111",
  27424=>"000000000",
  27425=>"000011111",
  27426=>"000000001",
  27427=>"000000000",
  27428=>"111110111",
  27429=>"111111111",
  27430=>"011000000",
  27431=>"001111111",
  27432=>"010011011",
  27433=>"000000000",
  27434=>"111111111",
  27435=>"111111011",
  27436=>"000000000",
  27437=>"100111111",
  27438=>"110111000",
  27439=>"110111000",
  27440=>"000000000",
  27441=>"000010001",
  27442=>"010111100",
  27443=>"110000000",
  27444=>"000000000",
  27445=>"001000000",
  27446=>"111111100",
  27447=>"111111111",
  27448=>"111111000",
  27449=>"111111111",
  27450=>"111111111",
  27451=>"100111111",
  27452=>"111111111",
  27453=>"000000010",
  27454=>"000111111",
  27455=>"110100000",
  27456=>"111111100",
  27457=>"000011011",
  27458=>"100110100",
  27459=>"111111111",
  27460=>"000000010",
  27461=>"111111111",
  27462=>"010000100",
  27463=>"011011000",
  27464=>"000000000",
  27465=>"111011111",
  27466=>"011001000",
  27467=>"101000000",
  27468=>"000000000",
  27469=>"100000000",
  27470=>"000000000",
  27471=>"001101111",
  27472=>"111011011",
  27473=>"000001100",
  27474=>"111011111",
  27475=>"100000000",
  27476=>"111111000",
  27477=>"011011011",
  27478=>"111111010",
  27479=>"111111111",
  27480=>"110111111",
  27481=>"111110111",
  27482=>"110110110",
  27483=>"001001010",
  27484=>"001000000",
  27485=>"000000000",
  27486=>"001111111",
  27487=>"111001000",
  27488=>"110110111",
  27489=>"111111101",
  27490=>"000000111",
  27491=>"111111111",
  27492=>"110111000",
  27493=>"111111111",
  27494=>"111000000",
  27495=>"110100000",
  27496=>"001011011",
  27497=>"010000000",
  27498=>"000000000",
  27499=>"010000000",
  27500=>"000000000",
  27501=>"000000000",
  27502=>"111111111",
  27503=>"010110110",
  27504=>"111010010",
  27505=>"100000000",
  27506=>"000000000",
  27507=>"111111111",
  27508=>"111100000",
  27509=>"111111100",
  27510=>"000000000",
  27511=>"000000000",
  27512=>"111000000",
  27513=>"011111000",
  27514=>"001111111",
  27515=>"000000000",
  27516=>"111111111",
  27517=>"000000000",
  27518=>"001000101",
  27519=>"101101111",
  27520=>"111111101",
  27521=>"100000000",
  27522=>"111111111",
  27523=>"111111111",
  27524=>"011011000",
  27525=>"110100110",
  27526=>"011111111",
  27527=>"010000000",
  27528=>"000000000",
  27529=>"111100100",
  27530=>"111111001",
  27531=>"111100000",
  27532=>"111111111",
  27533=>"010011000",
  27534=>"000000000",
  27535=>"110110000",
  27536=>"000000010",
  27537=>"110111111",
  27538=>"000000000",
  27539=>"111111111",
  27540=>"000000000",
  27541=>"000010010",
  27542=>"001000000",
  27543=>"100001000",
  27544=>"000000000",
  27545=>"000000000",
  27546=>"000000110",
  27547=>"110000000",
  27548=>"111111111",
  27549=>"111111110",
  27550=>"001001100",
  27551=>"001000000",
  27552=>"100010010",
  27553=>"001000011",
  27554=>"000000000",
  27555=>"100101111",
  27556=>"111111111",
  27557=>"111111010",
  27558=>"011000000",
  27559=>"000000111",
  27560=>"100111111",
  27561=>"100100111",
  27562=>"001001011",
  27563=>"011000101",
  27564=>"000000000",
  27565=>"000000000",
  27566=>"111111111",
  27567=>"111111111",
  27568=>"111111001",
  27569=>"000000000",
  27570=>"010110000",
  27571=>"011111111",
  27572=>"000000000",
  27573=>"101000001",
  27574=>"110110000",
  27575=>"011011111",
  27576=>"000000111",
  27577=>"000000000",
  27578=>"000000000",
  27579=>"100111111",
  27580=>"111001111",
  27581=>"100000000",
  27582=>"111111101",
  27583=>"110110010",
  27584=>"110000000",
  27585=>"100000000",
  27586=>"000000000",
  27587=>"111111110",
  27588=>"101000001",
  27589=>"110000100",
  27590=>"011001000",
  27591=>"000000000",
  27592=>"011001110",
  27593=>"000000000",
  27594=>"000100000",
  27595=>"111111000",
  27596=>"000000000",
  27597=>"111101100",
  27598=>"000000111",
  27599=>"000000000",
  27600=>"100000100",
  27601=>"000000000",
  27602=>"000000000",
  27603=>"010010110",
  27604=>"111111011",
  27605=>"001000011",
  27606=>"000000000",
  27607=>"000001111",
  27608=>"000000000",
  27609=>"111000001",
  27610=>"111111111",
  27611=>"011001101",
  27612=>"000000000",
  27613=>"101001000",
  27614=>"000000000",
  27615=>"011111111",
  27616=>"000000110",
  27617=>"000111111",
  27618=>"111111111",
  27619=>"000000000",
  27620=>"011111111",
  27621=>"000000000",
  27622=>"011000000",
  27623=>"000001011",
  27624=>"000000000",
  27625=>"000001001",
  27626=>"000100100",
  27627=>"010100000",
  27628=>"000000000",
  27629=>"000100110",
  27630=>"111111111",
  27631=>"000100111",
  27632=>"000000000",
  27633=>"111101111",
  27634=>"110000000",
  27635=>"000001000",
  27636=>"111111111",
  27637=>"000000000",
  27638=>"111111111",
  27639=>"000000100",
  27640=>"111111011",
  27641=>"001001100",
  27642=>"000111110",
  27643=>"100100110",
  27644=>"000000111",
  27645=>"000011111",
  27646=>"000011111",
  27647=>"111111111",
  27648=>"001001001",
  27649=>"111111111",
  27650=>"111111111",
  27651=>"111111000",
  27652=>"110110000",
  27653=>"001000001",
  27654=>"001001011",
  27655=>"111111111",
  27656=>"111111110",
  27657=>"111100101",
  27658=>"101001101",
  27659=>"111101111",
  27660=>"011011111",
  27661=>"111111111",
  27662=>"100100000",
  27663=>"000111111",
  27664=>"000000000",
  27665=>"111110110",
  27666=>"011001001",
  27667=>"000000101",
  27668=>"111111001",
  27669=>"000000000",
  27670=>"000000000",
  27671=>"111111111",
  27672=>"001001111",
  27673=>"011011001",
  27674=>"000111111",
  27675=>"001111101",
  27676=>"010000000",
  27677=>"111111111",
  27678=>"000000100",
  27679=>"000000000",
  27680=>"100100101",
  27681=>"111000000",
  27682=>"001001001",
  27683=>"001000000",
  27684=>"000000000",
  27685=>"110111110",
  27686=>"111101001",
  27687=>"111111100",
  27688=>"000000000",
  27689=>"000000000",
  27690=>"111011000",
  27691=>"000000000",
  27692=>"100000000",
  27693=>"111000000",
  27694=>"110110110",
  27695=>"101101101",
  27696=>"111111100",
  27697=>"000100000",
  27698=>"011000000",
  27699=>"011111111",
  27700=>"010101000",
  27701=>"100000000",
  27702=>"001101101",
  27703=>"000010110",
  27704=>"111111010",
  27705=>"000000000",
  27706=>"111111010",
  27707=>"010010000",
  27708=>"000001111",
  27709=>"111100000",
  27710=>"011111111",
  27711=>"111100100",
  27712=>"011011101",
  27713=>"010000000",
  27714=>"101000000",
  27715=>"000000000",
  27716=>"000001001",
  27717=>"111110110",
  27718=>"111111101",
  27719=>"100000000",
  27720=>"001011111",
  27721=>"001001111",
  27722=>"111111111",
  27723=>"111111111",
  27724=>"100000001",
  27725=>"111111111",
  27726=>"000000000",
  27727=>"000000000",
  27728=>"110111111",
  27729=>"011011010",
  27730=>"000000000",
  27731=>"111001100",
  27732=>"111111001",
  27733=>"011000000",
  27734=>"111101111",
  27735=>"111010111",
  27736=>"000101000",
  27737=>"000000000",
  27738=>"111110000",
  27739=>"110100100",
  27740=>"000110000",
  27741=>"001111111",
  27742=>"011111111",
  27743=>"000000000",
  27744=>"000000000",
  27745=>"000000001",
  27746=>"000000001",
  27747=>"000000000",
  27748=>"001111010",
  27749=>"011111111",
  27750=>"110100110",
  27751=>"111101001",
  27752=>"100111000",
  27753=>"111111111",
  27754=>"101000000",
  27755=>"111000000",
  27756=>"011110110",
  27757=>"110111111",
  27758=>"000000000",
  27759=>"100101100",
  27760=>"111111010",
  27761=>"111100000",
  27762=>"000001000",
  27763=>"011011011",
  27764=>"101001000",
  27765=>"001001000",
  27766=>"000000000",
  27767=>"111111101",
  27768=>"000101111",
  27769=>"111111101",
  27770=>"000000000",
  27771=>"111111111",
  27772=>"110010000",
  27773=>"111111010",
  27774=>"001110001",
  27775=>"001001011",
  27776=>"101111000",
  27777=>"000000111",
  27778=>"110000000",
  27779=>"100111111",
  27780=>"111111111",
  27781=>"000000100",
  27782=>"111111100",
  27783=>"001100111",
  27784=>"001111111",
  27785=>"000000000",
  27786=>"000000000",
  27787=>"110000000",
  27788=>"100000000",
  27789=>"111111110",
  27790=>"111111111",
  27791=>"111111011",
  27792=>"000000010",
  27793=>"111111111",
  27794=>"000000000",
  27795=>"000000000",
  27796=>"000100100",
  27797=>"000000111",
  27798=>"111111111",
  27799=>"100000000",
  27800=>"100000001",
  27801=>"111110111",
  27802=>"000000100",
  27803=>"001001000",
  27804=>"101111111",
  27805=>"000000000",
  27806=>"111111111",
  27807=>"001001001",
  27808=>"100111110",
  27809=>"111100000",
  27810=>"111111111",
  27811=>"110111011",
  27812=>"001001001",
  27813=>"011000000",
  27814=>"111111111",
  27815=>"011011001",
  27816=>"000000001",
  27817=>"000000001",
  27818=>"111000000",
  27819=>"111111111",
  27820=>"100100000",
  27821=>"111110110",
  27822=>"111111111",
  27823=>"000100000",
  27824=>"010010010",
  27825=>"100100000",
  27826=>"111111011",
  27827=>"111111111",
  27828=>"110110110",
  27829=>"100100101",
  27830=>"000000000",
  27831=>"010010111",
  27832=>"011000000",
  27833=>"111111111",
  27834=>"000000001",
  27835=>"111111111",
  27836=>"000000100",
  27837=>"000000000",
  27838=>"000000000",
  27839=>"000000000",
  27840=>"111111111",
  27841=>"001000000",
  27842=>"010000000",
  27843=>"001001000",
  27844=>"001001111",
  27845=>"000101111",
  27846=>"000001001",
  27847=>"101111001",
  27848=>"110110110",
  27849=>"000000001",
  27850=>"001000000",
  27851=>"111111111",
  27852=>"011111111",
  27853=>"000000110",
  27854=>"000000000",
  27855=>"111000000",
  27856=>"000000111",
  27857=>"000000000",
  27858=>"111111111",
  27859=>"000001101",
  27860=>"000000000",
  27861=>"111111111",
  27862=>"000111111",
  27863=>"001000100",
  27864=>"000111111",
  27865=>"111110110",
  27866=>"001000111",
  27867=>"111111111",
  27868=>"010111000",
  27869=>"101101111",
  27870=>"000000000",
  27871=>"101001111",
  27872=>"000000000",
  27873=>"011011000",
  27874=>"000010000",
  27875=>"000001111",
  27876=>"100100100",
  27877=>"000000111",
  27878=>"110111111",
  27879=>"111111111",
  27880=>"000000000",
  27881=>"000001111",
  27882=>"111111100",
  27883=>"110000000",
  27884=>"000000000",
  27885=>"011000000",
  27886=>"101000000",
  27887=>"000011000",
  27888=>"000111111",
  27889=>"111111111",
  27890=>"011111111",
  27891=>"000000000",
  27892=>"000000111",
  27893=>"011000100",
  27894=>"100001101",
  27895=>"001011010",
  27896=>"111101100",
  27897=>"111111111",
  27898=>"111111111",
  27899=>"000000111",
  27900=>"110110100",
  27901=>"000000000",
  27902=>"000100111",
  27903=>"111111101",
  27904=>"000000101",
  27905=>"000110110",
  27906=>"111111111",
  27907=>"000111101",
  27908=>"000000000",
  27909=>"111010000",
  27910=>"001000000",
  27911=>"001000101",
  27912=>"010110000",
  27913=>"111111000",
  27914=>"001000000",
  27915=>"111111111",
  27916=>"111001111",
  27917=>"111101001",
  27918=>"000000000",
  27919=>"000000000",
  27920=>"000000000",
  27921=>"000000111",
  27922=>"101001111",
  27923=>"011011111",
  27924=>"011000000",
  27925=>"111111010",
  27926=>"110000000",
  27927=>"111111111",
  27928=>"111111110",
  27929=>"100010011",
  27930=>"001000000",
  27931=>"111111111",
  27932=>"110100000",
  27933=>"000000111",
  27934=>"100000110",
  27935=>"000100111",
  27936=>"100001011",
  27937=>"111111111",
  27938=>"111001001",
  27939=>"111111111",
  27940=>"001000000",
  27941=>"001001101",
  27942=>"111100000",
  27943=>"000000001",
  27944=>"000000000",
  27945=>"111111001",
  27946=>"100000000",
  27947=>"111111000",
  27948=>"101000000",
  27949=>"000100111",
  27950=>"111111111",
  27951=>"111111000",
  27952=>"001001111",
  27953=>"111011001",
  27954=>"101000000",
  27955=>"000000000",
  27956=>"000000000",
  27957=>"000100111",
  27958=>"000000000",
  27959=>"011110100",
  27960=>"000000100",
  27961=>"111100100",
  27962=>"111101101",
  27963=>"000000111",
  27964=>"110110100",
  27965=>"111111010",
  27966=>"010000000",
  27967=>"110001111",
  27968=>"000000000",
  27969=>"000111111",
  27970=>"001101111",
  27971=>"000000000",
  27972=>"000000001",
  27973=>"111101111",
  27974=>"110111110",
  27975=>"101000001",
  27976=>"000000000",
  27977=>"000110111",
  27978=>"111111111",
  27979=>"000100100",
  27980=>"000100110",
  27981=>"000000100",
  27982=>"000000000",
  27983=>"000001001",
  27984=>"001011011",
  27985=>"111100100",
  27986=>"111001000",
  27987=>"111111111",
  27988=>"000000101",
  27989=>"011011011",
  27990=>"000110111",
  27991=>"000000000",
  27992=>"000000111",
  27993=>"000000000",
  27994=>"000011000",
  27995=>"110110111",
  27996=>"000100000",
  27997=>"111111111",
  27998=>"111000001",
  27999=>"101000100",
  28000=>"110110111",
  28001=>"111111110",
  28002=>"011011011",
  28003=>"101000001",
  28004=>"000000001",
  28005=>"000000000",
  28006=>"101001000",
  28007=>"000001111",
  28008=>"000000000",
  28009=>"000000000",
  28010=>"011111111",
  28011=>"010010011",
  28012=>"110110100",
  28013=>"000000100",
  28014=>"100000100",
  28015=>"011011011",
  28016=>"011001001",
  28017=>"010111111",
  28018=>"111111111",
  28019=>"000000100",
  28020=>"000011001",
  28021=>"000110111",
  28022=>"011110111",
  28023=>"000001000",
  28024=>"000000000",
  28025=>"111110000",
  28026=>"111001111",
  28027=>"000110000",
  28028=>"111010000",
  28029=>"111111110",
  28030=>"000111111",
  28031=>"111001111",
  28032=>"001000000",
  28033=>"100111001",
  28034=>"111001111",
  28035=>"000100001",
  28036=>"000000100",
  28037=>"111111011",
  28038=>"111111111",
  28039=>"001000000",
  28040=>"000000000",
  28041=>"010111111",
  28042=>"000000001",
  28043=>"110111111",
  28044=>"000000000",
  28045=>"011001001",
  28046=>"001100000",
  28047=>"000000000",
  28048=>"110110000",
  28049=>"111111111",
  28050=>"101110111",
  28051=>"011111010",
  28052=>"111000001",
  28053=>"000000000",
  28054=>"000000000",
  28055=>"111111000",
  28056=>"000111100",
  28057=>"000000000",
  28058=>"111111111",
  28059=>"111111111",
  28060=>"000100101",
  28061=>"000000000",
  28062=>"111110100",
  28063=>"000000000",
  28064=>"000001111",
  28065=>"001001000",
  28066=>"111001001",
  28067=>"111000000",
  28068=>"001000100",
  28069=>"111111001",
  28070=>"001111111",
  28071=>"001100111",
  28072=>"000000000",
  28073=>"000000101",
  28074=>"111110111",
  28075=>"111100100",
  28076=>"000000000",
  28077=>"110110110",
  28078=>"000000111",
  28079=>"100000101",
  28080=>"000000000",
  28081=>"000000000",
  28082=>"000000000",
  28083=>"111000110",
  28084=>"100000000",
  28085=>"111000000",
  28086=>"110111111",
  28087=>"001000000",
  28088=>"001001000",
  28089=>"101000100",
  28090=>"010010101",
  28091=>"111111100",
  28092=>"011101100",
  28093=>"101111111",
  28094=>"000000000",
  28095=>"110100000",
  28096=>"101111111",
  28097=>"000000000",
  28098=>"111111111",
  28099=>"000000000",
  28100=>"111001111",
  28101=>"000000100",
  28102=>"101101111",
  28103=>"001000000",
  28104=>"011001101",
  28105=>"100000000",
  28106=>"001000000",
  28107=>"111111111",
  28108=>"111111111",
  28109=>"110111010",
  28110=>"000000010",
  28111=>"001001000",
  28112=>"000000110",
  28113=>"000000100",
  28114=>"001011000",
  28115=>"000000000",
  28116=>"111111000",
  28117=>"111110100",
  28118=>"000100111",
  28119=>"100110110",
  28120=>"111111111",
  28121=>"111111101",
  28122=>"000000010",
  28123=>"010000110",
  28124=>"111000000",
  28125=>"000000101",
  28126=>"100000101",
  28127=>"110110000",
  28128=>"001000000",
  28129=>"101000000",
  28130=>"011000000",
  28131=>"010010011",
  28132=>"000000000",
  28133=>"000101101",
  28134=>"000001111",
  28135=>"000000000",
  28136=>"111110110",
  28137=>"000000111",
  28138=>"000000000",
  28139=>"111001001",
  28140=>"111111111",
  28141=>"111111011",
  28142=>"000011000",
  28143=>"110111111",
  28144=>"111111111",
  28145=>"000001001",
  28146=>"011111111",
  28147=>"001000000",
  28148=>"111100110",
  28149=>"100110110",
  28150=>"001000000",
  28151=>"011110111",
  28152=>"000000000",
  28153=>"001000000",
  28154=>"001000000",
  28155=>"000000010",
  28156=>"000100000",
  28157=>"111111111",
  28158=>"000000000",
  28159=>"101001111",
  28160=>"101111111",
  28161=>"110111111",
  28162=>"100100111",
  28163=>"000000000",
  28164=>"100001000",
  28165=>"000001111",
  28166=>"000000000",
  28167=>"101000000",
  28168=>"000000000",
  28169=>"000000000",
  28170=>"000100111",
  28171=>"111111111",
  28172=>"111110000",
  28173=>"111011000",
  28174=>"000000111",
  28175=>"001001111",
  28176=>"001000000",
  28177=>"010000011",
  28178=>"111111111",
  28179=>"011000000",
  28180=>"000000111",
  28181=>"111111111",
  28182=>"000100110",
  28183=>"010000110",
  28184=>"000011011",
  28185=>"111111111",
  28186=>"110111111",
  28187=>"111001100",
  28188=>"000000000",
  28189=>"110000000",
  28190=>"110000111",
  28191=>"000000111",
  28192=>"110111111",
  28193=>"111110000",
  28194=>"001001111",
  28195=>"000101100",
  28196=>"001111111",
  28197=>"111111011",
  28198=>"000000101",
  28199=>"000000111",
  28200=>"110000000",
  28201=>"111000000",
  28202=>"111111111",
  28203=>"000001111",
  28204=>"000101100",
  28205=>"110111111",
  28206=>"000010000",
  28207=>"000111111",
  28208=>"001101101",
  28209=>"111000000",
  28210=>"011000000",
  28211=>"000000000",
  28212=>"011000011",
  28213=>"110100000",
  28214=>"000111101",
  28215=>"000100001",
  28216=>"001111000",
  28217=>"110111111",
  28218=>"000000000",
  28219=>"111111000",
  28220=>"111110000",
  28221=>"000000000",
  28222=>"101001001",
  28223=>"000000101",
  28224=>"111110100",
  28225=>"111000000",
  28226=>"101101000",
  28227=>"000001001",
  28228=>"011111111",
  28229=>"011001000",
  28230=>"101000010",
  28231=>"111111111",
  28232=>"111100100",
  28233=>"000000000",
  28234=>"111111111",
  28235=>"110000001",
  28236=>"000000000",
  28237=>"100100000",
  28238=>"010000000",
  28239=>"111011111",
  28240=>"000001000",
  28241=>"111111011",
  28242=>"111011010",
  28243=>"000000001",
  28244=>"000000000",
  28245=>"111000000",
  28246=>"110111011",
  28247=>"000000000",
  28248=>"011111111",
  28249=>"000000000",
  28250=>"001111111",
  28251=>"111110100",
  28252=>"000000011",
  28253=>"111100100",
  28254=>"111001000",
  28255=>"001000000",
  28256=>"000000000",
  28257=>"000000010",
  28258=>"000110111",
  28259=>"000000110",
  28260=>"001000000",
  28261=>"000000000",
  28262=>"111111000",
  28263=>"110000100",
  28264=>"111111111",
  28265=>"100100111",
  28266=>"111111011",
  28267=>"111100000",
  28268=>"000000000",
  28269=>"001101111",
  28270=>"111000000",
  28271=>"100000000",
  28272=>"110111111",
  28273=>"111110000",
  28274=>"010111011",
  28275=>"100100000",
  28276=>"000000000",
  28277=>"001101111",
  28278=>"111111001",
  28279=>"111000000",
  28280=>"111110000",
  28281=>"111111000",
  28282=>"100001101",
  28283=>"111111000",
  28284=>"100000100",
  28285=>"000111111",
  28286=>"100100100",
  28287=>"111111111",
  28288=>"000000000",
  28289=>"000000000",
  28290=>"111011101",
  28291=>"000000111",
  28292=>"111111110",
  28293=>"111100000",
  28294=>"000001111",
  28295=>"111000000",
  28296=>"000000000",
  28297=>"000001111",
  28298=>"000000000",
  28299=>"001000000",
  28300=>"000000000",
  28301=>"111111101",
  28302=>"111111000",
  28303=>"011000000",
  28304=>"000111001",
  28305=>"000111111",
  28306=>"000000111",
  28307=>"000000000",
  28308=>"111000000",
  28309=>"111111111",
  28310=>"100000000",
  28311=>"000100111",
  28312=>"000001001",
  28313=>"000110100",
  28314=>"111111111",
  28315=>"111000000",
  28316=>"000101111",
  28317=>"000000111",
  28318=>"111000000",
  28319=>"111000000",
  28320=>"110000000",
  28321=>"001000000",
  28322=>"000000101",
  28323=>"111011101",
  28324=>"100100100",
  28325=>"000000111",
  28326=>"111111111",
  28327=>"111101001",
  28328=>"110111000",
  28329=>"000000111",
  28330=>"000111100",
  28331=>"110101000",
  28332=>"111101000",
  28333=>"110100101",
  28334=>"100111111",
  28335=>"000000111",
  28336=>"000000000",
  28337=>"110111111",
  28338=>"111110111",
  28339=>"011000111",
  28340=>"000000000",
  28341=>"101111111",
  28342=>"000000000",
  28343=>"000001001",
  28344=>"111100000",
  28345=>"000000000",
  28346=>"110111001",
  28347=>"111111111",
  28348=>"111111000",
  28349=>"000000011",
  28350=>"111110111",
  28351=>"111111000",
  28352=>"000001000",
  28353=>"000111010",
  28354=>"101001001",
  28355=>"011111010",
  28356=>"000000000",
  28357=>"000000111",
  28358=>"111111000",
  28359=>"100000000",
  28360=>"000000000",
  28361=>"111111111",
  28362=>"111111110",
  28363=>"111111011",
  28364=>"111110011",
  28365=>"110000000",
  28366=>"111001111",
  28367=>"000000000",
  28368=>"100111111",
  28369=>"100100111",
  28370=>"100000000",
  28371=>"000000000",
  28372=>"000000000",
  28373=>"101001000",
  28374=>"111110000",
  28375=>"111000000",
  28376=>"000000000",
  28377=>"000001001",
  28378=>"000000000",
  28379=>"000000000",
  28380=>"000001000",
  28381=>"111111111",
  28382=>"011111111",
  28383=>"101100000",
  28384=>"001000111",
  28385=>"001011110",
  28386=>"111111000",
  28387=>"111111101",
  28388=>"000000000",
  28389=>"010011111",
  28390=>"111111010",
  28391=>"110110011",
  28392=>"000111111",
  28393=>"111110111",
  28394=>"111111101",
  28395=>"101001111",
  28396=>"000000001",
  28397=>"000000000",
  28398=>"111111111",
  28399=>"010000000",
  28400=>"000000000",
  28401=>"000000000",
  28402=>"101100110",
  28403=>"010000000",
  28404=>"111001001",
  28405=>"111000000",
  28406=>"110111100",
  28407=>"100100000",
  28408=>"000101111",
  28409=>"010110000",
  28410=>"001001001",
  28411=>"000001000",
  28412=>"100100100",
  28413=>"111101111",
  28414=>"111111000",
  28415=>"101100100",
  28416=>"101001001",
  28417=>"111100000",
  28418=>"111001101",
  28419=>"000111111",
  28420=>"111111000",
  28421=>"001000000",
  28422=>"110111111",
  28423=>"000000111",
  28424=>"100000001",
  28425=>"111011000",
  28426=>"111111111",
  28427=>"000000001",
  28428=>"111111111",
  28429=>"111000000",
  28430=>"110111111",
  28431=>"000000000",
  28432=>"000000000",
  28433=>"000000001",
  28434=>"000000000",
  28435=>"100100100",
  28436=>"010000000",
  28437=>"001111111",
  28438=>"111110000",
  28439=>"101111111",
  28440=>"001011011",
  28441=>"101001101",
  28442=>"000000111",
  28443=>"101111111",
  28444=>"000101111",
  28445=>"001000000",
  28446=>"100111110",
  28447=>"000011111",
  28448=>"000000001",
  28449=>"000000001",
  28450=>"000001000",
  28451=>"110111111",
  28452=>"001001000",
  28453=>"011011111",
  28454=>"001001000",
  28455=>"010111011",
  28456=>"000000000",
  28457=>"111111111",
  28458=>"100111101",
  28459=>"000101111",
  28460=>"011001000",
  28461=>"100111000",
  28462=>"000000000",
  28463=>"000000111",
  28464=>"001001101",
  28465=>"000000000",
  28466=>"110000000",
  28467=>"111000110",
  28468=>"110101000",
  28469=>"111000001",
  28470=>"111000000",
  28471=>"000000000",
  28472=>"000000000",
  28473=>"111001000",
  28474=>"000101000",
  28475=>"111100111",
  28476=>"111101000",
  28477=>"001001000",
  28478=>"000000000",
  28479=>"000010000",
  28480=>"000111111",
  28481=>"101001100",
  28482=>"111001101",
  28483=>"111111000",
  28484=>"000000101",
  28485=>"111100000",
  28486=>"110111110",
  28487=>"000011111",
  28488=>"111000111",
  28489=>"000000000",
  28490=>"000111000",
  28491=>"000011111",
  28492=>"000000111",
  28493=>"000111111",
  28494=>"000000000",
  28495=>"011011001",
  28496=>"000101111",
  28497=>"100100101",
  28498=>"100111111",
  28499=>"000111101",
  28500=>"110110100",
  28501=>"011011011",
  28502=>"110000000",
  28503=>"000000000",
  28504=>"111111111",
  28505=>"111100111",
  28506=>"001001000",
  28507=>"000101101",
  28508=>"111111111",
  28509=>"111111111",
  28510=>"111111111",
  28511=>"000000100",
  28512=>"000111111",
  28513=>"000010011",
  28514=>"110000011",
  28515=>"111111111",
  28516=>"111111011",
  28517=>"000100000",
  28518=>"000000111",
  28519=>"100101111",
  28520=>"100100111",
  28521=>"000000111",
  28522=>"000000000",
  28523=>"000100101",
  28524=>"000011011",
  28525=>"111100000",
  28526=>"000000111",
  28527=>"000000000",
  28528=>"101101001",
  28529=>"111100100",
  28530=>"111010010",
  28531=>"001111110",
  28532=>"011001101",
  28533=>"100111111",
  28534=>"000000011",
  28535=>"001111111",
  28536=>"111000000",
  28537=>"111000001",
  28538=>"000000000",
  28539=>"000111000",
  28540=>"000000000",
  28541=>"111001000",
  28542=>"000100111",
  28543=>"111111111",
  28544=>"100101001",
  28545=>"000101100",
  28546=>"111100000",
  28547=>"000000000",
  28548=>"000000011",
  28549=>"111111111",
  28550=>"111000000",
  28551=>"000000000",
  28552=>"000000000",
  28553=>"010111111",
  28554=>"111011111",
  28555=>"110000000",
  28556=>"001000111",
  28557=>"000000111",
  28558=>"100111111",
  28559=>"000000110",
  28560=>"111000000",
  28561=>"100110111",
  28562=>"111000000",
  28563=>"111111101",
  28564=>"000000000",
  28565=>"000010000",
  28566=>"110110100",
  28567=>"100100100",
  28568=>"000011111",
  28569=>"000000101",
  28570=>"000000101",
  28571=>"000111111",
  28572=>"000000000",
  28573=>"111111111",
  28574=>"000000000",
  28575=>"001000000",
  28576=>"100111101",
  28577=>"101111111",
  28578=>"000000000",
  28579=>"000000111",
  28580=>"100110000",
  28581=>"000000000",
  28582=>"111110110",
  28583=>"000000111",
  28584=>"000000001",
  28585=>"100100110",
  28586=>"000000011",
  28587=>"000111010",
  28588=>"000000011",
  28589=>"111111001",
  28590=>"111100000",
  28591=>"111111111",
  28592=>"000111111",
  28593=>"111000000",
  28594=>"111110110",
  28595=>"010000000",
  28596=>"111111010",
  28597=>"100001000",
  28598=>"111101101",
  28599=>"000000000",
  28600=>"001000000",
  28601=>"111111111",
  28602=>"101001001",
  28603=>"001011001",
  28604=>"111101000",
  28605=>"000100110",
  28606=>"000111111",
  28607=>"110100111",
  28608=>"000000100",
  28609=>"110110010",
  28610=>"000000010",
  28611=>"000000000",
  28612=>"111111000",
  28613=>"110000000",
  28614=>"111111100",
  28615=>"000111111",
  28616=>"111001001",
  28617=>"000100111",
  28618=>"110000001",
  28619=>"000001000",
  28620=>"011000000",
  28621=>"000000111",
  28622=>"000100110",
  28623=>"001000000",
  28624=>"000000000",
  28625=>"111111111",
  28626=>"111111111",
  28627=>"111111111",
  28628=>"100100111",
  28629=>"111111000",
  28630=>"111001111",
  28631=>"110010011",
  28632=>"110000000",
  28633=>"110010110",
  28634=>"000000110",
  28635=>"000100111",
  28636=>"110110111",
  28637=>"011111111",
  28638=>"110000000",
  28639=>"100100000",
  28640=>"000000111",
  28641=>"000011111",
  28642=>"000000000",
  28643=>"011000000",
  28644=>"000000100",
  28645=>"101001000",
  28646=>"111011111",
  28647=>"000000001",
  28648=>"000001001",
  28649=>"111101111",
  28650=>"000111111",
  28651=>"000111111",
  28652=>"000000100",
  28653=>"001001101",
  28654=>"000111111",
  28655=>"111001000",
  28656=>"001111000",
  28657=>"000100011",
  28658=>"110000000",
  28659=>"000110110",
  28660=>"111101000",
  28661=>"001111111",
  28662=>"000000111",
  28663=>"101001011",
  28664=>"011111000",
  28665=>"111000110",
  28666=>"000000001",
  28667=>"111111011",
  28668=>"111111001",
  28669=>"111111001",
  28670=>"110000000",
  28671=>"111001000",
  28672=>"111111111",
  28673=>"111100110",
  28674=>"001101111",
  28675=>"111000000",
  28676=>"000000001",
  28677=>"111111111",
  28678=>"010010000",
  28679=>"111111111",
  28680=>"111111111",
  28681=>"111111111",
  28682=>"111000000",
  28683=>"000000000",
  28684=>"100111110",
  28685=>"000000110",
  28686=>"111111000",
  28687=>"000000001",
  28688=>"000000000",
  28689=>"000111111",
  28690=>"011011011",
  28691=>"000000000",
  28692=>"000000000",
  28693=>"110000100",
  28694=>"111111110",
  28695=>"111111000",
  28696=>"000000000",
  28697=>"010110100",
  28698=>"000100100",
  28699=>"100101111",
  28700=>"000100000",
  28701=>"000000001",
  28702=>"110110110",
  28703=>"010000011",
  28704=>"110110000",
  28705=>"010010110",
  28706=>"111111111",
  28707=>"111101111",
  28708=>"000000000",
  28709=>"000000000",
  28710=>"000110111",
  28711=>"000000111",
  28712=>"000000000",
  28713=>"000000000",
  28714=>"010110110",
  28715=>"111111111",
  28716=>"110000001",
  28717=>"111111111",
  28718=>"111101100",
  28719=>"000000000",
  28720=>"111011001",
  28721=>"000000000",
  28722=>"000111110",
  28723=>"000010010",
  28724=>"000000001",
  28725=>"000000000",
  28726=>"111011000",
  28727=>"001000000",
  28728=>"000000000",
  28729=>"111110111",
  28730=>"111111111",
  28731=>"111101111",
  28732=>"000000000",
  28733=>"000000000",
  28734=>"000000100",
  28735=>"111100100",
  28736=>"000110111",
  28737=>"000001000",
  28738=>"000100000",
  28739=>"000011000",
  28740=>"000000100",
  28741=>"100000000",
  28742=>"111111110",
  28743=>"111111010",
  28744=>"001011111",
  28745=>"000110111",
  28746=>"000000000",
  28747=>"001111110",
  28748=>"000000001",
  28749=>"000000101",
  28750=>"100000000",
  28751=>"000110100",
  28752=>"111111111",
  28753=>"101001000",
  28754=>"000000000",
  28755=>"111111111",
  28756=>"111110110",
  28757=>"000000111",
  28758=>"111100101",
  28759=>"110100111",
  28760=>"110000000",
  28761=>"111101111",
  28762=>"111111111",
  28763=>"110100000",
  28764=>"000101111",
  28765=>"000000001",
  28766=>"000000000",
  28767=>"000000000",
  28768=>"000111111",
  28769=>"111111111",
  28770=>"000000000",
  28771=>"111111111",
  28772=>"110000000",
  28773=>"110111111",
  28774=>"001001011",
  28775=>"001010011",
  28776=>"001000000",
  28777=>"111101001",
  28778=>"111111111",
  28779=>"101000000",
  28780=>"111111111",
  28781=>"000000000",
  28782=>"111111001",
  28783=>"000000000",
  28784=>"000000000",
  28785=>"000000000",
  28786=>"101101000",
  28787=>"111111001",
  28788=>"111111110",
  28789=>"110100100",
  28790=>"000000000",
  28791=>"000110000",
  28792=>"010110100",
  28793=>"000000001",
  28794=>"101100000",
  28795=>"000000000",
  28796=>"000000000",
  28797=>"000000000",
  28798=>"110110010",
  28799=>"000111111",
  28800=>"111011010",
  28801=>"000000000",
  28802=>"101101111",
  28803=>"111111111",
  28804=>"011111010",
  28805=>"000000000",
  28806=>"110000101",
  28807=>"000000110",
  28808=>"111111111",
  28809=>"000000000",
  28810=>"000000000",
  28811=>"110111010",
  28812=>"111111111",
  28813=>"111111111",
  28814=>"101110010",
  28815=>"000000000",
  28816=>"111000100",
  28817=>"111111111",
  28818=>"000000100",
  28819=>"011000000",
  28820=>"000000000",
  28821=>"000000000",
  28822=>"011011111",
  28823=>"111000000",
  28824=>"001000000",
  28825=>"111111000",
  28826=>"111111111",
  28827=>"000000101",
  28828=>"111111111",
  28829=>"110000000",
  28830=>"111101000",
  28831=>"001011011",
  28832=>"111111111",
  28833=>"111100000",
  28834=>"111000000",
  28835=>"001011111",
  28836=>"111111011",
  28837=>"000000010",
  28838=>"111101111",
  28839=>"110110000",
  28840=>"011110111",
  28841=>"000000000",
  28842=>"111001111",
  28843=>"000000000",
  28844=>"000000110",
  28845=>"101001111",
  28846=>"111101111",
  28847=>"100111111",
  28848=>"000000000",
  28849=>"000001000",
  28850=>"110111110",
  28851=>"111100111",
  28852=>"000000000",
  28853=>"000000000",
  28854=>"010110111",
  28855=>"111111111",
  28856=>"111110110",
  28857=>"111111111",
  28858=>"000000000",
  28859=>"111110111",
  28860=>"111111111",
  28861=>"111111010",
  28862=>"000101000",
  28863=>"100110011",
  28864=>"111100111",
  28865=>"100100100",
  28866=>"000000000",
  28867=>"000000000",
  28868=>"000111111",
  28869=>"011001110",
  28870=>"000000000",
  28871=>"110110111",
  28872=>"001000010",
  28873=>"000000100",
  28874=>"000101111",
  28875=>"000000001",
  28876=>"011011011",
  28877=>"001111001",
  28878=>"000000000",
  28879=>"010000010",
  28880=>"111111111",
  28881=>"001101111",
  28882=>"000100110",
  28883=>"000000110",
  28884=>"001000000",
  28885=>"001001000",
  28886=>"101000100",
  28887=>"000000110",
  28888=>"110111111",
  28889=>"000000000",
  28890=>"111111111",
  28891=>"010010111",
  28892=>"011011111",
  28893=>"110110100",
  28894=>"111110000",
  28895=>"111110111",
  28896=>"111001001",
  28897=>"000001011",
  28898=>"110000101",
  28899=>"000000000",
  28900=>"111011000",
  28901=>"110010000",
  28902=>"000000000",
  28903=>"110000000",
  28904=>"000001001",
  28905=>"111010001",
  28906=>"000000000",
  28907=>"010000010",
  28908=>"011001000",
  28909=>"111111111",
  28910=>"000111111",
  28911=>"111100100",
  28912=>"001011011",
  28913=>"101100000",
  28914=>"100000010",
  28915=>"110100000",
  28916=>"000000000",
  28917=>"100000000",
  28918=>"000000100",
  28919=>"111000000",
  28920=>"000000000",
  28921=>"111111111",
  28922=>"001000001",
  28923=>"111111111",
  28924=>"111111111",
  28925=>"111000000",
  28926=>"000000000",
  28927=>"000010000",
  28928=>"000000000",
  28929=>"000000000",
  28930=>"000000000",
  28931=>"111111111",
  28932=>"110110111",
  28933=>"000000000",
  28934=>"111111111",
  28935=>"011111111",
  28936=>"111111111",
  28937=>"000000000",
  28938=>"000000000",
  28939=>"111111111",
  28940=>"100000000",
  28941=>"111101111",
  28942=>"110111111",
  28943=>"111111000",
  28944=>"111111111",
  28945=>"001100100",
  28946=>"000000100",
  28947=>"000000000",
  28948=>"011111010",
  28949=>"000111011",
  28950=>"111111111",
  28951=>"111111111",
  28952=>"111111111",
  28953=>"011011000",
  28954=>"100110111",
  28955=>"000000000",
  28956=>"111111110",
  28957=>"110111111",
  28958=>"000010111",
  28959=>"011100000",
  28960=>"010100000",
  28961=>"000000000",
  28962=>"111111111",
  28963=>"111000000",
  28964=>"000000000",
  28965=>"111100000",
  28966=>"111111111",
  28967=>"111111000",
  28968=>"000000000",
  28969=>"000000000",
  28970=>"101100100",
  28971=>"000001000",
  28972=>"111101000",
  28973=>"001001001",
  28974=>"000000011",
  28975=>"000000001",
  28976=>"110100000",
  28977=>"000010000",
  28978=>"000000001",
  28979=>"000000010",
  28980=>"001101111",
  28981=>"111111111",
  28982=>"000000000",
  28983=>"111000100",
  28984=>"000111000",
  28985=>"111001000",
  28986=>"111000100",
  28987=>"111111111",
  28988=>"100110000",
  28989=>"100000100",
  28990=>"110010000",
  28991=>"111010000",
  28992=>"110111111",
  28993=>"111111111",
  28994=>"000000000",
  28995=>"000000000",
  28996=>"000000111",
  28997=>"111111011",
  28998=>"000010000",
  28999=>"111111010",
  29000=>"000000010",
  29001=>"011111111",
  29002=>"111111101",
  29003=>"100100110",
  29004=>"000000010",
  29005=>"000000011",
  29006=>"111000000",
  29007=>"111011011",
  29008=>"100110100",
  29009=>"010000000",
  29010=>"111111011",
  29011=>"000000000",
  29012=>"011111000",
  29013=>"011001011",
  29014=>"010000000",
  29015=>"100101111",
  29016=>"110101000",
  29017=>"101001111",
  29018=>"100100000",
  29019=>"000000111",
  29020=>"000000100",
  29021=>"000111111",
  29022=>"000000000",
  29023=>"110000000",
  29024=>"111111111",
  29025=>"111101111",
  29026=>"111111111",
  29027=>"100101000",
  29028=>"111011110",
  29029=>"000000000",
  29030=>"111011111",
  29031=>"111110110",
  29032=>"101101111",
  29033=>"000000000",
  29034=>"110110110",
  29035=>"000000000",
  29036=>"111111101",
  29037=>"111101001",
  29038=>"011001111",
  29039=>"000000000",
  29040=>"111111011",
  29041=>"000000000",
  29042=>"100110000",
  29043=>"000001001",
  29044=>"000000000",
  29045=>"111111111",
  29046=>"000000000",
  29047=>"010011000",
  29048=>"000000000",
  29049=>"000000111",
  29050=>"111110110",
  29051=>"111111110",
  29052=>"000000000",
  29053=>"000100111",
  29054=>"000000000",
  29055=>"111101111",
  29056=>"101111111",
  29057=>"111111111",
  29058=>"101001111",
  29059=>"010111111",
  29060=>"000000000",
  29061=>"111111111",
  29062=>"111000010",
  29063=>"000000000",
  29064=>"010000001",
  29065=>"000000000",
  29066=>"111111111",
  29067=>"111111011",
  29068=>"000000101",
  29069=>"110100000",
  29070=>"111111111",
  29071=>"000000010",
  29072=>"111111111",
  29073=>"110000000",
  29074=>"111111101",
  29075=>"011101000",
  29076=>"111111111",
  29077=>"000000000",
  29078=>"111111111",
  29079=>"010001000",
  29080=>"000000100",
  29081=>"111110110",
  29082=>"011010000",
  29083=>"111111111",
  29084=>"111010000",
  29085=>"000000000",
  29086=>"001000000",
  29087=>"111111111",
  29088=>"000000101",
  29089=>"111111100",
  29090=>"010000000",
  29091=>"010001000",
  29092=>"001000000",
  29093=>"111000000",
  29094=>"111111111",
  29095=>"111111011",
  29096=>"111111111",
  29097=>"000110111",
  29098=>"010011010",
  29099=>"000000000",
  29100=>"000000111",
  29101=>"110010000",
  29102=>"100100111",
  29103=>"111111111",
  29104=>"000000011",
  29105=>"110111010",
  29106=>"000111111",
  29107=>"000000000",
  29108=>"100100000",
  29109=>"000000010",
  29110=>"110110000",
  29111=>"010111010",
  29112=>"110111110",
  29113=>"111110111",
  29114=>"100000000",
  29115=>"011011001",
  29116=>"000000000",
  29117=>"110010110",
  29118=>"100100101",
  29119=>"100100100",
  29120=>"001101000",
  29121=>"000000000",
  29122=>"111111111",
  29123=>"100100100",
  29124=>"001000000",
  29125=>"000000010",
  29126=>"000000110",
  29127=>"001001101",
  29128=>"000000000",
  29129=>"000000000",
  29130=>"111110000",
  29131=>"000000000",
  29132=>"100111000",
  29133=>"000000010",
  29134=>"000000110",
  29135=>"000000100",
  29136=>"000000000",
  29137=>"000001001",
  29138=>"011000000",
  29139=>"000000000",
  29140=>"011001111",
  29141=>"100110011",
  29142=>"000000000",
  29143=>"111111111",
  29144=>"000000111",
  29145=>"111111011",
  29146=>"000100100",
  29147=>"000000000",
  29148=>"011111111",
  29149=>"111111101",
  29150=>"100000001",
  29151=>"001000001",
  29152=>"010000000",
  29153=>"000000000",
  29154=>"001101000",
  29155=>"111111011",
  29156=>"011010110",
  29157=>"111000010",
  29158=>"001101000",
  29159=>"010000000",
  29160=>"111111110",
  29161=>"111110010",
  29162=>"010010010",
  29163=>"111111011",
  29164=>"111111111",
  29165=>"111010011",
  29166=>"001000000",
  29167=>"000000110",
  29168=>"100000000",
  29169=>"111111111",
  29170=>"000000000",
  29171=>"000000111",
  29172=>"000000000",
  29173=>"111111010",
  29174=>"000000000",
  29175=>"000000111",
  29176=>"000000000",
  29177=>"000010010",
  29178=>"000100000",
  29179=>"000100000",
  29180=>"110010000",
  29181=>"110110110",
  29182=>"110111111",
  29183=>"111111110",
  29184=>"111111000",
  29185=>"000000111",
  29186=>"111000000",
  29187=>"010000000",
  29188=>"111100000",
  29189=>"111111110",
  29190=>"110110111",
  29191=>"000111111",
  29192=>"000001000",
  29193=>"100100100",
  29194=>"000000000",
  29195=>"010011111",
  29196=>"000100110",
  29197=>"000001111",
  29198=>"001001011",
  29199=>"011010000",
  29200=>"101000110",
  29201=>"111111101",
  29202=>"111110111",
  29203=>"000100000",
  29204=>"001000000",
  29205=>"000000000",
  29206=>"011001000",
  29207=>"011000011",
  29208=>"011111110",
  29209=>"101100111",
  29210=>"111111111",
  29211=>"000001001",
  29212=>"001111111",
  29213=>"001000111",
  29214=>"111001011",
  29215=>"111000000",
  29216=>"000111111",
  29217=>"111111111",
  29218=>"001001111",
  29219=>"101001111",
  29220=>"100100110",
  29221=>"000100111",
  29222=>"110110111",
  29223=>"011111101",
  29224=>"000011111",
  29225=>"111111111",
  29226=>"110111111",
  29227=>"000000000",
  29228=>"000000000",
  29229=>"111111100",
  29230=>"111101101",
  29231=>"001000111",
  29232=>"000000000",
  29233=>"111111111",
  29234=>"011011011",
  29235=>"101111111",
  29236=>"111110000",
  29237=>"111011011",
  29238=>"000011011",
  29239=>"110000001",
  29240=>"000000101",
  29241=>"010000000",
  29242=>"100000000",
  29243=>"000111111",
  29244=>"000000111",
  29245=>"010010000",
  29246=>"011001000",
  29247=>"110010010",
  29248=>"000100111",
  29249=>"000000000",
  29250=>"111000000",
  29251=>"011100111",
  29252=>"101100000",
  29253=>"111111101",
  29254=>"110111000",
  29255=>"111111111",
  29256=>"000001010",
  29257=>"000000000",
  29258=>"000000000",
  29259=>"100001001",
  29260=>"000100000",
  29261=>"000111101",
  29262=>"000010000",
  29263=>"111111111",
  29264=>"000011011",
  29265=>"011011111",
  29266=>"010111111",
  29267=>"110011001",
  29268=>"000000000",
  29269=>"111111100",
  29270=>"111111111",
  29271=>"000000000",
  29272=>"000000000",
  29273=>"100111111",
  29274=>"000111111",
  29275=>"001011110",
  29276=>"111111111",
  29277=>"000100111",
  29278=>"100100000",
  29279=>"111110110",
  29280=>"010000000",
  29281=>"001000001",
  29282=>"111111000",
  29283=>"111111111",
  29284=>"111000001",
  29285=>"000001111",
  29286=>"000000000",
  29287=>"100100100",
  29288=>"111111111",
  29289=>"110011001",
  29290=>"110110011",
  29291=>"001001101",
  29292=>"111100000",
  29293=>"111111111",
  29294=>"111111111",
  29295=>"111000000",
  29296=>"000100100",
  29297=>"001000001",
  29298=>"000000000",
  29299=>"111101101",
  29300=>"000000010",
  29301=>"111111011",
  29302=>"101000000",
  29303=>"101001001",
  29304=>"000000000",
  29305=>"111110110",
  29306=>"111111111",
  29307=>"000000100",
  29308=>"011001011",
  29309=>"100100100",
  29310=>"110111111",
  29311=>"000100111",
  29312=>"110000000",
  29313=>"001001000",
  29314=>"111000000",
  29315=>"111110110",
  29316=>"010000000",
  29317=>"111101111",
  29318=>"000000011",
  29319=>"011001001",
  29320=>"000010110",
  29321=>"101100001",
  29322=>"000001111",
  29323=>"111111111",
  29324=>"111000000",
  29325=>"000000111",
  29326=>"001000000",
  29327=>"111101111",
  29328=>"111111111",
  29329=>"000000000",
  29330=>"111111111",
  29331=>"111111111",
  29332=>"111101001",
  29333=>"111111010",
  29334=>"000000000",
  29335=>"000101000",
  29336=>"000000111",
  29337=>"111111111",
  29338=>"011011011",
  29339=>"111000000",
  29340=>"011011000",
  29341=>"000000111",
  29342=>"110110111",
  29343=>"111111110",
  29344=>"111111111",
  29345=>"110100100",
  29346=>"000000101",
  29347=>"001011011",
  29348=>"001001011",
  29349=>"111111111",
  29350=>"110100111",
  29351=>"011000000",
  29352=>"000000000",
  29353=>"000000100",
  29354=>"000000000",
  29355=>"010100111",
  29356=>"001000100",
  29357=>"000101001",
  29358=>"000000000",
  29359=>"011001111",
  29360=>"000000000",
  29361=>"011111111",
  29362=>"111111111",
  29363=>"101000000",
  29364=>"000110111",
  29365=>"000000000",
  29366=>"111111111",
  29367=>"111111111",
  29368=>"111111100",
  29369=>"111111111",
  29370=>"000001000",
  29371=>"111111111",
  29372=>"110110000",
  29373=>"000111001",
  29374=>"111111111",
  29375=>"000111111",
  29376=>"111111000",
  29377=>"000000000",
  29378=>"111110110",
  29379=>"000101000",
  29380=>"000000000",
  29381=>"000000000",
  29382=>"011001000",
  29383=>"111111000",
  29384=>"000011111",
  29385=>"000000000",
  29386=>"000000000",
  29387=>"111111111",
  29388=>"000000000",
  29389=>"111111001",
  29390=>"111111111",
  29391=>"111000000",
  29392=>"100100000",
  29393=>"000000000",
  29394=>"100000000",
  29395=>"111111000",
  29396=>"111111111",
  29397=>"001101111",
  29398=>"000001000",
  29399=>"110110000",
  29400=>"111100000",
  29401=>"101111111",
  29402=>"000000000",
  29403=>"010111111",
  29404=>"111110110",
  29405=>"000001111",
  29406=>"111101111",
  29407=>"000000000",
  29408=>"111111000",
  29409=>"011000000",
  29410=>"000000000",
  29411=>"000000000",
  29412=>"111001111",
  29413=>"011000001",
  29414=>"001111111",
  29415=>"000000110",
  29416=>"000000111",
  29417=>"000111111",
  29418=>"111011111",
  29419=>"001111111",
  29420=>"111111011",
  29421=>"000000000",
  29422=>"111001000",
  29423=>"100111111",
  29424=>"111011011",
  29425=>"000000111",
  29426=>"100100100",
  29427=>"001011011",
  29428=>"111111001",
  29429=>"111001000",
  29430=>"011100111",
  29431=>"001000000",
  29432=>"111111011",
  29433=>"000000000",
  29434=>"000000001",
  29435=>"100100100",
  29436=>"000000110",
  29437=>"100001000",
  29438=>"011000000",
  29439=>"100100101",
  29440=>"111101111",
  29441=>"010010000",
  29442=>"000000000",
  29443=>"101100100",
  29444=>"000000000",
  29445=>"001000000",
  29446=>"111111111",
  29447=>"111111111",
  29448=>"000110000",
  29449=>"101111111",
  29450=>"000000000",
  29451=>"001000100",
  29452=>"111111111",
  29453=>"111111111",
  29454=>"001001111",
  29455=>"000000111",
  29456=>"000000010",
  29457=>"110000010",
  29458=>"000000000",
  29459=>"000001111",
  29460=>"000000000",
  29461=>"111100100",
  29462=>"111011011",
  29463=>"011111111",
  29464=>"111111111",
  29465=>"111111111",
  29466=>"000000000",
  29467=>"111010000",
  29468=>"100100000",
  29469=>"101111111",
  29470=>"000000000",
  29471=>"000011111",
  29472=>"111111111",
  29473=>"000000000",
  29474=>"000100111",
  29475=>"010011010",
  29476=>"000000010",
  29477=>"111111011",
  29478=>"000000010",
  29479=>"100000111",
  29480=>"111100000",
  29481=>"000000111",
  29482=>"101000111",
  29483=>"001111111",
  29484=>"110110000",
  29485=>"100101101",
  29486=>"000000000",
  29487=>"000000000",
  29488=>"000000000",
  29489=>"000010011",
  29490=>"001111111",
  29491=>"001001001",
  29492=>"000000000",
  29493=>"000000100",
  29494=>"000100100",
  29495=>"111101000",
  29496=>"101001111",
  29497=>"100100111",
  29498=>"111111111",
  29499=>"111111111",
  29500=>"001100000",
  29501=>"000000101",
  29502=>"000000000",
  29503=>"111111110",
  29504=>"111111111",
  29505=>"000000001",
  29506=>"000001000",
  29507=>"111111100",
  29508=>"111110000",
  29509=>"010011001",
  29510=>"000000000",
  29511=>"111110000",
  29512=>"001011011",
  29513=>"000000000",
  29514=>"001111110",
  29515=>"001000001",
  29516=>"001000101",
  29517=>"001111000",
  29518=>"000000000",
  29519=>"111001001",
  29520=>"111001001",
  29521=>"111111111",
  29522=>"100100111",
  29523=>"000000000",
  29524=>"000000010",
  29525=>"111001111",
  29526=>"000100101",
  29527=>"010110111",
  29528=>"010010000",
  29529=>"110111110",
  29530=>"011111111",
  29531=>"001101111",
  29532=>"000000000",
  29533=>"111000000",
  29534=>"101100000",
  29535=>"111111111",
  29536=>"001000100",
  29537=>"010100111",
  29538=>"111100100",
  29539=>"100111111",
  29540=>"100001011",
  29541=>"000000000",
  29542=>"000000000",
  29543=>"111111101",
  29544=>"111100100",
  29545=>"111001001",
  29546=>"111111110",
  29547=>"101101111",
  29548=>"001111100",
  29549=>"111101000",
  29550=>"111111000",
  29551=>"000010111",
  29552=>"000000000",
  29553=>"111111111",
  29554=>"000000000",
  29555=>"111111111",
  29556=>"110110111",
  29557=>"000000000",
  29558=>"001111001",
  29559=>"000000000",
  29560=>"111111000",
  29561=>"000011101",
  29562=>"000000000",
  29563=>"011111100",
  29564=>"100100111",
  29565=>"000000000",
  29566=>"100100000",
  29567=>"110100000",
  29568=>"000111111",
  29569=>"001101111",
  29570=>"111000000",
  29571=>"000000000",
  29572=>"000100100",
  29573=>"110110000",
  29574=>"010111111",
  29575=>"100110110",
  29576=>"000000000",
  29577=>"100100111",
  29578=>"001001111",
  29579=>"110110000",
  29580=>"111000010",
  29581=>"110100000",
  29582=>"000100110",
  29583=>"111111111",
  29584=>"000000000",
  29585=>"111111001",
  29586=>"100101111",
  29587=>"000000000",
  29588=>"111111111",
  29589=>"001001001",
  29590=>"001011000",
  29591=>"000010010",
  29592=>"111111111",
  29593=>"111101111",
  29594=>"111000000",
  29595=>"111111111",
  29596=>"000000000",
  29597=>"000000000",
  29598=>"000000000",
  29599=>"110000110",
  29600=>"111111111",
  29601=>"010110010",
  29602=>"001011001",
  29603=>"000110000",
  29604=>"000000000",
  29605=>"110100000",
  29606=>"111110000",
  29607=>"011111000",
  29608=>"001000000",
  29609=>"100100000",
  29610=>"000000000",
  29611=>"111111000",
  29612=>"111111111",
  29613=>"000100100",
  29614=>"000000000",
  29615=>"111111111",
  29616=>"000000111",
  29617=>"100000000",
  29618=>"010010110",
  29619=>"000111111",
  29620=>"000000101",
  29621=>"111111111",
  29622=>"001111111",
  29623=>"000000000",
  29624=>"100101111",
  29625=>"100111111",
  29626=>"111111100",
  29627=>"000000000",
  29628=>"101100111",
  29629=>"111111010",
  29630=>"000000000",
  29631=>"111011001",
  29632=>"001011000",
  29633=>"101001000",
  29634=>"111111110",
  29635=>"001001001",
  29636=>"111111000",
  29637=>"111000101",
  29638=>"000110111",
  29639=>"000000000",
  29640=>"000000110",
  29641=>"110111111",
  29642=>"000110000",
  29643=>"100100111",
  29644=>"000000111",
  29645=>"000000000",
  29646=>"111110100",
  29647=>"111111011",
  29648=>"000000100",
  29649=>"000111000",
  29650=>"100111111",
  29651=>"011111111",
  29652=>"000001000",
  29653=>"110110000",
  29654=>"010000000",
  29655=>"100100100",
  29656=>"011111001",
  29657=>"000000000",
  29658=>"000111111",
  29659=>"100111110",
  29660=>"000000010",
  29661=>"111111111",
  29662=>"001011000",
  29663=>"110000000",
  29664=>"011111111",
  29665=>"111011000",
  29666=>"110000111",
  29667=>"000000000",
  29668=>"100100100",
  29669=>"001001111",
  29670=>"111101101",
  29671=>"111111011",
  29672=>"110110111",
  29673=>"000011011",
  29674=>"011111111",
  29675=>"111011111",
  29676=>"000000000",
  29677=>"110100111",
  29678=>"001001000",
  29679=>"111111110",
  29680=>"111111111",
  29681=>"100000000",
  29682=>"111101001",
  29683=>"010111111",
  29684=>"111111111",
  29685=>"000000000",
  29686=>"000000000",
  29687=>"111100111",
  29688=>"111111001",
  29689=>"111001001",
  29690=>"111001000",
  29691=>"000000000",
  29692=>"111111111",
  29693=>"000000000",
  29694=>"000010000",
  29695=>"111011111",
  29696=>"110110110",
  29697=>"000000110",
  29698=>"011011011",
  29699=>"000000000",
  29700=>"100110110",
  29701=>"001001101",
  29702=>"000001000",
  29703=>"111111111",
  29704=>"101101111",
  29705=>"000011011",
  29706=>"111111110",
  29707=>"100100100",
  29708=>"001001011",
  29709=>"111111010",
  29710=>"010011000",
  29711=>"010010110",
  29712=>"110111111",
  29713=>"000000000",
  29714=>"000000100",
  29715=>"000110010",
  29716=>"000000000",
  29717=>"000001101",
  29718=>"000100110",
  29719=>"111111111",
  29720=>"000000111",
  29721=>"000000001",
  29722=>"101000111",
  29723=>"011011111",
  29724=>"001001000",
  29725=>"000000000",
  29726=>"110111111",
  29727=>"000000000",
  29728=>"000000000",
  29729=>"000000000",
  29730=>"001001101",
  29731=>"000000101",
  29732=>"110110000",
  29733=>"110010000",
  29734=>"110111111",
  29735=>"011001000",
  29736=>"111111001",
  29737=>"000011001",
  29738=>"011000000",
  29739=>"111000101",
  29740=>"000000101",
  29741=>"111111000",
  29742=>"101000000",
  29743=>"011111111",
  29744=>"110110110",
  29745=>"111110010",
  29746=>"000001001",
  29747=>"000001011",
  29748=>"000000001",
  29749=>"001001000",
  29750=>"000000000",
  29751=>"001000001",
  29752=>"000111100",
  29753=>"111111011",
  29754=>"111011001",
  29755=>"111111111",
  29756=>"000000000",
  29757=>"111111111",
  29758=>"010111010",
  29759=>"001001001",
  29760=>"000000001",
  29761=>"000000000",
  29762=>"001000000",
  29763=>"111100000",
  29764=>"100100100",
  29765=>"000000110",
  29766=>"111111001",
  29767=>"001111111",
  29768=>"100100100",
  29769=>"111001011",
  29770=>"110010110",
  29771=>"000001000",
  29772=>"001101111",
  29773=>"010000000",
  29774=>"000011011",
  29775=>"110111110",
  29776=>"000000100",
  29777=>"000001000",
  29778=>"100000001",
  29779=>"110110000",
  29780=>"110110000",
  29781=>"000001111",
  29782=>"000000000",
  29783=>"000000000",
  29784=>"000000110",
  29785=>"111001111",
  29786=>"000101100",
  29787=>"000011000",
  29788=>"000001011",
  29789=>"111111111",
  29790=>"111001000",
  29791=>"011111110",
  29792=>"000000010",
  29793=>"111010000",
  29794=>"000000010",
  29795=>"001101101",
  29796=>"100000101",
  29797=>"000000100",
  29798=>"000001110",
  29799=>"111111000",
  29800=>"001111111",
  29801=>"101101111",
  29802=>"111111001",
  29803=>"000000000",
  29804=>"110110110",
  29805=>"111111111",
  29806=>"001001000",
  29807=>"111111111",
  29808=>"000000101",
  29809=>"110110000",
  29810=>"000000001",
  29811=>"000001111",
  29812=>"110000010",
  29813=>"110010010",
  29814=>"001001101",
  29815=>"001000001",
  29816=>"001000000",
  29817=>"001000010",
  29818=>"000000001",
  29819=>"111101000",
  29820=>"100110100",
  29821=>"100111000",
  29822=>"000000001",
  29823=>"000000000",
  29824=>"001001001",
  29825=>"000100110",
  29826=>"000000110",
  29827=>"011011000",
  29828=>"000001001",
  29829=>"000000000",
  29830=>"110110000",
  29831=>"000000000",
  29832=>"000100010",
  29833=>"000001001",
  29834=>"000001000",
  29835=>"000000111",
  29836=>"100100000",
  29837=>"001000000",
  29838=>"000101001",
  29839=>"000000000",
  29840=>"001100100",
  29841=>"110110000",
  29842=>"000000110",
  29843=>"111011111",
  29844=>"111001000",
  29845=>"111110111",
  29846=>"100100110",
  29847=>"000101101",
  29848=>"001111111",
  29849=>"111111111",
  29850=>"000001001",
  29851=>"000000000",
  29852=>"110000000",
  29853=>"011010110",
  29854=>"100000001",
  29855=>"000001001",
  29856=>"011001000",
  29857=>"000110111",
  29858=>"000001111",
  29859=>"000001101",
  29860=>"000001001",
  29861=>"000011001",
  29862=>"000000000",
  29863=>"100110000",
  29864=>"111111000",
  29865=>"000100000",
  29866=>"111111111",
  29867=>"000000000",
  29868=>"010011011",
  29869=>"000010111",
  29870=>"100101101",
  29871=>"000000111",
  29872=>"010110110",
  29873=>"010000100",
  29874=>"111111111",
  29875=>"000000000",
  29876=>"100000011",
  29877=>"000100111",
  29878=>"001101111",
  29879=>"000001001",
  29880=>"001101111",
  29881=>"010010011",
  29882=>"001001001",
  29883=>"100001000",
  29884=>"100111111",
  29885=>"001000000",
  29886=>"001001001",
  29887=>"011111111",
  29888=>"000000100",
  29889=>"000000100",
  29890=>"111111111",
  29891=>"000000000",
  29892=>"111111111",
  29893=>"000011000",
  29894=>"100110110",
  29895=>"000000101",
  29896=>"000000110",
  29897=>"100100111",
  29898=>"100000000",
  29899=>"001111100",
  29900=>"101101111",
  29901=>"011110111",
  29902=>"111111111",
  29903=>"000000010",
  29904=>"000000011",
  29905=>"000110111",
  29906=>"000010010",
  29907=>"101101101",
  29908=>"011001000",
  29909=>"111111111",
  29910=>"111111111",
  29911=>"110111000",
  29912=>"010001111",
  29913=>"111111111",
  29914=>"111000000",
  29915=>"000000111",
  29916=>"000100000",
  29917=>"100100111",
  29918=>"100101101",
  29919=>"000011011",
  29920=>"000000000",
  29921=>"000111111",
  29922=>"000000110",
  29923=>"010000000",
  29924=>"111110100",
  29925=>"111001000",
  29926=>"111000000",
  29927=>"111111110",
  29928=>"000000110",
  29929=>"000010111",
  29930=>"000101111",
  29931=>"110111111",
  29932=>"000000110",
  29933=>"001100000",
  29934=>"000000111",
  29935=>"000000001",
  29936=>"000000101",
  29937=>"111110000",
  29938=>"111111111",
  29939=>"000000000",
  29940=>"110111110",
  29941=>"000000001",
  29942=>"000000001",
  29943=>"111111111",
  29944=>"000000000",
  29945=>"000000010",
  29946=>"000010011",
  29947=>"000010010",
  29948=>"001001000",
  29949=>"000000001",
  29950=>"110110111",
  29951=>"101100001",
  29952=>"000111111",
  29953=>"111001101",
  29954=>"111101111",
  29955=>"000000000",
  29956=>"001001111",
  29957=>"110111111",
  29958=>"110101111",
  29959=>"000000111",
  29960=>"110111111",
  29961=>"000000000",
  29962=>"000000000",
  29963=>"100100000",
  29964=>"011001001",
  29965=>"000000000",
  29966=>"000000000",
  29967=>"011010000",
  29968=>"010100100",
  29969=>"000110111",
  29970=>"001001101",
  29971=>"000110111",
  29972=>"000000000",
  29973=>"011010000",
  29974=>"101101111",
  29975=>"111111101",
  29976=>"110110011",
  29977=>"111111110",
  29978=>"001011111",
  29979=>"000000111",
  29980=>"001101110",
  29981=>"000100110",
  29982=>"111001000",
  29983=>"000110110",
  29984=>"011011000",
  29985=>"000000001",
  29986=>"000011100",
  29987=>"111111011",
  29988=>"010010110",
  29989=>"100000101",
  29990=>"011001000",
  29991=>"110110000",
  29992=>"001001100",
  29993=>"110110010",
  29994=>"111111001",
  29995=>"011011011",
  29996=>"111111110",
  29997=>"100000001",
  29998=>"000000000",
  29999=>"100101101",
  30000=>"100011111",
  30001=>"000000110",
  30002=>"111111111",
  30003=>"100000111",
  30004=>"111000001",
  30005=>"010110010",
  30006=>"000011111",
  30007=>"111111111",
  30008=>"111001011",
  30009=>"111101001",
  30010=>"001111111",
  30011=>"100100111",
  30012=>"111001111",
  30013=>"001001001",
  30014=>"110110110",
  30015=>"110111000",
  30016=>"000000111",
  30017=>"000111111",
  30018=>"111111111",
  30019=>"111111000",
  30020=>"110111110",
  30021=>"000101111",
  30022=>"010000000",
  30023=>"000000000",
  30024=>"000000100",
  30025=>"000000000",
  30026=>"000000000",
  30027=>"000000100",
  30028=>"111111111",
  30029=>"000101111",
  30030=>"111111010",
  30031=>"110111111",
  30032=>"011111101",
  30033=>"111111111",
  30034=>"111111111",
  30035=>"000001111",
  30036=>"000011010",
  30037=>"011011001",
  30038=>"110110000",
  30039=>"000000001",
  30040=>"001000101",
  30041=>"000110000",
  30042=>"000000000",
  30043=>"111001101",
  30044=>"010010010",
  30045=>"000000000",
  30046=>"111111111",
  30047=>"111111111",
  30048=>"110000100",
  30049=>"110110000",
  30050=>"111111111",
  30051=>"000000010",
  30052=>"111111011",
  30053=>"000000000",
  30054=>"111111111",
  30055=>"001011111",
  30056=>"100010011",
  30057=>"111111111",
  30058=>"000000111",
  30059=>"000110110",
  30060=>"110110000",
  30061=>"001011000",
  30062=>"111111111",
  30063=>"000000000",
  30064=>"101100100",
  30065=>"000000000",
  30066=>"110111111",
  30067=>"000100111",
  30068=>"011011000",
  30069=>"101111111",
  30070=>"011011100",
  30071=>"100001111",
  30072=>"111111111",
  30073=>"010111110",
  30074=>"110110110",
  30075=>"000000000",
  30076=>"000000000",
  30077=>"110110010",
  30078=>"101101111",
  30079=>"000000101",
  30080=>"110110111",
  30081=>"110110100",
  30082=>"000000111",
  30083=>"101001011",
  30084=>"000000000",
  30085=>"111011000",
  30086=>"111011000",
  30087=>"111110110",
  30088=>"111101111",
  30089=>"000111111",
  30090=>"111111011",
  30091=>"000010111",
  30092=>"110010111",
  30093=>"000110011",
  30094=>"100000111",
  30095=>"000000111",
  30096=>"110010010",
  30097=>"110110000",
  30098=>"111111111",
  30099=>"100100110",
  30100=>"111111010",
  30101=>"000011000",
  30102=>"010000000",
  30103=>"000000000",
  30104=>"000000111",
  30105=>"111111111",
  30106=>"000000000",
  30107=>"110111000",
  30108=>"000100111",
  30109=>"000010000",
  30110=>"000000100",
  30111=>"000000100",
  30112=>"000110110",
  30113=>"000011000",
  30114=>"110111111",
  30115=>"101100100",
  30116=>"110111111",
  30117=>"000000000",
  30118=>"111111011",
  30119=>"000011110",
  30120=>"111101111",
  30121=>"111111001",
  30122=>"000000000",
  30123=>"101101001",
  30124=>"000000111",
  30125=>"110111101",
  30126=>"000000111",
  30127=>"111111111",
  30128=>"101001101",
  30129=>"111111000",
  30130=>"110111111",
  30131=>"010111001",
  30132=>"000000101",
  30133=>"100001001",
  30134=>"111111111",
  30135=>"001000000",
  30136=>"111000111",
  30137=>"110110010",
  30138=>"010000101",
  30139=>"110101111",
  30140=>"000001111",
  30141=>"111000000",
  30142=>"000000111",
  30143=>"101111001",
  30144=>"000000100",
  30145=>"111111111",
  30146=>"000000000",
  30147=>"000101111",
  30148=>"110011011",
  30149=>"010000011",
  30150=>"111011001",
  30151=>"000100000",
  30152=>"000001001",
  30153=>"000011011",
  30154=>"101001101",
  30155=>"101100111",
  30156=>"111111000",
  30157=>"110110000",
  30158=>"000000000",
  30159=>"001111011",
  30160=>"001001000",
  30161=>"100100111",
  30162=>"000011111",
  30163=>"000101000",
  30164=>"111111000",
  30165=>"111000000",
  30166=>"001000000",
  30167=>"100110100",
  30168=>"000000111",
  30169=>"010100100",
  30170=>"000000110",
  30171=>"111111111",
  30172=>"000010000",
  30173=>"110110000",
  30174=>"011000111",
  30175=>"111110101",
  30176=>"101101111",
  30177=>"000110111",
  30178=>"100000000",
  30179=>"010000010",
  30180=>"111101001",
  30181=>"100000111",
  30182=>"000111111",
  30183=>"111111000",
  30184=>"110010001",
  30185=>"000000000",
  30186=>"111111111",
  30187=>"001001001",
  30188=>"000000000",
  30189=>"100100000",
  30190=>"000000001",
  30191=>"110111111",
  30192=>"000000001",
  30193=>"000001101",
  30194=>"000001011",
  30195=>"100000000",
  30196=>"100001001",
  30197=>"111110010",
  30198=>"111111111",
  30199=>"000000000",
  30200=>"001000111",
  30201=>"111001111",
  30202=>"001001011",
  30203=>"001111111",
  30204=>"111111001",
  30205=>"110110110",
  30206=>"111101001",
  30207=>"000000111",
  30208=>"001011001",
  30209=>"000111111",
  30210=>"111101111",
  30211=>"100000000",
  30212=>"111111000",
  30213=>"000000000",
  30214=>"111001011",
  30215=>"111111111",
  30216=>"111111111",
  30217=>"001001000",
  30218=>"000000000",
  30219=>"000100000",
  30220=>"111111111",
  30221=>"000000000",
  30222=>"110100000",
  30223=>"000000000",
  30224=>"111111111",
  30225=>"111111111",
  30226=>"110111111",
  30227=>"000000000",
  30228=>"111111111",
  30229=>"111101000",
  30230=>"000000000",
  30231=>"001000100",
  30232=>"110111110",
  30233=>"111101101",
  30234=>"000101111",
  30235=>"111000000",
  30236=>"100000000",
  30237=>"111111111",
  30238=>"001111110",
  30239=>"000110100",
  30240=>"001001000",
  30241=>"111101100",
  30242=>"111111110",
  30243=>"100001001",
  30244=>"000000000",
  30245=>"111111001",
  30246=>"000010010",
  30247=>"111111110",
  30248=>"111000111",
  30249=>"000000000",
  30250=>"000000000",
  30251=>"101111111",
  30252=>"111111111",
  30253=>"000000000",
  30254=>"101101100",
  30255=>"000000100",
  30256=>"000010000",
  30257=>"001000000",
  30258=>"010110110",
  30259=>"000000000",
  30260=>"000000100",
  30261=>"111011101",
  30262=>"111111111",
  30263=>"101001111",
  30264=>"100111000",
  30265=>"000000000",
  30266=>"111111010",
  30267=>"111111111",
  30268=>"000101100",
  30269=>"110111111",
  30270=>"110000111",
  30271=>"111100000",
  30272=>"111110010",
  30273=>"000000000",
  30274=>"111111101",
  30275=>"001011011",
  30276=>"000100100",
  30277=>"001001100",
  30278=>"000111111",
  30279=>"111101111",
  30280=>"101110000",
  30281=>"000000000",
  30282=>"000000000",
  30283=>"000000001",
  30284=>"000110000",
  30285=>"000000000",
  30286=>"100111111",
  30287=>"110110110",
  30288=>"000000000",
  30289=>"111111001",
  30290=>"000010000",
  30291=>"001001001",
  30292=>"000000000",
  30293=>"000000111",
  30294=>"000000010",
  30295=>"111111111",
  30296=>"101001000",
  30297=>"000000000",
  30298=>"000000111",
  30299=>"000000111",
  30300=>"111011000",
  30301=>"111111111",
  30302=>"001000110",
  30303=>"000000100",
  30304=>"001001111",
  30305=>"001111011",
  30306=>"110110000",
  30307=>"111000111",
  30308=>"001000000",
  30309=>"101111111",
  30310=>"000000000",
  30311=>"000000000",
  30312=>"000000000",
  30313=>"111111000",
  30314=>"000110111",
  30315=>"110010000",
  30316=>"111011010",
  30317=>"111111110",
  30318=>"001001001",
  30319=>"000100111",
  30320=>"000111011",
  30321=>"111111000",
  30322=>"000000000",
  30323=>"111111110",
  30324=>"011111110",
  30325=>"011001111",
  30326=>"000111111",
  30327=>"000000000",
  30328=>"000000000",
  30329=>"000000011",
  30330=>"000000000",
  30331=>"000001011",
  30332=>"100100100",
  30333=>"111111111",
  30334=>"110110110",
  30335=>"110000000",
  30336=>"111111000",
  30337=>"100100110",
  30338=>"001001111",
  30339=>"110110110",
  30340=>"100111100",
  30341=>"001101111",
  30342=>"000000000",
  30343=>"100101111",
  30344=>"111001101",
  30345=>"000000000",
  30346=>"001111001",
  30347=>"111111111",
  30348=>"111111000",
  30349=>"110111111",
  30350=>"111111111",
  30351=>"000000000",
  30352=>"011111111",
  30353=>"000000000",
  30354=>"000000000",
  30355=>"111100000",
  30356=>"001011000",
  30357=>"110000000",
  30358=>"000000000",
  30359=>"111111111",
  30360=>"110111111",
  30361=>"111111000",
  30362=>"111011001",
  30363=>"000000000",
  30364=>"101111111",
  30365=>"111000010",
  30366=>"111111111",
  30367=>"000000000",
  30368=>"111011111",
  30369=>"110111111",
  30370=>"111111110",
  30371=>"111111110",
  30372=>"111111010",
  30373=>"111111111",
  30374=>"111111010",
  30375=>"110110110",
  30376=>"000000000",
  30377=>"000100111",
  30378=>"111111000",
  30379=>"111111000",
  30380=>"000010111",
  30381=>"100111111",
  30382=>"111000000",
  30383=>"001111011",
  30384=>"000000000",
  30385=>"111111111",
  30386=>"110110110",
  30387=>"111111011",
  30388=>"000000010",
  30389=>"001000000",
  30390=>"000001111",
  30391=>"111111111",
  30392=>"111011011",
  30393=>"111111111",
  30394=>"111111000",
  30395=>"111111111",
  30396=>"000000000",
  30397=>"000000101",
  30398=>"011111111",
  30399=>"111111111",
  30400=>"110111010",
  30401=>"001001000",
  30402=>"000001000",
  30403=>"111111111",
  30404=>"000000100",
  30405=>"000000000",
  30406=>"001000001",
  30407=>"000000000",
  30408=>"111111111",
  30409=>"000000000",
  30410=>"000000011",
  30411=>"000000000",
  30412=>"110111111",
  30413=>"100100011",
  30414=>"000000110",
  30415=>"111111111",
  30416=>"000111000",
  30417=>"111111000",
  30418=>"000100010",
  30419=>"000000000",
  30420=>"101110100",
  30421=>"111111111",
  30422=>"001001000",
  30423=>"111111111",
  30424=>"000000000",
  30425=>"111111111",
  30426=>"111101101",
  30427=>"000000010",
  30428=>"000000110",
  30429=>"010000000",
  30430=>"111111000",
  30431=>"000000000",
  30432=>"111101001",
  30433=>"100000000",
  30434=>"000000000",
  30435=>"111111011",
  30436=>"111111111",
  30437=>"000000110",
  30438=>"111111111",
  30439=>"000111111",
  30440=>"001001111",
  30441=>"111100000",
  30442=>"000000001",
  30443=>"001111010",
  30444=>"011111111",
  30445=>"000000000",
  30446=>"111111101",
  30447=>"000111111",
  30448=>"111110111",
  30449=>"111111111",
  30450=>"010000000",
  30451=>"010000000",
  30452=>"100100100",
  30453=>"100000011",
  30454=>"000100000",
  30455=>"110111111",
  30456=>"000000000",
  30457=>"000110111",
  30458=>"000000000",
  30459=>"111101101",
  30460=>"000000000",
  30461=>"100101000",
  30462=>"111111110",
  30463=>"000000000",
  30464=>"111111101",
  30465=>"000000000",
  30466=>"111111111",
  30467=>"101100110",
  30468=>"110111000",
  30469=>"111011001",
  30470=>"000000000",
  30471=>"000000000",
  30472=>"000000000",
  30473=>"000000000",
  30474=>"000000000",
  30475=>"000101000",
  30476=>"111100111",
  30477=>"111111111",
  30478=>"111111111",
  30479=>"001111001",
  30480=>"111111111",
  30481=>"001111111",
  30482=>"111111111",
  30483=>"000000000",
  30484=>"111011001",
  30485=>"000110110",
  30486=>"111111111",
  30487=>"111111111",
  30488=>"001001011",
  30489=>"000000000",
  30490=>"000000000",
  30491=>"000000000",
  30492=>"111111110",
  30493=>"001111111",
  30494=>"111111111",
  30495=>"101111001",
  30496=>"100000000",
  30497=>"111111000",
  30498=>"000000000",
  30499=>"110100110",
  30500=>"111111111",
  30501=>"000000100",
  30502=>"111111111",
  30503=>"000000000",
  30504=>"111111111",
  30505=>"110110010",
  30506=>"000111000",
  30507=>"000000000",
  30508=>"111111111",
  30509=>"110000000",
  30510=>"111111111",
  30511=>"000000100",
  30512=>"111001000",
  30513=>"111111111",
  30514=>"111111111",
  30515=>"100111111",
  30516=>"111101111",
  30517=>"110111111",
  30518=>"000000000",
  30519=>"001000000",
  30520=>"000100000",
  30521=>"000000000",
  30522=>"111111111",
  30523=>"111000101",
  30524=>"001000000",
  30525=>"001111110",
  30526=>"111011000",
  30527=>"000000110",
  30528=>"000000001",
  30529=>"000000111",
  30530=>"000000000",
  30531=>"111111111",
  30532=>"100100000",
  30533=>"110111111",
  30534=>"111011010",
  30535=>"111111111",
  30536=>"000000000",
  30537=>"000000111",
  30538=>"000111111",
  30539=>"000000000",
  30540=>"000100110",
  30541=>"000100010",
  30542=>"010000100",
  30543=>"000000000",
  30544=>"111000000",
  30545=>"000000000",
  30546=>"111111110",
  30547=>"011111111",
  30548=>"000000000",
  30549=>"001001011",
  30550=>"111011000",
  30551=>"011001001",
  30552=>"110000101",
  30553=>"000011000",
  30554=>"111111111",
  30555=>"010110111",
  30556=>"111111101",
  30557=>"111111110",
  30558=>"001011010",
  30559=>"101000000",
  30560=>"000000000",
  30561=>"000000000",
  30562=>"110111111",
  30563=>"001101111",
  30564=>"111110110",
  30565=>"000000001",
  30566=>"000000000",
  30567=>"000001111",
  30568=>"001000001",
  30569=>"111111000",
  30570=>"111011000",
  30571=>"000000000",
  30572=>"100100100",
  30573=>"000111110",
  30574=>"000000111",
  30575=>"000110000",
  30576=>"110110111",
  30577=>"000011111",
  30578=>"100100000",
  30579=>"000000000",
  30580=>"111111111",
  30581=>"000000000",
  30582=>"111111010",
  30583=>"000000011",
  30584=>"000000000",
  30585=>"000111111",
  30586=>"000001111",
  30587=>"000000000",
  30588=>"110111111",
  30589=>"000000000",
  30590=>"000111100",
  30591=>"000000000",
  30592=>"000101111",
  30593=>"000000000",
  30594=>"111111000",
  30595=>"111111001",
  30596=>"000000000",
  30597=>"111001000",
  30598=>"100000000",
  30599=>"110010111",
  30600=>"111111011",
  30601=>"111111110",
  30602=>"000000000",
  30603=>"000000001",
  30604=>"000000000",
  30605=>"111000000",
  30606=>"000111111",
  30607=>"000000000",
  30608=>"000000010",
  30609=>"000000100",
  30610=>"000000000",
  30611=>"001001001",
  30612=>"111011000",
  30613=>"000000000",
  30614=>"100100000",
  30615=>"111111110",
  30616=>"111111111",
  30617=>"111111111",
  30618=>"011111001",
  30619=>"101111111",
  30620=>"011000000",
  30621=>"100110000",
  30622=>"011001000",
  30623=>"111111111",
  30624=>"000000000",
  30625=>"111111000",
  30626=>"001000101",
  30627=>"000011111",
  30628=>"001111111",
  30629=>"011011111",
  30630=>"000000000",
  30631=>"001001111",
  30632=>"000101111",
  30633=>"110110111",
  30634=>"111111111",
  30635=>"000000000",
  30636=>"111111111",
  30637=>"000000000",
  30638=>"000000000",
  30639=>"100100000",
  30640=>"011000000",
  30641=>"000000000",
  30642=>"111111000",
  30643=>"010111111",
  30644=>"111111111",
  30645=>"110000000",
  30646=>"111111111",
  30647=>"111000000",
  30648=>"000111111",
  30649=>"111111111",
  30650=>"000000110",
  30651=>"100000010",
  30652=>"111111001",
  30653=>"000111111",
  30654=>"111111001",
  30655=>"101100110",
  30656=>"010111011",
  30657=>"111101111",
  30658=>"111111111",
  30659=>"111111011",
  30660=>"000000000",
  30661=>"001000000",
  30662=>"000000000",
  30663=>"111001001",
  30664=>"111000000",
  30665=>"000000000",
  30666=>"000000000",
  30667=>"000000000",
  30668=>"010111000",
  30669=>"000000000",
  30670=>"000001000",
  30671=>"000001000",
  30672=>"001000001",
  30673=>"111111111",
  30674=>"010000010",
  30675=>"000000000",
  30676=>"001000000",
  30677=>"000000100",
  30678=>"000000000",
  30679=>"111001111",
  30680=>"000001100",
  30681=>"111111001",
  30682=>"000000000",
  30683=>"111111111",
  30684=>"000100000",
  30685=>"000001101",
  30686=>"100000000",
  30687=>"000100110",
  30688=>"101000000",
  30689=>"111111111",
  30690=>"111000111",
  30691=>"111111111",
  30692=>"111111111",
  30693=>"000000100",
  30694=>"111110000",
  30695=>"000000000",
  30696=>"111111111",
  30697=>"000000111",
  30698=>"000000000",
  30699=>"000000000",
  30700=>"111110000",
  30701=>"011111110",
  30702=>"111111100",
  30703=>"000000000",
  30704=>"111111111",
  30705=>"001111111",
  30706=>"000111111",
  30707=>"000000000",
  30708=>"111111111",
  30709=>"000000000",
  30710=>"111111100",
  30711=>"100100111",
  30712=>"110101101",
  30713=>"101001000",
  30714=>"001111011",
  30715=>"000000000",
  30716=>"111111111",
  30717=>"110110000",
  30718=>"001011111",
  30719=>"111000000",
  30720=>"111110100",
  30721=>"011010000",
  30722=>"011111111",
  30723=>"000000100",
  30724=>"001011011",
  30725=>"110110001",
  30726=>"000000000",
  30727=>"111100110",
  30728=>"000000111",
  30729=>"000000000",
  30730=>"110000000",
  30731=>"000001101",
  30732=>"001101110",
  30733=>"111100100",
  30734=>"010100100",
  30735=>"111111111",
  30736=>"111111110",
  30737=>"010110111",
  30738=>"100111101",
  30739=>"010000000",
  30740=>"111010111",
  30741=>"111111000",
  30742=>"101111111",
  30743=>"011001000",
  30744=>"111110111",
  30745=>"001001101",
  30746=>"000000000",
  30747=>"111111100",
  30748=>"010111011",
  30749=>"110000000",
  30750=>"001001000",
  30751=>"100100110",
  30752=>"110000000",
  30753=>"110110110",
  30754=>"001001011",
  30755=>"001000101",
  30756=>"111011010",
  30757=>"010111110",
  30758=>"001101001",
  30759=>"000100110",
  30760=>"100000000",
  30761=>"001001111",
  30762=>"110111111",
  30763=>"111001001",
  30764=>"011000110",
  30765=>"111010011",
  30766=>"000001000",
  30767=>"111110010",
  30768=>"111111111",
  30769=>"001001101",
  30770=>"011011001",
  30771=>"110111110",
  30772=>"110110000",
  30773=>"000000000",
  30774=>"111111111",
  30775=>"000101111",
  30776=>"110111111",
  30777=>"000001100",
  30778=>"000000000",
  30779=>"000000000",
  30780=>"101100101",
  30781=>"100000000",
  30782=>"011011011",
  30783=>"000000111",
  30784=>"111111000",
  30785=>"011011110",
  30786=>"101000000",
  30787=>"001001001",
  30788=>"101111100",
  30789=>"001001001",
  30790=>"000000110",
  30791=>"111111111",
  30792=>"001011011",
  30793=>"000000001",
  30794=>"111111110",
  30795=>"100000000",
  30796=>"000110000",
  30797=>"111110110",
  30798=>"000000111",
  30799=>"001000000",
  30800=>"101000000",
  30801=>"011111010",
  30802=>"100000000",
  30803=>"000000000",
  30804=>"000000000",
  30805=>"000000011",
  30806=>"000000000",
  30807=>"000101010",
  30808=>"110110010",
  30809=>"000000000",
  30810=>"001000000",
  30811=>"110010110",
  30812=>"000010010",
  30813=>"111000100",
  30814=>"001000101",
  30815=>"000000011",
  30816=>"000000110",
  30817=>"001101101",
  30818=>"101110110",
  30819=>"111101111",
  30820=>"110111100",
  30821=>"111101101",
  30822=>"101001111",
  30823=>"001000101",
  30824=>"111111111",
  30825=>"000000010",
  30826=>"000000111",
  30827=>"000000010",
  30828=>"110111101",
  30829=>"100000000",
  30830=>"110010000",
  30831=>"111111111",
  30832=>"111110010",
  30833=>"111001011",
  30834=>"001000000",
  30835=>"001000010",
  30836=>"111111111",
  30837=>"000000000",
  30838=>"110111010",
  30839=>"111111101",
  30840=>"000101101",
  30841=>"001001001",
  30842=>"001001001",
  30843=>"110010000",
  30844=>"100100100",
  30845=>"001001000",
  30846=>"001100100",
  30847=>"010011000",
  30848=>"000000000",
  30849=>"000001001",
  30850=>"000000000",
  30851=>"000001011",
  30852=>"010000001",
  30853=>"000000000",
  30854=>"111111100",
  30855=>"001101101",
  30856=>"000000000",
  30857=>"000000000",
  30858=>"111101101",
  30859=>"010010000",
  30860=>"000000000",
  30861=>"111111010",
  30862=>"101111001",
  30863=>"111000000",
  30864=>"000000001",
  30865=>"111111010",
  30866=>"010010011",
  30867=>"010110000",
  30868=>"001001101",
  30869=>"000100110",
  30870=>"000000000",
  30871=>"111111111",
  30872=>"101100111",
  30873=>"001010011",
  30874=>"111111111",
  30875=>"001001000",
  30876=>"000000000",
  30877=>"100110101",
  30878=>"110111101",
  30879=>"001101000",
  30880=>"111011000",
  30881=>"000000000",
  30882=>"000000011",
  30883=>"000000101",
  30884=>"001001001",
  30885=>"111111100",
  30886=>"110111111",
  30887=>"001100100",
  30888=>"111101111",
  30889=>"000000001",
  30890=>"011000000",
  30891=>"110110000",
  30892=>"000001111",
  30893=>"110110110",
  30894=>"001001000",
  30895=>"111111111",
  30896=>"111111000",
  30897=>"111111110",
  30898=>"111111111",
  30899=>"010000000",
  30900=>"111111110",
  30901=>"111111110",
  30902=>"000000000",
  30903=>"000100000",
  30904=>"000111111",
  30905=>"001101001",
  30906=>"101001000",
  30907=>"001000000",
  30908=>"111111111",
  30909=>"010000000",
  30910=>"000000000",
  30911=>"110110110",
  30912=>"000110000",
  30913=>"110110000",
  30914=>"110110110",
  30915=>"111111111",
  30916=>"000000100",
  30917=>"111111111",
  30918=>"011010010",
  30919=>"111111000",
  30920=>"000000000",
  30921=>"000100011",
  30922=>"000000101",
  30923=>"111101000",
  30924=>"001111111",
  30925=>"000011111",
  30926=>"000000110",
  30927=>"000000000",
  30928=>"010010000",
  30929=>"001000010",
  30930=>"010110010",
  30931=>"000000000",
  30932=>"110011010",
  30933=>"001001011",
  30934=>"111101111",
  30935=>"100100111",
  30936=>"000000110",
  30937=>"111111010",
  30938=>"101100111",
  30939=>"101111111",
  30940=>"000000000",
  30941=>"000111101",
  30942=>"111111101",
  30943=>"010000000",
  30944=>"001011111",
  30945=>"111011011",
  30946=>"111110110",
  30947=>"011111110",
  30948=>"111111111",
  30949=>"100001001",
  30950=>"000001111",
  30951=>"000111110",
  30952=>"010111111",
  30953=>"110110110",
  30954=>"101000000",
  30955=>"101101111",
  30956=>"000101111",
  30957=>"000000111",
  30958=>"111011000",
  30959=>"111101100",
  30960=>"000000001",
  30961=>"000000110",
  30962=>"010000111",
  30963=>"101000000",
  30964=>"000110100",
  30965=>"000100110",
  30966=>"011011001",
  30967=>"100111000",
  30968=>"111110101",
  30969=>"111111111",
  30970=>"101111000",
  30971=>"010010010",
  30972=>"000000001",
  30973=>"111110001",
  30974=>"000000100",
  30975=>"111110110",
  30976=>"001000001",
  30977=>"100110000",
  30978=>"111111000",
  30979=>"000000000",
  30980=>"111101001",
  30981=>"000110000",
  30982=>"011111111",
  30983=>"110110110",
  30984=>"000000001",
  30985=>"101101100",
  30986=>"111111111",
  30987=>"000000100",
  30988=>"111101111",
  30989=>"010011000",
  30990=>"110111110",
  30991=>"010111010",
  30992=>"011111000",
  30993=>"000000010",
  30994=>"000000000",
  30995=>"110110011",
  30996=>"000000000",
  30997=>"000000000",
  30998=>"001001000",
  30999=>"111111110",
  31000=>"000000000",
  31001=>"111111011",
  31002=>"000100100",
  31003=>"111110000",
  31004=>"100110110",
  31005=>"000110111",
  31006=>"000000000",
  31007=>"111111111",
  31008=>"011111000",
  31009=>"000100000",
  31010=>"011111100",
  31011=>"000000110",
  31012=>"011000000",
  31013=>"111101001",
  31014=>"100110111",
  31015=>"111110000",
  31016=>"101000000",
  31017=>"100111011",
  31018=>"001000011",
  31019=>"011011010",
  31020=>"000010010",
  31021=>"110110110",
  31022=>"110010111",
  31023=>"101001101",
  31024=>"100111111",
  31025=>"010111011",
  31026=>"101001000",
  31027=>"011000000",
  31028=>"010000010",
  31029=>"011111000",
  31030=>"010000000",
  31031=>"000000000",
  31032=>"000000000",
  31033=>"000000000",
  31034=>"000000101",
  31035=>"101101000",
  31036=>"000000000",
  31037=>"001001101",
  31038=>"111101101",
  31039=>"111111100",
  31040=>"011111110",
  31041=>"111100100",
  31042=>"000011001",
  31043=>"101000000",
  31044=>"111001000",
  31045=>"111111111",
  31046=>"101111111",
  31047=>"000100000",
  31048=>"111101101",
  31049=>"010000000",
  31050=>"000000000",
  31051=>"011011011",
  31052=>"001011000",
  31053=>"001011111",
  31054=>"111001111",
  31055=>"001001001",
  31056=>"011011011",
  31057=>"001000000",
  31058=>"111110111",
  31059=>"100001101",
  31060=>"001001100",
  31061=>"111011001",
  31062=>"000000000",
  31063=>"001101111",
  31064=>"110110000",
  31065=>"111111111",
  31066=>"001000000",
  31067=>"111111101",
  31068=>"000000100",
  31069=>"111110100",
  31070=>"101001000",
  31071=>"011111111",
  31072=>"111011111",
  31073=>"000000000",
  31074=>"000000000",
  31075=>"101000000",
  31076=>"110100100",
  31077=>"000000000",
  31078=>"111111111",
  31079=>"000010010",
  31080=>"100100110",
  31081=>"111001110",
  31082=>"000000000",
  31083=>"000110110",
  31084=>"100100000",
  31085=>"001000011",
  31086=>"000000000",
  31087=>"111001001",
  31088=>"000000000",
  31089=>"000000000",
  31090=>"101111110",
  31091=>"110100110",
  31092=>"011001000",
  31093=>"000000100",
  31094=>"000001111",
  31095=>"111111000",
  31096=>"111101100",
  31097=>"111110111",
  31098=>"000000110",
  31099=>"000000010",
  31100=>"000000111",
  31101=>"111111111",
  31102=>"111111000",
  31103=>"000000001",
  31104=>"001010000",
  31105=>"101101101",
  31106=>"000000000",
  31107=>"000000111",
  31108=>"000000111",
  31109=>"000011010",
  31110=>"000111111",
  31111=>"000111111",
  31112=>"000000000",
  31113=>"100111011",
  31114=>"101000001",
  31115=>"111101000",
  31116=>"101111111",
  31117=>"110101011",
  31118=>"000000000",
  31119=>"000000000",
  31120=>"010111111",
  31121=>"110000000",
  31122=>"000100000",
  31123=>"000000000",
  31124=>"000111111",
  31125=>"000000000",
  31126=>"000010011",
  31127=>"111111010",
  31128=>"111111011",
  31129=>"110110100",
  31130=>"000000001",
  31131=>"000000111",
  31132=>"000000101",
  31133=>"111111111",
  31134=>"000000000",
  31135=>"000111111",
  31136=>"111111111",
  31137=>"011011001",
  31138=>"111111000",
  31139=>"011001000",
  31140=>"101110000",
  31141=>"111111111",
  31142=>"111101111",
  31143=>"111110110",
  31144=>"011110010",
  31145=>"100110000",
  31146=>"001001000",
  31147=>"000000110",
  31148=>"001000000",
  31149=>"101101101",
  31150=>"001101111",
  31151=>"111111011",
  31152=>"111011000",
  31153=>"000000001",
  31154=>"011101000",
  31155=>"111111010",
  31156=>"001111111",
  31157=>"111111111",
  31158=>"011000100",
  31159=>"000000000",
  31160=>"000001000",
  31161=>"011111011",
  31162=>"111101100",
  31163=>"001001111",
  31164=>"010110110",
  31165=>"000000000",
  31166=>"000000000",
  31167=>"001000110",
  31168=>"000000111",
  31169=>"100110111",
  31170=>"111101111",
  31171=>"100101111",
  31172=>"111111111",
  31173=>"011001101",
  31174=>"110001001",
  31175=>"111000000",
  31176=>"101101111",
  31177=>"101100100",
  31178=>"000000000",
  31179=>"000100000",
  31180=>"011010110",
  31181=>"000110100",
  31182=>"110110010",
  31183=>"000000000",
  31184=>"000000000",
  31185=>"101101100",
  31186=>"100100001",
  31187=>"001001101",
  31188=>"101000101",
  31189=>"001000000",
  31190=>"001000000",
  31191=>"000001011",
  31192=>"100000100",
  31193=>"110000000",
  31194=>"000000000",
  31195=>"111110000",
  31196=>"011111111",
  31197=>"111111111",
  31198=>"111011011",
  31199=>"100100100",
  31200=>"001000110",
  31201=>"000000001",
  31202=>"000000000",
  31203=>"111101000",
  31204=>"000000110",
  31205=>"101001111",
  31206=>"111110110",
  31207=>"000000000",
  31208=>"110110110",
  31209=>"111111001",
  31210=>"000000001",
  31211=>"000011001",
  31212=>"010111010",
  31213=>"111111010",
  31214=>"111111011",
  31215=>"110111111",
  31216=>"100001101",
  31217=>"000101111",
  31218=>"011111011",
  31219=>"011111110",
  31220=>"101100000",
  31221=>"110111111",
  31222=>"001000100",
  31223=>"110110110",
  31224=>"111111100",
  31225=>"000001001",
  31226=>"001000000",
  31227=>"010110000",
  31228=>"111111101",
  31229=>"110100110",
  31230=>"000000000",
  31231=>"110000110",
  31232=>"000010110",
  31233=>"000000000",
  31234=>"000000000",
  31235=>"111000000",
  31236=>"001111111",
  31237=>"111111111",
  31238=>"111101000",
  31239=>"011111111",
  31240=>"001111111",
  31241=>"111111001",
  31242=>"000000111",
  31243=>"000000111",
  31244=>"111111111",
  31245=>"111000000",
  31246=>"111111000",
  31247=>"000111111",
  31248=>"000000000",
  31249=>"000111111",
  31250=>"110000000",
  31251=>"000000111",
  31252=>"000111111",
  31253=>"000001011",
  31254=>"111101000",
  31255=>"000000100",
  31256=>"100110111",
  31257=>"001011000",
  31258=>"111101111",
  31259=>"011010110",
  31260=>"000000111",
  31261=>"111111000",
  31262=>"111011111",
  31263=>"010100111",
  31264=>"000111111",
  31265=>"110000000",
  31266=>"000000000",
  31267=>"111111111",
  31268=>"111000000",
  31269=>"100000000",
  31270=>"111111111",
  31271=>"111111110",
  31272=>"010010000",
  31273=>"101000000",
  31274=>"000111111",
  31275=>"111000100",
  31276=>"000110111",
  31277=>"111111011",
  31278=>"110101101",
  31279=>"000000111",
  31280=>"111000000",
  31281=>"011111111",
  31282=>"000000000",
  31283=>"000000110",
  31284=>"111000000",
  31285=>"110000000",
  31286=>"000000000",
  31287=>"000001011",
  31288=>"000000111",
  31289=>"101000000",
  31290=>"000000000",
  31291=>"000000111",
  31292=>"111111000",
  31293=>"110000000",
  31294=>"111110111",
  31295=>"000000000",
  31296=>"111000100",
  31297=>"111000000",
  31298=>"111111110",
  31299=>"101000000",
  31300=>"000000000",
  31301=>"000000101",
  31302=>"110110100",
  31303=>"000000000",
  31304=>"111011110",
  31305=>"000000000",
  31306=>"000101001",
  31307=>"000100100",
  31308=>"000110111",
  31309=>"110111111",
  31310=>"000000000",
  31311=>"111110100",
  31312=>"000000000",
  31313=>"111111111",
  31314=>"111011001",
  31315=>"100000000",
  31316=>"000000000",
  31317=>"100100000",
  31318=>"000111110",
  31319=>"001000000",
  31320=>"000000000",
  31321=>"001000000",
  31322=>"000101111",
  31323=>"001111111",
  31324=>"101000000",
  31325=>"000000101",
  31326=>"000000001",
  31327=>"000001000",
  31328=>"111000000",
  31329=>"110000000",
  31330=>"000010111",
  31331=>"111111111",
  31332=>"001111111",
  31333=>"111111001",
  31334=>"111011000",
  31335=>"000000000",
  31336=>"101111001",
  31337=>"000000101",
  31338=>"100000110",
  31339=>"000000000",
  31340=>"111111000",
  31341=>"111011101",
  31342=>"000000000",
  31343=>"000000000",
  31344=>"000000000",
  31345=>"111100000",
  31346=>"111001000",
  31347=>"000100101",
  31348=>"000000111",
  31349=>"011011001",
  31350=>"000000000",
  31351=>"000111000",
  31352=>"111111000",
  31353=>"000110000",
  31354=>"111111000",
  31355=>"111110000",
  31356=>"000000011",
  31357=>"111000111",
  31358=>"000000111",
  31359=>"001000000",
  31360=>"000000100",
  31361=>"000010110",
  31362=>"001011000",
  31363=>"111111000",
  31364=>"000000000",
  31365=>"111000101",
  31366=>"011011001",
  31367=>"111000111",
  31368=>"000000000",
  31369=>"001101111",
  31370=>"000000000",
  31371=>"111111000",
  31372=>"111000110",
  31373=>"001011000",
  31374=>"111011000",
  31375=>"000111111",
  31376=>"000000111",
  31377=>"000000110",
  31378=>"000111000",
  31379=>"000000000",
  31380=>"000000111",
  31381=>"001111111",
  31382=>"000000000",
  31383=>"000000111",
  31384=>"000000001",
  31385=>"000110110",
  31386=>"111101101",
  31387=>"000000111",
  31388=>"000000000",
  31389=>"111111000",
  31390=>"000000000",
  31391=>"010011001",
  31392=>"000000101",
  31393=>"111000000",
  31394=>"000000000",
  31395=>"010000000",
  31396=>"111111000",
  31397=>"111111010",
  31398=>"111111111",
  31399=>"011110000",
  31400=>"110000000",
  31401=>"111001000",
  31402=>"000000000",
  31403=>"111111110",
  31404=>"110101000",
  31405=>"000000001",
  31406=>"111111111",
  31407=>"111111110",
  31408=>"011111110",
  31409=>"111110000",
  31410=>"111101111",
  31411=>"111101100",
  31412=>"111000010",
  31413=>"000101101",
  31414=>"000000000",
  31415=>"111110000",
  31416=>"110111100",
  31417=>"111111000",
  31418=>"000000000",
  31419=>"000111111",
  31420=>"000000000",
  31421=>"001000000",
  31422=>"111111011",
  31423=>"000001001",
  31424=>"000000111",
  31425=>"000001111",
  31426=>"000011001",
  31427=>"001001111",
  31428=>"111111000",
  31429=>"100111101",
  31430=>"111111000",
  31431=>"000111111",
  31432=>"111011000",
  31433=>"100000001",
  31434=>"111111111",
  31435=>"000000111",
  31436=>"001000000",
  31437=>"001000100",
  31438=>"111111111",
  31439=>"010111000",
  31440=>"111101110",
  31441=>"111111001",
  31442=>"100000000",
  31443=>"011000000",
  31444=>"000000000",
  31445=>"000110011",
  31446=>"100000000",
  31447=>"111011010",
  31448=>"111000000",
  31449=>"000000111",
  31450=>"111111000",
  31451=>"000011001",
  31452=>"000111111",
  31453=>"001011111",
  31454=>"000000100",
  31455=>"111111000",
  31456=>"111111010",
  31457=>"101111111",
  31458=>"111111111",
  31459=>"000010110",
  31460=>"111000010",
  31461=>"000011111",
  31462=>"000000011",
  31463=>"000000000",
  31464=>"111000000",
  31465=>"100111111",
  31466=>"110111111",
  31467=>"000000111",
  31468=>"000101100",
  31469=>"110111000",
  31470=>"011001001",
  31471=>"111110000",
  31472=>"011000000",
  31473=>"110111110",
  31474=>"111100000",
  31475=>"000111111",
  31476=>"010001001",
  31477=>"000000000",
  31478=>"001011111",
  31479=>"000001110",
  31480=>"111111111",
  31481=>"000000100",
  31482=>"111110000",
  31483=>"000101000",
  31484=>"100000001",
  31485=>"011000011",
  31486=>"000111111",
  31487=>"000000000",
  31488=>"111001000",
  31489=>"000000000",
  31490=>"010010000",
  31491=>"111111111",
  31492=>"000000100",
  31493=>"111000000",
  31494=>"000000111",
  31495=>"000111000",
  31496=>"000000101",
  31497=>"000111011",
  31498=>"111000011",
  31499=>"000001101",
  31500=>"000000111",
  31501=>"000000111",
  31502=>"000000000",
  31503=>"001001111",
  31504=>"000000000",
  31505=>"111111000",
  31506=>"111000000",
  31507=>"000000000",
  31508=>"110000000",
  31509=>"000000111",
  31510=>"100100110",
  31511=>"111111101",
  31512=>"111111001",
  31513=>"000010111",
  31514=>"001000000",
  31515=>"000000111",
  31516=>"000000000",
  31517=>"111111111",
  31518=>"111111111",
  31519=>"110110111",
  31520=>"000000110",
  31521=>"000110111",
  31522=>"000000111",
  31523=>"110110111",
  31524=>"001101111",
  31525=>"111000000",
  31526=>"000000001",
  31527=>"000000111",
  31528=>"111111100",
  31529=>"111000000",
  31530=>"000011011",
  31531=>"111111111",
  31532=>"001111111",
  31533=>"000110111",
  31534=>"000000000",
  31535=>"101111000",
  31536=>"000000010",
  31537=>"110110100",
  31538=>"001111110",
  31539=>"000000000",
  31540=>"111111111",
  31541=>"000001001",
  31542=>"111000100",
  31543=>"111001001",
  31544=>"111111111",
  31545=>"111111111",
  31546=>"000111111",
  31547=>"111111111",
  31548=>"011000000",
  31549=>"000000111",
  31550=>"000000000",
  31551=>"110011111",
  31552=>"000101101",
  31553=>"111110110",
  31554=>"110111011",
  31555=>"111111100",
  31556=>"011111111",
  31557=>"001000000",
  31558=>"000000000",
  31559=>"111111111",
  31560=>"111111111",
  31561=>"111000011",
  31562=>"111111110",
  31563=>"000000110",
  31564=>"101100000",
  31565=>"000000100",
  31566=>"000111111",
  31567=>"100000000",
  31568=>"000011011",
  31569=>"111011000",
  31570=>"000000010",
  31571=>"111111111",
  31572=>"111101000",
  31573=>"011000010",
  31574=>"100100000",
  31575=>"100000001",
  31576=>"000000000",
  31577=>"111111111",
  31578=>"000010111",
  31579=>"111000001",
  31580=>"000101100",
  31581=>"101000000",
  31582=>"111001000",
  31583=>"111110010",
  31584=>"111111000",
  31585=>"000000111",
  31586=>"111100100",
  31587=>"011001001",
  31588=>"111000000",
  31589=>"000000001",
  31590=>"111111000",
  31591=>"000000000",
  31592=>"000000010",
  31593=>"111111010",
  31594=>"001001000",
  31595=>"111111001",
  31596=>"000000001",
  31597=>"100111111",
  31598=>"010000000",
  31599=>"000000000",
  31600=>"111000000",
  31601=>"000000100",
  31602=>"000000000",
  31603=>"111111100",
  31604=>"111111000",
  31605=>"111011111",
  31606=>"000110111",
  31607=>"000000010",
  31608=>"111001011",
  31609=>"111111100",
  31610=>"000010001",
  31611=>"111111111",
  31612=>"000000111",
  31613=>"111000000",
  31614=>"111111000",
  31615=>"111001111",
  31616=>"000010011",
  31617=>"001001111",
  31618=>"000110111",
  31619=>"000000111",
  31620=>"000101111",
  31621=>"111111111",
  31622=>"111000000",
  31623=>"110000111",
  31624=>"111000000",
  31625=>"011011110",
  31626=>"111111111",
  31627=>"111111000",
  31628=>"111001001",
  31629=>"111111000",
  31630=>"110100111",
  31631=>"000000001",
  31632=>"001001100",
  31633=>"000111101",
  31634=>"111111010",
  31635=>"000000000",
  31636=>"000101111",
  31637=>"000011010",
  31638=>"111111111",
  31639=>"000000000",
  31640=>"111111111",
  31641=>"011101111",
  31642=>"111000000",
  31643=>"000000000",
  31644=>"101000000",
  31645=>"001111000",
  31646=>"100000000",
  31647=>"000101111",
  31648=>"111000111",
  31649=>"010010000",
  31650=>"000001001",
  31651=>"001000000",
  31652=>"111110110",
  31653=>"011011111",
  31654=>"111111111",
  31655=>"000010111",
  31656=>"101111111",
  31657=>"111001000",
  31658=>"111111111",
  31659=>"000000111",
  31660=>"000100100",
  31661=>"001001000",
  31662=>"000001000",
  31663=>"000111111",
  31664=>"000000000",
  31665=>"101001000",
  31666=>"100100000",
  31667=>"000000001",
  31668=>"101000000",
  31669=>"111111000",
  31670=>"000110100",
  31671=>"110100111",
  31672=>"000000001",
  31673=>"000111111",
  31674=>"011001001",
  31675=>"010000000",
  31676=>"111111001",
  31677=>"111110111",
  31678=>"000000000",
  31679=>"100110100",
  31680=>"111100111",
  31681=>"111001111",
  31682=>"111111000",
  31683=>"111101000",
  31684=>"000111011",
  31685=>"110111011",
  31686=>"100000000",
  31687=>"111101000",
  31688=>"000000101",
  31689=>"000000111",
  31690=>"001001000",
  31691=>"001000111",
  31692=>"111111011",
  31693=>"000111000",
  31694=>"100101000",
  31695=>"111111110",
  31696=>"110000000",
  31697=>"000000000",
  31698=>"001101111",
  31699=>"000000100",
  31700=>"100000100",
  31701=>"000000000",
  31702=>"111111100",
  31703=>"111110000",
  31704=>"000111110",
  31705=>"000000000",
  31706=>"000000111",
  31707=>"000111111",
  31708=>"111111111",
  31709=>"001000011",
  31710=>"001111111",
  31711=>"000010110",
  31712=>"101111111",
  31713=>"110000110",
  31714=>"000000100",
  31715=>"001011000",
  31716=>"000000111",
  31717=>"000001000",
  31718=>"110111111",
  31719=>"110000000",
  31720=>"111100000",
  31721=>"000110111",
  31722=>"111111000",
  31723=>"000000111",
  31724=>"111111001",
  31725=>"011000000",
  31726=>"101101111",
  31727=>"111110001",
  31728=>"100111000",
  31729=>"111111111",
  31730=>"111101001",
  31731=>"111111100",
  31732=>"111110000",
  31733=>"011000000",
  31734=>"000111111",
  31735=>"111001000",
  31736=>"111111111",
  31737=>"011011011",
  31738=>"111111111",
  31739=>"000000000",
  31740=>"000001111",
  31741=>"111000001",
  31742=>"001001111",
  31743=>"001001111",
  31744=>"111000000",
  31745=>"000000010",
  31746=>"000000000",
  31747=>"111011111",
  31748=>"111000110",
  31749=>"010000000",
  31750=>"001000100",
  31751=>"000000000",
  31752=>"101000001",
  31753=>"111111111",
  31754=>"000001111",
  31755=>"111111111",
  31756=>"111000000",
  31757=>"101111111",
  31758=>"111001001",
  31759=>"111111111",
  31760=>"000100101",
  31761=>"010001001",
  31762=>"111001000",
  31763=>"000000000",
  31764=>"000000000",
  31765=>"111111011",
  31766=>"010000000",
  31767=>"000000100",
  31768=>"110111110",
  31769=>"000000011",
  31770=>"111011111",
  31771=>"000011001",
  31772=>"000000000",
  31773=>"111111000",
  31774=>"011001001",
  31775=>"111111111",
  31776=>"111111110",
  31777=>"000111001",
  31778=>"001001111",
  31779=>"000101101",
  31780=>"111111111",
  31781=>"000000101",
  31782=>"000000000",
  31783=>"100100111",
  31784=>"000000000",
  31785=>"000000000",
  31786=>"000111111",
  31787=>"000000000",
  31788=>"111111111",
  31789=>"110110000",
  31790=>"100000000",
  31791=>"111111111",
  31792=>"111111111",
  31793=>"111001000",
  31794=>"111110111",
  31795=>"100110000",
  31796=>"111110110",
  31797=>"111000000",
  31798=>"000111110",
  31799=>"000111111",
  31800=>"000000000",
  31801=>"000000110",
  31802=>"000000110",
  31803=>"000000001",
  31804=>"111111111",
  31805=>"000110000",
  31806=>"111111111",
  31807=>"111111111",
  31808=>"111110000",
  31809=>"111111110",
  31810=>"000001111",
  31811=>"100111111",
  31812=>"110111111",
  31813=>"001001001",
  31814=>"000101111",
  31815=>"111111111",
  31816=>"011011011",
  31817=>"111101111",
  31818=>"000111111",
  31819=>"010110111",
  31820=>"110100000",
  31821=>"000000001",
  31822=>"111111110",
  31823=>"000001111",
  31824=>"000111111",
  31825=>"111111111",
  31826=>"000000000",
  31827=>"000100111",
  31828=>"000000000",
  31829=>"000000000",
  31830=>"000011001",
  31831=>"000000000",
  31832=>"010110010",
  31833=>"001001101",
  31834=>"001011111",
  31835=>"000100100",
  31836=>"000000000",
  31837=>"111111111",
  31838=>"000111000",
  31839=>"111110001",
  31840=>"100000000",
  31841=>"000000000",
  31842=>"010010000",
  31843=>"111110110",
  31844=>"110111110",
  31845=>"000000000",
  31846=>"000000000",
  31847=>"011011001",
  31848=>"111111101",
  31849=>"001001001",
  31850=>"110110000",
  31851=>"000000001",
  31852=>"110110110",
  31853=>"111111110",
  31854=>"000000001",
  31855=>"010010010",
  31856=>"000110010",
  31857=>"000111111",
  31858=>"111111110",
  31859=>"000000010",
  31860=>"010000000",
  31861=>"011001011",
  31862=>"000000000",
  31863=>"101101100",
  31864=>"111110000",
  31865=>"001000010",
  31866=>"111000101",
  31867=>"000000000",
  31868=>"110111110",
  31869=>"111111111",
  31870=>"001111100",
  31871=>"111111111",
  31872=>"000000000",
  31873=>"000000101",
  31874=>"111111101",
  31875=>"000000001",
  31876=>"111000000",
  31877=>"101001111",
  31878=>"110111111",
  31879=>"111101111",
  31880=>"000000000",
  31881=>"101000000",
  31882=>"111111100",
  31883=>"111010000",
  31884=>"111001001",
  31885=>"111111000",
  31886=>"001011110",
  31887=>"000000000",
  31888=>"000000000",
  31889=>"110100000",
  31890=>"011001001",
  31891=>"110100110",
  31892=>"011011111",
  31893=>"111111111",
  31894=>"011011000",
  31895=>"111100000",
  31896=>"000000111",
  31897=>"111001000",
  31898=>"000000100",
  31899=>"000000000",
  31900=>"000011111",
  31901=>"000000111",
  31902=>"000001001",
  31903=>"110100110",
  31904=>"111111110",
  31905=>"000111111",
  31906=>"000000000",
  31907=>"000000000",
  31908=>"011000000",
  31909=>"111111110",
  31910=>"001111110",
  31911=>"111111011",
  31912=>"010111101",
  31913=>"111111111",
  31914=>"000000000",
  31915=>"000000000",
  31916=>"000111111",
  31917=>"011000100",
  31918=>"111111111",
  31919=>"110110110",
  31920=>"000000000",
  31921=>"100111011",
  31922=>"010000110",
  31923=>"000000000",
  31924=>"111111110",
  31925=>"111111111",
  31926=>"111000000",
  31927=>"111010000",
  31928=>"111100110",
  31929=>"000000000",
  31930=>"000000011",
  31931=>"000000000",
  31932=>"111111010",
  31933=>"100100111",
  31934=>"100000000",
  31935=>"111000000",
  31936=>"111111111",
  31937=>"000000110",
  31938=>"111100111",
  31939=>"000000000",
  31940=>"110111111",
  31941=>"111111111",
  31942=>"000001111",
  31943=>"010000000",
  31944=>"000000111",
  31945=>"111111111",
  31946=>"000000000",
  31947=>"111111111",
  31948=>"000000111",
  31949=>"000000000",
  31950=>"000000011",
  31951=>"111111000",
  31952=>"111111011",
  31953=>"011010111",
  31954=>"001001100",
  31955=>"111111101",
  31956=>"100000000",
  31957=>"001011000",
  31958=>"000000000",
  31959=>"100000000",
  31960=>"000000000",
  31961=>"000111101",
  31962=>"000000000",
  31963=>"111111111",
  31964=>"111111111",
  31965=>"000000111",
  31966=>"101001000",
  31967=>"111011000",
  31968=>"001000000",
  31969=>"000111100",
  31970=>"111011001",
  31971=>"111111111",
  31972=>"001001000",
  31973=>"000001011",
  31974=>"111111111",
  31975=>"111111011",
  31976=>"111111101",
  31977=>"110110111",
  31978=>"000000111",
  31979=>"000000100",
  31980=>"111111111",
  31981=>"101001010",
  31982=>"111001011",
  31983=>"111011111",
  31984=>"000110110",
  31985=>"100100000",
  31986=>"100000001",
  31987=>"000000111",
  31988=>"000111111",
  31989=>"111111000",
  31990=>"011011111",
  31991=>"111010000",
  31992=>"111111111",
  31993=>"111100111",
  31994=>"001100111",
  31995=>"110111111",
  31996=>"110110100",
  31997=>"111011000",
  31998=>"100111100",
  31999=>"011111011",
  32000=>"000101111",
  32001=>"111011111",
  32002=>"111111111",
  32003=>"101000000",
  32004=>"100000000",
  32005=>"000000000",
  32006=>"001001111",
  32007=>"000000110",
  32008=>"000100000",
  32009=>"000000000",
  32010=>"000000100",
  32011=>"001101111",
  32012=>"111000000",
  32013=>"000000001",
  32014=>"000011000",
  32015=>"111111111",
  32016=>"000000000",
  32017=>"000111111",
  32018=>"111001000",
  32019=>"111111111",
  32020=>"111110110",
  32021=>"111111011",
  32022=>"001000100",
  32023=>"111111110",
  32024=>"000000000",
  32025=>"000000000",
  32026=>"110000011",
  32027=>"111000000",
  32028=>"111001001",
  32029=>"000000000",
  32030=>"000000000",
  32031=>"111101111",
  32032=>"000110111",
  32033=>"000000010",
  32034=>"001101111",
  32035=>"111111111",
  32036=>"110000000",
  32037=>"111111111",
  32038=>"001101101",
  32039=>"000000111",
  32040=>"011011111",
  32041=>"000000000",
  32042=>"010010010",
  32043=>"111111110",
  32044=>"000001000",
  32045=>"000000000",
  32046=>"111000110",
  32047=>"111111010",
  32048=>"000000100",
  32049=>"000000000",
  32050=>"000000100",
  32051=>"000111000",
  32052=>"100100000",
  32053=>"111100111",
  32054=>"000000000",
  32055=>"111001011",
  32056=>"111111111",
  32057=>"010011111",
  32058=>"111111111",
  32059=>"100001000",
  32060=>"111111111",
  32061=>"000000101",
  32062=>"000010111",
  32063=>"000010000",
  32064=>"000111110",
  32065=>"111111000",
  32066=>"111111111",
  32067=>"111111110",
  32068=>"111111111",
  32069=>"001011111",
  32070=>"000111100",
  32071=>"111111011",
  32072=>"000000000",
  32073=>"000000000",
  32074=>"111111111",
  32075=>"111111100",
  32076=>"000000000",
  32077=>"111110111",
  32078=>"000001000",
  32079=>"110100000",
  32080=>"111111000",
  32081=>"000000000",
  32082=>"111111111",
  32083=>"111111111",
  32084=>"111000010",
  32085=>"011011011",
  32086=>"000000110",
  32087=>"110100000",
  32088=>"000001111",
  32089=>"111111111",
  32090=>"000010011",
  32091=>"001011110",
  32092=>"000000111",
  32093=>"100000000",
  32094=>"111111100",
  32095=>"110110111",
  32096=>"111000000",
  32097=>"000000000",
  32098=>"110100000",
  32099=>"000000000",
  32100=>"000000100",
  32101=>"111111111",
  32102=>"000000100",
  32103=>"000000101",
  32104=>"011111111",
  32105=>"111111111",
  32106=>"110111000",
  32107=>"111111110",
  32108=>"000000000",
  32109=>"000011001",
  32110=>"010000100",
  32111=>"000000011",
  32112=>"000000000",
  32113=>"000000000",
  32114=>"111001000",
  32115=>"110110111",
  32116=>"000000111",
  32117=>"111001000",
  32118=>"111111111",
  32119=>"000000011",
  32120=>"000000000",
  32121=>"000000111",
  32122=>"000000110",
  32123=>"110110110",
  32124=>"000000111",
  32125=>"000000000",
  32126=>"111000000",
  32127=>"001001111",
  32128=>"111111100",
  32129=>"111010110",
  32130=>"010000000",
  32131=>"100000011",
  32132=>"111111111",
  32133=>"001111111",
  32134=>"000000111",
  32135=>"111111000",
  32136=>"111111111",
  32137=>"111011001",
  32138=>"111101000",
  32139=>"101101111",
  32140=>"000101111",
  32141=>"000001011",
  32142=>"000001000",
  32143=>"111110100",
  32144=>"100111000",
  32145=>"000000000",
  32146=>"000000111",
  32147=>"111111110",
  32148=>"011001001",
  32149=>"010110000",
  32150=>"111111100",
  32151=>"000000100",
  32152=>"011111100",
  32153=>"000000010",
  32154=>"111111010",
  32155=>"000001000",
  32156=>"111111001",
  32157=>"111111111",
  32158=>"111111111",
  32159=>"110110000",
  32160=>"011111111",
  32161=>"000000011",
  32162=>"011000100",
  32163=>"000001111",
  32164=>"000111000",
  32165=>"111110001",
  32166=>"000000000",
  32167=>"001000000",
  32168=>"100011111",
  32169=>"000011000",
  32170=>"000001001",
  32171=>"111111001",
  32172=>"001000000",
  32173=>"001001000",
  32174=>"000000111",
  32175=>"111100101",
  32176=>"111111111",
  32177=>"111111111",
  32178=>"000000110",
  32179=>"110010000",
  32180=>"110111111",
  32181=>"111101000",
  32182=>"000110111",
  32183=>"000111111",
  32184=>"000001111",
  32185=>"111111001",
  32186=>"000000100",
  32187=>"000111111",
  32188=>"110110110",
  32189=>"000000000",
  32190=>"111111111",
  32191=>"111001011",
  32192=>"100111111",
  32193=>"111000101",
  32194=>"000000000",
  32195=>"000111010",
  32196=>"000000000",
  32197=>"110000100",
  32198=>"110010100",
  32199=>"101001000",
  32200=>"000001011",
  32201=>"111101000",
  32202=>"111111111",
  32203=>"000000000",
  32204=>"100110000",
  32205=>"000011111",
  32206=>"000111110",
  32207=>"111111111",
  32208=>"000000000",
  32209=>"111111111",
  32210=>"110110110",
  32211=>"101000000",
  32212=>"000000000",
  32213=>"000000010",
  32214=>"000000011",
  32215=>"100100100",
  32216=>"011000111",
  32217=>"110100101",
  32218=>"000000010",
  32219=>"110110100",
  32220=>"000111111",
  32221=>"111001111",
  32222=>"111111111",
  32223=>"100000000",
  32224=>"011010111",
  32225=>"000111111",
  32226=>"000000011",
  32227=>"111101100",
  32228=>"000111000",
  32229=>"001111000",
  32230=>"111111111",
  32231=>"000000000",
  32232=>"010000010",
  32233=>"101001100",
  32234=>"000011111",
  32235=>"111111111",
  32236=>"111111111",
  32237=>"000000000",
  32238=>"001000110",
  32239=>"111111011",
  32240=>"001000111",
  32241=>"111010110",
  32242=>"011111001",
  32243=>"111111111",
  32244=>"111111111",
  32245=>"101111111",
  32246=>"000000000",
  32247=>"110000111",
  32248=>"101101111",
  32249=>"100100100",
  32250=>"110110100",
  32251=>"111111110",
  32252=>"111111111",
  32253=>"111100100",
  32254=>"000000011",
  32255=>"111111101",
  32256=>"111000001",
  32257=>"000000010",
  32258=>"000001111",
  32259=>"000000000",
  32260=>"001000000",
  32261=>"000010000",
  32262=>"100000100",
  32263=>"111111111",
  32264=>"010000100",
  32265=>"110111000",
  32266=>"111111110",
  32267=>"111111111",
  32268=>"111110000",
  32269=>"111111110",
  32270=>"111111000",
  32271=>"000000000",
  32272=>"111011111",
  32273=>"111010000",
  32274=>"000111111",
  32275=>"000111111",
  32276=>"000000111",
  32277=>"000111111",
  32278=>"000000000",
  32279=>"000111111",
  32280=>"000000000",
  32281=>"101111110",
  32282=>"110000000",
  32283=>"101110000",
  32284=>"000000111",
  32285=>"100111111",
  32286=>"100110110",
  32287=>"100110111",
  32288=>"001000110",
  32289=>"111101001",
  32290=>"000000110",
  32291=>"111111011",
  32292=>"000111111",
  32293=>"011111111",
  32294=>"010000001",
  32295=>"010000000",
  32296=>"011111100",
  32297=>"000000000",
  32298=>"111000000",
  32299=>"110111111",
  32300=>"111111000",
  32301=>"111111011",
  32302=>"000111001",
  32303=>"111111111",
  32304=>"000000000",
  32305=>"110111110",
  32306=>"000000001",
  32307=>"111100000",
  32308=>"111000000",
  32309=>"000001111",
  32310=>"111111100",
  32311=>"011011111",
  32312=>"111000000",
  32313=>"111111000",
  32314=>"000000000",
  32315=>"111100111",
  32316=>"111101100",
  32317=>"110000011",
  32318=>"111101111",
  32319=>"001111001",
  32320=>"111100011",
  32321=>"000100000",
  32322=>"111111000",
  32323=>"111111001",
  32324=>"110110000",
  32325=>"111110111",
  32326=>"000000000",
  32327=>"111111100",
  32328=>"001001000",
  32329=>"000000111",
  32330=>"101000000",
  32331=>"111100001",
  32332=>"110110110",
  32333=>"101000111",
  32334=>"000000000",
  32335=>"001000000",
  32336=>"111001000",
  32337=>"111010000",
  32338=>"000000111",
  32339=>"111000000",
  32340=>"111110110",
  32341=>"000001011",
  32342=>"111001001",
  32343=>"100111111",
  32344=>"111111111",
  32345=>"000000000",
  32346=>"100111111",
  32347=>"001111000",
  32348=>"101001111",
  32349=>"010011000",
  32350=>"111000001",
  32351=>"110000010",
  32352=>"000000000",
  32353=>"000111000",
  32354=>"111100000",
  32355=>"000001110",
  32356=>"110000001",
  32357=>"000000100",
  32358=>"111111000",
  32359=>"111111101",
  32360=>"100000111",
  32361=>"100111111",
  32362=>"110000001",
  32363=>"111111111",
  32364=>"111001000",
  32365=>"000000001",
  32366=>"111000111",
  32367=>"000000011",
  32368=>"111111000",
  32369=>"111111000",
  32370=>"011011000",
  32371=>"000000101",
  32372=>"000000111",
  32373=>"001011000",
  32374=>"000000000",
  32375=>"000000000",
  32376=>"100100000",
  32377=>"000000001",
  32378=>"000000000",
  32379=>"000101001",
  32380=>"000101111",
  32381=>"000001111",
  32382=>"001011011",
  32383=>"110110010",
  32384=>"111111111",
  32385=>"111110010",
  32386=>"111000000",
  32387=>"000100000",
  32388=>"101111111",
  32389=>"111000111",
  32390=>"111111000",
  32391=>"000000000",
  32392=>"000111111",
  32393=>"000000000",
  32394=>"111000000",
  32395=>"000000100",
  32396=>"111000000",
  32397=>"100111111",
  32398=>"000101111",
  32399=>"000000000",
  32400=>"111111000",
  32401=>"010000000",
  32402=>"001000010",
  32403=>"100000000",
  32404=>"111111001",
  32405=>"111111000",
  32406=>"000000010",
  32407=>"000000000",
  32408=>"000111111",
  32409=>"111111111",
  32410=>"000001011",
  32411=>"000010001",
  32412=>"111001000",
  32413=>"000000000",
  32414=>"111100000",
  32415=>"111111000",
  32416=>"100000111",
  32417=>"001111101",
  32418=>"111111000",
  32419=>"111000100",
  32420=>"111100110",
  32421=>"100111111",
  32422=>"010111110",
  32423=>"101000000",
  32424=>"111011011",
  32425=>"111011000",
  32426=>"111110000",
  32427=>"111111100",
  32428=>"111000000",
  32429=>"111011001",
  32430=>"111000111",
  32431=>"010100111",
  32432=>"111100000",
  32433=>"111101001",
  32434=>"111111110",
  32435=>"110111011",
  32436=>"100100111",
  32437=>"000001011",
  32438=>"110110000",
  32439=>"111000010",
  32440=>"111111101",
  32441=>"001011111",
  32442=>"111101101",
  32443=>"000000010",
  32444=>"111000000",
  32445=>"000000001",
  32446=>"000111111",
  32447=>"000001101",
  32448=>"000000011",
  32449=>"111111000",
  32450=>"000000010",
  32451=>"111111111",
  32452=>"000000011",
  32453=>"000111111",
  32454=>"001000000",
  32455=>"111000000",
  32456=>"111000010",
  32457=>"110111000",
  32458=>"000111110",
  32459=>"000000001",
  32460=>"111000000",
  32461=>"111111000",
  32462=>"111000000",
  32463=>"111000010",
  32464=>"100000000",
  32465=>"010000100",
  32466=>"111010000",
  32467=>"111011001",
  32468=>"001100100",
  32469=>"000001000",
  32470=>"000000011",
  32471=>"001000000",
  32472=>"000001000",
  32473=>"000111111",
  32474=>"000000000",
  32475=>"000010111",
  32476=>"111110000",
  32477=>"000111111",
  32478=>"001000000",
  32479=>"101000001",
  32480=>"011000000",
  32481=>"000000010",
  32482=>"110111000",
  32483=>"111011111",
  32484=>"110111111",
  32485=>"100100100",
  32486=>"111111000",
  32487=>"000000000",
  32488=>"000000100",
  32489=>"110100000",
  32490=>"111111001",
  32491=>"111100000",
  32492=>"100000000",
  32493=>"000000000",
  32494=>"111100000",
  32495=>"000000000",
  32496=>"000011111",
  32497=>"011000000",
  32498=>"111111100",
  32499=>"111111001",
  32500=>"000000001",
  32501=>"111000000",
  32502=>"110110110",
  32503=>"000000000",
  32504=>"110010000",
  32505=>"110000000",
  32506=>"000000111",
  32507=>"000000011",
  32508=>"000100110",
  32509=>"111111111",
  32510=>"100000000",
  32511=>"000111111",
  32512=>"000001011",
  32513=>"001001001",
  32514=>"100111000",
  32515=>"000000000",
  32516=>"000001111",
  32517=>"000111111",
  32518=>"111000000",
  32519=>"101100000",
  32520=>"000011000",
  32521=>"000111111",
  32522=>"000000011",
  32523=>"000000111",
  32524=>"110000000",
  32525=>"111111000",
  32526=>"000011011",
  32527=>"111111000",
  32528=>"000111110",
  32529=>"000000000",
  32530=>"000000000",
  32531=>"111000011",
  32532=>"000111111",
  32533=>"000000000",
  32534=>"000111111",
  32535=>"000000111",
  32536=>"011111111",
  32537=>"000000001",
  32538=>"111111110",
  32539=>"000011111",
  32540=>"000000000",
  32541=>"000000111",
  32542=>"111111011",
  32543=>"111111000",
  32544=>"110111001",
  32545=>"110111111",
  32546=>"100111111",
  32547=>"101001001",
  32548=>"000011111",
  32549=>"000000001",
  32550=>"000111010",
  32551=>"000101111",
  32552=>"110111111",
  32553=>"111111111",
  32554=>"000000000",
  32555=>"111000000",
  32556=>"000000000",
  32557=>"000110100",
  32558=>"001000110",
  32559=>"000000000",
  32560=>"111111001",
  32561=>"000000001",
  32562=>"000011000",
  32563=>"111111110",
  32564=>"000000000",
  32565=>"010000100",
  32566=>"000000011",
  32567=>"000000000",
  32568=>"000000000",
  32569=>"011011011",
  32570=>"111000110",
  32571=>"010000000",
  32572=>"000111111",
  32573=>"111100000",
  32574=>"000111111",
  32575=>"000000111",
  32576=>"111000000",
  32577=>"101111100",
  32578=>"000000001",
  32579=>"000101111",
  32580=>"111011100",
  32581=>"000110111",
  32582=>"000000000",
  32583=>"100100000",
  32584=>"111000000",
  32585=>"000000000",
  32586=>"001000111",
  32587=>"100110000",
  32588=>"001000010",
  32589=>"100000000",
  32590=>"111011000",
  32591=>"000000111",
  32592=>"110110110",
  32593=>"000111111",
  32594=>"111000000",
  32595=>"101000000",
  32596=>"101111110",
  32597=>"001000111",
  32598=>"111111011",
  32599=>"110000000",
  32600=>"001111111",
  32601=>"111001000",
  32602=>"001000000",
  32603=>"000011011",
  32604=>"000000000",
  32605=>"111111001",
  32606=>"000000111",
  32607=>"001111000",
  32608=>"110111111",
  32609=>"111111000",
  32610=>"001110000",
  32611=>"000001000",
  32612=>"000100100",
  32613=>"000000000",
  32614=>"110111111",
  32615=>"111101001",
  32616=>"111111110",
  32617=>"000000000",
  32618=>"110111111",
  32619=>"001000001",
  32620=>"111100000",
  32621=>"111000000",
  32622=>"000000100",
  32623=>"000100111",
  32624=>"111111000",
  32625=>"010111111",
  32626=>"000111111",
  32627=>"100100100",
  32628=>"111100000",
  32629=>"000000000",
  32630=>"101000100",
  32631=>"110111111",
  32632=>"000011001",
  32633=>"000000100",
  32634=>"000000110",
  32635=>"111011111",
  32636=>"001001001",
  32637=>"001000000",
  32638=>"111111111",
  32639=>"111100100",
  32640=>"001001000",
  32641=>"000001101",
  32642=>"111011111",
  32643=>"000011011",
  32644=>"100100110",
  32645=>"011011001",
  32646=>"000111111",
  32647=>"111000000",
  32648=>"110000000",
  32649=>"111100111",
  32650=>"100111111",
  32651=>"000001011",
  32652=>"111111111",
  32653=>"110111111",
  32654=>"100110000",
  32655=>"000000011",
  32656=>"111000000",
  32657=>"111001001",
  32658=>"110111000",
  32659=>"000110110",
  32660=>"000000110",
  32661=>"000001000",
  32662=>"100111111",
  32663=>"111100100",
  32664=>"000000000",
  32665=>"111000000",
  32666=>"000111101",
  32667=>"100101000",
  32668=>"000000110",
  32669=>"000010011",
  32670=>"001000011",
  32671=>"111111001",
  32672=>"011001110",
  32673=>"000001111",
  32674=>"000000000",
  32675=>"111111111",
  32676=>"111111111",
  32677=>"000000000",
  32678=>"111100111",
  32679=>"111111111",
  32680=>"001000000",
  32681=>"000011000",
  32682=>"111000111",
  32683=>"000000000",
  32684=>"000000110",
  32685=>"100000000",
  32686=>"111000101",
  32687=>"110100100",
  32688=>"111010000",
  32689=>"000111111",
  32690=>"001001100",
  32691=>"011011111",
  32692=>"000000000",
  32693=>"100110110",
  32694=>"111111111",
  32695=>"101000000",
  32696=>"000000000",
  32697=>"111010000",
  32698=>"111000000",
  32699=>"011001000",
  32700=>"000000011",
  32701=>"001111111",
  32702=>"000011111",
  32703=>"011001001",
  32704=>"011011000",
  32705=>"111001111",
  32706=>"000000000",
  32707=>"111111111",
  32708=>"111000001",
  32709=>"100000000",
  32710=>"000000001",
  32711=>"000000000",
  32712=>"100001001",
  32713=>"111111111",
  32714=>"000000000",
  32715=>"000000000",
  32716=>"111100000",
  32717=>"100000000",
  32718=>"111110000",
  32719=>"000111111",
  32720=>"000111111",
  32721=>"110100100",
  32722=>"111000000",
  32723=>"000000111",
  32724=>"100100011",
  32725=>"111001100",
  32726=>"000000000",
  32727=>"011000000",
  32728=>"000000000",
  32729=>"000000000",
  32730=>"100000000",
  32731=>"100100110",
  32732=>"000100000",
  32733=>"000000111",
  32734=>"111111000",
  32735=>"100111000",
  32736=>"111010010",
  32737=>"111000111",
  32738=>"000000000",
  32739=>"111111011",
  32740=>"111111110",
  32741=>"111000000",
  32742=>"101111111",
  32743=>"000000111",
  32744=>"111000001",
  32745=>"000000101",
  32746=>"000000000",
  32747=>"100100000",
  32748=>"111000000",
  32749=>"111111000",
  32750=>"111110011",
  32751=>"011010000",
  32752=>"000000000",
  32753=>"000001000",
  32754=>"011000101",
  32755=>"111000000",
  32756=>"111011111",
  32757=>"000000111",
  32758=>"100000110",
  32759=>"000100111",
  32760=>"111000000",
  32761=>"000111010",
  32762=>"111000000",
  32763=>"000001111",
  32764=>"011010111",
  32765=>"001000000",
  32766=>"000000000",
  32767=>"001111111",
  32768=>"001000000",
  32769=>"011111001",
  32770=>"000010111",
  32771=>"011010111",
  32772=>"000000111",
  32773=>"111000000",
  32774=>"000000000",
  32775=>"000000000",
  32776=>"111111111",
  32777=>"011000000",
  32778=>"111111111",
  32779=>"000100000",
  32780=>"000000000",
  32781=>"000000011",
  32782=>"001111111",
  32783=>"000000000",
  32784=>"000000000",
  32785=>"000000000",
  32786=>"000000000",
  32787=>"111111111",
  32788=>"000000100",
  32789=>"111111110",
  32790=>"000101111",
  32791=>"111111000",
  32792=>"000000101",
  32793=>"000001011",
  32794=>"000110111",
  32795=>"110100100",
  32796=>"111111111",
  32797=>"000000000",
  32798=>"001000000",
  32799=>"000000000",
  32800=>"111100100",
  32801=>"111111111",
  32802=>"001001000",
  32803=>"111111111",
  32804=>"111110111",
  32805=>"000000001",
  32806=>"111111111",
  32807=>"000111111",
  32808=>"101000000",
  32809=>"111111111",
  32810=>"111101000",
  32811=>"000000001",
  32812=>"111111111",
  32813=>"000000000",
  32814=>"111111111",
  32815=>"110110000",
  32816=>"001011111",
  32817=>"100100000",
  32818=>"111111101",
  32819=>"011100100",
  32820=>"000000001",
  32821=>"011011000",
  32822=>"100101111",
  32823=>"000000011",
  32824=>"111111111",
  32825=>"000000000",
  32826=>"000000101",
  32827=>"000000000",
  32828=>"111001011",
  32829=>"000000000",
  32830=>"111111111",
  32831=>"111100100",
  32832=>"111111111",
  32833=>"001000000",
  32834=>"000000111",
  32835=>"000000000",
  32836=>"011111011",
  32837=>"100100110",
  32838=>"111001000",
  32839=>"000100100",
  32840=>"011111001",
  32841=>"110100111",
  32842=>"000000000",
  32843=>"000000000",
  32844=>"000000001",
  32845=>"000000010",
  32846=>"000000000",
  32847=>"000100111",
  32848=>"000000000",
  32849=>"100111100",
  32850=>"001001111",
  32851=>"110100111",
  32852=>"001111111",
  32853=>"000110111",
  32854=>"111111000",
  32855=>"111111111",
  32856=>"000001111",
  32857=>"000000000",
  32858=>"000010000",
  32859=>"110111110",
  32860=>"001001000",
  32861=>"000000000",
  32862=>"111111111",
  32863=>"000000000",
  32864=>"000000000",
  32865=>"001000000",
  32866=>"110111001",
  32867=>"000000111",
  32868=>"111000111",
  32869=>"001111111",
  32870=>"000000000",
  32871=>"000111111",
  32872=>"000000000",
  32873=>"111000000",
  32874=>"110110011",
  32875=>"100100000",
  32876=>"011011111",
  32877=>"000000000",
  32878=>"000000000",
  32879=>"000000111",
  32880=>"111111111",
  32881=>"000000000",
  32882=>"111111111",
  32883=>"000110100",
  32884=>"111111111",
  32885=>"000000111",
  32886=>"111111100",
  32887=>"111111100",
  32888=>"000100111",
  32889=>"000000000",
  32890=>"000000000",
  32891=>"000000000",
  32892=>"000000000",
  32893=>"000011010",
  32894=>"000000000",
  32895=>"001100100",
  32896=>"111111111",
  32897=>"000000000",
  32898=>"000000000",
  32899=>"111111111",
  32900=>"000000000",
  32901=>"000000000",
  32902=>"000000110",
  32903=>"110000000",
  32904=>"111111111",
  32905=>"111111111",
  32906=>"000000111",
  32907=>"111111111",
  32908=>"100000000",
  32909=>"000000111",
  32910=>"111111000",
  32911=>"111101000",
  32912=>"000000000",
  32913=>"111111111",
  32914=>"100001000",
  32915=>"000000000",
  32916=>"111010000",
  32917=>"011011111",
  32918=>"000000000",
  32919=>"111111111",
  32920=>"001101101",
  32921=>"100110111",
  32922=>"000111111",
  32923=>"101100111",
  32924=>"001011111",
  32925=>"111111111",
  32926=>"000000000",
  32927=>"111111011",
  32928=>"111111000",
  32929=>"111011001",
  32930=>"111001111",
  32931=>"111011111",
  32932=>"110110111",
  32933=>"000000011",
  32934=>"111111111",
  32935=>"000000001",
  32936=>"000001111",
  32937=>"000000000",
  32938=>"000000000",
  32939=>"011000000",
  32940=>"010000000",
  32941=>"100110000",
  32942=>"111111111",
  32943=>"000000000",
  32944=>"000000000",
  32945=>"111111111",
  32946=>"111111111",
  32947=>"111111111",
  32948=>"110111111",
  32949=>"000001000",
  32950=>"111111110",
  32951=>"111000001",
  32952=>"000011111",
  32953=>"100010000",
  32954=>"000000000",
  32955=>"010000000",
  32956=>"111111011",
  32957=>"000000000",
  32958=>"000000101",
  32959=>"000000000",
  32960=>"111111111",
  32961=>"000001111",
  32962=>"010000000",
  32963=>"111111101",
  32964=>"000000000",
  32965=>"000000110",
  32966=>"111011111",
  32967=>"111111111",
  32968=>"010111111",
  32969=>"111111110",
  32970=>"000000000",
  32971=>"111101101",
  32972=>"111111000",
  32973=>"000000000",
  32974=>"100111111",
  32975=>"000000000",
  32976=>"011111111",
  32977=>"101100000",
  32978=>"000000111",
  32979=>"000000000",
  32980=>"000110110",
  32981=>"000000001",
  32982=>"111011001",
  32983=>"101100101",
  32984=>"110000000",
  32985=>"011011111",
  32986=>"111100000",
  32987=>"000000110",
  32988=>"111111111",
  32989=>"111110111",
  32990=>"100000000",
  32991=>"000100110",
  32992=>"001111111",
  32993=>"111111111",
  32994=>"000000000",
  32995=>"000010111",
  32996=>"011001101",
  32997=>"111111011",
  32998=>"000000011",
  32999=>"111111101",
  33000=>"011001111",
  33001=>"001111111",
  33002=>"111111111",
  33003=>"000000000",
  33004=>"000000000",
  33005=>"000000000",
  33006=>"000000000",
  33007=>"111000000",
  33008=>"100000011",
  33009=>"000000101",
  33010=>"100000010",
  33011=>"011001001",
  33012=>"110111011",
  33013=>"110110000",
  33014=>"000000110",
  33015=>"100111111",
  33016=>"000000001",
  33017=>"000000000",
  33018=>"000111111",
  33019=>"100001001",
  33020=>"100100000",
  33021=>"111100000",
  33022=>"111110000",
  33023=>"111111111",
  33024=>"000000001",
  33025=>"111110100",
  33026=>"011011001",
  33027=>"000000000",
  33028=>"100100100",
  33029=>"111000001",
  33030=>"000000111",
  33031=>"101101100",
  33032=>"111111101",
  33033=>"111010000",
  33034=>"000111100",
  33035=>"001100111",
  33036=>"000000100",
  33037=>"110010000",
  33038=>"000000001",
  33039=>"110100100",
  33040=>"000000000",
  33041=>"111111001",
  33042=>"111111010",
  33043=>"111011000",
  33044=>"111111101",
  33045=>"000000000",
  33046=>"000000100",
  33047=>"111001000",
  33048=>"100000000",
  33049=>"001001111",
  33050=>"111111111",
  33051=>"001000000",
  33052=>"111111111",
  33053=>"100000000",
  33054=>"000000000",
  33055=>"111111001",
  33056=>"111100000",
  33057=>"011110111",
  33058=>"101111000",
  33059=>"000000000",
  33060=>"001001001",
  33061=>"111111111",
  33062=>"111111111",
  33063=>"111111111",
  33064=>"111110111",
  33065=>"000000000",
  33066=>"011000000",
  33067=>"111111110",
  33068=>"001001000",
  33069=>"110111111",
  33070=>"000000110",
  33071=>"000000001",
  33072=>"000001001",
  33073=>"111000000",
  33074=>"111111111",
  33075=>"100000000",
  33076=>"111111111",
  33077=>"001111101",
  33078=>"111101011",
  33079=>"000111111",
  33080=>"000000000",
  33081=>"111111111",
  33082=>"010111000",
  33083=>"000000000",
  33084=>"000000000",
  33085=>"110110111",
  33086=>"000000000",
  33087=>"111111111",
  33088=>"110111111",
  33089=>"100111111",
  33090=>"111111111",
  33091=>"111111111",
  33092=>"000011111",
  33093=>"111111111",
  33094=>"000000001",
  33095=>"111111111",
  33096=>"111101111",
  33097=>"111111111",
  33098=>"111111111",
  33099=>"011100111",
  33100=>"000011001",
  33101=>"000000011",
  33102=>"111000000",
  33103=>"011011011",
  33104=>"000001010",
  33105=>"000000000",
  33106=>"000000000",
  33107=>"001000000",
  33108=>"000000000",
  33109=>"110110111",
  33110=>"110111111",
  33111=>"111111111",
  33112=>"111111111",
  33113=>"000000000",
  33114=>"000111011",
  33115=>"101111000",
  33116=>"000000000",
  33117=>"000000001",
  33118=>"010111111",
  33119=>"000000001",
  33120=>"001101111",
  33121=>"000001111",
  33122=>"001001000",
  33123=>"111111001",
  33124=>"000000110",
  33125=>"111001000",
  33126=>"111001101",
  33127=>"111111111",
  33128=>"000011000",
  33129=>"100000000",
  33130=>"111111111",
  33131=>"111111111",
  33132=>"011001001",
  33133=>"000011001",
  33134=>"111111111",
  33135=>"101101101",
  33136=>"011111111",
  33137=>"111111111",
  33138=>"111111111",
  33139=>"100110100",
  33140=>"111111011",
  33141=>"000000001",
  33142=>"111010000",
  33143=>"100111111",
  33144=>"111011010",
  33145=>"000000000",
  33146=>"000000101",
  33147=>"110000000",
  33148=>"111110000",
  33149=>"111000000",
  33150=>"011001001",
  33151=>"000000001",
  33152=>"111111111",
  33153=>"000000000",
  33154=>"001011011",
  33155=>"000000000",
  33156=>"000000000",
  33157=>"111111111",
  33158=>"111111000",
  33159=>"011111111",
  33160=>"111110111",
  33161=>"010010100",
  33162=>"001000000",
  33163=>"111111111",
  33164=>"110000000",
  33165=>"110111100",
  33166=>"000111100",
  33167=>"010110010",
  33168=>"000000000",
  33169=>"111100010",
  33170=>"001001111",
  33171=>"000000000",
  33172=>"100000000",
  33173=>"100110000",
  33174=>"111011111",
  33175=>"000110000",
  33176=>"000000000",
  33177=>"111110111",
  33178=>"000100111",
  33179=>"000000000",
  33180=>"111110100",
  33181=>"000000001",
  33182=>"100100000",
  33183=>"100110000",
  33184=>"011111000",
  33185=>"000110110",
  33186=>"111010000",
  33187=>"000000000",
  33188=>"000000000",
  33189=>"111110010",
  33190=>"000000000",
  33191=>"111111111",
  33192=>"100101111",
  33193=>"000101111",
  33194=>"000000000",
  33195=>"010010111",
  33196=>"000000000",
  33197=>"110110111",
  33198=>"111111111",
  33199=>"001001111",
  33200=>"111111111",
  33201=>"000000000",
  33202=>"001111111",
  33203=>"111111111",
  33204=>"000000000",
  33205=>"011001101",
  33206=>"001111001",
  33207=>"011010111",
  33208=>"000000000",
  33209=>"011001000",
  33210=>"000000000",
  33211=>"111111111",
  33212=>"110110110",
  33213=>"111000001",
  33214=>"001000100",
  33215=>"111000000",
  33216=>"000000110",
  33217=>"110111111",
  33218=>"111111111",
  33219=>"000010000",
  33220=>"111110111",
  33221=>"000000001",
  33222=>"000000000",
  33223=>"111111000",
  33224=>"111111111",
  33225=>"111111000",
  33226=>"000000000",
  33227=>"010011000",
  33228=>"000000000",
  33229=>"000000000",
  33230=>"000000000",
  33231=>"000010111",
  33232=>"000000000",
  33233=>"010000001",
  33234=>"000000000",
  33235=>"111111111",
  33236=>"100111111",
  33237=>"111111110",
  33238=>"111101000",
  33239=>"100000000",
  33240=>"111111111",
  33241=>"011110110",
  33242=>"011000001",
  33243=>"111111111",
  33244=>"011000000",
  33245=>"000000111",
  33246=>"000110111",
  33247=>"010000000",
  33248=>"111111111",
  33249=>"111111111",
  33250=>"100000000",
  33251=>"000000000",
  33252=>"111000000",
  33253=>"000001001",
  33254=>"000110110",
  33255=>"000000000",
  33256=>"111111111",
  33257=>"111111111",
  33258=>"000000000",
  33259=>"000000001",
  33260=>"000001011",
  33261=>"001101011",
  33262=>"110111111",
  33263=>"100110111",
  33264=>"000000001",
  33265=>"000000000",
  33266=>"111111111",
  33267=>"101111100",
  33268=>"000001001",
  33269=>"000000011",
  33270=>"111111001",
  33271=>"000111111",
  33272=>"111111111",
  33273=>"000001000",
  33274=>"001001111",
  33275=>"010110011",
  33276=>"111111111",
  33277=>"100110110",
  33278=>"111111001",
  33279=>"000000011",
  33280=>"011110110",
  33281=>"110111111",
  33282=>"111111110",
  33283=>"101111110",
  33284=>"110110000",
  33285=>"001000000",
  33286=>"111111010",
  33287=>"000001111",
  33288=>"111000100",
  33289=>"110110111",
  33290=>"101001001",
  33291=>"000110110",
  33292=>"100110100",
  33293=>"000000000",
  33294=>"100100111",
  33295=>"111011010",
  33296=>"000000000",
  33297=>"111111110",
  33298=>"000000000",
  33299=>"111111111",
  33300=>"111111111",
  33301=>"010000000",
  33302=>"101001001",
  33303=>"001000000",
  33304=>"101101100",
  33305=>"011001000",
  33306=>"000000000",
  33307=>"100100100",
  33308=>"111111111",
  33309=>"111000000",
  33310=>"111000000",
  33311=>"111011011",
  33312=>"111111111",
  33313=>"111111001",
  33314=>"001000101",
  33315=>"101101111",
  33316=>"111111111",
  33317=>"100001101",
  33318=>"000001111",
  33319=>"000000000",
  33320=>"000000000",
  33321=>"000000000",
  33322=>"000000000",
  33323=>"110110000",
  33324=>"001000000",
  33325=>"000111000",
  33326=>"001001101",
  33327=>"001001111",
  33328=>"000010000",
  33329=>"111111011",
  33330=>"100111111",
  33331=>"000001001",
  33332=>"001011000",
  33333=>"110110010",
  33334=>"000000101",
  33335=>"000000000",
  33336=>"000100000",
  33337=>"000000000",
  33338=>"110110010",
  33339=>"111111111",
  33340=>"100000000",
  33341=>"010111010",
  33342=>"111111111",
  33343=>"110000000",
  33344=>"011001001",
  33345=>"000010000",
  33346=>"000111111",
  33347=>"000000000",
  33348=>"110110110",
  33349=>"000000000",
  33350=>"000000000",
  33351=>"001001001",
  33352=>"011111111",
  33353=>"000000111",
  33354=>"111111010",
  33355=>"001000000",
  33356=>"000110111",
  33357=>"000010000",
  33358=>"110110110",
  33359=>"000100100",
  33360=>"101000001",
  33361=>"011010000",
  33362=>"000001111",
  33363=>"110110000",
  33364=>"011011000",
  33365=>"000000000",
  33366=>"000000000",
  33367=>"011111110",
  33368=>"000110010",
  33369=>"000001111",
  33370=>"000100110",
  33371=>"110110110",
  33372=>"000000000",
  33373=>"000000000",
  33374=>"000000001",
  33375=>"101001001",
  33376=>"000111111",
  33377=>"101011000",
  33378=>"000000000",
  33379=>"000000110",
  33380=>"100000000",
  33381=>"000000111",
  33382=>"000000110",
  33383=>"111100000",
  33384=>"100011000",
  33385=>"000101111",
  33386=>"111111010",
  33387=>"000010010",
  33388=>"110111100",
  33389=>"111111111",
  33390=>"101111111",
  33391=>"010010011",
  33392=>"111010110",
  33393=>"001001101",
  33394=>"111111000",
  33395=>"000000111",
  33396=>"000000000",
  33397=>"111111110",
  33398=>"000000000",
  33399=>"111111111",
  33400=>"000000111",
  33401=>"101111000",
  33402=>"100101100",
  33403=>"001000000",
  33404=>"111111100",
  33405=>"111111111",
  33406=>"000000000",
  33407=>"111110000",
  33408=>"111111111",
  33409=>"111111110",
  33410=>"000001111",
  33411=>"011111000",
  33412=>"110000100",
  33413=>"111101101",
  33414=>"101100100",
  33415=>"000001000",
  33416=>"010010010",
  33417=>"001001111",
  33418=>"000000000",
  33419=>"100000000",
  33420=>"001001111",
  33421=>"000000001",
  33422=>"100000000",
  33423=>"111111110",
  33424=>"101101111",
  33425=>"011011000",
  33426=>"010111111",
  33427=>"100100111",
  33428=>"010000000",
  33429=>"111110010",
  33430=>"000011001",
  33431=>"001001000",
  33432=>"000000100",
  33433=>"100111111",
  33434=>"111000000",
  33435=>"000000000",
  33436=>"100000001",
  33437=>"011001001",
  33438=>"100000001",
  33439=>"111111000",
  33440=>"111111011",
  33441=>"100111100",
  33442=>"000110010",
  33443=>"110100111",
  33444=>"000100100",
  33445=>"001001101",
  33446=>"111111101",
  33447=>"111100000",
  33448=>"000000101",
  33449=>"000000001",
  33450=>"111001001",
  33451=>"000000000",
  33452=>"101101000",
  33453=>"000010010",
  33454=>"001000000",
  33455=>"000001111",
  33456=>"000111000",
  33457=>"111111001",
  33458=>"111111110",
  33459=>"101101000",
  33460=>"111000001",
  33461=>"000000000",
  33462=>"000011010",
  33463=>"000000000",
  33464=>"001000101",
  33465=>"111111111",
  33466=>"101001001",
  33467=>"000000000",
  33468=>"000000111",
  33469=>"111111111",
  33470=>"000000111",
  33471=>"000000000",
  33472=>"010010100",
  33473=>"111111111",
  33474=>"111111111",
  33475=>"000000111",
  33476=>"000101111",
  33477=>"000100010",
  33478=>"110110000",
  33479=>"000000000",
  33480=>"000000001",
  33481=>"101001001",
  33482=>"000000001",
  33483=>"111000000",
  33484=>"000100100",
  33485=>"000000000",
  33486=>"000111111",
  33487=>"000111001",
  33488=>"100000000",
  33489=>"101000111",
  33490=>"110000001",
  33491=>"101001101",
  33492=>"111000000",
  33493=>"000000000",
  33494=>"110110110",
  33495=>"111110110",
  33496=>"110100110",
  33497=>"000110111",
  33498=>"111011011",
  33499=>"111111000",
  33500=>"110100000",
  33501=>"000100111",
  33502=>"111111010",
  33503=>"001001001",
  33504=>"000000110",
  33505=>"000000000",
  33506=>"111111010",
  33507=>"000000001",
  33508=>"111111111",
  33509=>"101111111",
  33510=>"000000101",
  33511=>"100111111",
  33512=>"000000111",
  33513=>"001001100",
  33514=>"110110010",
  33515=>"110111100",
  33516=>"111111001",
  33517=>"000101000",
  33518=>"000000000",
  33519=>"000000111",
  33520=>"101111111",
  33521=>"000000001",
  33522=>"101101001",
  33523=>"000000000",
  33524=>"111111011",
  33525=>"000100110",
  33526=>"010111010",
  33527=>"000110111",
  33528=>"010110110",
  33529=>"111111111",
  33530=>"000010000",
  33531=>"100100110",
  33532=>"001011011",
  33533=>"000000001",
  33534=>"011000000",
  33535=>"111100110",
  33536=>"000000001",
  33537=>"000001011",
  33538=>"000000101",
  33539=>"000001001",
  33540=>"111111110",
  33541=>"111100111",
  33542=>"000000111",
  33543=>"001001001",
  33544=>"100110010",
  33545=>"110000000",
  33546=>"000001101",
  33547=>"110111010",
  33548=>"000000100",
  33549=>"111001101",
  33550=>"010110011",
  33551=>"111111111",
  33552=>"111110011",
  33553=>"001000001",
  33554=>"111001000",
  33555=>"101110111",
  33556=>"111100101",
  33557=>"111111111",
  33558=>"100110000",
  33559=>"101111110",
  33560=>"111111000",
  33561=>"000111101",
  33562=>"111111010",
  33563=>"111000000",
  33564=>"001001011",
  33565=>"000000000",
  33566=>"001000000",
  33567=>"001011111",
  33568=>"100000000",
  33569=>"000000000",
  33570=>"010110111",
  33571=>"111111010",
  33572=>"110101101",
  33573=>"111111111",
  33574=>"000000000",
  33575=>"111111111",
  33576=>"110001101",
  33577=>"110000000",
  33578=>"011111110",
  33579=>"011011010",
  33580=>"000000000",
  33581=>"010010010",
  33582=>"111000111",
  33583=>"110000010",
  33584=>"110110110",
  33585=>"000000000",
  33586=>"110111111",
  33587=>"111110000",
  33588=>"000000011",
  33589=>"000000001",
  33590=>"001011000",
  33591=>"000000101",
  33592=>"010010000",
  33593=>"101000101",
  33594=>"111111111",
  33595=>"111111000",
  33596=>"000001111",
  33597=>"000000000",
  33598=>"111111111",
  33599=>"111111111",
  33600=>"000000000",
  33601=>"111111011",
  33602=>"001011011",
  33603=>"000001111",
  33604=>"000000110",
  33605=>"000000100",
  33606=>"111000000",
  33607=>"001011111",
  33608=>"000000000",
  33609=>"000000111",
  33610=>"000000001",
  33611=>"011011000",
  33612=>"111000010",
  33613=>"001000000",
  33614=>"110111111",
  33615=>"111100000",
  33616=>"111010000",
  33617=>"100000001",
  33618=>"001001000",
  33619=>"000000101",
  33620=>"000110111",
  33621=>"001001000",
  33622=>"010110000",
  33623=>"111011000",
  33624=>"011111111",
  33625=>"001111111",
  33626=>"011000000",
  33627=>"000000001",
  33628=>"000110110",
  33629=>"010011110",
  33630=>"010000000",
  33631=>"000001101",
  33632=>"111001000",
  33633=>"000000000",
  33634=>"111001000",
  33635=>"000000000",
  33636=>"001001000",
  33637=>"011110000",
  33638=>"000010010",
  33639=>"000000000",
  33640=>"111011000",
  33641=>"110000011",
  33642=>"100000000",
  33643=>"110110010",
  33644=>"110110110",
  33645=>"000001111",
  33646=>"111111111",
  33647=>"001001101",
  33648=>"111111111",
  33649=>"001000000",
  33650=>"010111111",
  33651=>"100100000",
  33652=>"000110000",
  33653=>"101001101",
  33654=>"000000000",
  33655=>"111110000",
  33656=>"000000001",
  33657=>"111110010",
  33658=>"101001111",
  33659=>"000000000",
  33660=>"100100111",
  33661=>"111111111",
  33662=>"111011000",
  33663=>"000000101",
  33664=>"110010000",
  33665=>"100110111",
  33666=>"110001000",
  33667=>"111101111",
  33668=>"111110111",
  33669=>"000001111",
  33670=>"111111100",
  33671=>"111101001",
  33672=>"000000010",
  33673=>"000000010",
  33674=>"000101111",
  33675=>"000100100",
  33676=>"000110111",
  33677=>"110100000",
  33678=>"000000010",
  33679=>"110110000",
  33680=>"011001001",
  33681=>"111111111",
  33682=>"111111110",
  33683=>"000111111",
  33684=>"000000000",
  33685=>"010010000",
  33686=>"000000000",
  33687=>"110110000",
  33688=>"111100000",
  33689=>"000100100",
  33690=>"010010010",
  33691=>"110110010",
  33692=>"000010110",
  33693=>"010110110",
  33694=>"111101001",
  33695=>"111111111",
  33696=>"100000000",
  33697=>"111011001",
  33698=>"000000000",
  33699=>"100000000",
  33700=>"111101111",
  33701=>"000010010",
  33702=>"000010111",
  33703=>"000000000",
  33704=>"001001000",
  33705=>"001001000",
  33706=>"010110111",
  33707=>"001011000",
  33708=>"011001111",
  33709=>"000000101",
  33710=>"000111111",
  33711=>"110111110",
  33712=>"000000111",
  33713=>"000000000",
  33714=>"000000000",
  33715=>"010000000",
  33716=>"001000101",
  33717=>"000000000",
  33718=>"111111111",
  33719=>"111111000",
  33720=>"111000000",
  33721=>"000010111",
  33722=>"111100000",
  33723=>"111111111",
  33724=>"000000000",
  33725=>"101000000",
  33726=>"111011010",
  33727=>"110110000",
  33728=>"000000001",
  33729=>"000110111",
  33730=>"000110111",
  33731=>"001000011",
  33732=>"110110010",
  33733=>"100100000",
  33734=>"010010000",
  33735=>"011111100",
  33736=>"111001000",
  33737=>"111111111",
  33738=>"001001111",
  33739=>"000001001",
  33740=>"010010000",
  33741=>"111111111",
  33742=>"101000111",
  33743=>"110010000",
  33744=>"100110000",
  33745=>"110110010",
  33746=>"000100111",
  33747=>"100110010",
  33748=>"000000001",
  33749=>"000000000",
  33750=>"111111111",
  33751=>"011011010",
  33752=>"000001111",
  33753=>"000001001",
  33754=>"111000111",
  33755=>"111001101",
  33756=>"000000000",
  33757=>"111111110",
  33758=>"111011101",
  33759=>"100100000",
  33760=>"000011000",
  33761=>"010110110",
  33762=>"011000001",
  33763=>"110110010",
  33764=>"111010110",
  33765=>"000111111",
  33766=>"111011000",
  33767=>"000000000",
  33768=>"110111010",
  33769=>"111111001",
  33770=>"000000000",
  33771=>"111111111",
  33772=>"111111111",
  33773=>"011111000",
  33774=>"001000000",
  33775=>"111000001",
  33776=>"101001000",
  33777=>"000000101",
  33778=>"101001101",
  33779=>"011000010",
  33780=>"100000101",
  33781=>"111111000",
  33782=>"110111111",
  33783=>"000000000",
  33784=>"000010010",
  33785=>"111111000",
  33786=>"111000000",
  33787=>"000000000",
  33788=>"000000111",
  33789=>"000000000",
  33790=>"111111111",
  33791=>"000000111",
  33792=>"111111111",
  33793=>"111000000",
  33794=>"111111101",
  33795=>"000000100",
  33796=>"011111111",
  33797=>"111110000",
  33798=>"111001111",
  33799=>"111001001",
  33800=>"000000111",
  33801=>"111011000",
  33802=>"111111111",
  33803=>"001000101",
  33804=>"110010000",
  33805=>"000001111",
  33806=>"101100000",
  33807=>"100000000",
  33808=>"011101101",
  33809=>"010000000",
  33810=>"110110110",
  33811=>"111111111",
  33812=>"000000111",
  33813=>"000000000",
  33814=>"000000110",
  33815=>"011111111",
  33816=>"111111111",
  33817=>"110110011",
  33818=>"011011000",
  33819=>"100001000",
  33820=>"000000000",
  33821=>"000000001",
  33822=>"111011000",
  33823=>"001000000",
  33824=>"001000000",
  33825=>"110110110",
  33826=>"000111010",
  33827=>"111000000",
  33828=>"000110010",
  33829=>"000000000",
  33830=>"000000000",
  33831=>"111111111",
  33832=>"111111111",
  33833=>"010111010",
  33834=>"111110111",
  33835=>"010111100",
  33836=>"000000111",
  33837=>"001100111",
  33838=>"111000000",
  33839=>"111000110",
  33840=>"100111000",
  33841=>"101000100",
  33842=>"000000000",
  33843=>"011111111",
  33844=>"000011111",
  33845=>"011111111",
  33846=>"111001000",
  33847=>"000001010",
  33848=>"000001111",
  33849=>"010010000",
  33850=>"101000000",
  33851=>"000000000",
  33852=>"111001100",
  33853=>"111101001",
  33854=>"110110111",
  33855=>"000000000",
  33856=>"101000000",
  33857=>"000001101",
  33858=>"111000100",
  33859=>"010000111",
  33860=>"010001001",
  33861=>"001001000",
  33862=>"000000000",
  33863=>"000000000",
  33864=>"000000110",
  33865=>"101000001",
  33866=>"000111111",
  33867=>"111111000",
  33868=>"110000101",
  33869=>"000000000",
  33870=>"000001011",
  33871=>"111111111",
  33872=>"000000000",
  33873=>"111101000",
  33874=>"000000000",
  33875=>"000000100",
  33876=>"111001111",
  33877=>"111111111",
  33878=>"000000000",
  33879=>"111111111",
  33880=>"111000011",
  33881=>"111000000",
  33882=>"111110000",
  33883=>"000000001",
  33884=>"110111111",
  33885=>"110000000",
  33886=>"111111111",
  33887=>"000100111",
  33888=>"100101100",
  33889=>"111111111",
  33890=>"000000000",
  33891=>"101101111",
  33892=>"110000000",
  33893=>"001000101",
  33894=>"000001111",
  33895=>"110100100",
  33896=>"100101111",
  33897=>"101111000",
  33898=>"010110010",
  33899=>"101000101",
  33900=>"111111001",
  33901=>"000111111",
  33902=>"100110111",
  33903=>"000100100",
  33904=>"111111110",
  33905=>"111111010",
  33906=>"000111111",
  33907=>"111111111",
  33908=>"110000000",
  33909=>"000111010",
  33910=>"111101111",
  33911=>"111111001",
  33912=>"001000100",
  33913=>"111111111",
  33914=>"000000000",
  33915=>"000000001",
  33916=>"110110000",
  33917=>"000010000",
  33918=>"000000000",
  33919=>"000000000",
  33920=>"000000111",
  33921=>"000000111",
  33922=>"111111111",
  33923=>"000011111",
  33924=>"000000111",
  33925=>"111100101",
  33926=>"010110110",
  33927=>"111011001",
  33928=>"000000001",
  33929=>"011111111",
  33930=>"000000001",
  33931=>"111111111",
  33932=>"101001001",
  33933=>"000000000",
  33934=>"011001001",
  33935=>"000000001",
  33936=>"111111111",
  33937=>"000001111",
  33938=>"111111111",
  33939=>"110111111",
  33940=>"111111111",
  33941=>"000000000",
  33942=>"110000111",
  33943=>"000000111",
  33944=>"000001110",
  33945=>"111111011",
  33946=>"000000000",
  33947=>"001000001",
  33948=>"111111111",
  33949=>"011000000",
  33950=>"111111111",
  33951=>"000000000",
  33952=>"000110101",
  33953=>"111011011",
  33954=>"011111000",
  33955=>"111000000",
  33956=>"111101100",
  33957=>"111111101",
  33958=>"111111000",
  33959=>"111111111",
  33960=>"010111111",
  33961=>"000000000",
  33962=>"111111111",
  33963=>"111111111",
  33964=>"000000000",
  33965=>"000000000",
  33966=>"111110000",
  33967=>"011001000",
  33968=>"111111111",
  33969=>"011001011",
  33970=>"110111110",
  33971=>"000001111",
  33972=>"000000111",
  33973=>"000000000",
  33974=>"111110000",
  33975=>"000100111",
  33976=>"001001000",
  33977=>"000000001",
  33978=>"101001001",
  33979=>"000000001",
  33980=>"110111111",
  33981=>"000000000",
  33982=>"100000100",
  33983=>"000000001",
  33984=>"001000000",
  33985=>"000000000",
  33986=>"000000000",
  33987=>"110111010",
  33988=>"000000111",
  33989=>"111110111",
  33990=>"110100111",
  33991=>"000100100",
  33992=>"000000000",
  33993=>"101000101",
  33994=>"100000100",
  33995=>"000000010",
  33996=>"000000000",
  33997=>"001001000",
  33998=>"111000000",
  33999=>"000100111",
  34000=>"001001001",
  34001=>"100110110",
  34002=>"000010000",
  34003=>"111100111",
  34004=>"001100100",
  34005=>"001000001",
  34006=>"000000000",
  34007=>"001111111",
  34008=>"100111000",
  34009=>"111111111",
  34010=>"000000000",
  34011=>"111111111",
  34012=>"000000111",
  34013=>"000000000",
  34014=>"010111111",
  34015=>"100100101",
  34016=>"011001111",
  34017=>"000000000",
  34018=>"000101110",
  34019=>"111001001",
  34020=>"111011011",
  34021=>"011001101",
  34022=>"111111111",
  34023=>"111111111",
  34024=>"001000110",
  34025=>"000000010",
  34026=>"011011000",
  34027=>"000000011",
  34028=>"010000000",
  34029=>"000111110",
  34030=>"111111101",
  34031=>"000000000",
  34032=>"000000000",
  34033=>"001111111",
  34034=>"111111101",
  34035=>"000000000",
  34036=>"000011111",
  34037=>"000000001",
  34038=>"011111111",
  34039=>"010111110",
  34040=>"000000111",
  34041=>"000000000",
  34042=>"000000000",
  34043=>"111001001",
  34044=>"101000000",
  34045=>"110000100",
  34046=>"111111111",
  34047=>"001001000",
  34048=>"000000000",
  34049=>"000011011",
  34050=>"000000000",
  34051=>"000000000",
  34052=>"111111111",
  34053=>"111000000",
  34054=>"000101101",
  34055=>"010000000",
  34056=>"000001011",
  34057=>"111100000",
  34058=>"111111111",
  34059=>"111111111",
  34060=>"010111111",
  34061=>"000000000",
  34062=>"111110111",
  34063=>"011011111",
  34064=>"111111111",
  34065=>"011110010",
  34066=>"000000000",
  34067=>"000000100",
  34068=>"111000000",
  34069=>"000100000",
  34070=>"110110110",
  34071=>"001000111",
  34072=>"011111111",
  34073=>"111110100",
  34074=>"000000000",
  34075=>"000000010",
  34076=>"000000011",
  34077=>"000000000",
  34078=>"111001111",
  34079=>"011001001",
  34080=>"000100111",
  34081=>"111110110",
  34082=>"100100100",
  34083=>"111111111",
  34084=>"010111111",
  34085=>"000000001",
  34086=>"101101111",
  34087=>"110110000",
  34088=>"110011001",
  34089=>"000000100",
  34090=>"111101000",
  34091=>"000100101",
  34092=>"100000000",
  34093=>"110100111",
  34094=>"011011000",
  34095=>"000000100",
  34096=>"100111110",
  34097=>"000000000",
  34098=>"111001001",
  34099=>"100000110",
  34100=>"100111111",
  34101=>"110110111",
  34102=>"000000011",
  34103=>"101000000",
  34104=>"000000111",
  34105=>"000000000",
  34106=>"000000100",
  34107=>"000111111",
  34108=>"111111011",
  34109=>"110000110",
  34110=>"110000000",
  34111=>"000000001",
  34112=>"001000000",
  34113=>"111111110",
  34114=>"111011111",
  34115=>"000000000",
  34116=>"000000000",
  34117=>"011000110",
  34118=>"000000000",
  34119=>"110111111",
  34120=>"000111111",
  34121=>"000000000",
  34122=>"111111111",
  34123=>"000100110",
  34124=>"000000000",
  34125=>"110110000",
  34126=>"000000000",
  34127=>"010000000",
  34128=>"011111000",
  34129=>"111011000",
  34130=>"111110101",
  34131=>"000000001",
  34132=>"000000000",
  34133=>"001000001",
  34134=>"010110000",
  34135=>"111011000",
  34136=>"111111000",
  34137=>"111111111",
  34138=>"011001001",
  34139=>"011111111",
  34140=>"111111111",
  34141=>"111000001",
  34142=>"000000000",
  34143=>"011111111",
  34144=>"001001111",
  34145=>"111111111",
  34146=>"110110110",
  34147=>"111111111",
  34148=>"011011111",
  34149=>"001000000",
  34150=>"000111111",
  34151=>"010110010",
  34152=>"100010111",
  34153=>"111111010",
  34154=>"001001001",
  34155=>"011111111",
  34156=>"111001000",
  34157=>"111111111",
  34158=>"101000111",
  34159=>"100000001",
  34160=>"000001000",
  34161=>"010001011",
  34162=>"001001100",
  34163=>"111001000",
  34164=>"111111000",
  34165=>"001000000",
  34166=>"011111010",
  34167=>"000010000",
  34168=>"000000100",
  34169=>"000111111",
  34170=>"000000000",
  34171=>"000110000",
  34172=>"000000100",
  34173=>"111110000",
  34174=>"111110110",
  34175=>"111111111",
  34176=>"001001001",
  34177=>"000000100",
  34178=>"100000001",
  34179=>"111111111",
  34180=>"011111011",
  34181=>"111111110",
  34182=>"000000000",
  34183=>"000000110",
  34184=>"101000000",
  34185=>"100100000",
  34186=>"101000000",
  34187=>"000111000",
  34188=>"011111111",
  34189=>"001001100",
  34190=>"001011111",
  34191=>"110100100",
  34192=>"010111000",
  34193=>"111111000",
  34194=>"000010000",
  34195=>"110111111",
  34196=>"000000000",
  34197=>"000000000",
  34198=>"111101101",
  34199=>"001000010",
  34200=>"111100010",
  34201=>"000000001",
  34202=>"000101001",
  34203=>"001000100",
  34204=>"001000000",
  34205=>"000011111",
  34206=>"000000110",
  34207=>"000100111",
  34208=>"100000100",
  34209=>"011111001",
  34210=>"000101111",
  34211=>"000000000",
  34212=>"111001111",
  34213=>"000001001",
  34214=>"111111111",
  34215=>"111111111",
  34216=>"000000000",
  34217=>"000000000",
  34218=>"000000010",
  34219=>"000000011",
  34220=>"000111000",
  34221=>"111111111",
  34222=>"110000000",
  34223=>"111011001",
  34224=>"011011000",
  34225=>"000110110",
  34226=>"001011011",
  34227=>"000011111",
  34228=>"010011010",
  34229=>"111111101",
  34230=>"110111111",
  34231=>"001000000",
  34232=>"010000011",
  34233=>"111111110",
  34234=>"000000011",
  34235=>"101000101",
  34236=>"000000010",
  34237=>"001001111",
  34238=>"000000000",
  34239=>"000010001",
  34240=>"111111011",
  34241=>"000111111",
  34242=>"111111111",
  34243=>"000001001",
  34244=>"111011111",
  34245=>"110100000",
  34246=>"111010000",
  34247=>"000000101",
  34248=>"011000000",
  34249=>"111111000",
  34250=>"000000000",
  34251=>"000000000",
  34252=>"000000000",
  34253=>"000000000",
  34254=>"000000001",
  34255=>"111001001",
  34256=>"111111111",
  34257=>"100111111",
  34258=>"111111110",
  34259=>"000111111",
  34260=>"100100000",
  34261=>"111001000",
  34262=>"000000100",
  34263=>"100100001",
  34264=>"011001111",
  34265=>"111111111",
  34266=>"000000000",
  34267=>"110100110",
  34268=>"100001001",
  34269=>"000000111",
  34270=>"000000111",
  34271=>"100100110",
  34272=>"110111111",
  34273=>"111111111",
  34274=>"111111111",
  34275=>"101000001",
  34276=>"111111111",
  34277=>"000111111",
  34278=>"100110000",
  34279=>"000111111",
  34280=>"111101000",
  34281=>"111110111",
  34282=>"110111000",
  34283=>"000000000",
  34284=>"000011111",
  34285=>"001001000",
  34286=>"000111110",
  34287=>"000101100",
  34288=>"000000001",
  34289=>"111111111",
  34290=>"111111111",
  34291=>"000000001",
  34292=>"011011111",
  34293=>"111000000",
  34294=>"111101000",
  34295=>"111010111",
  34296=>"010000111",
  34297=>"001001001",
  34298=>"000000000",
  34299=>"000100111",
  34300=>"111111110",
  34301=>"000111011",
  34302=>"010000011",
  34303=>"111001101",
  34304=>"001111011",
  34305=>"000000000",
  34306=>"000101111",
  34307=>"000110111",
  34308=>"110111111",
  34309=>"011001111",
  34310=>"000000000",
  34311=>"111111111",
  34312=>"111111111",
  34313=>"100110111",
  34314=>"001110111",
  34315=>"000001011",
  34316=>"001001011",
  34317=>"000111111",
  34318=>"000000000",
  34319=>"110010000",
  34320=>"111101101",
  34321=>"101000000",
  34322=>"111111001",
  34323=>"000000100",
  34324=>"000000000",
  34325=>"011101101",
  34326=>"111111000",
  34327=>"111000000",
  34328=>"011000000",
  34329=>"010000001",
  34330=>"000000000",
  34331=>"111111100",
  34332=>"000000000",
  34333=>"111111001",
  34334=>"100000100",
  34335=>"000000010",
  34336=>"111111111",
  34337=>"000000000",
  34338=>"000000001",
  34339=>"010000000",
  34340=>"010010111",
  34341=>"110111111",
  34342=>"111101101",
  34343=>"011111111",
  34344=>"011111111",
  34345=>"000000000",
  34346=>"110110000",
  34347=>"110111111",
  34348=>"111111111",
  34349=>"000000000",
  34350=>"100000000",
  34351=>"111111111",
  34352=>"000000000",
  34353=>"000000000",
  34354=>"100100111",
  34355=>"001111000",
  34356=>"001001001",
  34357=>"111111111",
  34358=>"010000000",
  34359=>"110110001",
  34360=>"000000100",
  34361=>"111110111",
  34362=>"111111111",
  34363=>"111001000",
  34364=>"001111111",
  34365=>"111111111",
  34366=>"000110011",
  34367=>"111111111",
  34368=>"000000000",
  34369=>"001001000",
  34370=>"000000000",
  34371=>"001000011",
  34372=>"111000000",
  34373=>"111111110",
  34374=>"111011011",
  34375=>"111000111",
  34376=>"111110110",
  34377=>"000000000",
  34378=>"011011011",
  34379=>"111111111",
  34380=>"000100111",
  34381=>"111111111",
  34382=>"111111111",
  34383=>"000000000",
  34384=>"111111000",
  34385=>"001000000",
  34386=>"010111110",
  34387=>"011111110",
  34388=>"111101101",
  34389=>"000000000",
  34390=>"000000000",
  34391=>"110110000",
  34392=>"000111111",
  34393=>"000000000",
  34394=>"010000111",
  34395=>"111111111",
  34396=>"000000001",
  34397=>"000110010",
  34398=>"000011000",
  34399=>"000000000",
  34400=>"000111001",
  34401=>"110110110",
  34402=>"000000000",
  34403=>"111111111",
  34404=>"000111111",
  34405=>"010110000",
  34406=>"111110110",
  34407=>"111111111",
  34408=>"001001111",
  34409=>"000000000",
  34410=>"011011011",
  34411=>"011001000",
  34412=>"110100110",
  34413=>"000100110",
  34414=>"111111111",
  34415=>"000111111",
  34416=>"101000000",
  34417=>"001000110",
  34418=>"100001001",
  34419=>"110110110",
  34420=>"111100100",
  34421=>"111111110",
  34422=>"000000000",
  34423=>"111101000",
  34424=>"111101100",
  34425=>"000111111",
  34426=>"010010000",
  34427=>"011000101",
  34428=>"010010110",
  34429=>"000010110",
  34430=>"000000000",
  34431=>"000000000",
  34432=>"000000000",
  34433=>"000000000",
  34434=>"110100100",
  34435=>"000000000",
  34436=>"000000011",
  34437=>"001000000",
  34438=>"111111111",
  34439=>"001000011",
  34440=>"000001000",
  34441=>"011000011",
  34442=>"111101111",
  34443=>"111100000",
  34444=>"111011001",
  34445=>"001000000",
  34446=>"101000000",
  34447=>"111011111",
  34448=>"000000001",
  34449=>"111101101",
  34450=>"011100100",
  34451=>"001001111",
  34452=>"000000000",
  34453=>"100100100",
  34454=>"110110000",
  34455=>"111011000",
  34456=>"000000000",
  34457=>"010010111",
  34458=>"000000000",
  34459=>"111111110",
  34460=>"010010000",
  34461=>"000000000",
  34462=>"111111000",
  34463=>"001000111",
  34464=>"000000000",
  34465=>"111111011",
  34466=>"001000010",
  34467=>"111111111",
  34468=>"111111110",
  34469=>"111111111",
  34470=>"001000000",
  34471=>"111101001",
  34472=>"110111110",
  34473=>"100000000",
  34474=>"010010000",
  34475=>"000001111",
  34476=>"011010111",
  34477=>"100100100",
  34478=>"011000000",
  34479=>"000000001",
  34480=>"000111111",
  34481=>"111100100",
  34482=>"011001011",
  34483=>"011000000",
  34484=>"111111110",
  34485=>"100100000",
  34486=>"110111111",
  34487=>"000010111",
  34488=>"111000000",
  34489=>"001000000",
  34490=>"010111110",
  34491=>"010111000",
  34492=>"111111110",
  34493=>"000111111",
  34494=>"001100000",
  34495=>"000000110",
  34496=>"001000111",
  34497=>"011000000",
  34498=>"011011110",
  34499=>"000000000",
  34500=>"011111000",
  34501=>"000000000",
  34502=>"000011110",
  34503=>"111111111",
  34504=>"000111111",
  34505=>"001000000",
  34506=>"100110111",
  34507=>"111111111",
  34508=>"001001001",
  34509=>"001111010",
  34510=>"111011011",
  34511=>"000000110",
  34512=>"111111111",
  34513=>"000000101",
  34514=>"000001111",
  34515=>"111101101",
  34516=>"000100001",
  34517=>"000001011",
  34518=>"000000000",
  34519=>"000000000",
  34520=>"000100100",
  34521=>"000000101",
  34522=>"010111111",
  34523=>"000000100",
  34524=>"110111111",
  34525=>"000000000",
  34526=>"001000111",
  34527=>"111111000",
  34528=>"000000000",
  34529=>"001000000",
  34530=>"111111111",
  34531=>"111000000",
  34532=>"110110110",
  34533=>"011111111",
  34534=>"111111110",
  34535=>"111111000",
  34536=>"101000000",
  34537=>"101111000",
  34538=>"111111011",
  34539=>"111000000",
  34540=>"000000000",
  34541=>"010000000",
  34542=>"111101000",
  34543=>"000000000",
  34544=>"000000000",
  34545=>"111000000",
  34546=>"000001010",
  34547=>"000000000",
  34548=>"010000100",
  34549=>"110000000",
  34550=>"011011111",
  34551=>"000000000",
  34552=>"111110011",
  34553=>"001111111",
  34554=>"111111111",
  34555=>"100111111",
  34556=>"100000001",
  34557=>"111111110",
  34558=>"111111111",
  34559=>"111111110",
  34560=>"000100000",
  34561=>"001101101",
  34562=>"000000000",
  34563=>"100000001",
  34564=>"111111111",
  34565=>"000000111",
  34566=>"111111000",
  34567=>"001011000",
  34568=>"000000000",
  34569=>"000000111",
  34570=>"111111111",
  34571=>"110011011",
  34572=>"111111111",
  34573=>"111101111",
  34574=>"000000111",
  34575=>"111111111",
  34576=>"010000000",
  34577=>"000000101",
  34578=>"000000000",
  34579=>"001001000",
  34580=>"000000000",
  34581=>"111000011",
  34582=>"110100100",
  34583=>"101101001",
  34584=>"000000000",
  34585=>"000000100",
  34586=>"000000001",
  34587=>"111110000",
  34588=>"111110110",
  34589=>"000000110",
  34590=>"010011111",
  34591=>"111000011",
  34592=>"110111111",
  34593=>"000000000",
  34594=>"001111111",
  34595=>"000001001",
  34596=>"111110110",
  34597=>"111111111",
  34598=>"001101101",
  34599=>"001000000",
  34600=>"010000000",
  34601=>"000000000",
  34602=>"111111111",
  34603=>"001001100",
  34604=>"000000001",
  34605=>"100100000",
  34606=>"000000000",
  34607=>"000000001",
  34608=>"000001000",
  34609=>"111000001",
  34610=>"111100101",
  34611=>"000000110",
  34612=>"111001001",
  34613=>"000000001",
  34614=>"110010000",
  34615=>"000011111",
  34616=>"111000111",
  34617=>"000000011",
  34618=>"010000001",
  34619=>"111111111",
  34620=>"000000000",
  34621=>"111111111",
  34622=>"010000000",
  34623=>"010000000",
  34624=>"000000000",
  34625=>"111101011",
  34626=>"000111111",
  34627=>"001000000",
  34628=>"000000000",
  34629=>"000001001",
  34630=>"110000000",
  34631=>"111101001",
  34632=>"111111101",
  34633=>"111111111",
  34634=>"000000000",
  34635=>"011001001",
  34636=>"110111000",
  34637=>"011011011",
  34638=>"011111000",
  34639=>"000100110",
  34640=>"000100100",
  34641=>"000000000",
  34642=>"110110111",
  34643=>"000100110",
  34644=>"111111000",
  34645=>"011011011",
  34646=>"010000000",
  34647=>"110110110",
  34648=>"111000000",
  34649=>"011011001",
  34650=>"111100100",
  34651=>"011000000",
  34652=>"000000100",
  34653=>"001011111",
  34654=>"111111011",
  34655=>"111111100",
  34656=>"101100100",
  34657=>"000000000",
  34658=>"111001000",
  34659=>"000001111",
  34660=>"100111101",
  34661=>"011111011",
  34662=>"001111111",
  34663=>"111111111",
  34664=>"111111000",
  34665=>"100000000",
  34666=>"100100111",
  34667=>"000000100",
  34668=>"011000000",
  34669=>"000000000",
  34670=>"000000100",
  34671=>"111100111",
  34672=>"000000101",
  34673=>"111100000",
  34674=>"011111111",
  34675=>"100000100",
  34676=>"110110100",
  34677=>"100000000",
  34678=>"000000000",
  34679=>"000001001",
  34680=>"110110110",
  34681=>"000110010",
  34682=>"000000000",
  34683=>"111111111",
  34684=>"111111111",
  34685=>"001001000",
  34686=>"111011000",
  34687=>"000000000",
  34688=>"100100000",
  34689=>"110111101",
  34690=>"111111111",
  34691=>"100100110",
  34692=>"000110111",
  34693=>"001000000",
  34694=>"110110110",
  34695=>"000011111",
  34696=>"000000000",
  34697=>"100000010",
  34698=>"001000000",
  34699=>"111000000",
  34700=>"111111111",
  34701=>"100110111",
  34702=>"111001001",
  34703=>"011111011",
  34704=>"111111111",
  34705=>"000000000",
  34706=>"111111011",
  34707=>"000000111",
  34708=>"111111110",
  34709=>"000010000",
  34710=>"110000000",
  34711=>"111001001",
  34712=>"111111111",
  34713=>"110110110",
  34714=>"000010010",
  34715=>"000011111",
  34716=>"000111011",
  34717=>"111111111",
  34718=>"000000000",
  34719=>"000000000",
  34720=>"110000000",
  34721=>"111111011",
  34722=>"111111111",
  34723=>"000000111",
  34724=>"000010011",
  34725=>"000000000",
  34726=>"000000000",
  34727=>"101111111",
  34728=>"011011011",
  34729=>"111111011",
  34730=>"000000100",
  34731=>"000000000",
  34732=>"000000000",
  34733=>"000000100",
  34734=>"000000000",
  34735=>"111111111",
  34736=>"000000000",
  34737=>"111111111",
  34738=>"000000001",
  34739=>"110110110",
  34740=>"111000000",
  34741=>"000000000",
  34742=>"011111111",
  34743=>"000000111",
  34744=>"011011010",
  34745=>"111101111",
  34746=>"111000000",
  34747=>"100110100",
  34748=>"001001001",
  34749=>"000010110",
  34750=>"001000000",
  34751=>"100100000",
  34752=>"111111001",
  34753=>"100111111",
  34754=>"000000000",
  34755=>"111111011",
  34756=>"100110110",
  34757=>"000000111",
  34758=>"000000000",
  34759=>"001001111",
  34760=>"111000000",
  34761=>"000000000",
  34762=>"000000000",
  34763=>"000000010",
  34764=>"111001111",
  34765=>"000000000",
  34766=>"111111111",
  34767=>"000000000",
  34768=>"001000010",
  34769=>"001001000",
  34770=>"111111111",
  34771=>"000000000",
  34772=>"111011011",
  34773=>"110010111",
  34774=>"111111111",
  34775=>"000000000",
  34776=>"000100111",
  34777=>"111101100",
  34778=>"100010110",
  34779=>"111110000",
  34780=>"011011111",
  34781=>"010000000",
  34782=>"000001000",
  34783=>"111111101",
  34784=>"011101101",
  34785=>"111010010",
  34786=>"000001111",
  34787=>"110111111",
  34788=>"111110110",
  34789=>"000010110",
  34790=>"000100111",
  34791=>"000000000",
  34792=>"011010010",
  34793=>"100100000",
  34794=>"100000111",
  34795=>"000000001",
  34796=>"000000000",
  34797=>"111001001",
  34798=>"111111111",
  34799=>"001000000",
  34800=>"001001101",
  34801=>"100000000",
  34802=>"111111011",
  34803=>"000000000",
  34804=>"110111010",
  34805=>"000000000",
  34806=>"000000000",
  34807=>"110110010",
  34808=>"011111111",
  34809=>"011010011",
  34810=>"111110111",
  34811=>"001111110",
  34812=>"000100101",
  34813=>"011000000",
  34814=>"111111100",
  34815=>"001011111",
  34816=>"111001000",
  34817=>"110111111",
  34818=>"111111111",
  34819=>"111111111",
  34820=>"001000000",
  34821=>"101000000",
  34822=>"000011011",
  34823=>"111111111",
  34824=>"001001001",
  34825=>"111111001",
  34826=>"000000000",
  34827=>"000110110",
  34828=>"110100000",
  34829=>"110100000",
  34830=>"000000100",
  34831=>"001001001",
  34832=>"010000111",
  34833=>"000111101",
  34834=>"111111111",
  34835=>"111111111",
  34836=>"111001000",
  34837=>"111110110",
  34838=>"110111100",
  34839=>"011111001",
  34840=>"111111110",
  34841=>"111110111",
  34842=>"000000000",
  34843=>"010010111",
  34844=>"110110111",
  34845=>"110110111",
  34846=>"111110111",
  34847=>"110110000",
  34848=>"011000111",
  34849=>"111111111",
  34850=>"000000110",
  34851=>"111000011",
  34852=>"111111000",
  34853=>"111101111",
  34854=>"001000000",
  34855=>"111110000",
  34856=>"111000000",
  34857=>"000000000",
  34858=>"000000111",
  34859=>"111101111",
  34860=>"011111111",
  34861=>"011011011",
  34862=>"000000111",
  34863=>"001001000",
  34864=>"000000000",
  34865=>"111111111",
  34866=>"111111001",
  34867=>"001100111",
  34868=>"011111111",
  34869=>"111110110",
  34870=>"100000111",
  34871=>"110111011",
  34872=>"000000000",
  34873=>"000000111",
  34874=>"111110111",
  34875=>"001000000",
  34876=>"100000000",
  34877=>"011000000",
  34878=>"111111111",
  34879=>"000000000",
  34880=>"011111011",
  34881=>"000000000",
  34882=>"111111011",
  34883=>"000011000",
  34884=>"001000110",
  34885=>"111111111",
  34886=>"111111000",
  34887=>"000000000",
  34888=>"011000000",
  34889=>"110100111",
  34890=>"011111111",
  34891=>"011111111",
  34892=>"110100000",
  34893=>"111111111",
  34894=>"110000000",
  34895=>"100101011",
  34896=>"111010000",
  34897=>"000000111",
  34898=>"000000100",
  34899=>"111111111",
  34900=>"000000000",
  34901=>"111111111",
  34902=>"001011111",
  34903=>"100110100",
  34904=>"111111111",
  34905=>"010000000",
  34906=>"011111111",
  34907=>"000110000",
  34908=>"000000000",
  34909=>"000000000",
  34910=>"111100100",
  34911=>"111011001",
  34912=>"111111111",
  34913=>"101111101",
  34914=>"010110010",
  34915=>"000111111",
  34916=>"000000011",
  34917=>"011001000",
  34918=>"110000100",
  34919=>"000100110",
  34920=>"111100000",
  34921=>"000000000",
  34922=>"111111111",
  34923=>"111111000",
  34924=>"111110111",
  34925=>"111111111",
  34926=>"110000001",
  34927=>"111111111",
  34928=>"111110110",
  34929=>"000000100",
  34930=>"000000111",
  34931=>"010000000",
  34932=>"000000000",
  34933=>"110110110",
  34934=>"011111110",
  34935=>"111001001",
  34936=>"111111111",
  34937=>"111001101",
  34938=>"000001011",
  34939=>"111111111",
  34940=>"010110111",
  34941=>"111111011",
  34942=>"000000110",
  34943=>"001001001",
  34944=>"000001111",
  34945=>"000000011",
  34946=>"111100000",
  34947=>"111111111",
  34948=>"110110111",
  34949=>"010111111",
  34950=>"001101111",
  34951=>"111011000",
  34952=>"111111010",
  34953=>"000001111",
  34954=>"100000000",
  34955=>"011111111",
  34956=>"000000000",
  34957=>"100001101",
  34958=>"111111111",
  34959=>"000000100",
  34960=>"000011011",
  34961=>"011001000",
  34962=>"000111011",
  34963=>"111001001",
  34964=>"011111000",
  34965=>"001001000",
  34966=>"111111111",
  34967=>"000000000",
  34968=>"111010011",
  34969=>"011000000",
  34970=>"111111111",
  34971=>"000000000",
  34972=>"111001001",
  34973=>"101100101",
  34974=>"000000000",
  34975=>"000000000",
  34976=>"000000000",
  34977=>"011000001",
  34978=>"000110000",
  34979=>"000000000",
  34980=>"110111100",
  34981=>"111000000",
  34982=>"000000000",
  34983=>"100111111",
  34984=>"111000000",
  34985=>"000000000",
  34986=>"111111111",
  34987=>"000000000",
  34988=>"111100100",
  34989=>"011001000",
  34990=>"000001111",
  34991=>"111111101",
  34992=>"000000000",
  34993=>"101011111",
  34994=>"000000000",
  34995=>"111111111",
  34996=>"000000000",
  34997=>"001111111",
  34998=>"000100001",
  34999=>"111111001",
  35000=>"111100101",
  35001=>"000000000",
  35002=>"001001001",
  35003=>"001000000",
  35004=>"100110111",
  35005=>"110111000",
  35006=>"111000111",
  35007=>"000000000",
  35008=>"111110000",
  35009=>"011111110",
  35010=>"000000000",
  35011=>"111111111",
  35012=>"111111111",
  35013=>"000000000",
  35014=>"110101111",
  35015=>"010010011",
  35016=>"111100111",
  35017=>"000000000",
  35018=>"111011000",
  35019=>"111011111",
  35020=>"000000000",
  35021=>"111000000",
  35022=>"111111111",
  35023=>"111100011",
  35024=>"111111111",
  35025=>"000100111",
  35026=>"111110110",
  35027=>"000000000",
  35028=>"110001001",
  35029=>"111111110",
  35030=>"000000000",
  35031=>"111000001",
  35032=>"011111111",
  35033=>"000000000",
  35034=>"000001111",
  35035=>"000000000",
  35036=>"101111111",
  35037=>"111110110",
  35038=>"000000000",
  35039=>"001001011",
  35040=>"000000000",
  35041=>"000000000",
  35042=>"111110000",
  35043=>"001000011",
  35044=>"100000000",
  35045=>"101100100",
  35046=>"011000000",
  35047=>"001000000",
  35048=>"111111111",
  35049=>"111111111",
  35050=>"111010001",
  35051=>"000000111",
  35052=>"111111111",
  35053=>"001000000",
  35054=>"111011111",
  35055=>"000000000",
  35056=>"000100000",
  35057=>"111111111",
  35058=>"101000000",
  35059=>"011001000",
  35060=>"011111111",
  35061=>"111110110",
  35062=>"111111110",
  35063=>"000100100",
  35064=>"000110111",
  35065=>"111111110",
  35066=>"010010000",
  35067=>"000001001",
  35068=>"100001110",
  35069=>"000000000",
  35070=>"111001011",
  35071=>"101000000",
  35072=>"111111111",
  35073=>"111101000",
  35074=>"111111111",
  35075=>"110010111",
  35076=>"111011011",
  35077=>"111100100",
  35078=>"000000011",
  35079=>"110000000",
  35080=>"011000000",
  35081=>"000100000",
  35082=>"000000000",
  35083=>"011010111",
  35084=>"100110000",
  35085=>"001000101",
  35086=>"111111111",
  35087=>"000000111",
  35088=>"000100111",
  35089=>"100000011",
  35090=>"110110101",
  35091=>"100100110",
  35092=>"110111111",
  35093=>"000100000",
  35094=>"100100100",
  35095=>"110110000",
  35096=>"101101111",
  35097=>"000011011",
  35098=>"000000000",
  35099=>"111111111",
  35100=>"010010000",
  35101=>"111111111",
  35102=>"111111111",
  35103=>"000000000",
  35104=>"111001001",
  35105=>"011001000",
  35106=>"111111111",
  35107=>"100100111",
  35108=>"111111111",
  35109=>"000000000",
  35110=>"000000111",
  35111=>"000001000",
  35112=>"000101111",
  35113=>"100100111",
  35114=>"000000000",
  35115=>"111000000",
  35116=>"111001001",
  35117=>"101010111",
  35118=>"111010111",
  35119=>"111111111",
  35120=>"100100000",
  35121=>"000000101",
  35122=>"000000000",
  35123=>"000000000",
  35124=>"000000000",
  35125=>"100110110",
  35126=>"010111111",
  35127=>"100111100",
  35128=>"000000000",
  35129=>"000000000",
  35130=>"111111000",
  35131=>"000000000",
  35132=>"111111111",
  35133=>"110000000",
  35134=>"100000100",
  35135=>"111111111",
  35136=>"000000000",
  35137=>"111111100",
  35138=>"111111111",
  35139=>"000000110",
  35140=>"011010000",
  35141=>"000000111",
  35142=>"100100100",
  35143=>"110111111",
  35144=>"111111111",
  35145=>"000000000",
  35146=>"111010000",
  35147=>"011111011",
  35148=>"111100111",
  35149=>"110111111",
  35150=>"000000110",
  35151=>"111110100",
  35152=>"100001000",
  35153=>"010000000",
  35154=>"000000000",
  35155=>"111111000",
  35156=>"111100100",
  35157=>"000000000",
  35158=>"111110000",
  35159=>"000000000",
  35160=>"111001010",
  35161=>"000000000",
  35162=>"000000000",
  35163=>"000000000",
  35164=>"000000011",
  35165=>"110111111",
  35166=>"110111111",
  35167=>"111111111",
  35168=>"111111111",
  35169=>"111101000",
  35170=>"110011111",
  35171=>"111111111",
  35172=>"100100111",
  35173=>"100000100",
  35174=>"000100000",
  35175=>"000000000",
  35176=>"100000000",
  35177=>"011111111",
  35178=>"000000000",
  35179=>"100111001",
  35180=>"100000000",
  35181=>"011000000",
  35182=>"100000000",
  35183=>"000100000",
  35184=>"000000000",
  35185=>"001001000",
  35186=>"000000110",
  35187=>"001000001",
  35188=>"111000100",
  35189=>"000000111",
  35190=>"111100100",
  35191=>"000000000",
  35192=>"111111111",
  35193=>"000000000",
  35194=>"111111111",
  35195=>"001111100",
  35196=>"111001000",
  35197=>"111111111",
  35198=>"000000000",
  35199=>"111111001",
  35200=>"111100110",
  35201=>"111111111",
  35202=>"111111111",
  35203=>"011000000",
  35204=>"101000000",
  35205=>"000000000",
  35206=>"111101101",
  35207=>"000000000",
  35208=>"000000000",
  35209=>"000000000",
  35210=>"011110011",
  35211=>"000000000",
  35212=>"000000000",
  35213=>"110110110",
  35214=>"111100111",
  35215=>"000000000",
  35216=>"000010111",
  35217=>"000001000",
  35218=>"111111111",
  35219=>"111111110",
  35220=>"011000000",
  35221=>"001111111",
  35222=>"001000000",
  35223=>"010010100",
  35224=>"111111111",
  35225=>"111001000",
  35226=>"001000000",
  35227=>"101101111",
  35228=>"011111111",
  35229=>"111001000",
  35230=>"001011111",
  35231=>"000000000",
  35232=>"011111000",
  35233=>"000000011",
  35234=>"001110100",
  35235=>"001011011",
  35236=>"111111111",
  35237=>"111111111",
  35238=>"000010000",
  35239=>"100111111",
  35240=>"111111110",
  35241=>"111111000",
  35242=>"100111110",
  35243=>"000000001",
  35244=>"111111111",
  35245=>"000000001",
  35246=>"111111111",
  35247=>"111011001",
  35248=>"000000000",
  35249=>"111111111",
  35250=>"001000000",
  35251=>"111111111",
  35252=>"001001001",
  35253=>"000000000",
  35254=>"111100110",
  35255=>"111000000",
  35256=>"111111111",
  35257=>"111111011",
  35258=>"000000101",
  35259=>"110110100",
  35260=>"000000000",
  35261=>"111111111",
  35262=>"000000000",
  35263=>"110111111",
  35264=>"000001001",
  35265=>"111001001",
  35266=>"111111111",
  35267=>"111111011",
  35268=>"111010010",
  35269=>"111001000",
  35270=>"011000000",
  35271=>"000010001",
  35272=>"011111111",
  35273=>"011011000",
  35274=>"011000000",
  35275=>"000000111",
  35276=>"011111111",
  35277=>"000000000",
  35278=>"000000000",
  35279=>"011000000",
  35280=>"111111111",
  35281=>"001111111",
  35282=>"011010111",
  35283=>"100000000",
  35284=>"110100110",
  35285=>"111111111",
  35286=>"000000010",
  35287=>"011111111",
  35288=>"001000000",
  35289=>"101100110",
  35290=>"111111101",
  35291=>"001001110",
  35292=>"111100000",
  35293=>"001001001",
  35294=>"001001010",
  35295=>"111111111",
  35296=>"000001000",
  35297=>"000000000",
  35298=>"101001000",
  35299=>"101101000",
  35300=>"111111111",
  35301=>"100111111",
  35302=>"111000100",
  35303=>"001001001",
  35304=>"000110100",
  35305=>"101000000",
  35306=>"001111111",
  35307=>"000110000",
  35308=>"000000101",
  35309=>"000000001",
  35310=>"000000111",
  35311=>"111111111",
  35312=>"001000000",
  35313=>"000111111",
  35314=>"011001000",
  35315=>"010110010",
  35316=>"111110111",
  35317=>"000000110",
  35318=>"111111110",
  35319=>"101101111",
  35320=>"000000000",
  35321=>"111101001",
  35322=>"100110111",
  35323=>"000000000",
  35324=>"000000100",
  35325=>"111111111",
  35326=>"000000111",
  35327=>"000000000",
  35328=>"000000000",
  35329=>"111110111",
  35330=>"000000000",
  35331=>"111111111",
  35332=>"110001001",
  35333=>"000011011",
  35334=>"000000100",
  35335=>"000000000",
  35336=>"110110100",
  35337=>"001001001",
  35338=>"110000000",
  35339=>"111000110",
  35340=>"001000001",
  35341=>"000000000",
  35342=>"001011111",
  35343=>"111111111",
  35344=>"000100101",
  35345=>"000010000",
  35346=>"000000111",
  35347=>"100111111",
  35348=>"011111111",
  35349=>"000000001",
  35350=>"110110000",
  35351=>"111111111",
  35352=>"000000000",
  35353=>"100100101",
  35354=>"111111111",
  35355=>"100100111",
  35356=>"111010100",
  35357=>"000000000",
  35358=>"010000000",
  35359=>"110000000",
  35360=>"101111111",
  35361=>"110100000",
  35362=>"000001100",
  35363=>"001000000",
  35364=>"000000000",
  35365=>"111011101",
  35366=>"011111111",
  35367=>"110110100",
  35368=>"111111111",
  35369=>"100101110",
  35370=>"000000000",
  35371=>"000000000",
  35372=>"000000000",
  35373=>"100111111",
  35374=>"001000000",
  35375=>"111110101",
  35376=>"111110000",
  35377=>"000000011",
  35378=>"111101111",
  35379=>"111111111",
  35380=>"011111111",
  35381=>"111111001",
  35382=>"111000111",
  35383=>"111111101",
  35384=>"000100100",
  35385=>"000000000",
  35386=>"110111111",
  35387=>"110000000",
  35388=>"000000000",
  35389=>"110110000",
  35390=>"010001000",
  35391=>"000000000",
  35392=>"010000110",
  35393=>"001111011",
  35394=>"111100000",
  35395=>"111110110",
  35396=>"111001011",
  35397=>"110110110",
  35398=>"000000000",
  35399=>"111111110",
  35400=>"011000111",
  35401=>"000000000",
  35402=>"000000000",
  35403=>"001001101",
  35404=>"000000000",
  35405=>"111011000",
  35406=>"000001011",
  35407=>"111111111",
  35408=>"000000100",
  35409=>"000110110",
  35410=>"111111111",
  35411=>"001001000",
  35412=>"111111000",
  35413=>"100000110",
  35414=>"111101110",
  35415=>"001000000",
  35416=>"000001111",
  35417=>"010010000",
  35418=>"101000001",
  35419=>"111011001",
  35420=>"100001001",
  35421=>"000000000",
  35422=>"000000000",
  35423=>"110110110",
  35424=>"111111111",
  35425=>"111111111",
  35426=>"101000111",
  35427=>"111111111",
  35428=>"111111111",
  35429=>"111110000",
  35430=>"000000000",
  35431=>"000000000",
  35432=>"000000000",
  35433=>"111111111",
  35434=>"101110100",
  35435=>"111111110",
  35436=>"001001000",
  35437=>"000000001",
  35438=>"000000000",
  35439=>"000000000",
  35440=>"111111111",
  35441=>"001000111",
  35442=>"001001011",
  35443=>"101000000",
  35444=>"000000000",
  35445=>"111101111",
  35446=>"000011010",
  35447=>"000001000",
  35448=>"001000000",
  35449=>"000000100",
  35450=>"000000010",
  35451=>"111111011",
  35452=>"000000000",
  35453=>"110111110",
  35454=>"000000000",
  35455=>"000001111",
  35456=>"111111111",
  35457=>"111111111",
  35458=>"000101000",
  35459=>"100100100",
  35460=>"101111111",
  35461=>"110111111",
  35462=>"000000000",
  35463=>"111111010",
  35464=>"111111001",
  35465=>"000000110",
  35466=>"110000111",
  35467=>"000000100",
  35468=>"000101111",
  35469=>"111111111",
  35470=>"001001100",
  35471=>"100010011",
  35472=>"000000000",
  35473=>"001001001",
  35474=>"111111111",
  35475=>"111111111",
  35476=>"000000000",
  35477=>"000000101",
  35478=>"000000000",
  35479=>"111000000",
  35480=>"001101101",
  35481=>"111111111",
  35482=>"000100000",
  35483=>"000000111",
  35484=>"000000100",
  35485=>"111111111",
  35486=>"111111111",
  35487=>"000111000",
  35488=>"110111011",
  35489=>"000000000",
  35490=>"111111111",
  35491=>"111111111",
  35492=>"000100110",
  35493=>"111111111",
  35494=>"111111111",
  35495=>"011011001",
  35496=>"111111111",
  35497=>"000000001",
  35498=>"110111111",
  35499=>"000000000",
  35500=>"111111110",
  35501=>"111111111",
  35502=>"000111111",
  35503=>"001000111",
  35504=>"010110000",
  35505=>"111111001",
  35506=>"100000000",
  35507=>"000000000",
  35508=>"000000000",
  35509=>"000000000",
  35510=>"110111111",
  35511=>"000000000",
  35512=>"101111011",
  35513=>"000000000",
  35514=>"000000000",
  35515=>"100111111",
  35516=>"001000100",
  35517=>"000110111",
  35518=>"000000000",
  35519=>"111111111",
  35520=>"111000000",
  35521=>"100000100",
  35522=>"000000000",
  35523=>"111111001",
  35524=>"000000001",
  35525=>"000000000",
  35526=>"000001110",
  35527=>"000000000",
  35528=>"000111010",
  35529=>"000000111",
  35530=>"111000000",
  35531=>"000000011",
  35532=>"000000111",
  35533=>"000000000",
  35534=>"111110111",
  35535=>"110000010",
  35536=>"000101101",
  35537=>"001101111",
  35538=>"111000000",
  35539=>"110110111",
  35540=>"000000000",
  35541=>"011011111",
  35542=>"000000111",
  35543=>"111001111",
  35544=>"000000111",
  35545=>"111111111",
  35546=>"111111111",
  35547=>"111111111",
  35548=>"111111111",
  35549=>"111111111",
  35550=>"111100100",
  35551=>"000000000",
  35552=>"110011010",
  35553=>"000000011",
  35554=>"111111010",
  35555=>"101111111",
  35556=>"000000100",
  35557=>"110110111",
  35558=>"111110111",
  35559=>"000110111",
  35560=>"111111111",
  35561=>"111111000",
  35562=>"101100111",
  35563=>"001000111",
  35564=>"000000111",
  35565=>"000011111",
  35566=>"000000111",
  35567=>"000000000",
  35568=>"111011011",
  35569=>"111111111",
  35570=>"000101101",
  35571=>"000000001",
  35572=>"000111111",
  35573=>"111000001",
  35574=>"000000000",
  35575=>"111011000",
  35576=>"000000000",
  35577=>"000000000",
  35578=>"111111111",
  35579=>"111001000",
  35580=>"111111111",
  35581=>"010000111",
  35582=>"110111111",
  35583=>"100100010",
  35584=>"011001001",
  35585=>"001001001",
  35586=>"111111111",
  35587=>"000011011",
  35588=>"111100000",
  35589=>"000100100",
  35590=>"100000000",
  35591=>"111111100",
  35592=>"000000001",
  35593=>"000000000",
  35594=>"000000000",
  35595=>"110111111",
  35596=>"110111111",
  35597=>"010000000",
  35598=>"011111111",
  35599=>"000000000",
  35600=>"100011111",
  35601=>"000000000",
  35602=>"000000000",
  35603=>"000111001",
  35604=>"111111111",
  35605=>"111000000",
  35606=>"111111111",
  35607=>"011000000",
  35608=>"000000000",
  35609=>"111111000",
  35610=>"000000100",
  35611=>"000100111",
  35612=>"110110111",
  35613=>"111111111",
  35614=>"000000000",
  35615=>"000000000",
  35616=>"001000000",
  35617=>"000000000",
  35618=>"001111111",
  35619=>"000000000",
  35620=>"111000101",
  35621=>"000000100",
  35622=>"100101101",
  35623=>"000000000",
  35624=>"000000000",
  35625=>"010000000",
  35626=>"111000000",
  35627=>"111101000",
  35628=>"001000111",
  35629=>"000100000",
  35630=>"000000000",
  35631=>"011001000",
  35632=>"000000000",
  35633=>"100000000",
  35634=>"111111111",
  35635=>"000000000",
  35636=>"000001111",
  35637=>"000000011",
  35638=>"100111000",
  35639=>"000000100",
  35640=>"000000000",
  35641=>"000000000",
  35642=>"000000000",
  35643=>"111111000",
  35644=>"000000000",
  35645=>"100000101",
  35646=>"000000000",
  35647=>"101100000",
  35648=>"000000110",
  35649=>"111110110",
  35650=>"000000000",
  35651=>"111111111",
  35652=>"000000110",
  35653=>"111111111",
  35654=>"000111111",
  35655=>"000000111",
  35656=>"110000111",
  35657=>"000000100",
  35658=>"111000101",
  35659=>"111001101",
  35660=>"000110110",
  35661=>"000100000",
  35662=>"000111111",
  35663=>"111111111",
  35664=>"010000000",
  35665=>"100100100",
  35666=>"111011011",
  35667=>"000000000",
  35668=>"001000000",
  35669=>"000000000",
  35670=>"111111010",
  35671=>"001000111",
  35672=>"011111111",
  35673=>"111110110",
  35674=>"001111111",
  35675=>"000000000",
  35676=>"001001000",
  35677=>"000000000",
  35678=>"110100110",
  35679=>"000000000",
  35680=>"000000111",
  35681=>"000000000",
  35682=>"001001001",
  35683=>"001001111",
  35684=>"111111111",
  35685=>"000000000",
  35686=>"000000000",
  35687=>"011111111",
  35688=>"111010000",
  35689=>"111110111",
  35690=>"000000011",
  35691=>"000000000",
  35692=>"000111111",
  35693=>"000111101",
  35694=>"011011110",
  35695=>"000000001",
  35696=>"000000111",
  35697=>"000000000",
  35698=>"011011001",
  35699=>"011111111",
  35700=>"110110110",
  35701=>"110110111",
  35702=>"011011001",
  35703=>"001111111",
  35704=>"000000000",
  35705=>"111111111",
  35706=>"010011111",
  35707=>"111111111",
  35708=>"000000100",
  35709=>"111111111",
  35710=>"111111001",
  35711=>"000000000",
  35712=>"000000000",
  35713=>"001111111",
  35714=>"111100100",
  35715=>"111110000",
  35716=>"000000111",
  35717=>"000000000",
  35718=>"000001101",
  35719=>"110110110",
  35720=>"100000000",
  35721=>"000000100",
  35722=>"000000001",
  35723=>"010000000",
  35724=>"111111111",
  35725=>"101111111",
  35726=>"000000100",
  35727=>"011011111",
  35728=>"000000000",
  35729=>"111111111",
  35730=>"000000000",
  35731=>"000000000",
  35732=>"111111111",
  35733=>"000110110",
  35734=>"000000000",
  35735=>"000000001",
  35736=>"000001111",
  35737=>"111111111",
  35738=>"000000000",
  35739=>"000000000",
  35740=>"100110111",
  35741=>"000000111",
  35742=>"011011010",
  35743=>"111111111",
  35744=>"011111100",
  35745=>"011011001",
  35746=>"001000000",
  35747=>"110111111",
  35748=>"001001111",
  35749=>"111111111",
  35750=>"110111111",
  35751=>"100011111",
  35752=>"001001001",
  35753=>"000000000",
  35754=>"111111111",
  35755=>"010001001",
  35756=>"111001001",
  35757=>"000000000",
  35758=>"000000100",
  35759=>"100000101",
  35760=>"000000000",
  35761=>"000000000",
  35762=>"100010000",
  35763=>"111000000",
  35764=>"000000001",
  35765=>"111111011",
  35766=>"110000000",
  35767=>"111111111",
  35768=>"000000111",
  35769=>"100110000",
  35770=>"111111111",
  35771=>"111111111",
  35772=>"110001111",
  35773=>"001000101",
  35774=>"111100111",
  35775=>"001001001",
  35776=>"001000110",
  35777=>"000000000",
  35778=>"000000000",
  35779=>"000000000",
  35780=>"001000000",
  35781=>"000000000",
  35782=>"111111010",
  35783=>"001101101",
  35784=>"010011010",
  35785=>"000000000",
  35786=>"001000101",
  35787=>"110111111",
  35788=>"000000100",
  35789=>"000000111",
  35790=>"000001001",
  35791=>"011001000",
  35792=>"111101001",
  35793=>"011011011",
  35794=>"000000000",
  35795=>"111111111",
  35796=>"111111111",
  35797=>"111111111",
  35798=>"011011000",
  35799=>"111000000",
  35800=>"000000000",
  35801=>"010000000",
  35802=>"001000100",
  35803=>"000001000",
  35804=>"000000000",
  35805=>"111000000",
  35806=>"000100011",
  35807=>"000000001",
  35808=>"001000000",
  35809=>"011111000",
  35810=>"111111111",
  35811=>"111011000",
  35812=>"111001001",
  35813=>"111110111",
  35814=>"111111111",
  35815=>"000000111",
  35816=>"111111111",
  35817=>"000000000",
  35818=>"101000000",
  35819=>"111111111",
  35820=>"001000110",
  35821=>"000110111",
  35822=>"011011011",
  35823=>"001011001",
  35824=>"000000110",
  35825=>"011111111",
  35826=>"000000100",
  35827=>"000000000",
  35828=>"000100111",
  35829=>"000000000",
  35830=>"001011111",
  35831=>"110100000",
  35832=>"001000000",
  35833=>"010010110",
  35834=>"100000000",
  35835=>"000000111",
  35836=>"011011111",
  35837=>"111000011",
  35838=>"000000010",
  35839=>"111111111",
  35840=>"111100000",
  35841=>"000011011",
  35842=>"000000000",
  35843=>"000000111",
  35844=>"000110111",
  35845=>"001110110",
  35846=>"111111111",
  35847=>"000111111",
  35848=>"000111000",
  35849=>"000000001",
  35850=>"000000000",
  35851=>"111001001",
  35852=>"111111111",
  35853=>"000000111",
  35854=>"111011011",
  35855=>"000011110",
  35856=>"000100000",
  35857=>"111110110",
  35858=>"111101111",
  35859=>"000000111",
  35860=>"100000000",
  35861=>"111111111",
  35862=>"111111111",
  35863=>"000000000",
  35864=>"000000000",
  35865=>"111111111",
  35866=>"000000000",
  35867=>"000000000",
  35868=>"110110000",
  35869=>"111101000",
  35870=>"110111011",
  35871=>"000001111",
  35872=>"110000000",
  35873=>"011000000",
  35874=>"000011111",
  35875=>"100000000",
  35876=>"111000000",
  35877=>"111101100",
  35878=>"111111111",
  35879=>"111111111",
  35880=>"000000000",
  35881=>"000001111",
  35882=>"000000000",
  35883=>"011000100",
  35884=>"000000000",
  35885=>"100001111",
  35886=>"001101101",
  35887=>"111111111",
  35888=>"011110010",
  35889=>"000000100",
  35890=>"111110000",
  35891=>"111111111",
  35892=>"111101101",
  35893=>"110010000",
  35894=>"000000000",
  35895=>"100000001",
  35896=>"000000001",
  35897=>"000000000",
  35898=>"111111111",
  35899=>"100111001",
  35900=>"011111111",
  35901=>"000000000",
  35902=>"000000001",
  35903=>"011000000",
  35904=>"000000000",
  35905=>"010010010",
  35906=>"110111111",
  35907=>"000110011",
  35908=>"000000111",
  35909=>"111011110",
  35910=>"111011111",
  35911=>"111111001",
  35912=>"111111011",
  35913=>"000010000",
  35914=>"111111111",
  35915=>"111111000",
  35916=>"111111111",
  35917=>"010100100",
  35918=>"011111000",
  35919=>"000000101",
  35920=>"111111111",
  35921=>"011010000",
  35922=>"000110010",
  35923=>"000000000",
  35924=>"110000000",
  35925=>"000011111",
  35926=>"000000000",
  35927=>"001000000",
  35928=>"111111110",
  35929=>"001001001",
  35930=>"111111011",
  35931=>"000000111",
  35932=>"111111111",
  35933=>"111111111",
  35934=>"000001001",
  35935=>"111101111",
  35936=>"000000000",
  35937=>"011011111",
  35938=>"000000000",
  35939=>"000000000",
  35940=>"111111001",
  35941=>"110111011",
  35942=>"000000001",
  35943=>"111101111",
  35944=>"111110000",
  35945=>"000000000",
  35946=>"111110111",
  35947=>"111000000",
  35948=>"000000000",
  35949=>"000000000",
  35950=>"001001000",
  35951=>"111111111",
  35952=>"101111111",
  35953=>"011111111",
  35954=>"000000100",
  35955=>"100100110",
  35956=>"000000000",
  35957=>"000000001",
  35958=>"000000000",
  35959=>"110110100",
  35960=>"001100110",
  35961=>"111111111",
  35962=>"110110010",
  35963=>"001111111",
  35964=>"000000100",
  35965=>"000000000",
  35966=>"110010000",
  35967=>"000100001",
  35968=>"000000000",
  35969=>"111111111",
  35970=>"001001111",
  35971=>"000000000",
  35972=>"100000000",
  35973=>"011111111",
  35974=>"111111011",
  35975=>"111100100",
  35976=>"001000001",
  35977=>"111111111",
  35978=>"000111111",
  35979=>"000000110",
  35980=>"000000000",
  35981=>"111111111",
  35982=>"011000000",
  35983=>"111111111",
  35984=>"000000100",
  35985=>"100100000",
  35986=>"111111000",
  35987=>"000000110",
  35988=>"111000000",
  35989=>"011111110",
  35990=>"111111111",
  35991=>"000000000",
  35992=>"000000000",
  35993=>"000000000",
  35994=>"110111111",
  35995=>"110101000",
  35996=>"000100110",
  35997=>"001111111",
  35998=>"111111001",
  35999=>"000100111",
  36000=>"110100000",
  36001=>"111111111",
  36002=>"110110101",
  36003=>"000000000",
  36004=>"110110110",
  36005=>"100101011",
  36006=>"000000101",
  36007=>"110111111",
  36008=>"111011000",
  36009=>"000000100",
  36010=>"111111111",
  36011=>"000000000",
  36012=>"000001011",
  36013=>"010010110",
  36014=>"111111111",
  36015=>"011111111",
  36016=>"111111111",
  36017=>"111111111",
  36018=>"011111111",
  36019=>"111111111",
  36020=>"000110110",
  36021=>"000000000",
  36022=>"001000000",
  36023=>"111111000",
  36024=>"001001111",
  36025=>"111111110",
  36026=>"011111000",
  36027=>"001110001",
  36028=>"110010010",
  36029=>"000001010",
  36030=>"111111111",
  36031=>"110110110",
  36032=>"000000000",
  36033=>"111111111",
  36034=>"000000000",
  36035=>"000000000",
  36036=>"111111011",
  36037=>"000000011",
  36038=>"100000000",
  36039=>"111111110",
  36040=>"000000000",
  36041=>"001001000",
  36042=>"111111111",
  36043=>"111111111",
  36044=>"011001101",
  36045=>"011001001",
  36046=>"111111110",
  36047=>"011000000",
  36048=>"000000000",
  36049=>"100000000",
  36050=>"000000111",
  36051=>"111111010",
  36052=>"111101101",
  36053=>"110111111",
  36054=>"000000000",
  36055=>"000010101",
  36056=>"000011001",
  36057=>"000000001",
  36058=>"000000000",
  36059=>"111111111",
  36060=>"111111111",
  36061=>"000000000",
  36062=>"100110100",
  36063=>"010011001",
  36064=>"000000010",
  36065=>"000000000",
  36066=>"000000011",
  36067=>"001111111",
  36068=>"010010011",
  36069=>"001001001",
  36070=>"111111111",
  36071=>"111011111",
  36072=>"000000000",
  36073=>"111110000",
  36074=>"111011111",
  36075=>"000000000",
  36076=>"000000000",
  36077=>"000011111",
  36078=>"111111000",
  36079=>"111111111",
  36080=>"111110000",
  36081=>"010000000",
  36082=>"000100000",
  36083=>"011111100",
  36084=>"010111111",
  36085=>"111111111",
  36086=>"000000000",
  36087=>"111011111",
  36088=>"111111111",
  36089=>"000000000",
  36090=>"011111111",
  36091=>"110110001",
  36092=>"111111101",
  36093=>"010011001",
  36094=>"001001000",
  36095=>"100100111",
  36096=>"000011111",
  36097=>"100100110",
  36098=>"011001000",
  36099=>"000100000",
  36100=>"000001010",
  36101=>"100100100",
  36102=>"000000111",
  36103=>"000000000",
  36104=>"000000001",
  36105=>"110111000",
  36106=>"111111111",
  36107=>"110110110",
  36108=>"111111011",
  36109=>"001000000",
  36110=>"111111111",
  36111=>"000000000",
  36112=>"110100010",
  36113=>"011011001",
  36114=>"000001000",
  36115=>"001000000",
  36116=>"001001000",
  36117=>"111010111",
  36118=>"001111111",
  36119=>"011001000",
  36120=>"111100100",
  36121=>"111111111",
  36122=>"000000000",
  36123=>"000000100",
  36124=>"110001111",
  36125=>"111111111",
  36126=>"000000001",
  36127=>"111100000",
  36128=>"110110110",
  36129=>"111111111",
  36130=>"111111111",
  36131=>"111111001",
  36132=>"011011001",
  36133=>"011000000",
  36134=>"111111111",
  36135=>"111110000",
  36136=>"001000000",
  36137=>"111111111",
  36138=>"001000000",
  36139=>"110111011",
  36140=>"000000000",
  36141=>"000010010",
  36142=>"011111000",
  36143=>"111001001",
  36144=>"000000111",
  36145=>"110110110",
  36146=>"011000000",
  36147=>"000000000",
  36148=>"000000000",
  36149=>"000101001",
  36150=>"101110110",
  36151=>"101101111",
  36152=>"000000000",
  36153=>"000000000",
  36154=>"000000000",
  36155=>"000000111",
  36156=>"100111111",
  36157=>"000100111",
  36158=>"011111111",
  36159=>"111111000",
  36160=>"000111111",
  36161=>"111111111",
  36162=>"000000001",
  36163=>"000000000",
  36164=>"111100001",
  36165=>"100110000",
  36166=>"011111111",
  36167=>"111110111",
  36168=>"000000000",
  36169=>"000000000",
  36170=>"100000100",
  36171=>"100110010",
  36172=>"100111111",
  36173=>"111111111",
  36174=>"000001001",
  36175=>"001111111",
  36176=>"000001000",
  36177=>"001111111",
  36178=>"011011110",
  36179=>"000010010",
  36180=>"110111111",
  36181=>"111111011",
  36182=>"000000000",
  36183=>"111111111",
  36184=>"000000000",
  36185=>"111111000",
  36186=>"111111110",
  36187=>"000100100",
  36188=>"000000000",
  36189=>"100101111",
  36190=>"111111101",
  36191=>"111011001",
  36192=>"111111111",
  36193=>"011111111",
  36194=>"110100100",
  36195=>"111111011",
  36196=>"001001010",
  36197=>"000000000",
  36198=>"111111111",
  36199=>"110111111",
  36200=>"001011011",
  36201=>"110011001",
  36202=>"111100000",
  36203=>"000111111",
  36204=>"111111111",
  36205=>"001110110",
  36206=>"111000000",
  36207=>"000000100",
  36208=>"000000000",
  36209=>"000101111",
  36210=>"001001101",
  36211=>"100110111",
  36212=>"000000000",
  36213=>"000000000",
  36214=>"000000000",
  36215=>"000000001",
  36216=>"011011111",
  36217=>"000000000",
  36218=>"000000000",
  36219=>"000000000",
  36220=>"110100000",
  36221=>"000000001",
  36222=>"111111111",
  36223=>"111111101",
  36224=>"111011010",
  36225=>"111011011",
  36226=>"111111111",
  36227=>"000000000",
  36228=>"111011000",
  36229=>"000001000",
  36230=>"001111111",
  36231=>"011000000",
  36232=>"000000000",
  36233=>"110110100",
  36234=>"001001000",
  36235=>"000000000",
  36236=>"111111111",
  36237=>"001111111",
  36238=>"111111111",
  36239=>"000111111",
  36240=>"000000000",
  36241=>"000000000",
  36242=>"111111111",
  36243=>"001011111",
  36244=>"111111111",
  36245=>"000000000",
  36246=>"000000000",
  36247=>"010010000",
  36248=>"111110000",
  36249=>"010111000",
  36250=>"000011011",
  36251=>"011000000",
  36252=>"001000001",
  36253=>"110000010",
  36254=>"011001001",
  36255=>"000000000",
  36256=>"111101111",
  36257=>"111111110",
  36258=>"111110110",
  36259=>"011000011",
  36260=>"000011001",
  36261=>"000000111",
  36262=>"111001000",
  36263=>"000110010",
  36264=>"111111110",
  36265=>"000000000",
  36266=>"001011111",
  36267=>"101100100",
  36268=>"000000000",
  36269=>"001001001",
  36270=>"000000100",
  36271=>"111111111",
  36272=>"111111111",
  36273=>"111010011",
  36274=>"000000000",
  36275=>"000000000",
  36276=>"101111111",
  36277=>"000000000",
  36278=>"000111111",
  36279=>"000011111",
  36280=>"111000000",
  36281=>"000000000",
  36282=>"111101111",
  36283=>"111111110",
  36284=>"000000000",
  36285=>"100100011",
  36286=>"000100111",
  36287=>"100101101",
  36288=>"000111111",
  36289=>"000000000",
  36290=>"111111111",
  36291=>"000000000",
  36292=>"000000000",
  36293=>"011111111",
  36294=>"111111111",
  36295=>"000101001",
  36296=>"001000000",
  36297=>"000000000",
  36298=>"111011001",
  36299=>"111111111",
  36300=>"000000000",
  36301=>"000001000",
  36302=>"111111111",
  36303=>"000010010",
  36304=>"110110111",
  36305=>"001000000",
  36306=>"110110110",
  36307=>"111111011",
  36308=>"000000000",
  36309=>"111000001",
  36310=>"000011011",
  36311=>"110111111",
  36312=>"111111111",
  36313=>"101101001",
  36314=>"000000000",
  36315=>"000000000",
  36316=>"111110000",
  36317=>"000000000",
  36318=>"111111111",
  36319=>"100100101",
  36320=>"011110111",
  36321=>"111111001",
  36322=>"010110110",
  36323=>"000000000",
  36324=>"110111111",
  36325=>"000000000",
  36326=>"000000001",
  36327=>"000000000",
  36328=>"001001001",
  36329=>"001001111",
  36330=>"111100100",
  36331=>"000000100",
  36332=>"110111110",
  36333=>"111110110",
  36334=>"001001000",
  36335=>"000000000",
  36336=>"011111111",
  36337=>"111110110",
  36338=>"011011000",
  36339=>"010000000",
  36340=>"111111011",
  36341=>"000000000",
  36342=>"000000011",
  36343=>"001000000",
  36344=>"001111111",
  36345=>"001001001",
  36346=>"000000000",
  36347=>"001000000",
  36348=>"110000000",
  36349=>"011111111",
  36350=>"000100000",
  36351=>"111111111",
  36352=>"000000111",
  36353=>"000000010",
  36354=>"111101000",
  36355=>"111001000",
  36356=>"000000110",
  36357=>"111101000",
  36358=>"000000000",
  36359=>"110111111",
  36360=>"001001011",
  36361=>"010000000",
  36362=>"100000000",
  36363=>"100111111",
  36364=>"000000100",
  36365=>"001000000",
  36366=>"000010000",
  36367=>"101000000",
  36368=>"111111110",
  36369=>"000000010",
  36370=>"000000111",
  36371=>"111110000",
  36372=>"011011010",
  36373=>"000000101",
  36374=>"000000000",
  36375=>"001100001",
  36376=>"110110100",
  36377=>"101001001",
  36378=>"011011101",
  36379=>"100000000",
  36380=>"111111111",
  36381=>"100000101",
  36382=>"001001001",
  36383=>"100110000",
  36384=>"000000000",
  36385=>"000000000",
  36386=>"000000001",
  36387=>"110110110",
  36388=>"000000001",
  36389=>"000001001",
  36390=>"000000111",
  36391=>"111111011",
  36392=>"000000000",
  36393=>"000100110",
  36394=>"111111111",
  36395=>"000000000",
  36396=>"000001011",
  36397=>"000000000",
  36398=>"111111111",
  36399=>"111111111",
  36400=>"111001000",
  36401=>"000000111",
  36402=>"001000000",
  36403=>"111111011",
  36404=>"110010000",
  36405=>"001101111",
  36406=>"100110110",
  36407=>"000000000",
  36408=>"111111000",
  36409=>"111101101",
  36410=>"111111100",
  36411=>"110110100",
  36412=>"111001111",
  36413=>"110111111",
  36414=>"111111111",
  36415=>"111111111",
  36416=>"111100001",
  36417=>"111111111",
  36418=>"110000000",
  36419=>"111111001",
  36420=>"100000000",
  36421=>"101110111",
  36422=>"110100101",
  36423=>"111111111",
  36424=>"111111000",
  36425=>"000000111",
  36426=>"000100000",
  36427=>"011111111",
  36428=>"101101111",
  36429=>"000011110",
  36430=>"001000000",
  36431=>"000000000",
  36432=>"101111111",
  36433=>"110110100",
  36434=>"000000000",
  36435=>"000000000",
  36436=>"000000000",
  36437=>"111111111",
  36438=>"111100101",
  36439=>"111111111",
  36440=>"000000100",
  36441=>"000000000",
  36442=>"011111111",
  36443=>"011111111",
  36444=>"001111111",
  36445=>"000000000",
  36446=>"110011001",
  36447=>"111111111",
  36448=>"110000101",
  36449=>"000000000",
  36450=>"011111101",
  36451=>"000000101",
  36452=>"001000000",
  36453=>"101101111",
  36454=>"101101101",
  36455=>"000000000",
  36456=>"111111111",
  36457=>"000000111",
  36458=>"111100011",
  36459=>"001011011",
  36460=>"011111100",
  36461=>"001111111",
  36462=>"111111111",
  36463=>"110110110",
  36464=>"000000011",
  36465=>"000000000",
  36466=>"011000000",
  36467=>"111100100",
  36468=>"001101001",
  36469=>"001000000",
  36470=>"011001111",
  36471=>"101101001",
  36472=>"000000000",
  36473=>"101000000",
  36474=>"111110100",
  36475=>"011000000",
  36476=>"001001000",
  36477=>"110111000",
  36478=>"000111111",
  36479=>"000000000",
  36480=>"000000101",
  36481=>"010111011",
  36482=>"111111011",
  36483=>"000011000",
  36484=>"001001001",
  36485=>"111111111",
  36486=>"001001001",
  36487=>"001111111",
  36488=>"000000100",
  36489=>"000100000",
  36490=>"000000100",
  36491=>"001000111",
  36492=>"000110110",
  36493=>"111111100",
  36494=>"011000010",
  36495=>"000101111",
  36496=>"110111111",
  36497=>"111000000",
  36498=>"110000100",
  36499=>"001001001",
  36500=>"111111111",
  36501=>"111111110",
  36502=>"000001000",
  36503=>"111000000",
  36504=>"111110010",
  36505=>"111110000",
  36506=>"111111111",
  36507=>"111111111",
  36508=>"000000000",
  36509=>"001000000",
  36510=>"111111110",
  36511=>"000000100",
  36512=>"111000111",
  36513=>"101101111",
  36514=>"111010000",
  36515=>"000000000",
  36516=>"111000101",
  36517=>"110000110",
  36518=>"000000000",
  36519=>"001001001",
  36520=>"000000000",
  36521=>"000000000",
  36522=>"111001000",
  36523=>"111111101",
  36524=>"111001111",
  36525=>"110110000",
  36526=>"100000000",
  36527=>"101111111",
  36528=>"000000000",
  36529=>"001111100",
  36530=>"111111011",
  36531=>"000010000",
  36532=>"000110110",
  36533=>"001111111",
  36534=>"001000000",
  36535=>"111111111",
  36536=>"111111111",
  36537=>"111000000",
  36538=>"000000111",
  36539=>"111011011",
  36540=>"010110110",
  36541=>"000000000",
  36542=>"000000110",
  36543=>"111111111",
  36544=>"000000100",
  36545=>"110111011",
  36546=>"101001101",
  36547=>"000000000",
  36548=>"011111111",
  36549=>"000101111",
  36550=>"111111110",
  36551=>"000000000",
  36552=>"000100000",
  36553=>"111000000",
  36554=>"000000000",
  36555=>"000110111",
  36556=>"111101001",
  36557=>"000001100",
  36558=>"011001000",
  36559=>"111101000",
  36560=>"010111111",
  36561=>"000000000",
  36562=>"000000000",
  36563=>"000000000",
  36564=>"001001001",
  36565=>"001001001",
  36566=>"000000000",
  36567=>"000001111",
  36568=>"101111101",
  36569=>"111111111",
  36570=>"000000111",
  36571=>"110000011",
  36572=>"000110110",
  36573=>"001001111",
  36574=>"111111111",
  36575=>"011000000",
  36576=>"000000000",
  36577=>"000000000",
  36578=>"000000000",
  36579=>"000000011",
  36580=>"000110110",
  36581=>"111100011",
  36582=>"111000000",
  36583=>"011001000",
  36584=>"111010000",
  36585=>"011111110",
  36586=>"110111111",
  36587=>"101101111",
  36588=>"111101100",
  36589=>"111111110",
  36590=>"111111111",
  36591=>"111001000",
  36592=>"111111111",
  36593=>"111111111",
  36594=>"000000000",
  36595=>"000000110",
  36596=>"000001111",
  36597=>"111110110",
  36598=>"111111111",
  36599=>"000000000",
  36600=>"111001000",
  36601=>"000000000",
  36602=>"000000000",
  36603=>"000011011",
  36604=>"000000100",
  36605=>"101111111",
  36606=>"111000001",
  36607=>"000111111",
  36608=>"100000001",
  36609=>"110000000",
  36610=>"000000000",
  36611=>"101001000",
  36612=>"000111110",
  36613=>"000000000",
  36614=>"111111111",
  36615=>"011011001",
  36616=>"110110111",
  36617=>"111111111",
  36618=>"111111110",
  36619=>"001011011",
  36620=>"111111111",
  36621=>"111000000",
  36622=>"111111111",
  36623=>"110110000",
  36624=>"111111111",
  36625=>"101001001",
  36626=>"011011000",
  36627=>"000000111",
  36628=>"111000000",
  36629=>"111111111",
  36630=>"110110110",
  36631=>"111110000",
  36632=>"111101111",
  36633=>"000111111",
  36634=>"111111011",
  36635=>"100000000",
  36636=>"000001000",
  36637=>"001000100",
  36638=>"000010111",
  36639=>"101110111",
  36640=>"000000000",
  36641=>"000110111",
  36642=>"110100101",
  36643=>"111111110",
  36644=>"111001001",
  36645=>"111011011",
  36646=>"001001001",
  36647=>"000000100",
  36648=>"001001001",
  36649=>"001000000",
  36650=>"100000100",
  36651=>"000000000",
  36652=>"111011011",
  36653=>"110000100",
  36654=>"111000111",
  36655=>"000000001",
  36656=>"100110111",
  36657=>"000000111",
  36658=>"000100111",
  36659=>"001111111",
  36660=>"111111110",
  36661=>"000001011",
  36662=>"001000000",
  36663=>"101000000",
  36664=>"000000000",
  36665=>"001000000",
  36666=>"111011011",
  36667=>"011111000",
  36668=>"101100111",
  36669=>"001001111",
  36670=>"101101001",
  36671=>"000000010",
  36672=>"000000111",
  36673=>"001000000",
  36674=>"000000110",
  36675=>"000000000",
  36676=>"001011001",
  36677=>"111000101",
  36678=>"000000000",
  36679=>"100111111",
  36680=>"111111111",
  36681=>"000010110",
  36682=>"001000000",
  36683=>"000000000",
  36684=>"111111111",
  36685=>"000100000",
  36686=>"111100111",
  36687=>"101101000",
  36688=>"001001011",
  36689=>"000000000",
  36690=>"001001000",
  36691=>"110000000",
  36692=>"111001101",
  36693=>"011011001",
  36694=>"001000000",
  36695=>"111111111",
  36696=>"001001011",
  36697=>"111111111",
  36698=>"111111111",
  36699=>"010000110",
  36700=>"111000000",
  36701=>"111111111",
  36702=>"101101101",
  36703=>"111110110",
  36704=>"000100111",
  36705=>"111111111",
  36706=>"101100110",
  36707=>"000000000",
  36708=>"000000111",
  36709=>"000101100",
  36710=>"000111111",
  36711=>"111111111",
  36712=>"000000010",
  36713=>"111111110",
  36714=>"011001001",
  36715=>"101101000",
  36716=>"100010000",
  36717=>"110110010",
  36718=>"000000000",
  36719=>"111001111",
  36720=>"000000000",
  36721=>"011001001",
  36722=>"000001111",
  36723=>"100111101",
  36724=>"001001001",
  36725=>"000111111",
  36726=>"000000000",
  36727=>"110110000",
  36728=>"011111111",
  36729=>"000001000",
  36730=>"000000000",
  36731=>"111111111",
  36732=>"110000100",
  36733=>"000000000",
  36734=>"000000000",
  36735=>"000000000",
  36736=>"100110100",
  36737=>"001001001",
  36738=>"111111011",
  36739=>"000111111",
  36740=>"000000000",
  36741=>"110110000",
  36742=>"000000000",
  36743=>"000001111",
  36744=>"000000000",
  36745=>"111111111",
  36746=>"111111111",
  36747=>"110110000",
  36748=>"100110111",
  36749=>"100110100",
  36750=>"110111110",
  36751=>"000000000",
  36752=>"000000000",
  36753=>"111111111",
  36754=>"111011010",
  36755=>"000000111",
  36756=>"111111111",
  36757=>"000010000",
  36758=>"000000001",
  36759=>"110111110",
  36760=>"001111111",
  36761=>"100111111",
  36762=>"000000000",
  36763=>"001000000",
  36764=>"011000000",
  36765=>"000000001",
  36766=>"000000000",
  36767=>"001001001",
  36768=>"110011011",
  36769=>"011111100",
  36770=>"000000100",
  36771=>"001001000",
  36772=>"000000111",
  36773=>"000000000",
  36774=>"000110011",
  36775=>"010111111",
  36776=>"000011101",
  36777=>"110100111",
  36778=>"110010010",
  36779=>"000000011",
  36780=>"000000000",
  36781=>"111111111",
  36782=>"101101101",
  36783=>"111111111",
  36784=>"111111111",
  36785=>"000001001",
  36786=>"000000000",
  36787=>"000011001",
  36788=>"100000000",
  36789=>"001001111",
  36790=>"111100100",
  36791=>"000000000",
  36792=>"111111111",
  36793=>"000011101",
  36794=>"011111111",
  36795=>"110010011",
  36796=>"011000000",
  36797=>"000010111",
  36798=>"000000000",
  36799=>"110100100",
  36800=>"101111011",
  36801=>"111111111",
  36802=>"000000000",
  36803=>"000000101",
  36804=>"111111111",
  36805=>"111001111",
  36806=>"000000101",
  36807=>"000000110",
  36808=>"111000110",
  36809=>"111001000",
  36810=>"101000000",
  36811=>"000010110",
  36812=>"111001000",
  36813=>"000000000",
  36814=>"000000000",
  36815=>"111111111",
  36816=>"111111011",
  36817=>"000000000",
  36818=>"000000001",
  36819=>"000000001",
  36820=>"110111111",
  36821=>"111111001",
  36822=>"001000111",
  36823=>"110000000",
  36824=>"000000000",
  36825=>"011111110",
  36826=>"111000111",
  36827=>"101111111",
  36828=>"000000000",
  36829=>"101111111",
  36830=>"000000111",
  36831=>"110111110",
  36832=>"001001100",
  36833=>"111111111",
  36834=>"111111111",
  36835=>"111011010",
  36836=>"111111111",
  36837=>"111111111",
  36838=>"110111111",
  36839=>"000001001",
  36840=>"100000100",
  36841=>"000000000",
  36842=>"111000100",
  36843=>"111111111",
  36844=>"111111111",
  36845=>"111111011",
  36846=>"000111111",
  36847=>"111111111",
  36848=>"000000000",
  36849=>"100000000",
  36850=>"111111011",
  36851=>"010111000",
  36852=>"111111011",
  36853=>"011011000",
  36854=>"001001101",
  36855=>"110111111",
  36856=>"011001011",
  36857=>"011001001",
  36858=>"100100100",
  36859=>"111000111",
  36860=>"110110111",
  36861=>"100000000",
  36862=>"100100110",
  36863=>"001111111",
  36864=>"111111111",
  36865=>"111111011",
  36866=>"101111111",
  36867=>"111111011",
  36868=>"011011011",
  36869=>"110011011",
  36870=>"000010111",
  36871=>"111010100",
  36872=>"000100111",
  36873=>"000000001",
  36874=>"111111111",
  36875=>"000000011",
  36876=>"000111111",
  36877=>"110000011",
  36878=>"111011011",
  36879=>"111010010",
  36880=>"000000000",
  36881=>"000000000",
  36882=>"000000000",
  36883=>"000000000",
  36884=>"011110100",
  36885=>"111001101",
  36886=>"101101001",
  36887=>"001001001",
  36888=>"000000100",
  36889=>"001001001",
  36890=>"011000000",
  36891=>"111111111",
  36892=>"100000000",
  36893=>"000001001",
  36894=>"000100111",
  36895=>"111110000",
  36896=>"100111000",
  36897=>"111000000",
  36898=>"100111111",
  36899=>"111111000",
  36900=>"010000000",
  36901=>"000000000",
  36902=>"000000111",
  36903=>"000000000",
  36904=>"001001011",
  36905=>"111111111",
  36906=>"001011111",
  36907=>"000000100",
  36908=>"110111110",
  36909=>"111000000",
  36910=>"111011000",
  36911=>"111001000",
  36912=>"000011011",
  36913=>"010111011",
  36914=>"000000010",
  36915=>"001011011",
  36916=>"011111000",
  36917=>"001101111",
  36918=>"000000000",
  36919=>"001001100",
  36920=>"111111111",
  36921=>"001011111",
  36922=>"011111111",
  36923=>"011000000",
  36924=>"001000000",
  36925=>"100100000",
  36926=>"111100101",
  36927=>"000000000",
  36928=>"000111111",
  36929=>"111111100",
  36930=>"011000000",
  36931=>"011011011",
  36932=>"100000000",
  36933=>"010011000",
  36934=>"110000110",
  36935=>"100100000",
  36936=>"100110111",
  36937=>"000000000",
  36938=>"111111111",
  36939=>"101111101",
  36940=>"101000000",
  36941=>"011010011",
  36942=>"000110110",
  36943=>"111011000",
  36944=>"110010000",
  36945=>"100000000",
  36946=>"011111111",
  36947=>"111110110",
  36948=>"001000000",
  36949=>"000010000",
  36950=>"000001001",
  36951=>"000000000",
  36952=>"000011000",
  36953=>"000000100",
  36954=>"000000000",
  36955=>"110110110",
  36956=>"111110110",
  36957=>"000000000",
  36958=>"000000000",
  36959=>"100100110",
  36960=>"101101101",
  36961=>"000000000",
  36962=>"011011011",
  36963=>"111101001",
  36964=>"000000010",
  36965=>"111110000",
  36966=>"111111111",
  36967=>"111111111",
  36968=>"001111111",
  36969=>"001011111",
  36970=>"111111111",
  36971=>"000000000",
  36972=>"111111000",
  36973=>"011111111",
  36974=>"001000000",
  36975=>"100111111",
  36976=>"001001000",
  36977=>"000000111",
  36978=>"111110110",
  36979=>"111111010",
  36980=>"000000000",
  36981=>"111111111",
  36982=>"000000100",
  36983=>"001011010",
  36984=>"110110110",
  36985=>"000011000",
  36986=>"111111111",
  36987=>"000000000",
  36988=>"000000000",
  36989=>"001001111",
  36990=>"011111111",
  36991=>"001001010",
  36992=>"001000000",
  36993=>"001001000",
  36994=>"000110000",
  36995=>"000001000",
  36996=>"111111111",
  36997=>"001101111",
  36998=>"001011001",
  36999=>"000000111",
  37000=>"111111111",
  37001=>"111111001",
  37002=>"111110110",
  37003=>"000000000",
  37004=>"101000010",
  37005=>"000001011",
  37006=>"111111111",
  37007=>"000000001",
  37008=>"111111111",
  37009=>"000000000",
  37010=>"000010000",
  37011=>"000100111",
  37012=>"011011011",
  37013=>"000000000",
  37014=>"111111111",
  37015=>"000000000",
  37016=>"111110111",
  37017=>"111111111",
  37018=>"000000110",
  37019=>"000000000",
  37020=>"011111111",
  37021=>"001000000",
  37022=>"111000000",
  37023=>"000000000",
  37024=>"111111111",
  37025=>"000001111",
  37026=>"001001000",
  37027=>"111110110",
  37028=>"011011010",
  37029=>"000010000",
  37030=>"111111111",
  37031=>"111011111",
  37032=>"000011000",
  37033=>"000000000",
  37034=>"011011000",
  37035=>"101001011",
  37036=>"000110000",
  37037=>"001001000",
  37038=>"000111111",
  37039=>"111111000",
  37040=>"111010000",
  37041=>"000100100",
  37042=>"111111111",
  37043=>"111111111",
  37044=>"001001000",
  37045=>"100000000",
  37046=>"000001011",
  37047=>"001000101",
  37048=>"111111110",
  37049=>"111111111",
  37050=>"110000000",
  37051=>"100111111",
  37052=>"111000000",
  37053=>"111111111",
  37054=>"111100001",
  37055=>"111001000",
  37056=>"010011111",
  37057=>"011000000",
  37058=>"001000000",
  37059=>"100000000",
  37060=>"110110010",
  37061=>"000000000",
  37062=>"000000100",
  37063=>"000000111",
  37064=>"111111111",
  37065=>"000000000",
  37066=>"000010011",
  37067=>"111111111",
  37068=>"100000000",
  37069=>"000110111",
  37070=>"011011011",
  37071=>"000000000",
  37072=>"000000000",
  37073=>"011011111",
  37074=>"000000000",
  37075=>"001011011",
  37076=>"101111011",
  37077=>"000000000",
  37078=>"000000001",
  37079=>"010111111",
  37080=>"111111111",
  37081=>"000000111",
  37082=>"000000000",
  37083=>"110110110",
  37084=>"000000001",
  37085=>"000000001",
  37086=>"111111111",
  37087=>"111111100",
  37088=>"000000000",
  37089=>"011011000",
  37090=>"000000000",
  37091=>"000001111",
  37092=>"000000000",
  37093=>"000111111",
  37094=>"000100111",
  37095=>"000000111",
  37096=>"111111111",
  37097=>"111111111",
  37098=>"000000000",
  37099=>"111000100",
  37100=>"110111111",
  37101=>"000110111",
  37102=>"101111111",
  37103=>"000000000",
  37104=>"100111100",
  37105=>"000000101",
  37106=>"000000000",
  37107=>"010111000",
  37108=>"001101111",
  37109=>"001001001",
  37110=>"100100100",
  37111=>"000001111",
  37112=>"111111001",
  37113=>"000000000",
  37114=>"000000010",
  37115=>"111111011",
  37116=>"000000000",
  37117=>"011001111",
  37118=>"000011001",
  37119=>"011111111",
  37120=>"111111011",
  37121=>"001001011",
  37122=>"111110111",
  37123=>"111011111",
  37124=>"001000110",
  37125=>"000110110",
  37126=>"111111111",
  37127=>"001011111",
  37128=>"000010010",
  37129=>"111110011",
  37130=>"000000001",
  37131=>"111111111",
  37132=>"111000000",
  37133=>"000000000",
  37134=>"000000111",
  37135=>"000000000",
  37136=>"000000010",
  37137=>"000000000",
  37138=>"000000000",
  37139=>"110000001",
  37140=>"011011011",
  37141=>"000100000",
  37142=>"000000111",
  37143=>"000110000",
  37144=>"111111011",
  37145=>"000000000",
  37146=>"000000000",
  37147=>"010000110",
  37148=>"011011000",
  37149=>"000000111",
  37150=>"001001001",
  37151=>"110000000",
  37152=>"101101111",
  37153=>"111111111",
  37154=>"000000000",
  37155=>"000000000",
  37156=>"111111111",
  37157=>"000110111",
  37158=>"000000000",
  37159=>"000010011",
  37160=>"000110011",
  37161=>"010000000",
  37162=>"000111011",
  37163=>"000101111",
  37164=>"000111111",
  37165=>"100001011",
  37166=>"000000100",
  37167=>"000000000",
  37168=>"011001000",
  37169=>"011000000",
  37170=>"111111111",
  37171=>"001000001",
  37172=>"000010000",
  37173=>"110111110",
  37174=>"000000001",
  37175=>"100100110",
  37176=>"111111000",
  37177=>"111010000",
  37178=>"111000011",
  37179=>"001000000",
  37180=>"110111111",
  37181=>"101000001",
  37182=>"011001000",
  37183=>"111111110",
  37184=>"000001101",
  37185=>"000000000",
  37186=>"100101110",
  37187=>"000000000",
  37188=>"011011011",
  37189=>"000000000",
  37190=>"000000000",
  37191=>"111111110",
  37192=>"110111111",
  37193=>"000000000",
  37194=>"011010010",
  37195=>"100101101",
  37196=>"100000100",
  37197=>"000000010",
  37198=>"000000000",
  37199=>"000100100",
  37200=>"111111111",
  37201=>"000000000",
  37202=>"000000000",
  37203=>"111001000",
  37204=>"001000000",
  37205=>"011011011",
  37206=>"000000010",
  37207=>"100000000",
  37208=>"000000000",
  37209=>"111111010",
  37210=>"000001001",
  37211=>"011111000",
  37212=>"000000000",
  37213=>"111111111",
  37214=>"000000000",
  37215=>"110111111",
  37216=>"100000000",
  37217=>"110111000",
  37218=>"110111111",
  37219=>"000000000",
  37220=>"110111111",
  37221=>"000000000",
  37222=>"000000000",
  37223=>"000011111",
  37224=>"100110110",
  37225=>"111111100",
  37226=>"000000000",
  37227=>"000001111",
  37228=>"001000000",
  37229=>"111011000",
  37230=>"011011111",
  37231=>"100100100",
  37232=>"000000000",
  37233=>"000111010",
  37234=>"111000000",
  37235=>"111001000",
  37236=>"111111111",
  37237=>"000000000",
  37238=>"000111111",
  37239=>"111111111",
  37240=>"111111111",
  37241=>"001110111",
  37242=>"000000000",
  37243=>"111111111",
  37244=>"000000010",
  37245=>"111001011",
  37246=>"000000000",
  37247=>"100111111",
  37248=>"000000000",
  37249=>"111111111",
  37250=>"011011011",
  37251=>"111001000",
  37252=>"000000000",
  37253=>"011111011",
  37254=>"100110111",
  37255=>"001000000",
  37256=>"111111111",
  37257=>"000000011",
  37258=>"010000000",
  37259=>"111000000",
  37260=>"000100101",
  37261=>"111011000",
  37262=>"000011010",
  37263=>"000010010",
  37264=>"000010010",
  37265=>"000100100",
  37266=>"000000000",
  37267=>"000001011",
  37268=>"111111100",
  37269=>"000000000",
  37270=>"011111110",
  37271=>"011011011",
  37272=>"111111111",
  37273=>"000000001",
  37274=>"011010110",
  37275=>"001001111",
  37276=>"000110110",
  37277=>"000101111",
  37278=>"000100111",
  37279=>"000000000",
  37280=>"000000000",
  37281=>"011011011",
  37282=>"111111111",
  37283=>"011111111",
  37284=>"101111110",
  37285=>"111111111",
  37286=>"000110010",
  37287=>"100110110",
  37288=>"110000000",
  37289=>"000000000",
  37290=>"111111100",
  37291=>"000000100",
  37292=>"000011011",
  37293=>"000010010",
  37294=>"000000000",
  37295=>"000010110",
  37296=>"000000100",
  37297=>"000000010",
  37298=>"000000111",
  37299=>"000000000",
  37300=>"111111111",
  37301=>"100000110",
  37302=>"001100100",
  37303=>"111111000",
  37304=>"111111111",
  37305=>"101101011",
  37306=>"011000011",
  37307=>"111110000",
  37308=>"111111011",
  37309=>"011011111",
  37310=>"000101100",
  37311=>"111101110",
  37312=>"000000000",
  37313=>"100111111",
  37314=>"111111111",
  37315=>"000110000",
  37316=>"000001000",
  37317=>"111101001",
  37318=>"000000000",
  37319=>"000100000",
  37320=>"100000000",
  37321=>"001000110",
  37322=>"000000000",
  37323=>"011010010",
  37324=>"111110000",
  37325=>"000100000",
  37326=>"111000001",
  37327=>"111111100",
  37328=>"000010111",
  37329=>"100100111",
  37330=>"100100100",
  37331=>"010110111",
  37332=>"111110110",
  37333=>"001011111",
  37334=>"011011011",
  37335=>"000101001",
  37336=>"000000000",
  37337=>"100000100",
  37338=>"111111111",
  37339=>"000111111",
  37340=>"111111111",
  37341=>"110100111",
  37342=>"111111111",
  37343=>"111111111",
  37344=>"111000000",
  37345=>"000000000",
  37346=>"111011011",
  37347=>"111101100",
  37348=>"111111011",
  37349=>"111111000",
  37350=>"101001111",
  37351=>"000000000",
  37352=>"010000000",
  37353=>"000000000",
  37354=>"000000000",
  37355=>"010011010",
  37356=>"000000110",
  37357=>"111111111",
  37358=>"111111111",
  37359=>"111111111",
  37360=>"110110001",
  37361=>"000000000",
  37362=>"000000000",
  37363=>"000011110",
  37364=>"111111011",
  37365=>"100000000",
  37366=>"000000100",
  37367=>"100110100",
  37368=>"000001111",
  37369=>"010011111",
  37370=>"111111011",
  37371=>"000001111",
  37372=>"100111111",
  37373=>"000000000",
  37374=>"100111010",
  37375=>"110111111",
  37376=>"111111111",
  37377=>"000000000",
  37378=>"000000000",
  37379=>"111000000",
  37380=>"110111111",
  37381=>"110111000",
  37382=>"011001111",
  37383=>"111111111",
  37384=>"111111111",
  37385=>"001101000",
  37386=>"001000000",
  37387=>"111100000",
  37388=>"000110100",
  37389=>"111111111",
  37390=>"000001111",
  37391=>"000011011",
  37392=>"000101000",
  37393=>"000000111",
  37394=>"001011011",
  37395=>"111111000",
  37396=>"100101000",
  37397=>"000000000",
  37398=>"001001000",
  37399=>"000100000",
  37400=>"000000100",
  37401=>"000100001",
  37402=>"000100111",
  37403=>"000000011",
  37404=>"000000111",
  37405=>"000000000",
  37406=>"000111110",
  37407=>"111111000",
  37408=>"101011011",
  37409=>"000100110",
  37410=>"000000100",
  37411=>"000011111",
  37412=>"111111110",
  37413=>"000000000",
  37414=>"011011000",
  37415=>"111111111",
  37416=>"001000000",
  37417=>"000000001",
  37418=>"001001000",
  37419=>"111111111",
  37420=>"111111111",
  37421=>"111011010",
  37422=>"001001011",
  37423=>"000000000",
  37424=>"000000000",
  37425=>"000010010",
  37426=>"100100001",
  37427=>"011001000",
  37428=>"000000000",
  37429=>"100100000",
  37430=>"111111011",
  37431=>"000101001",
  37432=>"111111111",
  37433=>"000000100",
  37434=>"000000000",
  37435=>"111111111",
  37436=>"000000000",
  37437=>"001111001",
  37438=>"111111011",
  37439=>"001111001",
  37440=>"000000000",
  37441=>"100111111",
  37442=>"111110100",
  37443=>"001000000",
  37444=>"111111111",
  37445=>"001011011",
  37446=>"000000111",
  37447=>"000011000",
  37448=>"000001111",
  37449=>"000000000",
  37450=>"000001001",
  37451=>"010000001",
  37452=>"111111111",
  37453=>"011011110",
  37454=>"000000000",
  37455=>"011000111",
  37456=>"000000001",
  37457=>"100111111",
  37458=>"000111111",
  37459=>"101001110",
  37460=>"001111111",
  37461=>"111000000",
  37462=>"000111011",
  37463=>"110101111",
  37464=>"000000000",
  37465=>"111111111",
  37466=>"111110000",
  37467=>"100100111",
  37468=>"000000000",
  37469=>"100100101",
  37470=>"111100100",
  37471=>"111111011",
  37472=>"111000000",
  37473=>"011000000",
  37474=>"111111111",
  37475=>"000000000",
  37476=>"110111100",
  37477=>"101000000",
  37478=>"111111111",
  37479=>"000001001",
  37480=>"001001000",
  37481=>"000000111",
  37482=>"001111111",
  37483=>"001111001",
  37484=>"111111100",
  37485=>"000000000",
  37486=>"000000000",
  37487=>"101000001",
  37488=>"111111111",
  37489=>"111111101",
  37490=>"000111111",
  37491=>"000000000",
  37492=>"001000000",
  37493=>"000000111",
  37494=>"100100111",
  37495=>"000010010",
  37496=>"010000000",
  37497=>"101100100",
  37498=>"000011000",
  37499=>"111000000",
  37500=>"000110110",
  37501=>"000000100",
  37502=>"011001011",
  37503=>"000100110",
  37504=>"000001001",
  37505=>"100000000",
  37506=>"000000111",
  37507=>"011111111",
  37508=>"000000000",
  37509=>"000000111",
  37510=>"111000000",
  37511=>"000000000",
  37512=>"000000000",
  37513=>"110000101",
  37514=>"000000000",
  37515=>"100111111",
  37516=>"111111101",
  37517=>"000001101",
  37518=>"000000000",
  37519=>"000000000",
  37520=>"111111000",
  37521=>"100111111",
  37522=>"111111111",
  37523=>"000000010",
  37524=>"100100111",
  37525=>"000000000",
  37526=>"111111111",
  37527=>"111000000",
  37528=>"000000100",
  37529=>"111111001",
  37530=>"001011011",
  37531=>"000000000",
  37532=>"111011111",
  37533=>"000000000",
  37534=>"000100000",
  37535=>"000000111",
  37536=>"001000111",
  37537=>"111111000",
  37538=>"000000001",
  37539=>"000000000",
  37540=>"100100000",
  37541=>"000000000",
  37542=>"000111111",
  37543=>"000000100",
  37544=>"111111111",
  37545=>"001000000",
  37546=>"000000000",
  37547=>"001111111",
  37548=>"000000101",
  37549=>"111111111",
  37550=>"111111111",
  37551=>"000000000",
  37552=>"000111111",
  37553=>"011011111",
  37554=>"111111111",
  37555=>"000100000",
  37556=>"111111011",
  37557=>"111011111",
  37558=>"111111111",
  37559=>"111000000",
  37560=>"000000000",
  37561=>"111111000",
  37562=>"000100100",
  37563=>"001010111",
  37564=>"111111100",
  37565=>"111111111",
  37566=>"111111011",
  37567=>"000000001",
  37568=>"001000000",
  37569=>"000110110",
  37570=>"000000001",
  37571=>"111111111",
  37572=>"110111010",
  37573=>"000000110",
  37574=>"000000000",
  37575=>"111111111",
  37576=>"111111100",
  37577=>"000000000",
  37578=>"001101001",
  37579=>"000000101",
  37580=>"000000000",
  37581=>"000000111",
  37582=>"000000000",
  37583=>"000000000",
  37584=>"001000000",
  37585=>"000000000",
  37586=>"001000011",
  37587=>"111111110",
  37588=>"110111101",
  37589=>"111111000",
  37590=>"110111111",
  37591=>"000000100",
  37592=>"000111011",
  37593=>"000110110",
  37594=>"000110100",
  37595=>"000000000",
  37596=>"111111001",
  37597=>"111111111",
  37598=>"000000000",
  37599=>"001001000",
  37600=>"000000000",
  37601=>"000000111",
  37602=>"111111111",
  37603=>"001111011",
  37604=>"000001011",
  37605=>"001000000",
  37606=>"111111111",
  37607=>"000000000",
  37608=>"000001000",
  37609=>"000000000",
  37610=>"101111111",
  37611=>"111001001",
  37612=>"000000001",
  37613=>"111111111",
  37614=>"110111111",
  37615=>"000001111",
  37616=>"011011001",
  37617=>"000000000",
  37618=>"000000000",
  37619=>"110100101",
  37620=>"111111111",
  37621=>"111110110",
  37622=>"000001000",
  37623=>"111111111",
  37624=>"111111111",
  37625=>"000000000",
  37626=>"000110110",
  37627=>"010000000",
  37628=>"111111000",
  37629=>"001111111",
  37630=>"111001001",
  37631=>"000100000",
  37632=>"110110110",
  37633=>"110100110",
  37634=>"011010110",
  37635=>"100000100",
  37636=>"111000000",
  37637=>"001001111",
  37638=>"111100000",
  37639=>"000001001",
  37640=>"000000100",
  37641=>"111000000",
  37642=>"001111011",
  37643=>"000000001",
  37644=>"000000000",
  37645=>"110110010",
  37646=>"111111111",
  37647=>"111111000",
  37648=>"000000000",
  37649=>"000001000",
  37650=>"100000000",
  37651=>"000000000",
  37652=>"111101111",
  37653=>"111111001",
  37654=>"110111111",
  37655=>"111111001",
  37656=>"000011111",
  37657=>"100111001",
  37658=>"011011000",
  37659=>"111111111",
  37660=>"001111111",
  37661=>"000111111",
  37662=>"111000000",
  37663=>"111111111",
  37664=>"111101000",
  37665=>"111111111",
  37666=>"111111000",
  37667=>"111101100",
  37668=>"000000000",
  37669=>"000000000",
  37670=>"000000000",
  37671=>"110000000",
  37672=>"000110110",
  37673=>"000000000",
  37674=>"000011111",
  37675=>"111000000",
  37676=>"000000000",
  37677=>"000011000",
  37678=>"101000111",
  37679=>"111111111",
  37680=>"000111101",
  37681=>"100111000",
  37682=>"001000111",
  37683=>"000110011",
  37684=>"111000000",
  37685=>"001000110",
  37686=>"000000000",
  37687=>"000000000",
  37688=>"111111111",
  37689=>"000101111",
  37690=>"001001000",
  37691=>"000000000",
  37692=>"111111111",
  37693=>"000000000",
  37694=>"111001001",
  37695=>"011001000",
  37696=>"111000000",
  37697=>"000000000",
  37698=>"110110010",
  37699=>"100100101",
  37700=>"000001000",
  37701=>"000000001",
  37702=>"000000000",
  37703=>"111101101",
  37704=>"000000000",
  37705=>"000000000",
  37706=>"111000000",
  37707=>"001011011",
  37708=>"100111111",
  37709=>"000000000",
  37710=>"000000110",
  37711=>"000110111",
  37712=>"111101101",
  37713=>"111111111",
  37714=>"111111111",
  37715=>"000000000",
  37716=>"000000000",
  37717=>"011111011",
  37718=>"000000000",
  37719=>"100100101",
  37720=>"001011001",
  37721=>"100000101",
  37722=>"111011000",
  37723=>"000000000",
  37724=>"110111000",
  37725=>"111111111",
  37726=>"111111011",
  37727=>"000100110",
  37728=>"111111000",
  37729=>"111001011",
  37730=>"101100000",
  37731=>"000111111",
  37732=>"111011011",
  37733=>"001001000",
  37734=>"000000000",
  37735=>"110110111",
  37736=>"000100100",
  37737=>"000000100",
  37738=>"000000000",
  37739=>"000001111",
  37740=>"100101110",
  37741=>"000000000",
  37742=>"111111110",
  37743=>"111111111",
  37744=>"101000000",
  37745=>"111000000",
  37746=>"100001101",
  37747=>"000000011",
  37748=>"000000000",
  37749=>"011011011",
  37750=>"110111111",
  37751=>"100000000",
  37752=>"000001001",
  37753=>"011100111",
  37754=>"000000000",
  37755=>"100100100",
  37756=>"011010011",
  37757=>"111000100",
  37758=>"000111111",
  37759=>"110111111",
  37760=>"000100100",
  37761=>"111111111",
  37762=>"111111010",
  37763=>"111111001",
  37764=>"000100111",
  37765=>"111111111",
  37766=>"100000001",
  37767=>"100010000",
  37768=>"111111001",
  37769=>"000000000",
  37770=>"111111101",
  37771=>"000000001",
  37772=>"111111111",
  37773=>"000001011",
  37774=>"000111000",
  37775=>"000000000",
  37776=>"111111111",
  37777=>"110100110",
  37778=>"100000000",
  37779=>"110110111",
  37780=>"111111111",
  37781=>"000000000",
  37782=>"110100000",
  37783=>"110100000",
  37784=>"111101001",
  37785=>"100100101",
  37786=>"000000001",
  37787=>"111111101",
  37788=>"000000000",
  37789=>"111111111",
  37790=>"101001001",
  37791=>"000000000",
  37792=>"000000001",
  37793=>"100101111",
  37794=>"111111111",
  37795=>"000000000",
  37796=>"000000000",
  37797=>"010111111",
  37798=>"000000000",
  37799=>"111111111",
  37800=>"100000000",
  37801=>"111000000",
  37802=>"000000000",
  37803=>"111111110",
  37804=>"000000000",
  37805=>"111111000",
  37806=>"010011011",
  37807=>"001000100",
  37808=>"100100000",
  37809=>"000000000",
  37810=>"000000000",
  37811=>"111110000",
  37812=>"111110000",
  37813=>"001101110",
  37814=>"100101111",
  37815=>"111110111",
  37816=>"000000001",
  37817=>"110111111",
  37818=>"000000000",
  37819=>"111000000",
  37820=>"000000000",
  37821=>"111111101",
  37822=>"000111010",
  37823=>"000101111",
  37824=>"111110100",
  37825=>"111000000",
  37826=>"100000000",
  37827=>"111111000",
  37828=>"110101000",
  37829=>"000000000",
  37830=>"000000000",
  37831=>"000000000",
  37832=>"111111111",
  37833=>"111111111",
  37834=>"100000111",
  37835=>"000000111",
  37836=>"000000000",
  37837=>"111111111",
  37838=>"111111111",
  37839=>"000000000",
  37840=>"000111000",
  37841=>"000000000",
  37842=>"000000000",
  37843=>"000000001",
  37844=>"011111111",
  37845=>"000111111",
  37846=>"001000000",
  37847=>"000000010",
  37848=>"000111111",
  37849=>"011000000",
  37850=>"110110000",
  37851=>"011010110",
  37852=>"111111001",
  37853=>"000000000",
  37854=>"000000000",
  37855=>"100100000",
  37856=>"000000000",
  37857=>"010000000",
  37858=>"111111010",
  37859=>"000100000",
  37860=>"110100100",
  37861=>"000000011",
  37862=>"010000000",
  37863=>"011111111",
  37864=>"000111111",
  37865=>"001000000",
  37866=>"000000100",
  37867=>"100110111",
  37868=>"100000000",
  37869=>"111110100",
  37870=>"111111000",
  37871=>"110001010",
  37872=>"111000000",
  37873=>"100010000",
  37874=>"000000001",
  37875=>"110111101",
  37876=>"011001000",
  37877=>"111111111",
  37878=>"000000101",
  37879=>"001001000",
  37880=>"111111111",
  37881=>"001001011",
  37882=>"001111000",
  37883=>"111000000",
  37884=>"100000110",
  37885=>"010111111",
  37886=>"111111111",
  37887=>"100100110",
  37888=>"000000000",
  37889=>"001000000",
  37890=>"111000001",
  37891=>"111111111",
  37892=>"000100111",
  37893=>"111010100",
  37894=>"111111001",
  37895=>"111111111",
  37896=>"111111110",
  37897=>"111000000",
  37898=>"001111111",
  37899=>"111001101",
  37900=>"000100110",
  37901=>"111001000",
  37902=>"000000000",
  37903=>"000000010",
  37904=>"100111111",
  37905=>"000000111",
  37906=>"010000100",
  37907=>"111000000",
  37908=>"000010000",
  37909=>"000100000",
  37910=>"111111001",
  37911=>"111100100",
  37912=>"100110110",
  37913=>"000001111",
  37914=>"000000000",
  37915=>"100100100",
  37916=>"111100111",
  37917=>"101111111",
  37918=>"000100100",
  37919=>"111111111",
  37920=>"000010000",
  37921=>"000001111",
  37922=>"110100000",
  37923=>"000111111",
  37924=>"111111110",
  37925=>"111011000",
  37926=>"111111101",
  37927=>"011101111",
  37928=>"111111111",
  37929=>"000101001",
  37930=>"111000000",
  37931=>"111111111",
  37932=>"111111000",
  37933=>"111111111",
  37934=>"000110100",
  37935=>"111111111",
  37936=>"111100010",
  37937=>"010111111",
  37938=>"000000001",
  37939=>"101001000",
  37940=>"011111111",
  37941=>"100111000",
  37942=>"100000011",
  37943=>"000100111",
  37944=>"000000000",
  37945=>"010000111",
  37946=>"000001000",
  37947=>"010110000",
  37948=>"111111111",
  37949=>"000000111",
  37950=>"000101111",
  37951=>"001001000",
  37952=>"111000000",
  37953=>"111011000",
  37954=>"000000000",
  37955=>"111000111",
  37956=>"100100110",
  37957=>"000000000",
  37958=>"000000000",
  37959=>"000000000",
  37960=>"011000001",
  37961=>"000000111",
  37962=>"111111000",
  37963=>"100000000",
  37964=>"000000000",
  37965=>"111111111",
  37966=>"000000000",
  37967=>"000000000",
  37968=>"000000001",
  37969=>"000110111",
  37970=>"011000000",
  37971=>"110110000",
  37972=>"000000011",
  37973=>"010010000",
  37974=>"000000111",
  37975=>"010000000",
  37976=>"000000000",
  37977=>"001000101",
  37978=>"000000000",
  37979=>"001111100",
  37980=>"000000000",
  37981=>"001000000",
  37982=>"011011000",
  37983=>"000000001",
  37984=>"111000111",
  37985=>"000000000",
  37986=>"000001000",
  37987=>"000100111",
  37988=>"000110100",
  37989=>"011001111",
  37990=>"000111111",
  37991=>"000001011",
  37992=>"010111000",
  37993=>"000000000",
  37994=>"001000000",
  37995=>"001001001",
  37996=>"111111100",
  37997=>"000000000",
  37998=>"000000010",
  37999=>"000111111",
  38000=>"001011011",
  38001=>"000000001",
  38002=>"000011011",
  38003=>"000111111",
  38004=>"111000000",
  38005=>"010111111",
  38006=>"110110110",
  38007=>"111111110",
  38008=>"111111111",
  38009=>"111100000",
  38010=>"010111111",
  38011=>"111111000",
  38012=>"000001111",
  38013=>"111111100",
  38014=>"111111111",
  38015=>"000000000",
  38016=>"111111111",
  38017=>"000000111",
  38018=>"001001000",
  38019=>"111111111",
  38020=>"111000000",
  38021=>"101000000",
  38022=>"101110000",
  38023=>"110111111",
  38024=>"111111000",
  38025=>"000000011",
  38026=>"000000000",
  38027=>"111011000",
  38028=>"000000110",
  38029=>"110000000",
  38030=>"101101101",
  38031=>"111111111",
  38032=>"111111111",
  38033=>"000001111",
  38034=>"000000000",
  38035=>"000000000",
  38036=>"111111111",
  38037=>"000010111",
  38038=>"001000000",
  38039=>"000011000",
  38040=>"111111000",
  38041=>"111001000",
  38042=>"110110000",
  38043=>"100111000",
  38044=>"000000000",
  38045=>"010110110",
  38046=>"111000000",
  38047=>"000000000",
  38048=>"000000000",
  38049=>"111011000",
  38050=>"110111111",
  38051=>"000110000",
  38052=>"000111111",
  38053=>"111101101",
  38054=>"000111000",
  38055=>"000111111",
  38056=>"110000111",
  38057=>"001000001",
  38058=>"111001000",
  38059=>"111100111",
  38060=>"111111111",
  38061=>"111101000",
  38062=>"111111101",
  38063=>"000000000",
  38064=>"111111111",
  38065=>"000000000",
  38066=>"111111110",
  38067=>"111111000",
  38068=>"111111101",
  38069=>"000000000",
  38070=>"000000000",
  38071=>"110110000",
  38072=>"111000000",
  38073=>"000000000",
  38074=>"000000110",
  38075=>"101001011",
  38076=>"111110100",
  38077=>"000001111",
  38078=>"111110000",
  38079=>"111000101",
  38080=>"110111111",
  38081=>"011111001",
  38082=>"011011000",
  38083=>"000111000",
  38084=>"111111111",
  38085=>"000000111",
  38086=>"100000100",
  38087=>"110111100",
  38088=>"000111111",
  38089=>"111010000",
  38090=>"111111111",
  38091=>"011000000",
  38092=>"000001001",
  38093=>"111111111",
  38094=>"111000000",
  38095=>"000011000",
  38096=>"000100111",
  38097=>"111111111",
  38098=>"000010110",
  38099=>"110111000",
  38100=>"000100111",
  38101=>"000111000",
  38102=>"000111110",
  38103=>"011000000",
  38104=>"111111111",
  38105=>"111111110",
  38106=>"111000110",
  38107=>"010111111",
  38108=>"111111101",
  38109=>"001000000",
  38110=>"000000110",
  38111=>"111111000",
  38112=>"000000000",
  38113=>"001000000",
  38114=>"000000001",
  38115=>"111111000",
  38116=>"011001000",
  38117=>"000000010",
  38118=>"000001111",
  38119=>"111110000",
  38120=>"111111110",
  38121=>"000111111",
  38122=>"111111111",
  38123=>"111000111",
  38124=>"110001010",
  38125=>"000111111",
  38126=>"000001111",
  38127=>"000000000",
  38128=>"100000000",
  38129=>"011000111",
  38130=>"111000101",
  38131=>"000010010",
  38132=>"001000111",
  38133=>"000000000",
  38134=>"000111111",
  38135=>"111101111",
  38136=>"111111111",
  38137=>"111111000",
  38138=>"101101101",
  38139=>"001011010",
  38140=>"000011000",
  38141=>"000010111",
  38142=>"000000111",
  38143=>"111101001",
  38144=>"000110100",
  38145=>"100100000",
  38146=>"100000101",
  38147=>"000000000",
  38148=>"111111111",
  38149=>"111000000",
  38150=>"111111000",
  38151=>"111001011",
  38152=>"100110111",
  38153=>"111000000",
  38154=>"111111110",
  38155=>"000001001",
  38156=>"001111111",
  38157=>"000000000",
  38158=>"111111111",
  38159=>"111011000",
  38160=>"010110110",
  38161=>"111111111",
  38162=>"000011111",
  38163=>"101111111",
  38164=>"111111110",
  38165=>"000111111",
  38166=>"100100000",
  38167=>"101011000",
  38168=>"100000000",
  38169=>"000111111",
  38170=>"000111111",
  38171=>"110110111",
  38172=>"100000100",
  38173=>"000000111",
  38174=>"011011111",
  38175=>"001000000",
  38176=>"000000111",
  38177=>"000111111",
  38178=>"000100010",
  38179=>"111000000",
  38180=>"000001001",
  38181=>"001011111",
  38182=>"000000000",
  38183=>"000000001",
  38184=>"000011010",
  38185=>"000000000",
  38186=>"011000111",
  38187=>"000000000",
  38188=>"000111000",
  38189=>"001001001",
  38190=>"000000000",
  38191=>"000000001",
  38192=>"110111100",
  38193=>"000000111",
  38194=>"000100111",
  38195=>"000111111",
  38196=>"100101101",
  38197=>"111000000",
  38198=>"111111110",
  38199=>"000000100",
  38200=>"101001111",
  38201=>"000000000",
  38202=>"000011000",
  38203=>"000000110",
  38204=>"000110111",
  38205=>"101111111",
  38206=>"010000000",
  38207=>"110100111",
  38208=>"101101111",
  38209=>"111111111",
  38210=>"111110000",
  38211=>"000000000",
  38212=>"000111111",
  38213=>"000111111",
  38214=>"000000000",
  38215=>"111111000",
  38216=>"000000000",
  38217=>"000000000",
  38218=>"111101100",
  38219=>"111111110",
  38220=>"110110111",
  38221=>"011111111",
  38222=>"111100000",
  38223=>"000100100",
  38224=>"110111111",
  38225=>"111111111",
  38226=>"000000000",
  38227=>"111111000",
  38228=>"000000000",
  38229=>"011011011",
  38230=>"111011110",
  38231=>"100000011",
  38232=>"000000000",
  38233=>"110000000",
  38234=>"000001001",
  38235=>"111111111",
  38236=>"000000000",
  38237=>"000000111",
  38238=>"000001000",
  38239=>"001001100",
  38240=>"100001111",
  38241=>"101000000",
  38242=>"011001000",
  38243=>"101111111",
  38244=>"111111111",
  38245=>"111111000",
  38246=>"100000011",
  38247=>"111000000",
  38248=>"111111111",
  38249=>"010111011",
  38250=>"111111111",
  38251=>"111111000",
  38252=>"110000000",
  38253=>"000100110",
  38254=>"010000000",
  38255=>"000000000",
  38256=>"011111111",
  38257=>"111111111",
  38258=>"000111110",
  38259=>"011111110",
  38260=>"110111111",
  38261=>"001000000",
  38262=>"111111000",
  38263=>"000000000",
  38264=>"000010111",
  38265=>"110011000",
  38266=>"111100111",
  38267=>"000010111",
  38268=>"110111111",
  38269=>"000001111",
  38270=>"000000000",
  38271=>"000000000",
  38272=>"000001001",
  38273=>"000000001",
  38274=>"000000000",
  38275=>"000000001",
  38276=>"000110111",
  38277=>"111000000",
  38278=>"000000000",
  38279=>"110000000",
  38280=>"000001001",
  38281=>"000111111",
  38282=>"010010000",
  38283=>"101111111",
  38284=>"111111111",
  38285=>"000100111",
  38286=>"001000000",
  38287=>"000111111",
  38288=>"000000000",
  38289=>"111110111",
  38290=>"110111111",
  38291=>"000100111",
  38292=>"111000000",
  38293=>"000010000",
  38294=>"000000111",
  38295=>"001111111",
  38296=>"000100111",
  38297=>"000111011",
  38298=>"100100111",
  38299=>"111111000",
  38300=>"111011000",
  38301=>"111001000",
  38302=>"000000000",
  38303=>"000000000",
  38304=>"000111111",
  38305=>"110111000",
  38306=>"110000001",
  38307=>"110101110",
  38308=>"111111011",
  38309=>"100000000",
  38310=>"000001000",
  38311=>"111100110",
  38312=>"011000000",
  38313=>"001001111",
  38314=>"100000000",
  38315=>"111110001",
  38316=>"110010011",
  38317=>"010010010",
  38318=>"011011000",
  38319=>"001100111",
  38320=>"111000000",
  38321=>"000000000",
  38322=>"000000000",
  38323=>"111011000",
  38324=>"011000000",
  38325=>"000001111",
  38326=>"111111001",
  38327=>"000000000",
  38328=>"000111111",
  38329=>"000000101",
  38330=>"000011111",
  38331=>"100111111",
  38332=>"111010010",
  38333=>"000001000",
  38334=>"001000000",
  38335=>"111111100",
  38336=>"000000000",
  38337=>"111000000",
  38338=>"000000000",
  38339=>"111000000",
  38340=>"111010111",
  38341=>"101111111",
  38342=>"111001001",
  38343=>"100100000",
  38344=>"111111010",
  38345=>"111000000",
  38346=>"000001111",
  38347=>"000000111",
  38348=>"111111111",
  38349=>"110010110",
  38350=>"100000000",
  38351=>"100111111",
  38352=>"111111111",
  38353=>"000000000",
  38354=>"111001111",
  38355=>"000000000",
  38356=>"111111011",
  38357=>"111000000",
  38358=>"100110110",
  38359=>"000000000",
  38360=>"111111111",
  38361=>"011000000",
  38362=>"010110111",
  38363=>"000111101",
  38364=>"000010110",
  38365=>"111111111",
  38366=>"011111111",
  38367=>"000110111",
  38368=>"111111011",
  38369=>"111111111",
  38370=>"111111100",
  38371=>"111011111",
  38372=>"111111111",
  38373=>"100110010",
  38374=>"000001111",
  38375=>"000000111",
  38376=>"111111000",
  38377=>"111000000",
  38378=>"001111111",
  38379=>"111111111",
  38380=>"111111110",
  38381=>"011111111",
  38382=>"111111000",
  38383=>"000000000",
  38384=>"000111111",
  38385=>"000111110",
  38386=>"000001010",
  38387=>"000000000",
  38388=>"111110110",
  38389=>"000100110",
  38390=>"010111000",
  38391=>"000001000",
  38392=>"011111101",
  38393=>"000000000",
  38394=>"000010110",
  38395=>"111000000",
  38396=>"000000000",
  38397=>"110111100",
  38398=>"111011010",
  38399=>"100000000",
  38400=>"100000000",
  38401=>"110001101",
  38402=>"111111111",
  38403=>"000000000",
  38404=>"000000100",
  38405=>"010010011",
  38406=>"000000000",
  38407=>"110111111",
  38408=>"111111111",
  38409=>"000000100",
  38410=>"000000000",
  38411=>"111111100",
  38412=>"011011000",
  38413=>"000000001",
  38414=>"001101001",
  38415=>"000100000",
  38416=>"110000011",
  38417=>"000001111",
  38418=>"101111111",
  38419=>"000000101",
  38420=>"000000111",
  38421=>"101101111",
  38422=>"000000000",
  38423=>"110110111",
  38424=>"111111111",
  38425=>"000100000",
  38426=>"000000101",
  38427=>"000000100",
  38428=>"111111111",
  38429=>"111011001",
  38430=>"000000000",
  38431=>"100100110",
  38432=>"111000000",
  38433=>"000000000",
  38434=>"111111111",
  38435=>"000000000",
  38436=>"110111010",
  38437=>"000000011",
  38438=>"000000000",
  38439=>"110100000",
  38440=>"101001111",
  38441=>"111111111",
  38442=>"000000001",
  38443=>"001001111",
  38444=>"000000000",
  38445=>"000000101",
  38446=>"000000000",
  38447=>"111111000",
  38448=>"110000000",
  38449=>"000001000",
  38450=>"000001001",
  38451=>"000000000",
  38452=>"000000000",
  38453=>"110111111",
  38454=>"111111111",
  38455=>"111111101",
  38456=>"000000000",
  38457=>"111111111",
  38458=>"111111111",
  38459=>"100100110",
  38460=>"000000001",
  38461=>"000001000",
  38462=>"000000000",
  38463=>"100110110",
  38464=>"111111101",
  38465=>"011011010",
  38466=>"000000000",
  38467=>"110111111",
  38468=>"111011001",
  38469=>"111111111",
  38470=>"010000100",
  38471=>"000000000",
  38472=>"000010000",
  38473=>"111111111",
  38474=>"111111111",
  38475=>"111100100",
  38476=>"000000000",
  38477=>"111111110",
  38478=>"010000100",
  38479=>"000000000",
  38480=>"101111111",
  38481=>"000000001",
  38482=>"000000010",
  38483=>"000001010",
  38484=>"000000000",
  38485=>"111111111",
  38486=>"111110111",
  38487=>"111111111",
  38488=>"110011111",
  38489=>"111111111",
  38490=>"000000111",
  38491=>"100000000",
  38492=>"000000000",
  38493=>"000000000",
  38494=>"001001000",
  38495=>"001000000",
  38496=>"000000000",
  38497=>"011001111",
  38498=>"111000000",
  38499=>"000000000",
  38500=>"000001011",
  38501=>"000000000",
  38502=>"000000000",
  38503=>"000000000",
  38504=>"111111111",
  38505=>"111111110",
  38506=>"111111111",
  38507=>"111100001",
  38508=>"000000000",
  38509=>"100000000",
  38510=>"111111111",
  38511=>"111111111",
  38512=>"000000000",
  38513=>"111011001",
  38514=>"000000000",
  38515=>"101100000",
  38516=>"110010000",
  38517=>"000000100",
  38518=>"111100000",
  38519=>"000000000",
  38520=>"000110110",
  38521=>"011000000",
  38522=>"000011111",
  38523=>"000000101",
  38524=>"110110110",
  38525=>"111111011",
  38526=>"000000000",
  38527=>"000000101",
  38528=>"111111111",
  38529=>"100100000",
  38530=>"111000000",
  38531=>"000000000",
  38532=>"000000000",
  38533=>"000000001",
  38534=>"111111001",
  38535=>"110100100",
  38536=>"111001001",
  38537=>"000000000",
  38538=>"000000000",
  38539=>"000000000",
  38540=>"111111111",
  38541=>"111111111",
  38542=>"010111000",
  38543=>"101001000",
  38544=>"000001001",
  38545=>"000000000",
  38546=>"000000000",
  38547=>"111110111",
  38548=>"000000000",
  38549=>"110100011",
  38550=>"111111111",
  38551=>"111111001",
  38552=>"100111101",
  38553=>"100110000",
  38554=>"100000000",
  38555=>"111101111",
  38556=>"000000000",
  38557=>"010010111",
  38558=>"111111111",
  38559=>"000011000",
  38560=>"000001000",
  38561=>"011111111",
  38562=>"111111111",
  38563=>"000000000",
  38564=>"000110010",
  38565=>"111111111",
  38566=>"111100000",
  38567=>"100000000",
  38568=>"011000000",
  38569=>"000000000",
  38570=>"111001001",
  38571=>"111111111",
  38572=>"101111111",
  38573=>"100000000",
  38574=>"000001111",
  38575=>"110110100",
  38576=>"111111111",
  38577=>"111110000",
  38578=>"111111111",
  38579=>"000000000",
  38580=>"000011011",
  38581=>"110100000",
  38582=>"000000000",
  38583=>"111111111",
  38584=>"111111111",
  38585=>"111011010",
  38586=>"111111001",
  38587=>"111111111",
  38588=>"000000000",
  38589=>"111111111",
  38590=>"000000000",
  38591=>"001001000",
  38592=>"100000111",
  38593=>"011001011",
  38594=>"111001010",
  38595=>"000000000",
  38596=>"111111111",
  38597=>"000011000",
  38598=>"011110110",
  38599=>"000000100",
  38600=>"111111111",
  38601=>"000000000",
  38602=>"001000000",
  38603=>"111111111",
  38604=>"111111111",
  38605=>"100100100",
  38606=>"000000001",
  38607=>"101101111",
  38608=>"000000100",
  38609=>"111111111",
  38610=>"000000000",
  38611=>"001011011",
  38612=>"001100000",
  38613=>"111111111",
  38614=>"000000000",
  38615=>"111111111",
  38616=>"100100000",
  38617=>"110111000",
  38618=>"111100000",
  38619=>"000101000",
  38620=>"000000000",
  38621=>"111111111",
  38622=>"000000111",
  38623=>"000000000",
  38624=>"000000100",
  38625=>"111011001",
  38626=>"000000000",
  38627=>"100000000",
  38628=>"000111100",
  38629=>"000000100",
  38630=>"000000000",
  38631=>"101110110",
  38632=>"111111111",
  38633=>"000000000",
  38634=>"111111111",
  38635=>"000000011",
  38636=>"000000000",
  38637=>"000000000",
  38638=>"001111111",
  38639=>"111010111",
  38640=>"000000000",
  38641=>"000100110",
  38642=>"111111111",
  38643=>"001000000",
  38644=>"111111111",
  38645=>"000000000",
  38646=>"100100100",
  38647=>"111111111",
  38648=>"111111111",
  38649=>"111000111",
  38650=>"111111111",
  38651=>"000000000",
  38652=>"001001001",
  38653=>"001001001",
  38654=>"110110000",
  38655=>"100100110",
  38656=>"000001000",
  38657=>"000001001",
  38658=>"000000001",
  38659=>"111111111",
  38660=>"111111000",
  38661=>"000000001",
  38662=>"000000000",
  38663=>"100100101",
  38664=>"000000001",
  38665=>"000000000",
  38666=>"111110111",
  38667=>"000001001",
  38668=>"000000000",
  38669=>"000000000",
  38670=>"101100111",
  38671=>"001111111",
  38672=>"011111111",
  38673=>"111111111",
  38674=>"000101111",
  38675=>"111011111",
  38676=>"111111111",
  38677=>"100000000",
  38678=>"000000000",
  38679=>"000000000",
  38680=>"000111110",
  38681=>"000000000",
  38682=>"111100101",
  38683=>"111111111",
  38684=>"000000000",
  38685=>"111100000",
  38686=>"000000000",
  38687=>"111001101",
  38688=>"001100000",
  38689=>"011111111",
  38690=>"111001000",
  38691=>"111111111",
  38692=>"011000101",
  38693=>"111111111",
  38694=>"111111111",
  38695=>"000000100",
  38696=>"000000011",
  38697=>"111101101",
  38698=>"111011001",
  38699=>"000000000",
  38700=>"111111111",
  38701=>"000001001",
  38702=>"111000111",
  38703=>"110111111",
  38704=>"000111111",
  38705=>"111111110",
  38706=>"001000111",
  38707=>"000000000",
  38708=>"111111111",
  38709=>"000000000",
  38710=>"110000000",
  38711=>"000000000",
  38712=>"110110110",
  38713=>"000000111",
  38714=>"011011000",
  38715=>"110111000",
  38716=>"001111011",
  38717=>"011110000",
  38718=>"000000000",
  38719=>"110111111",
  38720=>"011011000",
  38721=>"110000000",
  38722=>"111111111",
  38723=>"111111110",
  38724=>"011001000",
  38725=>"000000011",
  38726=>"110111111",
  38727=>"000000000",
  38728=>"110110000",
  38729=>"111010110",
  38730=>"111111111",
  38731=>"000100100",
  38732=>"000110110",
  38733=>"111111001",
  38734=>"111111111",
  38735=>"000000000",
  38736=>"000000000",
  38737=>"001000000",
  38738=>"001001001",
  38739=>"011000000",
  38740=>"111111111",
  38741=>"011011011",
  38742=>"000000001",
  38743=>"000001101",
  38744=>"100000000",
  38745=>"000000000",
  38746=>"000001001",
  38747=>"000000111",
  38748=>"000000010",
  38749=>"111100000",
  38750=>"000000111",
  38751=>"111111111",
  38752=>"000000000",
  38753=>"011111111",
  38754=>"001011111",
  38755=>"111111011",
  38756=>"101000000",
  38757=>"000000000",
  38758=>"000000101",
  38759=>"000000000",
  38760=>"110100100",
  38761=>"111111001",
  38762=>"010011000",
  38763=>"000000000",
  38764=>"011110110",
  38765=>"000011000",
  38766=>"111110110",
  38767=>"111001000",
  38768=>"111111111",
  38769=>"000001011",
  38770=>"000001000",
  38771=>"111001000",
  38772=>"110000000",
  38773=>"000000000",
  38774=>"011111000",
  38775=>"010111111",
  38776=>"111111001",
  38777=>"001000000",
  38778=>"000000000",
  38779=>"000111110",
  38780=>"111111000",
  38781=>"000000000",
  38782=>"111000000",
  38783=>"111001000",
  38784=>"111111101",
  38785=>"101101111",
  38786=>"111111111",
  38787=>"000000000",
  38788=>"000000110",
  38789=>"111111000",
  38790=>"010110110",
  38791=>"100000111",
  38792=>"011001101",
  38793=>"000000000",
  38794=>"000000000",
  38795=>"111111111",
  38796=>"011111011",
  38797=>"101000011",
  38798=>"000000000",
  38799=>"111111111",
  38800=>"111111011",
  38801=>"110000000",
  38802=>"101111111",
  38803=>"110110100",
  38804=>"001011111",
  38805=>"000000000",
  38806=>"111111110",
  38807=>"010010000",
  38808=>"111110110",
  38809=>"111000000",
  38810=>"000100100",
  38811=>"000001001",
  38812=>"111111001",
  38813=>"111111111",
  38814=>"000100010",
  38815=>"000000000",
  38816=>"111111111",
  38817=>"000000010",
  38818=>"111011111",
  38819=>"111001000",
  38820=>"111111111",
  38821=>"000001001",
  38822=>"001001000",
  38823=>"000100101",
  38824=>"000000000",
  38825=>"111111111",
  38826=>"111111111",
  38827=>"000000000",
  38828=>"111000111",
  38829=>"000001001",
  38830=>"000001011",
  38831=>"011011111",
  38832=>"000010101",
  38833=>"000000000",
  38834=>"100110101",
  38835=>"000000000",
  38836=>"111110111",
  38837=>"111111011",
  38838=>"111111111",
  38839=>"010111011",
  38840=>"000000000",
  38841=>"000111001",
  38842=>"000000000",
  38843=>"110010000",
  38844=>"111111111",
  38845=>"111111001",
  38846=>"000000000",
  38847=>"100101111",
  38848=>"111111111",
  38849=>"000000000",
  38850=>"000101111",
  38851=>"000001111",
  38852=>"000000111",
  38853=>"100100000",
  38854=>"000000000",
  38855=>"111111111",
  38856=>"000011000",
  38857=>"000011000",
  38858=>"111111111",
  38859=>"000011111",
  38860=>"000000000",
  38861=>"111111100",
  38862=>"101111111",
  38863=>"000000100",
  38864=>"000010110",
  38865=>"111111111",
  38866=>"000101000",
  38867=>"000000001",
  38868=>"111111001",
  38869=>"111011111",
  38870=>"000000111",
  38871=>"110110110",
  38872=>"101101101",
  38873=>"000000000",
  38874=>"000000001",
  38875=>"000001000",
  38876=>"111111111",
  38877=>"111101111",
  38878=>"000000000",
  38879=>"100000001",
  38880=>"000000000",
  38881=>"111111001",
  38882=>"000110111",
  38883=>"000000000",
  38884=>"000000000",
  38885=>"000000000",
  38886=>"001101101",
  38887=>"010000000",
  38888=>"000010110",
  38889=>"111000000",
  38890=>"110110000",
  38891=>"111111010",
  38892=>"000011111",
  38893=>"000000000",
  38894=>"000000000",
  38895=>"000000111",
  38896=>"000000000",
  38897=>"000000000",
  38898=>"111111111",
  38899=>"000000000",
  38900=>"111000100",
  38901=>"110110000",
  38902=>"111000000",
  38903=>"110010000",
  38904=>"000000000",
  38905=>"000010010",
  38906=>"111110000",
  38907=>"111111111",
  38908=>"000000000",
  38909=>"000110111",
  38910=>"011111111",
  38911=>"111111111",
  38912=>"001000000",
  38913=>"000000100",
  38914=>"000000000",
  38915=>"000000111",
  38916=>"000000000",
  38917=>"111001001",
  38918=>"000000000",
  38919=>"000111111",
  38920=>"111111111",
  38921=>"011011000",
  38922=>"000000000",
  38923=>"111111111",
  38924=>"110110100",
  38925=>"000000000",
  38926=>"111001000",
  38927=>"111111111",
  38928=>"111111111",
  38929=>"000111100",
  38930=>"000111000",
  38931=>"111111111",
  38932=>"000000000",
  38933=>"010111111",
  38934=>"000000000",
  38935=>"011011000",
  38936=>"111000000",
  38937=>"111111111",
  38938=>"000000001",
  38939=>"110100000",
  38940=>"000000000",
  38941=>"001001000",
  38942=>"000111111",
  38943=>"100111110",
  38944=>"000000111",
  38945=>"111111000",
  38946=>"111110110",
  38947=>"010000001",
  38948=>"000000000",
  38949=>"000000100",
  38950=>"000000111",
  38951=>"100000110",
  38952=>"000000011",
  38953=>"110110111",
  38954=>"111111111",
  38955=>"001001110",
  38956=>"111111110",
  38957=>"111111111",
  38958=>"001000000",
  38959=>"000000000",
  38960=>"111111111",
  38961=>"111111111",
  38962=>"001000001",
  38963=>"111111111",
  38964=>"000011011",
  38965=>"111111111",
  38966=>"101100111",
  38967=>"111110000",
  38968=>"000000000",
  38969=>"110111111",
  38970=>"000000000",
  38971=>"111110111",
  38972=>"111111111",
  38973=>"101101111",
  38974=>"000000001",
  38975=>"111111111",
  38976=>"000000000",
  38977=>"111111000",
  38978=>"111111111",
  38979=>"111111001",
  38980=>"011110110",
  38981=>"000000000",
  38982=>"111111110",
  38983=>"000000000",
  38984=>"011001011",
  38985=>"001001001",
  38986=>"000000000",
  38987=>"100000000",
  38988=>"111111111",
  38989=>"000000111",
  38990=>"000000110",
  38991=>"111111111",
  38992=>"010010011",
  38993=>"000000110",
  38994=>"100000110",
  38995=>"111111111",
  38996=>"111111110",
  38997=>"111001000",
  38998=>"110100000",
  38999=>"001000000",
  39000=>"111111111",
  39001=>"111110110",
  39002=>"000000000",
  39003=>"001001111",
  39004=>"011010010",
  39005=>"111111111",
  39006=>"001111111",
  39007=>"111111111",
  39008=>"000000000",
  39009=>"000000111",
  39010=>"110110110",
  39011=>"000000000",
  39012=>"000000000",
  39013=>"111000010",
  39014=>"001000010",
  39015=>"111111111",
  39016=>"100000000",
  39017=>"001000000",
  39018=>"111110000",
  39019=>"000001000",
  39020=>"000000000",
  39021=>"111111111",
  39022=>"011000111",
  39023=>"000000000",
  39024=>"010000111",
  39025=>"000000011",
  39026=>"011111111",
  39027=>"000000000",
  39028=>"111010000",
  39029=>"111111001",
  39030=>"111111110",
  39031=>"111111111",
  39032=>"111111111",
  39033=>"100000000",
  39034=>"000000000",
  39035=>"000000000",
  39036=>"100110000",
  39037=>"111001001",
  39038=>"000000000",
  39039=>"101101111",
  39040=>"011111111",
  39041=>"001000001",
  39042=>"111111111",
  39043=>"111111111",
  39044=>"110111111",
  39045=>"011111111",
  39046=>"000000000",
  39047=>"001000000",
  39048=>"110111000",
  39049=>"000000000",
  39050=>"100100010",
  39051=>"111111111",
  39052=>"111101000",
  39053=>"111111111",
  39054=>"000000000",
  39055=>"000000000",
  39056=>"111111111",
  39057=>"111111111",
  39058=>"000000000",
  39059=>"100001000",
  39060=>"010111011",
  39061=>"111111000",
  39062=>"011000000",
  39063=>"000000000",
  39064=>"011101111",
  39065=>"111111111",
  39066=>"001010110",
  39067=>"111111100",
  39068=>"111111111",
  39069=>"001000000",
  39070=>"111011111",
  39071=>"000000000",
  39072=>"000100111",
  39073=>"111011111",
  39074=>"111111111",
  39075=>"000000000",
  39076=>"000000000",
  39077=>"110111111",
  39078=>"111111111",
  39079=>"110110111",
  39080=>"000001000",
  39081=>"111111111",
  39082=>"111111011",
  39083=>"111101111",
  39084=>"111111111",
  39085=>"000000001",
  39086=>"111000011",
  39087=>"000000000",
  39088=>"111111000",
  39089=>"111111111",
  39090=>"010110110",
  39091=>"111111111",
  39092=>"011000000",
  39093=>"111111111",
  39094=>"000111111",
  39095=>"011001111",
  39096=>"111011111",
  39097=>"000001001",
  39098=>"001111111",
  39099=>"001000111",
  39100=>"111100101",
  39101=>"000000000",
  39102=>"000000000",
  39103=>"000000111",
  39104=>"100000000",
  39105=>"000000000",
  39106=>"111111111",
  39107=>"111111111",
  39108=>"011001111",
  39109=>"111111111",
  39110=>"001001101",
  39111=>"000000001",
  39112=>"011111111",
  39113=>"111111110",
  39114=>"000000000",
  39115=>"111111111",
  39116=>"000001101",
  39117=>"110000000",
  39118=>"111111111",
  39119=>"111111111",
  39120=>"111011101",
  39121=>"000000010",
  39122=>"000000010",
  39123=>"111111111",
  39124=>"001000000",
  39125=>"101111011",
  39126=>"001001011",
  39127=>"111111111",
  39128=>"111101110",
  39129=>"111111111",
  39130=>"000011011",
  39131=>"100000001",
  39132=>"000000000",
  39133=>"111100101",
  39134=>"100000000",
  39135=>"000000000",
  39136=>"000000000",
  39137=>"111111000",
  39138=>"000000000",
  39139=>"000000000",
  39140=>"000000000",
  39141=>"110100111",
  39142=>"111111111",
  39143=>"000000111",
  39144=>"000000110",
  39145=>"110110111",
  39146=>"001011111",
  39147=>"100110111",
  39148=>"111111111",
  39149=>"000000000",
  39150=>"110111000",
  39151=>"001010111",
  39152=>"101111111",
  39153=>"111111000",
  39154=>"001111111",
  39155=>"001000000",
  39156=>"000000000",
  39157=>"111111111",
  39158=>"101000000",
  39159=>"100100000",
  39160=>"111111111",
  39161=>"000000000",
  39162=>"111111011",
  39163=>"000000000",
  39164=>"001001011",
  39165=>"110000000",
  39166=>"000000111",
  39167=>"111000000",
  39168=>"000000000",
  39169=>"110110110",
  39170=>"100101111",
  39171=>"111111111",
  39172=>"111111111",
  39173=>"111111111",
  39174=>"000111111",
  39175=>"010000001",
  39176=>"000000000",
  39177=>"111111111",
  39178=>"111100100",
  39179=>"100110010",
  39180=>"100100000",
  39181=>"111111111",
  39182=>"000000000",
  39183=>"110111111",
  39184=>"000000000",
  39185=>"000000111",
  39186=>"011011111",
  39187=>"111001101",
  39188=>"111111111",
  39189=>"111111111",
  39190=>"011111111",
  39191=>"111111000",
  39192=>"000000000",
  39193=>"000000000",
  39194=>"111101111",
  39195=>"111011001",
  39196=>"111110111",
  39197=>"000010011",
  39198=>"111111011",
  39199=>"000000011",
  39200=>"011001000",
  39201=>"000000000",
  39202=>"000000001",
  39203=>"000111110",
  39204=>"111111111",
  39205=>"000000110",
  39206=>"011011011",
  39207=>"000000000",
  39208=>"101101101",
  39209=>"000000000",
  39210=>"001111111",
  39211=>"111111111",
  39212=>"111111111",
  39213=>"000000000",
  39214=>"000000111",
  39215=>"111111111",
  39216=>"000000000",
  39217=>"000010111",
  39218=>"111111011",
  39219=>"111111100",
  39220=>"111111000",
  39221=>"001001111",
  39222=>"111011011",
  39223=>"000000000",
  39224=>"001000010",
  39225=>"001101111",
  39226=>"111111111",
  39227=>"000000000",
  39228=>"111111111",
  39229=>"000000111",
  39230=>"000000000",
  39231=>"001000111",
  39232=>"101000000",
  39233=>"010010000",
  39234=>"000001111",
  39235=>"000000001",
  39236=>"000000000",
  39237=>"100100000",
  39238=>"000000000",
  39239=>"111110110",
  39240=>"111111111",
  39241=>"100000000",
  39242=>"000000111",
  39243=>"000000011",
  39244=>"000000000",
  39245=>"000011111",
  39246=>"100110111",
  39247=>"111001001",
  39248=>"111101101",
  39249=>"111111111",
  39250=>"111101111",
  39251=>"111111111",
  39252=>"111101111",
  39253=>"000000000",
  39254=>"111111111",
  39255=>"000000000",
  39256=>"111100011",
  39257=>"111111111",
  39258=>"010000011",
  39259=>"000011001",
  39260=>"111111011",
  39261=>"011000000",
  39262=>"111111111",
  39263=>"001111011",
  39264=>"000000000",
  39265=>"011001000",
  39266=>"000100001",
  39267=>"111111111",
  39268=>"001000010",
  39269=>"000000000",
  39270=>"000000000",
  39271=>"111111111",
  39272=>"000100111",
  39273=>"000000111",
  39274=>"111111111",
  39275=>"000011001",
  39276=>"100000100",
  39277=>"000011011",
  39278=>"111111000",
  39279=>"000000000",
  39280=>"111111111",
  39281=>"000000000",
  39282=>"011000011",
  39283=>"010111001",
  39284=>"111111111",
  39285=>"110111111",
  39286=>"000000010",
  39287=>"011111100",
  39288=>"110111111",
  39289=>"111111111",
  39290=>"000011011",
  39291=>"110100100",
  39292=>"111111110",
  39293=>"111111110",
  39294=>"000000111",
  39295=>"111111111",
  39296=>"010011111",
  39297=>"110111111",
  39298=>"000000000",
  39299=>"111111111",
  39300=>"111111000",
  39301=>"001000111",
  39302=>"111111011",
  39303=>"111111111",
  39304=>"011110111",
  39305=>"100100000",
  39306=>"111110000",
  39307=>"011000000",
  39308=>"000000000",
  39309=>"110100000",
  39310=>"000000000",
  39311=>"000000000",
  39312=>"011000000",
  39313=>"111111111",
  39314=>"011000001",
  39315=>"111111010",
  39316=>"000000000",
  39317=>"010111111",
  39318=>"000000000",
  39319=>"111010000",
  39320=>"001001000",
  39321=>"111111111",
  39322=>"000000000",
  39323=>"100111111",
  39324=>"000000000",
  39325=>"011000111",
  39326=>"000000000",
  39327=>"111110110",
  39328=>"100000101",
  39329=>"000010010",
  39330=>"000000110",
  39331=>"111111000",
  39332=>"111111111",
  39333=>"111111111",
  39334=>"111111111",
  39335=>"011111101",
  39336=>"000000000",
  39337=>"111111011",
  39338=>"000000000",
  39339=>"111111100",
  39340=>"101000000",
  39341=>"000000000",
  39342=>"100100101",
  39343=>"111111111",
  39344=>"000000000",
  39345=>"111000000",
  39346=>"000000111",
  39347=>"001000000",
  39348=>"000000001",
  39349=>"100100000",
  39350=>"000000001",
  39351=>"000111111",
  39352=>"111101111",
  39353=>"100100000",
  39354=>"000000000",
  39355=>"000000000",
  39356=>"000000000",
  39357=>"111111111",
  39358=>"111111111",
  39359=>"001001001",
  39360=>"111111000",
  39361=>"001001101",
  39362=>"111111111",
  39363=>"111111111",
  39364=>"111111111",
  39365=>"100000010",
  39366=>"111111000",
  39367=>"010011110",
  39368=>"000000101",
  39369=>"000001111",
  39370=>"110000100",
  39371=>"001001000",
  39372=>"000000000",
  39373=>"000000000",
  39374=>"111111111",
  39375=>"100100100",
  39376=>"000111111",
  39377=>"111111111",
  39378=>"111111111",
  39379=>"001000011",
  39380=>"111000000",
  39381=>"111111111",
  39382=>"101111111",
  39383=>"000001011",
  39384=>"000000000",
  39385=>"000000011",
  39386=>"000000001",
  39387=>"001000000",
  39388=>"000000000",
  39389=>"000100000",
  39390=>"000000000",
  39391=>"101101001",
  39392=>"000000000",
  39393=>"001100111",
  39394=>"000000000",
  39395=>"000000100",
  39396=>"111111111",
  39397=>"111111111",
  39398=>"111111101",
  39399=>"110000000",
  39400=>"000000101",
  39401=>"000000000",
  39402=>"000011111",
  39403=>"111101001",
  39404=>"101100000",
  39405=>"000000000",
  39406=>"000001111",
  39407=>"111111111",
  39408=>"000000000",
  39409=>"000000000",
  39410=>"111001001",
  39411=>"000111111",
  39412=>"000010000",
  39413=>"011111111",
  39414=>"000000000",
  39415=>"110110110",
  39416=>"000000111",
  39417=>"100101100",
  39418=>"111111111",
  39419=>"101000101",
  39420=>"000001111",
  39421=>"111111111",
  39422=>"000000000",
  39423=>"111111111",
  39424=>"111000000",
  39425=>"000010010",
  39426=>"111111111",
  39427=>"000000000",
  39428=>"000000000",
  39429=>"110110110",
  39430=>"000000000",
  39431=>"111111111",
  39432=>"100111100",
  39433=>"000111111",
  39434=>"000000110",
  39435=>"111011111",
  39436=>"011011111",
  39437=>"111100100",
  39438=>"011101111",
  39439=>"000000000",
  39440=>"111111111",
  39441=>"000000000",
  39442=>"111111111",
  39443=>"011111111",
  39444=>"111111111",
  39445=>"111111111",
  39446=>"110110000",
  39447=>"101001000",
  39448=>"000000000",
  39449=>"100000100",
  39450=>"101000000",
  39451=>"011011111",
  39452=>"111100000",
  39453=>"111000001",
  39454=>"000100100",
  39455=>"100100111",
  39456=>"111011011",
  39457=>"111111100",
  39458=>"001111001",
  39459=>"111111111",
  39460=>"001001011",
  39461=>"111111111",
  39462=>"111111101",
  39463=>"000000111",
  39464=>"111111111",
  39465=>"000000000",
  39466=>"000000000",
  39467=>"111101110",
  39468=>"000111111",
  39469=>"111111111",
  39470=>"000000000",
  39471=>"000000000",
  39472=>"010000111",
  39473=>"111111111",
  39474=>"100000000",
  39475=>"011011111",
  39476=>"001001001",
  39477=>"000011000",
  39478=>"110000000",
  39479=>"101111111",
  39480=>"000000000",
  39481=>"110000000",
  39482=>"000100000",
  39483=>"000000001",
  39484=>"000000000",
  39485=>"111111011",
  39486=>"111111111",
  39487=>"100100000",
  39488=>"111100000",
  39489=>"001000010",
  39490=>"000111111",
  39491=>"000000111",
  39492=>"101000100",
  39493=>"110000000",
  39494=>"101100000",
  39495=>"111111111",
  39496=>"000001000",
  39497=>"000000000",
  39498=>"111111011",
  39499=>"100001011",
  39500=>"000000000",
  39501=>"111111111",
  39502=>"111111111",
  39503=>"111111101",
  39504=>"011011011",
  39505=>"111111101",
  39506=>"111110000",
  39507=>"111011110",
  39508=>"011111011",
  39509=>"000000100",
  39510=>"110101001",
  39511=>"101111111",
  39512=>"011100110",
  39513=>"001000101",
  39514=>"010110110",
  39515=>"111101000",
  39516=>"000000000",
  39517=>"111111111",
  39518=>"100101001",
  39519=>"000000000",
  39520=>"100000000",
  39521=>"011000110",
  39522=>"000000000",
  39523=>"111111110",
  39524=>"000000000",
  39525=>"001001001",
  39526=>"000000111",
  39527=>"001000000",
  39528=>"100000000",
  39529=>"000101111",
  39530=>"100000001",
  39531=>"111111111",
  39532=>"010111100",
  39533=>"000000000",
  39534=>"001000001",
  39535=>"010000111",
  39536=>"111111111",
  39537=>"000000111",
  39538=>"000000000",
  39539=>"111100101",
  39540=>"000000000",
  39541=>"111101101",
  39542=>"000001011",
  39543=>"001000000",
  39544=>"001001000",
  39545=>"101000000",
  39546=>"111111111",
  39547=>"101000000",
  39548=>"111110110",
  39549=>"101111111",
  39550=>"000000001",
  39551=>"000000000",
  39552=>"100101111",
  39553=>"000111111",
  39554=>"000000000",
  39555=>"000101100",
  39556=>"000000001",
  39557=>"000000000",
  39558=>"000110110",
  39559=>"111111111",
  39560=>"111111111",
  39561=>"100100101",
  39562=>"000000100",
  39563=>"111111111",
  39564=>"000001001",
  39565=>"000111111",
  39566=>"111000000",
  39567=>"000000111",
  39568=>"000000000",
  39569=>"001001001",
  39570=>"111111111",
  39571=>"100000000",
  39572=>"011000000",
  39573=>"000100110",
  39574=>"000111111",
  39575=>"000000000",
  39576=>"000000000",
  39577=>"111111111",
  39578=>"000000000",
  39579=>"101111111",
  39580=>"100001000",
  39581=>"000000000",
  39582=>"000000111",
  39583=>"100111111",
  39584=>"110111111",
  39585=>"000000000",
  39586=>"000000000",
  39587=>"111111011",
  39588=>"111101111",
  39589=>"100100110",
  39590=>"111111111",
  39591=>"001110110",
  39592=>"001111111",
  39593=>"111111111",
  39594=>"000000001",
  39595=>"111111111",
  39596=>"000001001",
  39597=>"011111100",
  39598=>"111111111",
  39599=>"000000100",
  39600=>"111111000",
  39601=>"111111001",
  39602=>"000000000",
  39603=>"001000000",
  39604=>"000110100",
  39605=>"110111110",
  39606=>"000000000",
  39607=>"000000110",
  39608=>"111000000",
  39609=>"111000000",
  39610=>"111110110",
  39611=>"000001011",
  39612=>"001111111",
  39613=>"000001111",
  39614=>"111111111",
  39615=>"000111111",
  39616=>"111111111",
  39617=>"000000100",
  39618=>"101001001",
  39619=>"111111111",
  39620=>"100001000",
  39621=>"000110110",
  39622=>"001111000",
  39623=>"001001000",
  39624=>"000000000",
  39625=>"001000000",
  39626=>"111100100",
  39627=>"111111011",
  39628=>"111110110",
  39629=>"101101000",
  39630=>"000110111",
  39631=>"111001000",
  39632=>"000000000",
  39633=>"000001011",
  39634=>"111011000",
  39635=>"111101000",
  39636=>"100000100",
  39637=>"111111111",
  39638=>"000000000",
  39639=>"110110100",
  39640=>"000000000",
  39641=>"000100100",
  39642=>"111111111",
  39643=>"000000000",
  39644=>"000000001",
  39645=>"011111110",
  39646=>"000000000",
  39647=>"110111101",
  39648=>"000001001",
  39649=>"001100000",
  39650=>"100101111",
  39651=>"000011011",
  39652=>"111111111",
  39653=>"111111000",
  39654=>"111111111",
  39655=>"111111111",
  39656=>"111000000",
  39657=>"111001001",
  39658=>"101101001",
  39659=>"000000011",
  39660=>"000000000",
  39661=>"000000000",
  39662=>"000100100",
  39663=>"000000111",
  39664=>"001101000",
  39665=>"111111101",
  39666=>"111111001",
  39667=>"000001111",
  39668=>"000000000",
  39669=>"001001011",
  39670=>"000100110",
  39671=>"001111111",
  39672=>"000000000",
  39673=>"000001000",
  39674=>"100101101",
  39675=>"011010010",
  39676=>"000001001",
  39677=>"000000010",
  39678=>"110110100",
  39679=>"001000111",
  39680=>"000100111",
  39681=>"000000000",
  39682=>"000000000",
  39683=>"000010000",
  39684=>"110000000",
  39685=>"000110100",
  39686=>"000000000",
  39687=>"000111111",
  39688=>"111111111",
  39689=>"000000000",
  39690=>"111111110",
  39691=>"010000110",
  39692=>"000000100",
  39693=>"111000001",
  39694=>"000000001",
  39695=>"000000000",
  39696=>"011000000",
  39697=>"000000011",
  39698=>"000000000",
  39699=>"000111111",
  39700=>"111111111",
  39701=>"100000000",
  39702=>"111111111",
  39703=>"111111111",
  39704=>"111111111",
  39705=>"111111111",
  39706=>"000000000",
  39707=>"111111111",
  39708=>"000100000",
  39709=>"000000000",
  39710=>"110111111",
  39711=>"111001111",
  39712=>"001000000",
  39713=>"000000000",
  39714=>"000111011",
  39715=>"111111011",
  39716=>"100000000",
  39717=>"000000000",
  39718=>"000110011",
  39719=>"100101000",
  39720=>"001000000",
  39721=>"000000011",
  39722=>"010110111",
  39723=>"001001111",
  39724=>"011011011",
  39725=>"101000000",
  39726=>"100100000",
  39727=>"000000000",
  39728=>"111111111",
  39729=>"000111111",
  39730=>"000000000",
  39731=>"000000011",
  39732=>"111100100",
  39733=>"011011111",
  39734=>"111111111",
  39735=>"000000000",
  39736=>"000000010",
  39737=>"000000000",
  39738=>"111111111",
  39739=>"111111110",
  39740=>"000000000",
  39741=>"000111111",
  39742=>"000000000",
  39743=>"000000110",
  39744=>"000000000",
  39745=>"000000000",
  39746=>"101111111",
  39747=>"101001111",
  39748=>"000000000",
  39749=>"111110110",
  39750=>"111000100",
  39751=>"011011001",
  39752=>"000100100",
  39753=>"100100100",
  39754=>"100111111",
  39755=>"001110111",
  39756=>"111111111",
  39757=>"000010000",
  39758=>"000000100",
  39759=>"111111000",
  39760=>"000000000",
  39761=>"000100000",
  39762=>"101111001",
  39763=>"000000000",
  39764=>"111111101",
  39765=>"000000000",
  39766=>"110000000",
  39767=>"111111111",
  39768=>"001000000",
  39769=>"000001110",
  39770=>"000000011",
  39771=>"111111111",
  39772=>"100111111",
  39773=>"000000000",
  39774=>"000000011",
  39775=>"110110111",
  39776=>"111111110",
  39777=>"111111110",
  39778=>"111111011",
  39779=>"111111111",
  39780=>"011011001",
  39781=>"000000000",
  39782=>"001111111",
  39783=>"100111111",
  39784=>"100000000",
  39785=>"000000000",
  39786=>"000000000",
  39787=>"000000000",
  39788=>"000000000",
  39789=>"000001001",
  39790=>"000000000",
  39791=>"000000000",
  39792=>"000000000",
  39793=>"111110000",
  39794=>"111010111",
  39795=>"100100111",
  39796=>"010001001",
  39797=>"110001001",
  39798=>"000000000",
  39799=>"010010000",
  39800=>"011001111",
  39801=>"000001111",
  39802=>"110111111",
  39803=>"110111111",
  39804=>"111111110",
  39805=>"111111111",
  39806=>"000000111",
  39807=>"101111111",
  39808=>"111111001",
  39809=>"000000000",
  39810=>"011111111",
  39811=>"100100100",
  39812=>"000000000",
  39813=>"000000000",
  39814=>"100000000",
  39815=>"100000000",
  39816=>"100110100",
  39817=>"000000000",
  39818=>"111111111",
  39819=>"111111111",
  39820=>"000100111",
  39821=>"000110000",
  39822=>"111101111",
  39823=>"000110110",
  39824=>"111111000",
  39825=>"001111111",
  39826=>"000000000",
  39827=>"111111110",
  39828=>"001001000",
  39829=>"000000000",
  39830=>"000000000",
  39831=>"100100001",
  39832=>"000000000",
  39833=>"111000000",
  39834=>"111111111",
  39835=>"000010000",
  39836=>"000000000",
  39837=>"000000000",
  39838=>"111011000",
  39839=>"000000000",
  39840=>"110111111",
  39841=>"010011111",
  39842=>"000100101",
  39843=>"000001011",
  39844=>"101101111",
  39845=>"001011001",
  39846=>"111111111",
  39847=>"111110000",
  39848=>"000010000",
  39849=>"110100100",
  39850=>"000111111",
  39851=>"111000000",
  39852=>"000101110",
  39853=>"000000000",
  39854=>"000000000",
  39855=>"000000000",
  39856=>"100101000",
  39857=>"011111000",
  39858=>"000111001",
  39859=>"010111011",
  39860=>"111111111",
  39861=>"011001001",
  39862=>"001111001",
  39863=>"001001000",
  39864=>"000000111",
  39865=>"000000001",
  39866=>"000000111",
  39867=>"000000000",
  39868=>"001000111",
  39869=>"111000110",
  39870=>"110100101",
  39871=>"001011111",
  39872=>"000000000",
  39873=>"000000000",
  39874=>"111111111",
  39875=>"000000000",
  39876=>"000000000",
  39877=>"000001100",
  39878=>"000001011",
  39879=>"000000001",
  39880=>"000000001",
  39881=>"000000000",
  39882=>"000000101",
  39883=>"111000101",
  39884=>"001000000",
  39885=>"000000111",
  39886=>"000000001",
  39887=>"000110011",
  39888=>"011000000",
  39889=>"000000000",
  39890=>"111111111",
  39891=>"111011111",
  39892=>"000101101",
  39893=>"000000000",
  39894=>"000101111",
  39895=>"000000000",
  39896=>"100001010",
  39897=>"000111011",
  39898=>"000010110",
  39899=>"000000000",
  39900=>"111011110",
  39901=>"000000001",
  39902=>"000000000",
  39903=>"100100000",
  39904=>"001000001",
  39905=>"111111111",
  39906=>"000111111",
  39907=>"111111100",
  39908=>"001000011",
  39909=>"000111100",
  39910=>"000110100",
  39911=>"000111000",
  39912=>"000000111",
  39913=>"000101100",
  39914=>"000000011",
  39915=>"000000001",
  39916=>"000011111",
  39917=>"111111111",
  39918=>"001111111",
  39919=>"111111111",
  39920=>"111111111",
  39921=>"000000000",
  39922=>"100000001",
  39923=>"011011111",
  39924=>"000111001",
  39925=>"110111111",
  39926=>"111111111",
  39927=>"011111111",
  39928=>"111100000",
  39929=>"111111111",
  39930=>"101001011",
  39931=>"111111000",
  39932=>"000000000",
  39933=>"000101111",
  39934=>"110110000",
  39935=>"000000100",
  39936=>"100100000",
  39937=>"000000000",
  39938=>"111111000",
  39939=>"000000000",
  39940=>"000000000",
  39941=>"100000000",
  39942=>"011011111",
  39943=>"001000000",
  39944=>"111111111",
  39945=>"111111000",
  39946=>"000000000",
  39947=>"111011001",
  39948=>"111110100",
  39949=>"000000110",
  39950=>"110000100",
  39951=>"111111100",
  39952=>"000010000",
  39953=>"001111110",
  39954=>"100111111",
  39955=>"111001111",
  39956=>"000000110",
  39957=>"111111000",
  39958=>"000111111",
  39959=>"111111001",
  39960=>"000000110",
  39961=>"000000001",
  39962=>"001011111",
  39963=>"111111111",
  39964=>"111111111",
  39965=>"000000100",
  39966=>"100100101",
  39967=>"110111000",
  39968=>"001101000",
  39969=>"010000110",
  39970=>"000011011",
  39971=>"111111111",
  39972=>"000000001",
  39973=>"111101101",
  39974=>"000000000",
  39975=>"010000111",
  39976=>"000000000",
  39977=>"000000010",
  39978=>"111111001",
  39979=>"000011000",
  39980=>"000000000",
  39981=>"111111000",
  39982=>"111111111",
  39983=>"111110000",
  39984=>"110110111",
  39985=>"111011001",
  39986=>"111001001",
  39987=>"110000000",
  39988=>"000000001",
  39989=>"001001011",
  39990=>"000000000",
  39991=>"000000000",
  39992=>"011111100",
  39993=>"000000000",
  39994=>"000000000",
  39995=>"000001000",
  39996=>"001000001",
  39997=>"000000111",
  39998=>"000010000",
  39999=>"000000000",
  40000=>"110001000",
  40001=>"111011001",
  40002=>"111100111",
  40003=>"000000000",
  40004=>"000000000",
  40005=>"011000000",
  40006=>"110000000",
  40007=>"111111111",
  40008=>"011001000",
  40009=>"000100100",
  40010=>"111100010",
  40011=>"000000000",
  40012=>"111111000",
  40013=>"111111110",
  40014=>"010111111",
  40015=>"000000000",
  40016=>"000000000",
  40017=>"010000000",
  40018=>"000110111",
  40019=>"100100111",
  40020=>"110111110",
  40021=>"001111111",
  40022=>"111111000",
  40023=>"000000000",
  40024=>"111110111",
  40025=>"100111111",
  40026=>"111111100",
  40027=>"001001001",
  40028=>"111111111",
  40029=>"000000000",
  40030=>"111111000",
  40031=>"110111111",
  40032=>"000000000",
  40033=>"111111111",
  40034=>"100000000",
  40035=>"011011111",
  40036=>"111000000",
  40037=>"110110111",
  40038=>"000000110",
  40039=>"000000000",
  40040=>"000000000",
  40041=>"001011111",
  40042=>"000100111",
  40043=>"111100000",
  40044=>"000000010",
  40045=>"111111111",
  40046=>"000100111",
  40047=>"000000000",
  40048=>"010010000",
  40049=>"000000000",
  40050=>"111111111",
  40051=>"111001101",
  40052=>"111111111",
  40053=>"101111111",
  40054=>"010000000",
  40055=>"000000111",
  40056=>"111000000",
  40057=>"111000000",
  40058=>"100000000",
  40059=>"000000111",
  40060=>"111011011",
  40061=>"000110100",
  40062=>"111111111",
  40063=>"111011000",
  40064=>"100100000",
  40065=>"001011000",
  40066=>"000110111",
  40067=>"001000000",
  40068=>"001000001",
  40069=>"000000000",
  40070=>"111111111",
  40071=>"111111010",
  40072=>"111110111",
  40073=>"100100000",
  40074=>"111111111",
  40075=>"100100100",
  40076=>"101001000",
  40077=>"000000000",
  40078=>"111111100",
  40079=>"111111111",
  40080=>"000000111",
  40081=>"001000000",
  40082=>"000011011",
  40083=>"111011111",
  40084=>"111000000",
  40085=>"011000000",
  40086=>"000000000",
  40087=>"000000000",
  40088=>"111111011",
  40089=>"011111111",
  40090=>"111111111",
  40091=>"111000000",
  40092=>"000001001",
  40093=>"000000111",
  40094=>"100100000",
  40095=>"001000010",
  40096=>"000000001",
  40097=>"110110101",
  40098=>"111000000",
  40099=>"100111111",
  40100=>"011011111",
  40101=>"111011000",
  40102=>"111010110",
  40103=>"110100100",
  40104=>"111111111",
  40105=>"111000101",
  40106=>"111001001",
  40107=>"111000000",
  40108=>"000001100",
  40109=>"111011000",
  40110=>"000110011",
  40111=>"111111111",
  40112=>"011011000",
  40113=>"000001100",
  40114=>"111111110",
  40115=>"000000000",
  40116=>"000000000",
  40117=>"000011111",
  40118=>"111111111",
  40119=>"111111111",
  40120=>"110100000",
  40121=>"111111110",
  40122=>"111100100",
  40123=>"111111111",
  40124=>"000000000",
  40125=>"111110110",
  40126=>"111101111",
  40127=>"000001010",
  40128=>"000111111",
  40129=>"000110110",
  40130=>"001001000",
  40131=>"000000000",
  40132=>"111110000",
  40133=>"110100111",
  40134=>"001000001",
  40135=>"000000000",
  40136=>"111110111",
  40137=>"111000000",
  40138=>"101000111",
  40139=>"000111111",
  40140=>"000000111",
  40141=>"000111111",
  40142=>"000000100",
  40143=>"000000110",
  40144=>"111000000",
  40145=>"001000000",
  40146=>"011000000",
  40147=>"000000000",
  40148=>"000000111",
  40149=>"011111111",
  40150=>"110000000",
  40151=>"001010000",
  40152=>"000000111",
  40153=>"110000001",
  40154=>"000000111",
  40155=>"000000000",
  40156=>"111111111",
  40157=>"110100000",
  40158=>"111011000",
  40159=>"100110110",
  40160=>"000000000",
  40161=>"001000100",
  40162=>"111111111",
  40163=>"111100000",
  40164=>"111101101",
  40165=>"110111001",
  40166=>"111111111",
  40167=>"111111111",
  40168=>"001011111",
  40169=>"111111111",
  40170=>"000001111",
  40171=>"000001111",
  40172=>"010010000",
  40173=>"110111111",
  40174=>"111111111",
  40175=>"000000000",
  40176=>"111100101",
  40177=>"111101101",
  40178=>"000000000",
  40179=>"001111111",
  40180=>"000001111",
  40181=>"001101111",
  40182=>"000000000",
  40183=>"000000000",
  40184=>"111111111",
  40185=>"110111111",
  40186=>"000000000",
  40187=>"000011011",
  40188=>"111101001",
  40189=>"000000010",
  40190=>"000110111",
  40191=>"000000000",
  40192=>"011111100",
  40193=>"111011000",
  40194=>"011000110",
  40195=>"000100111",
  40196=>"000000000",
  40197=>"001111011",
  40198=>"000000000",
  40199=>"000101100",
  40200=>"000000000",
  40201=>"000111111",
  40202=>"111110000",
  40203=>"011001000",
  40204=>"111111111",
  40205=>"001001000",
  40206=>"111111111",
  40207=>"000000000",
  40208=>"000100111",
  40209=>"100010000",
  40210=>"000000111",
  40211=>"000000000",
  40212=>"000001010",
  40213=>"110111111",
  40214=>"111111111",
  40215=>"001000001",
  40216=>"011111111",
  40217=>"111000000",
  40218=>"110010000",
  40219=>"011000000",
  40220=>"011000000",
  40221=>"111101111",
  40222=>"111001000",
  40223=>"110100000",
  40224=>"111011100",
  40225=>"111111100",
  40226=>"111110100",
  40227=>"000000000",
  40228=>"110110111",
  40229=>"111100000",
  40230=>"001011001",
  40231=>"000101000",
  40232=>"110111110",
  40233=>"111011111",
  40234=>"000110110",
  40235=>"000000000",
  40236=>"000000000",
  40237=>"001001000",
  40238=>"100000000",
  40239=>"000000001",
  40240=>"000000000",
  40241=>"000000000",
  40242=>"000010111",
  40243=>"000000000",
  40244=>"000100111",
  40245=>"111000000",
  40246=>"000000000",
  40247=>"111111111",
  40248=>"000011011",
  40249=>"000000101",
  40250=>"110100111",
  40251=>"000000100",
  40252=>"110000000",
  40253=>"000000000",
  40254=>"111111101",
  40255=>"111111001",
  40256=>"111100000",
  40257=>"000100111",
  40258=>"100000010",
  40259=>"111111000",
  40260=>"011011111",
  40261=>"010001000",
  40262=>"000000110",
  40263=>"111111111",
  40264=>"111111111",
  40265=>"000000000",
  40266=>"111110100",
  40267=>"110110000",
  40268=>"101111100",
  40269=>"000000000",
  40270=>"010110110",
  40271=>"001001111",
  40272=>"000011011",
  40273=>"001011001",
  40274=>"000000001",
  40275=>"000000000",
  40276=>"101101111",
  40277=>"100100110",
  40278=>"111011000",
  40279=>"000000100",
  40280=>"110111111",
  40281=>"001001001",
  40282=>"111111111",
  40283=>"000000000",
  40284=>"000000000",
  40285=>"111111101",
  40286=>"001001111",
  40287=>"011111100",
  40288=>"111000000",
  40289=>"000000100",
  40290=>"011011111",
  40291=>"001000111",
  40292=>"001011011",
  40293=>"000000000",
  40294=>"000111111",
  40295=>"110111000",
  40296=>"001000000",
  40297=>"000000111",
  40298=>"011011001",
  40299=>"000001001",
  40300=>"000000000",
  40301=>"001000011",
  40302=>"011011111",
  40303=>"111111111",
  40304=>"110111111",
  40305=>"000011001",
  40306=>"000000011",
  40307=>"100100110",
  40308=>"111111111",
  40309=>"110100000",
  40310=>"111011011",
  40311=>"000000010",
  40312=>"111111111",
  40313=>"000100111",
  40314=>"100110000",
  40315=>"000000000",
  40316=>"000100111",
  40317=>"000000000",
  40318=>"110000000",
  40319=>"111111000",
  40320=>"011011111",
  40321=>"110110111",
  40322=>"000100111",
  40323=>"001000111",
  40324=>"000001001",
  40325=>"110000000",
  40326=>"101111111",
  40327=>"010000000",
  40328=>"111111111",
  40329=>"000000000",
  40330=>"001000000",
  40331=>"111100101",
  40332=>"111111110",
  40333=>"000100100",
  40334=>"000000000",
  40335=>"000010111",
  40336=>"000001011",
  40337=>"000000000",
  40338=>"110010111",
  40339=>"111110000",
  40340=>"110111111",
  40341=>"000000000",
  40342=>"101001000",
  40343=>"110110010",
  40344=>"111111111",
  40345=>"111111111",
  40346=>"011011111",
  40347=>"111100100",
  40348=>"000010000",
  40349=>"000000000",
  40350=>"000000111",
  40351=>"000000000",
  40352=>"111111111",
  40353=>"000100111",
  40354=>"000111000",
  40355=>"000000000",
  40356=>"111111100",
  40357=>"010000000",
  40358=>"111000001",
  40359=>"111111111",
  40360=>"011000000",
  40361=>"111100000",
  40362=>"111111001",
  40363=>"001001111",
  40364=>"000000000",
  40365=>"000000000",
  40366=>"000001111",
  40367=>"000000111",
  40368=>"110110111",
  40369=>"111000000",
  40370=>"000000111",
  40371=>"000000000",
  40372=>"000111111",
  40373=>"100110111",
  40374=>"111111111",
  40375=>"111000000",
  40376=>"000000110",
  40377=>"111111111",
  40378=>"000000000",
  40379=>"000000000",
  40380=>"000000000",
  40381=>"111011000",
  40382=>"100000000",
  40383=>"001000011",
  40384=>"000000000",
  40385=>"111101000",
  40386=>"111010010",
  40387=>"000001000",
  40388=>"000111111",
  40389=>"111101001",
  40390=>"000001001",
  40391=>"111000001",
  40392=>"000000100",
  40393=>"111111111",
  40394=>"000000000",
  40395=>"000000000",
  40396=>"110110110",
  40397=>"111111011",
  40398=>"111110000",
  40399=>"111111100",
  40400=>"111000001",
  40401=>"000011000",
  40402=>"110000110",
  40403=>"000000111",
  40404=>"111110110",
  40405=>"100000000",
  40406=>"000000000",
  40407=>"100000001",
  40408=>"001010111",
  40409=>"000000001",
  40410=>"111111111",
  40411=>"111100100",
  40412=>"101111111",
  40413=>"000000111",
  40414=>"000111000",
  40415=>"110000100",
  40416=>"011001011",
  40417=>"001011111",
  40418=>"000000000",
  40419=>"000000000",
  40420=>"000000000",
  40421=>"001000000",
  40422=>"111111001",
  40423=>"100100100",
  40424=>"000000000",
  40425=>"000111100",
  40426=>"000000101",
  40427=>"000000111",
  40428=>"000111111",
  40429=>"000100000",
  40430=>"111010000",
  40431=>"011111110",
  40432=>"111111111",
  40433=>"000000001",
  40434=>"111011011",
  40435=>"011001001",
  40436=>"111111111",
  40437=>"011000100",
  40438=>"111111111",
  40439=>"001011111",
  40440=>"011001000",
  40441=>"100101111",
  40442=>"000001111",
  40443=>"110001000",
  40444=>"000000000",
  40445=>"111111111",
  40446=>"000000000",
  40447=>"111011011",
  40448=>"000000000",
  40449=>"000000100",
  40450=>"000000000",
  40451=>"111111000",
  40452=>"000110111",
  40453=>"000000000",
  40454=>"000000001",
  40455=>"000111111",
  40456=>"111011011",
  40457=>"010000000",
  40458=>"000000000",
  40459=>"001000000",
  40460=>"110110111",
  40461=>"101101111",
  40462=>"000011011",
  40463=>"000000000",
  40464=>"011111000",
  40465=>"111000111",
  40466=>"110110000",
  40467=>"111111111",
  40468=>"000000100",
  40469=>"000000001",
  40470=>"000000000",
  40471=>"010011000",
  40472=>"001011111",
  40473=>"000000000",
  40474=>"111111111",
  40475=>"001101100",
  40476=>"000000000",
  40477=>"111110000",
  40478=>"011110100",
  40479=>"100100111",
  40480=>"011111000",
  40481=>"110111100",
  40482=>"010100101",
  40483=>"111111111",
  40484=>"000000000",
  40485=>"000000000",
  40486=>"001001000",
  40487=>"111011000",
  40488=>"010000001",
  40489=>"000000000",
  40490=>"111111111",
  40491=>"111111111",
  40492=>"111110110",
  40493=>"000000000",
  40494=>"000001010",
  40495=>"111111111",
  40496=>"000111100",
  40497=>"000011011",
  40498=>"000000000",
  40499=>"000011010",
  40500=>"111111111",
  40501=>"110110000",
  40502=>"000000000",
  40503=>"111101101",
  40504=>"000000000",
  40505=>"011111110",
  40506=>"011111111",
  40507=>"111011111",
  40508=>"000000100",
  40509=>"111110100",
  40510=>"001001001",
  40511=>"011111111",
  40512=>"011111110",
  40513=>"101101000",
  40514=>"111111110",
  40515=>"011011000",
  40516=>"011011111",
  40517=>"000000100",
  40518=>"111111111",
  40519=>"111111000",
  40520=>"111111011",
  40521=>"000000000",
  40522=>"000000000",
  40523=>"000000011",
  40524=>"011010110",
  40525=>"100000000",
  40526=>"011000110",
  40527=>"111111111",
  40528=>"001000000",
  40529=>"011000000",
  40530=>"000000000",
  40531=>"000011110",
  40532=>"010010011",
  40533=>"111111111",
  40534=>"010000000",
  40535=>"011111110",
  40536=>"111111001",
  40537=>"000000100",
  40538=>"100111111",
  40539=>"111101101",
  40540=>"111001111",
  40541=>"000000000",
  40542=>"001111100",
  40543=>"101011011",
  40544=>"001000000",
  40545=>"000000100",
  40546=>"011000000",
  40547=>"000000111",
  40548=>"000001000",
  40549=>"110110110",
  40550=>"101111111",
  40551=>"111111111",
  40552=>"111111111",
  40553=>"001000000",
  40554=>"001111111",
  40555=>"111000000",
  40556=>"000000000",
  40557=>"000000010",
  40558=>"000000000",
  40559=>"111111110",
  40560=>"000000110",
  40561=>"011001101",
  40562=>"011111111",
  40563=>"000111111",
  40564=>"100000000",
  40565=>"111010000",
  40566=>"111111111",
  40567=>"111111111",
  40568=>"000000000",
  40569=>"111111111",
  40570=>"111001000",
  40571=>"111111111",
  40572=>"000000000",
  40573=>"000101001",
  40574=>"011000000",
  40575=>"000000000",
  40576=>"111111111",
  40577=>"011000111",
  40578=>"100101000",
  40579=>"000001001",
  40580=>"111001001",
  40581=>"000000000",
  40582=>"000000000",
  40583=>"001000000",
  40584=>"111111111",
  40585=>"001000111",
  40586=>"001011000",
  40587=>"000000000",
  40588=>"011111100",
  40589=>"000000001",
  40590=>"011110100",
  40591=>"111110110",
  40592=>"100101111",
  40593=>"000000000",
  40594=>"100110111",
  40595=>"110111111",
  40596=>"000100000",
  40597=>"100000000",
  40598=>"000000101",
  40599=>"111111111",
  40600=>"001000100",
  40601=>"010111111",
  40602=>"011000000",
  40603=>"110111111",
  40604=>"000000000",
  40605=>"000000110",
  40606=>"111110110",
  40607=>"001111000",
  40608=>"000000000",
  40609=>"111111111",
  40610=>"111001000",
  40611=>"000000000",
  40612=>"110110110",
  40613=>"011111110",
  40614=>"000101111",
  40615=>"000000001",
  40616=>"111110111",
  40617=>"111111111",
  40618=>"110111111",
  40619=>"000000000",
  40620=>"001001001",
  40621=>"111111100",
  40622=>"010010011",
  40623=>"011011101",
  40624=>"111111000",
  40625=>"001111111",
  40626=>"111111111",
  40627=>"111111111",
  40628=>"000001001",
  40629=>"111000000",
  40630=>"111111111",
  40631=>"111111111",
  40632=>"010000000",
  40633=>"000111111",
  40634=>"000000000",
  40635=>"011111111",
  40636=>"100100101",
  40637=>"001000000",
  40638=>"000001101",
  40639=>"000000000",
  40640=>"111100100",
  40641=>"000000000",
  40642=>"110001000",
  40643=>"110110111",
  40644=>"000001111",
  40645=>"001111111",
  40646=>"111111111",
  40647=>"000000000",
  40648=>"001001000",
  40649=>"001000000",
  40650=>"000000100",
  40651=>"000000000",
  40652=>"011011100",
  40653=>"001011011",
  40654=>"111111001",
  40655=>"110100000",
  40656=>"111111111",
  40657=>"011000000",
  40658=>"011001101",
  40659=>"000111111",
  40660=>"001111111",
  40661=>"000000000",
  40662=>"000111111",
  40663=>"111111100",
  40664=>"111100000",
  40665=>"110101000",
  40666=>"111100100",
  40667=>"111010110",
  40668=>"111111000",
  40669=>"111111111",
  40670=>"110111111",
  40671=>"000000000",
  40672=>"110111000",
  40673=>"111011000",
  40674=>"111001111",
  40675=>"110010000",
  40676=>"100000000",
  40677=>"111111011",
  40678=>"111101000",
  40679=>"111111111",
  40680=>"111111111",
  40681=>"111110100",
  40682=>"110000100",
  40683=>"001111111",
  40684=>"000011111",
  40685=>"100111111",
  40686=>"100000001",
  40687=>"011000001",
  40688=>"111111000",
  40689=>"000000000",
  40690=>"100111100",
  40691=>"000110100",
  40692=>"000011011",
  40693=>"111111111",
  40694=>"011011011",
  40695=>"110010110",
  40696=>"011011000",
  40697=>"011011111",
  40698=>"111111111",
  40699=>"001001001",
  40700=>"011111111",
  40701=>"000010110",
  40702=>"111111111",
  40703=>"001000000",
  40704=>"000000111",
  40705=>"000000111",
  40706=>"111111111",
  40707=>"000111000",
  40708=>"100101111",
  40709=>"000000000",
  40710=>"000101111",
  40711=>"011001000",
  40712=>"111111111",
  40713=>"000000000",
  40714=>"111111111",
  40715=>"011011001",
  40716=>"101100100",
  40717=>"011000100",
  40718=>"000000000",
  40719=>"111110111",
  40720=>"000001111",
  40721=>"000000100",
  40722=>"000000000",
  40723=>"000000001",
  40724=>"111111111",
  40725=>"111111110",
  40726=>"000000001",
  40727=>"011011011",
  40728=>"111111110",
  40729=>"100010000",
  40730=>"000000001",
  40731=>"101101101",
  40732=>"000000000",
  40733=>"111111111",
  40734=>"101100000",
  40735=>"100000001",
  40736=>"011001011",
  40737=>"111111111",
  40738=>"111111011",
  40739=>"111101101",
  40740=>"111111111",
  40741=>"001001111",
  40742=>"001100110",
  40743=>"011011001",
  40744=>"110111000",
  40745=>"000000000",
  40746=>"111011111",
  40747=>"000000011",
  40748=>"010011001",
  40749=>"000110111",
  40750=>"111111111",
  40751=>"000000000",
  40752=>"100000000",
  40753=>"111101101",
  40754=>"001111111",
  40755=>"000000000",
  40756=>"000001111",
  40757=>"000000001",
  40758=>"111110111",
  40759=>"001001000",
  40760=>"000000000",
  40761=>"000000000",
  40762=>"110111011",
  40763=>"000011111",
  40764=>"111110100",
  40765=>"001000011",
  40766=>"000000000",
  40767=>"011011011",
  40768=>"000000111",
  40769=>"100111000",
  40770=>"011001000",
  40771=>"000000000",
  40772=>"000000100",
  40773=>"111111111",
  40774=>"000000000",
  40775=>"111111111",
  40776=>"000000000",
  40777=>"001000000",
  40778=>"001100110",
  40779=>"000000000",
  40780=>"111011011",
  40781=>"111000000",
  40782=>"011111000",
  40783=>"000110110",
  40784=>"110100000",
  40785=>"111101111",
  40786=>"000000000",
  40787=>"111111110",
  40788=>"000000000",
  40789=>"001001011",
  40790=>"000000100",
  40791=>"111111001",
  40792=>"000000000",
  40793=>"000000111",
  40794=>"000000000",
  40795=>"110011011",
  40796=>"000000001",
  40797=>"000000000",
  40798=>"011001111",
  40799=>"111111010",
  40800=>"011111111",
  40801=>"111001111",
  40802=>"011011011",
  40803=>"110111111",
  40804=>"111110111",
  40805=>"000000000",
  40806=>"111111111",
  40807=>"111111111",
  40808=>"001001101",
  40809=>"000000111",
  40810=>"111001000",
  40811=>"000011111",
  40812=>"100010000",
  40813=>"011011011",
  40814=>"111111111",
  40815=>"000011011",
  40816=>"111111111",
  40817=>"000000000",
  40818=>"011001001",
  40819=>"000000000",
  40820=>"000000000",
  40821=>"000000000",
  40822=>"000000000",
  40823=>"000000000",
  40824=>"000000000",
  40825=>"011000011",
  40826=>"100111111",
  40827=>"000000000",
  40828=>"111101101",
  40829=>"000000000",
  40830=>"001000000",
  40831=>"000000000",
  40832=>"000000000",
  40833=>"010000100",
  40834=>"000000000",
  40835=>"000000100",
  40836=>"000000000",
  40837=>"000111000",
  40838=>"101100000",
  40839=>"011111000",
  40840=>"001101101",
  40841=>"100100000",
  40842=>"100000000",
  40843=>"111111101",
  40844=>"101001111",
  40845=>"001101111",
  40846=>"001001101",
  40847=>"001001111",
  40848=>"000000000",
  40849=>"111111111",
  40850=>"010001000",
  40851=>"011011111",
  40852=>"111111000",
  40853=>"000001011",
  40854=>"000000000",
  40855=>"111010000",
  40856=>"000000000",
  40857=>"011011110",
  40858=>"000000000",
  40859=>"000000000",
  40860=>"100111101",
  40861=>"000000000",
  40862=>"000111111",
  40863=>"000101111",
  40864=>"110000000",
  40865=>"111111101",
  40866=>"001001101",
  40867=>"111000000",
  40868=>"001101000",
  40869=>"111111111",
  40870=>"001000111",
  40871=>"000000000",
  40872=>"111111111",
  40873=>"000000000",
  40874=>"110110111",
  40875=>"000000100",
  40876=>"111101111",
  40877=>"111001100",
  40878=>"110110111",
  40879=>"000000000",
  40880=>"000000000",
  40881=>"111111111",
  40882=>"111000000",
  40883=>"111110101",
  40884=>"000111111",
  40885=>"111111110",
  40886=>"000110111",
  40887=>"000101111",
  40888=>"000000110",
  40889=>"111111111",
  40890=>"011111011",
  40891=>"111111111",
  40892=>"111111010",
  40893=>"111000011",
  40894=>"111001011",
  40895=>"011011111",
  40896=>"111111111",
  40897=>"000000000",
  40898=>"000000001",
  40899=>"001001111",
  40900=>"000000000",
  40901=>"000000000",
  40902=>"111000000",
  40903=>"111111111",
  40904=>"111011110",
  40905=>"000111111",
  40906=>"111111111",
  40907=>"111111111",
  40908=>"011001000",
  40909=>"111111111",
  40910=>"100000000",
  40911=>"110000110",
  40912=>"010011110",
  40913=>"000000001",
  40914=>"001000000",
  40915=>"000000000",
  40916=>"011111111",
  40917=>"000000001",
  40918=>"111111111",
  40919=>"100100110",
  40920=>"000000100",
  40921=>"110110000",
  40922=>"110100000",
  40923=>"000001000",
  40924=>"000000000",
  40925=>"111111111",
  40926=>"000001001",
  40927=>"000001111",
  40928=>"000000110",
  40929=>"000000000",
  40930=>"100111110",
  40931=>"111111111",
  40932=>"110111111",
  40933=>"000000000",
  40934=>"000001001",
  40935=>"110100100",
  40936=>"010011100",
  40937=>"100000001",
  40938=>"000000100",
  40939=>"111111011",
  40940=>"100000000",
  40941=>"111111000",
  40942=>"000000000",
  40943=>"000000101",
  40944=>"111111011",
  40945=>"111111011",
  40946=>"000000000",
  40947=>"111111111",
  40948=>"011111111",
  40949=>"101101101",
  40950=>"000000000",
  40951=>"001100111",
  40952=>"010000001",
  40953=>"000010001",
  40954=>"000000110",
  40955=>"011111111",
  40956=>"111111010",
  40957=>"000100000",
  40958=>"000000000",
  40959=>"000000010",
  40960=>"000011000",
  40961=>"010110000",
  40962=>"000000101",
  40963=>"011111000",
  40964=>"001111111",
  40965=>"000001111",
  40966=>"000000000",
  40967=>"111111111",
  40968=>"111111000",
  40969=>"000100111",
  40970=>"111100110",
  40971=>"111111111",
  40972=>"000000000",
  40973=>"110010111",
  40974=>"111110100",
  40975=>"111111001",
  40976=>"011011011",
  40977=>"000000111",
  40978=>"111111111",
  40979=>"111111111",
  40980=>"110111000",
  40981=>"111000000",
  40982=>"001101100",
  40983=>"111100100",
  40984=>"110110000",
  40985=>"001001100",
  40986=>"111000111",
  40987=>"000001101",
  40988=>"101111000",
  40989=>"000000000",
  40990=>"111000000",
  40991=>"000000000",
  40992=>"001011000",
  40993=>"110010000",
  40994=>"010001001",
  40995=>"001001010",
  40996=>"011001011",
  40997=>"001111111",
  40998=>"111111111",
  40999=>"000100100",
  41000=>"000000000",
  41001=>"110110110",
  41002=>"000100110",
  41003=>"111111111",
  41004=>"111111001",
  41005=>"000001000",
  41006=>"000000010",
  41007=>"011000000",
  41008=>"111101000",
  41009=>"111111111",
  41010=>"110111000",
  41011=>"000110110",
  41012=>"000001000",
  41013=>"100111111",
  41014=>"001101111",
  41015=>"000110100",
  41016=>"110111111",
  41017=>"101111111",
  41018=>"000011111",
  41019=>"111110000",
  41020=>"001100110",
  41021=>"111101111",
  41022=>"000000000",
  41023=>"111000111",
  41024=>"110110000",
  41025=>"000011010",
  41026=>"000000010",
  41027=>"111111010",
  41028=>"000000000",
  41029=>"111111110",
  41030=>"100111000",
  41031=>"110010000",
  41032=>"000001011",
  41033=>"000001111",
  41034=>"000000100",
  41035=>"110111010",
  41036=>"000110101",
  41037=>"111110000",
  41038=>"100000011",
  41039=>"111111111",
  41040=>"110111111",
  41041=>"111000111",
  41042=>"000000000",
  41043=>"001011011",
  41044=>"101001000",
  41045=>"100100110",
  41046=>"111110011",
  41047=>"000000000",
  41048=>"101111111",
  41049=>"111101111",
  41050=>"010000000",
  41051=>"110110000",
  41052=>"110000011",
  41053=>"110111111",
  41054=>"000100111",
  41055=>"100000001",
  41056=>"010000110",
  41057=>"000000000",
  41058=>"111111111",
  41059=>"000000011",
  41060=>"000110010",
  41061=>"111111000",
  41062=>"010011011",
  41063=>"111000101",
  41064=>"000000000",
  41065=>"000000010",
  41066=>"011000001",
  41067=>"000000000",
  41068=>"000000111",
  41069=>"001001001",
  41070=>"000001111",
  41071=>"110000111",
  41072=>"000011111",
  41073=>"000111111",
  41074=>"000001001",
  41075=>"000000111",
  41076=>"011001100",
  41077=>"000100110",
  41078=>"010010110",
  41079=>"111110000",
  41080=>"000000000",
  41081=>"111101000",
  41082=>"000001000",
  41083=>"100000011",
  41084=>"000000000",
  41085=>"100110111",
  41086=>"000000000",
  41087=>"111111011",
  41088=>"000101100",
  41089=>"111111011",
  41090=>"111011011",
  41091=>"000001000",
  41092=>"001001001",
  41093=>"001000000",
  41094=>"100110000",
  41095=>"000011111",
  41096=>"111111011",
  41097=>"000000000",
  41098=>"000000000",
  41099=>"000111111",
  41100=>"111111101",
  41101=>"111111000",
  41102=>"111111110",
  41103=>"000001111",
  41104=>"000000000",
  41105=>"111111111",
  41106=>"000111111",
  41107=>"000100000",
  41108=>"000011001",
  41109=>"101001001",
  41110=>"100111111",
  41111=>"000011111",
  41112=>"000001111",
  41113=>"011111101",
  41114=>"110110110",
  41115=>"010011001",
  41116=>"111100100",
  41117=>"111000000",
  41118=>"111111111",
  41119=>"011111111",
  41120=>"111110110",
  41121=>"111011011",
  41122=>"111000111",
  41123=>"001000000",
  41124=>"000010001",
  41125=>"111000111",
  41126=>"010001111",
  41127=>"101101101",
  41128=>"110111000",
  41129=>"000111111",
  41130=>"110111000",
  41131=>"101000001",
  41132=>"000000111",
  41133=>"000001000",
  41134=>"111111111",
  41135=>"000011001",
  41136=>"110111111",
  41137=>"111010011",
  41138=>"011001011",
  41139=>"010111111",
  41140=>"111001011",
  41141=>"101100100",
  41142=>"100101111",
  41143=>"111111110",
  41144=>"001000000",
  41145=>"111111111",
  41146=>"000000000",
  41147=>"001001100",
  41148=>"100000000",
  41149=>"001111111",
  41150=>"111111100",
  41151=>"011111111",
  41152=>"001001000",
  41153=>"010000000",
  41154=>"000000111",
  41155=>"111111111",
  41156=>"100111111",
  41157=>"000111111",
  41158=>"010010000",
  41159=>"001111101",
  41160=>"010110111",
  41161=>"100111001",
  41162=>"000000111",
  41163=>"011001101",
  41164=>"100001011",
  41165=>"111110110",
  41166=>"000000010",
  41167=>"110000000",
  41168=>"110010110",
  41169=>"000000111",
  41170=>"000010111",
  41171=>"000000000",
  41172=>"000101111",
  41173=>"010000001",
  41174=>"000110110",
  41175=>"000100100",
  41176=>"111111101",
  41177=>"000000111",
  41178=>"000110110",
  41179=>"000111001",
  41180=>"010110111",
  41181=>"000000000",
  41182=>"000111001",
  41183=>"101001001",
  41184=>"000000000",
  41185=>"111111111",
  41186=>"000000111",
  41187=>"111110000",
  41188=>"000000000",
  41189=>"011011001",
  41190=>"000110111",
  41191=>"110110000",
  41192=>"101111111",
  41193=>"111110000",
  41194=>"100100100",
  41195=>"100111111",
  41196=>"111111111",
  41197=>"000010100",
  41198=>"111000000",
  41199=>"000001000",
  41200=>"110110000",
  41201=>"111000000",
  41202=>"100000111",
  41203=>"001011111",
  41204=>"000110110",
  41205=>"011001111",
  41206=>"000111111",
  41207=>"000000001",
  41208=>"000000011",
  41209=>"001000001",
  41210=>"000000100",
  41211=>"111111111",
  41212=>"100100000",
  41213=>"111001000",
  41214=>"111000000",
  41215=>"101000000",
  41216=>"001000100",
  41217=>"000100100",
  41218=>"011111000",
  41219=>"101000001",
  41220=>"000111110",
  41221=>"001111111",
  41222=>"111011000",
  41223=>"000111001",
  41224=>"110111101",
  41225=>"100100111",
  41226=>"010111001",
  41227=>"000011111",
  41228=>"001101111",
  41229=>"000000111",
  41230=>"000000101",
  41231=>"111110100",
  41232=>"111000000",
  41233=>"000000000",
  41234=>"100000000",
  41235=>"111111001",
  41236=>"000000111",
  41237=>"000000101",
  41238=>"000100100",
  41239=>"000001000",
  41240=>"001001100",
  41241=>"110110111",
  41242=>"001111111",
  41243=>"111111111",
  41244=>"001000000",
  41245=>"000000001",
  41246=>"111111111",
  41247=>"000000001",
  41248=>"000000000",
  41249=>"000001001",
  41250=>"000001001",
  41251=>"111111111",
  41252=>"010110110",
  41253=>"111111111",
  41254=>"001001001",
  41255=>"000110111",
  41256=>"111001000",
  41257=>"000010111",
  41258=>"000000000",
  41259=>"001111110",
  41260=>"000100110",
  41261=>"000000111",
  41262=>"000000111",
  41263=>"000001001",
  41264=>"100101001",
  41265=>"111000111",
  41266=>"011011000",
  41267=>"010110111",
  41268=>"011000000",
  41269=>"100000001",
  41270=>"111000011",
  41271=>"000011000",
  41272=>"011111000",
  41273=>"111100111",
  41274=>"111111110",
  41275=>"110101000",
  41276=>"011100000",
  41277=>"111101000",
  41278=>"111111111",
  41279=>"000001000",
  41280=>"000000000",
  41281=>"111000001",
  41282=>"100100000",
  41283=>"001001000",
  41284=>"000000000",
  41285=>"111100000",
  41286=>"110111111",
  41287=>"000001011",
  41288=>"111001000",
  41289=>"000010010",
  41290=>"110011001",
  41291=>"001011011",
  41292=>"110110100",
  41293=>"110101111",
  41294=>"100100110",
  41295=>"000111111",
  41296=>"111011000",
  41297=>"101111000",
  41298=>"001111111",
  41299=>"101001001",
  41300=>"000000000",
  41301=>"000001011",
  41302=>"000000000",
  41303=>"111100111",
  41304=>"111011011",
  41305=>"010000000",
  41306=>"110000000",
  41307=>"000000110",
  41308=>"000001001",
  41309=>"100110110",
  41310=>"000010111",
  41311=>"000111011",
  41312=>"001001001",
  41313=>"000000000",
  41314=>"110111111",
  41315=>"001111111",
  41316=>"000011011",
  41317=>"001001011",
  41318=>"111111111",
  41319=>"000001111",
  41320=>"000110110",
  41321=>"000010000",
  41322=>"111111000",
  41323=>"101000110",
  41324=>"001001011",
  41325=>"111011011",
  41326=>"001001000",
  41327=>"000000110",
  41328=>"000000111",
  41329=>"111100100",
  41330=>"111000000",
  41331=>"001000000",
  41332=>"111100100",
  41333=>"010000110",
  41334=>"111101000",
  41335=>"100110000",
  41336=>"011011011",
  41337=>"110110111",
  41338=>"000000001",
  41339=>"111010011",
  41340=>"000111111",
  41341=>"001111110",
  41342=>"111000000",
  41343=>"111111111",
  41344=>"000000000",
  41345=>"001001001",
  41346=>"100000011",
  41347=>"100111000",
  41348=>"100100110",
  41349=>"000000000",
  41350=>"000000110",
  41351=>"010110000",
  41352=>"010011000",
  41353=>"001101100",
  41354=>"000000111",
  41355=>"011011000",
  41356=>"111111111",
  41357=>"101101100",
  41358=>"011100001",
  41359=>"010000111",
  41360=>"000001001",
  41361=>"110010010",
  41362=>"111111000",
  41363=>"110000001",
  41364=>"101001111",
  41365=>"000110110",
  41366=>"011111110",
  41367=>"001001001",
  41368=>"110111110",
  41369=>"111010000",
  41370=>"101000000",
  41371=>"111111000",
  41372=>"000100000",
  41373=>"110000000",
  41374=>"000001111",
  41375=>"001001010",
  41376=>"111001000",
  41377=>"100100100",
  41378=>"000000000",
  41379=>"110100000",
  41380=>"000100000",
  41381=>"011011011",
  41382=>"110000011",
  41383=>"111111001",
  41384=>"000000011",
  41385=>"110111111",
  41386=>"000001100",
  41387=>"000011011",
  41388=>"110100100",
  41389=>"111000000",
  41390=>"100000101",
  41391=>"110111000",
  41392=>"110000011",
  41393=>"111111101",
  41394=>"011000001",
  41395=>"110111111",
  41396=>"000001001",
  41397=>"001000110",
  41398=>"000111110",
  41399=>"101011111",
  41400=>"111010101",
  41401=>"000011111",
  41402=>"000000100",
  41403=>"011000000",
  41404=>"111000000",
  41405=>"010011010",
  41406=>"000000000",
  41407=>"100100000",
  41408=>"000011000",
  41409=>"110111111",
  41410=>"000111111",
  41411=>"111111111",
  41412=>"111100000",
  41413=>"010000000",
  41414=>"000000001",
  41415=>"000000001",
  41416=>"000000100",
  41417=>"000100100",
  41418=>"000111001",
  41419=>"000000010",
  41420=>"000000000",
  41421=>"001001011",
  41422=>"000011001",
  41423=>"111111000",
  41424=>"000011011",
  41425=>"000001111",
  41426=>"000000001",
  41427=>"000111111",
  41428=>"000111111",
  41429=>"111000000",
  41430=>"000000110",
  41431=>"000000000",
  41432=>"100101101",
  41433=>"110000010",
  41434=>"000000111",
  41435=>"000100000",
  41436=>"011011000",
  41437=>"111001011",
  41438=>"011111001",
  41439=>"110100000",
  41440=>"000101000",
  41441=>"000111101",
  41442=>"001000111",
  41443=>"010111111",
  41444=>"110010111",
  41445=>"110110000",
  41446=>"011001001",
  41447=>"100100111",
  41448=>"111111001",
  41449=>"111001000",
  41450=>"011010111",
  41451=>"111111101",
  41452=>"000100111",
  41453=>"111111000",
  41454=>"001101000",
  41455=>"000111111",
  41456=>"001000000",
  41457=>"111111011",
  41458=>"100011111",
  41459=>"000011001",
  41460=>"000110111",
  41461=>"100000100",
  41462=>"001110111",
  41463=>"000000000",
  41464=>"010000000",
  41465=>"001001001",
  41466=>"000000111",
  41467=>"001001000",
  41468=>"000000000",
  41469=>"111111101",
  41470=>"000000000",
  41471=>"011111111",
  41472=>"111111001",
  41473=>"111110110",
  41474=>"001100100",
  41475=>"010010110",
  41476=>"011000001",
  41477=>"000001011",
  41478=>"010110110",
  41479=>"001000111",
  41480=>"000000000",
  41481=>"011001000",
  41482=>"111001001",
  41483=>"110000001",
  41484=>"111111011",
  41485=>"000000000",
  41486=>"000101111",
  41487=>"111110001",
  41488=>"111111100",
  41489=>"111011001",
  41490=>"000000111",
  41491=>"111101111",
  41492=>"110000000",
  41493=>"000000011",
  41494=>"001000000",
  41495=>"011001001",
  41496=>"110110100",
  41497=>"001011111",
  41498=>"111011011",
  41499=>"100000000",
  41500=>"111000000",
  41501=>"110000110",
  41502=>"001001011",
  41503=>"000000000",
  41504=>"010111010",
  41505=>"000001001",
  41506=>"000000000",
  41507=>"000000000",
  41508=>"000001001",
  41509=>"011011001",
  41510=>"000000111",
  41511=>"000000000",
  41512=>"111111000",
  41513=>"111011011",
  41514=>"001000000",
  41515=>"000001111",
  41516=>"001000000",
  41517=>"011111111",
  41518=>"011000000",
  41519=>"111111011",
  41520=>"001001001",
  41521=>"111111111",
  41522=>"111011111",
  41523=>"111111010",
  41524=>"111111111",
  41525=>"110110110",
  41526=>"110010001",
  41527=>"000000000",
  41528=>"100001111",
  41529=>"111111111",
  41530=>"110111111",
  41531=>"011000101",
  41532=>"111111111",
  41533=>"111000000",
  41534=>"110111010",
  41535=>"011111111",
  41536=>"111101111",
  41537=>"101101001",
  41538=>"111111111",
  41539=>"110010000",
  41540=>"000000100",
  41541=>"011010100",
  41542=>"111111000",
  41543=>"100100111",
  41544=>"000111011",
  41545=>"000000000",
  41546=>"000000000",
  41547=>"000110111",
  41548=>"110110110",
  41549=>"010000001",
  41550=>"101001000",
  41551=>"000000111",
  41552=>"000000000",
  41553=>"001001111",
  41554=>"100000110",
  41555=>"000000001",
  41556=>"111111111",
  41557=>"000100111",
  41558=>"001011111",
  41559=>"111000000",
  41560=>"001111111",
  41561=>"000000101",
  41562=>"000000000",
  41563=>"111111110",
  41564=>"000000100",
  41565=>"111111111",
  41566=>"000001101",
  41567=>"011011110",
  41568=>"001111111",
  41569=>"000000000",
  41570=>"111110010",
  41571=>"111111111",
  41572=>"000000000",
  41573=>"010110111",
  41574=>"001001000",
  41575=>"000000000",
  41576=>"111111111",
  41577=>"000000011",
  41578=>"000000000",
  41579=>"111111000",
  41580=>"001001000",
  41581=>"100100000",
  41582=>"000000001",
  41583=>"111111111",
  41584=>"101000111",
  41585=>"111101001",
  41586=>"111111011",
  41587=>"000001000",
  41588=>"000101111",
  41589=>"000000011",
  41590=>"111111110",
  41591=>"000101111",
  41592=>"011110110",
  41593=>"111011000",
  41594=>"100000000",
  41595=>"000000000",
  41596=>"001001001",
  41597=>"100110111",
  41598=>"000000110",
  41599=>"011111111",
  41600=>"001000110",
  41601=>"000000000",
  41602=>"111111001",
  41603=>"111111111",
  41604=>"100100110",
  41605=>"000110111",
  41606=>"100110110",
  41607=>"001001000",
  41608=>"000000000",
  41609=>"101101111",
  41610=>"000101111",
  41611=>"000000111",
  41612=>"111111000",
  41613=>"111111111",
  41614=>"111111111",
  41615=>"111101000",
  41616=>"100000000",
  41617=>"111001001",
  41618=>"111111111",
  41619=>"100000000",
  41620=>"000001111",
  41621=>"110010001",
  41622=>"000000001",
  41623=>"011001111",
  41624=>"001000100",
  41625=>"000000011",
  41626=>"111111000",
  41627=>"101101101",
  41628=>"110111111",
  41629=>"010000001",
  41630=>"110000000",
  41631=>"000111111",
  41632=>"011010000",
  41633=>"011111011",
  41634=>"111110111",
  41635=>"011111111",
  41636=>"111001000",
  41637=>"000000000",
  41638=>"001000000",
  41639=>"101000100",
  41640=>"000000110",
  41641=>"001000000",
  41642=>"111111000",
  41643=>"000000000",
  41644=>"000100100",
  41645=>"000001011",
  41646=>"000000111",
  41647=>"000100111",
  41648=>"000010111",
  41649=>"011000100",
  41650=>"011111111",
  41651=>"111111001",
  41652=>"010010111",
  41653=>"000100000",
  41654=>"000000000",
  41655=>"000000000",
  41656=>"111100111",
  41657=>"000111111",
  41658=>"111000000",
  41659=>"100000000",
  41660=>"000000000",
  41661=>"000101110",
  41662=>"000010000",
  41663=>"111111011",
  41664=>"111111111",
  41665=>"111111110",
  41666=>"000000000",
  41667=>"111111111",
  41668=>"000000000",
  41669=>"000000110",
  41670=>"110110000",
  41671=>"010110011",
  41672=>"000000111",
  41673=>"000100101",
  41674=>"001000000",
  41675=>"000111101",
  41676=>"100111100",
  41677=>"000100000",
  41678=>"111000110",
  41679=>"110000000",
  41680=>"000011111",
  41681=>"000000001",
  41682=>"100000111",
  41683=>"000111010",
  41684=>"111111111",
  41685=>"111001000",
  41686=>"001000000",
  41687=>"000001001",
  41688=>"011111111",
  41689=>"101111111",
  41690=>"000000000",
  41691=>"000000000",
  41692=>"110110111",
  41693=>"000000111",
  41694=>"000000111",
  41695=>"000101111",
  41696=>"000000001",
  41697=>"000000111",
  41698=>"001000010",
  41699=>"111000010",
  41700=>"110111111",
  41701=>"111111111",
  41702=>"000010110",
  41703=>"000000000",
  41704=>"111111111",
  41705=>"010010000",
  41706=>"011111111",
  41707=>"000000000",
  41708=>"111110100",
  41709=>"011000000",
  41710=>"111011001",
  41711=>"101000000",
  41712=>"000000000",
  41713=>"010000100",
  41714=>"101100100",
  41715=>"001101101",
  41716=>"111111111",
  41717=>"111101001",
  41718=>"111101111",
  41719=>"111111111",
  41720=>"000000000",
  41721=>"111111111",
  41722=>"000000001",
  41723=>"111111111",
  41724=>"000000000",
  41725=>"001000001",
  41726=>"000000000",
  41727=>"100111111",
  41728=>"100111111",
  41729=>"111111001",
  41730=>"111111111",
  41731=>"001000000",
  41732=>"000000111",
  41733=>"000111111",
  41734=>"011111100",
  41735=>"110111111",
  41736=>"100111111",
  41737=>"101101111",
  41738=>"111111000",
  41739=>"000000000",
  41740=>"000000111",
  41741=>"011001011",
  41742=>"111111001",
  41743=>"111000000",
  41744=>"111110000",
  41745=>"001000000",
  41746=>"000000000",
  41747=>"111100101",
  41748=>"000000100",
  41749=>"111000000",
  41750=>"111111111",
  41751=>"100110111",
  41752=>"111111111",
  41753=>"000000000",
  41754=>"011001001",
  41755=>"000010010",
  41756=>"000000000",
  41757=>"000000010",
  41758=>"010000000",
  41759=>"100000000",
  41760=>"000000000",
  41761=>"000000111",
  41762=>"011010000",
  41763=>"001001111",
  41764=>"000000000",
  41765=>"000000100",
  41766=>"011011001",
  41767=>"110000110",
  41768=>"000000000",
  41769=>"111111110",
  41770=>"000110000",
  41771=>"000110010",
  41772=>"100011111",
  41773=>"110100100",
  41774=>"111111000",
  41775=>"000000010",
  41776=>"000000000",
  41777=>"000011011",
  41778=>"011111110",
  41779=>"111011000",
  41780=>"000000000",
  41781=>"111111110",
  41782=>"111000110",
  41783=>"000111111",
  41784=>"000000010",
  41785=>"000111111",
  41786=>"110111101",
  41787=>"111010110",
  41788=>"110000000",
  41789=>"000000010",
  41790=>"111000000",
  41791=>"000110111",
  41792=>"111000110",
  41793=>"111111111",
  41794=>"111111111",
  41795=>"100110001",
  41796=>"000000111",
  41797=>"101111101",
  41798=>"000000000",
  41799=>"001001000",
  41800=>"000000001",
  41801=>"001000000",
  41802=>"001000000",
  41803=>"111110000",
  41804=>"000000000",
  41805=>"000000000",
  41806=>"010111000",
  41807=>"000000110",
  41808=>"000000110",
  41809=>"000000000",
  41810=>"111000000",
  41811=>"010010110",
  41812=>"111111011",
  41813=>"000000000",
  41814=>"111111000",
  41815=>"111101001",
  41816=>"111111111",
  41817=>"000001000",
  41818=>"101100110",
  41819=>"000000101",
  41820=>"011000000",
  41821=>"000001001",
  41822=>"111111111",
  41823=>"111110110",
  41824=>"000110111",
  41825=>"100000000",
  41826=>"111111100",
  41827=>"010111111",
  41828=>"001100111",
  41829=>"111111111",
  41830=>"000000000",
  41831=>"111111111",
  41832=>"001110111",
  41833=>"001000000",
  41834=>"011011111",
  41835=>"111111100",
  41836=>"110110000",
  41837=>"111111101",
  41838=>"000000100",
  41839=>"001101101",
  41840=>"111111111",
  41841=>"111111101",
  41842=>"111111110",
  41843=>"101111111",
  41844=>"111111111",
  41845=>"111111111",
  41846=>"000000000",
  41847=>"100111110",
  41848=>"010000000",
  41849=>"000000000",
  41850=>"111111111",
  41851=>"000110111",
  41852=>"101100000",
  41853=>"111111111",
  41854=>"000000111",
  41855=>"000000100",
  41856=>"111111110",
  41857=>"000111100",
  41858=>"110010011",
  41859=>"111111001",
  41860=>"000000000",
  41861=>"010000100",
  41862=>"001101001",
  41863=>"111001001",
  41864=>"111111000",
  41865=>"000000011",
  41866=>"000010000",
  41867=>"000000001",
  41868=>"001000101",
  41869=>"000000110",
  41870=>"111111111",
  41871=>"111111011",
  41872=>"111101101",
  41873=>"000111111",
  41874=>"000000000",
  41875=>"111011111",
  41876=>"111111011",
  41877=>"000000000",
  41878=>"111010000",
  41879=>"111111100",
  41880=>"111111111",
  41881=>"111100001",
  41882=>"010000000",
  41883=>"111110000",
  41884=>"000011000",
  41885=>"011010000",
  41886=>"000000111",
  41887=>"000000000",
  41888=>"000000000",
  41889=>"000000001",
  41890=>"011100101",
  41891=>"011011111",
  41892=>"111111111",
  41893=>"011011000",
  41894=>"101111001",
  41895=>"001001000",
  41896=>"111001000",
  41897=>"111011011",
  41898=>"111111010",
  41899=>"001000011",
  41900=>"111101001",
  41901=>"010001000",
  41902=>"000000000",
  41903=>"000000010",
  41904=>"100101111",
  41905=>"001011111",
  41906=>"111111111",
  41907=>"000000000",
  41908=>"111111111",
  41909=>"000000000",
  41910=>"100000001",
  41911=>"000011111",
  41912=>"001101111",
  41913=>"111111111",
  41914=>"111111010",
  41915=>"011011111",
  41916=>"111111111",
  41917=>"000000010",
  41918=>"000000000",
  41919=>"111111001",
  41920=>"111111001",
  41921=>"111111111",
  41922=>"111001111",
  41923=>"011001000",
  41924=>"111110101",
  41925=>"000110110",
  41926=>"110000000",
  41927=>"001001111",
  41928=>"000101111",
  41929=>"000001011",
  41930=>"000000011",
  41931=>"000010000",
  41932=>"001001000",
  41933=>"010000000",
  41934=>"011011111",
  41935=>"111110000",
  41936=>"111100100",
  41937=>"111111111",
  41938=>"010011000",
  41939=>"000000011",
  41940=>"111111011",
  41941=>"111111111",
  41942=>"000000010",
  41943=>"011011011",
  41944=>"000000000",
  41945=>"000000111",
  41946=>"000000000",
  41947=>"111111111",
  41948=>"110000000",
  41949=>"000100101",
  41950=>"111011001",
  41951=>"100011011",
  41952=>"111111111",
  41953=>"111000000",
  41954=>"111111111",
  41955=>"111111111",
  41956=>"111111111",
  41957=>"000010000",
  41958=>"000000001",
  41959=>"111110000",
  41960=>"111101101",
  41961=>"111000000",
  41962=>"000011010",
  41963=>"000000001",
  41964=>"101000111",
  41965=>"111110000",
  41966=>"111111111",
  41967=>"000000100",
  41968=>"111000000",
  41969=>"111011011",
  41970=>"001000001",
  41971=>"010000000",
  41972=>"000011111",
  41973=>"111000001",
  41974=>"111111100",
  41975=>"011111101",
  41976=>"000100111",
  41977=>"011000010",
  41978=>"110111110",
  41979=>"000000111",
  41980=>"100111111",
  41981=>"000000000",
  41982=>"100111111",
  41983=>"000000000",
  41984=>"000000100",
  41985=>"000110111",
  41986=>"000010000",
  41987=>"100100101",
  41988=>"111001001",
  41989=>"110000000",
  41990=>"111110110",
  41991=>"011111011",
  41992=>"000000000",
  41993=>"000001000",
  41994=>"111111001",
  41995=>"101111000",
  41996=>"000000111",
  41997=>"111111110",
  41998=>"000000111",
  41999=>"110000000",
  42000=>"100100100",
  42001=>"110110100",
  42002=>"101000011",
  42003=>"000001111",
  42004=>"000000100",
  42005=>"001001111",
  42006=>"100111111",
  42007=>"001000000",
  42008=>"111100100",
  42009=>"000100100",
  42010=>"001001101",
  42011=>"011011100",
  42012=>"000001100",
  42013=>"100100101",
  42014=>"001001011",
  42015=>"001000000",
  42016=>"111111111",
  42017=>"111111111",
  42018=>"111111001",
  42019=>"001000001",
  42020=>"001000000",
  42021=>"101000101",
  42022=>"101001000",
  42023=>"000000001",
  42024=>"111111111",
  42025=>"100111001",
  42026=>"110100000",
  42027=>"000000000",
  42028=>"000000011",
  42029=>"000111000",
  42030=>"000000101",
  42031=>"110000011",
  42032=>"101100000",
  42033=>"110111111",
  42034=>"000000011",
  42035=>"000000001",
  42036=>"000000000",
  42037=>"001000111",
  42038=>"101000000",
  42039=>"111011111",
  42040=>"000000111",
  42041=>"000101001",
  42042=>"111111111",
  42043=>"111111111",
  42044=>"100100110",
  42045=>"111111001",
  42046=>"111111001",
  42047=>"000101111",
  42048=>"000001011",
  42049=>"000100000",
  42050=>"011011000",
  42051=>"000111001",
  42052=>"001001101",
  42053=>"111111111",
  42054=>"000010000",
  42055=>"000000000",
  42056=>"011011011",
  42057=>"011001111",
  42058=>"111011001",
  42059=>"000000001",
  42060=>"000100101",
  42061=>"100100000",
  42062=>"000000000",
  42063=>"001001111",
  42064=>"101001000",
  42065=>"000000000",
  42066=>"000000011",
  42067=>"110111001",
  42068=>"100100000",
  42069=>"001111111",
  42070=>"000001001",
  42071=>"110010000",
  42072=>"100111000",
  42073=>"000000111",
  42074=>"111101111",
  42075=>"110100100",
  42076=>"111001111",
  42077=>"000000111",
  42078=>"100100111",
  42079=>"011001000",
  42080=>"010110010",
  42081=>"110111001",
  42082=>"111111111",
  42083=>"000110110",
  42084=>"000000111",
  42085=>"000000101",
  42086=>"110110100",
  42087=>"100100100",
  42088=>"111011000",
  42089=>"000000010",
  42090=>"011111111",
  42091=>"000110000",
  42092=>"000111111",
  42093=>"100111111",
  42094=>"001000100",
  42095=>"000100100",
  42096=>"000100100",
  42097=>"000110111",
  42098=>"010110000",
  42099=>"000000111",
  42100=>"000000000",
  42101=>"001101111",
  42102=>"111111110",
  42103=>"101100111",
  42104=>"000000111",
  42105=>"000000111",
  42106=>"000000000",
  42107=>"000000000",
  42108=>"000010110",
  42109=>"111111111",
  42110=>"111011000",
  42111=>"000000000",
  42112=>"001001111",
  42113=>"110100111",
  42114=>"110111110",
  42115=>"011011000",
  42116=>"110110000",
  42117=>"000000111",
  42118=>"000000011",
  42119=>"000000000",
  42120=>"111111010",
  42121=>"000001111",
  42122=>"111010001",
  42123=>"011011001",
  42124=>"000000000",
  42125=>"000011111",
  42126=>"111111000",
  42127=>"111111111",
  42128=>"000000000",
  42129=>"000000000",
  42130=>"000001000",
  42131=>"011011000",
  42132=>"001101110",
  42133=>"100100110",
  42134=>"111111111",
  42135=>"001001111",
  42136=>"000000101",
  42137=>"111101101",
  42138=>"111000000",
  42139=>"000100110",
  42140=>"111111100",
  42141=>"000001001",
  42142=>"110111011",
  42143=>"110111110",
  42144=>"100000000",
  42145=>"111111111",
  42146=>"111111010",
  42147=>"111111111",
  42148=>"000000000",
  42149=>"100100000",
  42150=>"000000000",
  42151=>"100100101",
  42152=>"011111111",
  42153=>"000000000",
  42154=>"011001000",
  42155=>"001000000",
  42156=>"111111111",
  42157=>"000000000",
  42158=>"000000001",
  42159=>"111111111",
  42160=>"000111111",
  42161=>"000000001",
  42162=>"010011000",
  42163=>"100101111",
  42164=>"111111000",
  42165=>"000111110",
  42166=>"111111111",
  42167=>"111111111",
  42168=>"101000111",
  42169=>"000000000",
  42170=>"000000111",
  42171=>"000000000",
  42172=>"101101111",
  42173=>"110111110",
  42174=>"000010000",
  42175=>"001111101",
  42176=>"110100011",
  42177=>"111111111",
  42178=>"111011111",
  42179=>"000000000",
  42180=>"011110110",
  42181=>"000000000",
  42182=>"000000000",
  42183=>"010010110",
  42184=>"000000000",
  42185=>"000000001",
  42186=>"001000000",
  42187=>"000000010",
  42188=>"110110000",
  42189=>"000000000",
  42190=>"001000111",
  42191=>"111010110",
  42192=>"001000000",
  42193=>"000000000",
  42194=>"100110111",
  42195=>"000000111",
  42196=>"000000000",
  42197=>"111111111",
  42198=>"001000000",
  42199=>"000000001",
  42200=>"111111111",
  42201=>"111111111",
  42202=>"100000000",
  42203=>"110111111",
  42204=>"000001101",
  42205=>"111111110",
  42206=>"111111111",
  42207=>"001000000",
  42208=>"000000000",
  42209=>"000111010",
  42210=>"111110110",
  42211=>"111011111",
  42212=>"001110100",
  42213=>"000000001",
  42214=>"010010000",
  42215=>"111110111",
  42216=>"000101111",
  42217=>"001001000",
  42218=>"000000101",
  42219=>"011000101",
  42220=>"111101111",
  42221=>"001001111",
  42222=>"000111111",
  42223=>"000000000",
  42224=>"000000000",
  42225=>"011011000",
  42226=>"001000000",
  42227=>"000000111",
  42228=>"111111111",
  42229=>"011001111",
  42230=>"111111011",
  42231=>"001001111",
  42232=>"110111110",
  42233=>"001001101",
  42234=>"000010000",
  42235=>"000100111",
  42236=>"001001111",
  42237=>"000000111",
  42238=>"101000000",
  42239=>"100000000",
  42240=>"001000111",
  42241=>"100110001",
  42242=>"111111111",
  42243=>"010111111",
  42244=>"110111110",
  42245=>"000000000",
  42246=>"001001111",
  42247=>"001111101",
  42248=>"001000011",
  42249=>"111111111",
  42250=>"100111110",
  42251=>"100100101",
  42252=>"110000010",
  42253=>"000000000",
  42254=>"111111011",
  42255=>"000100100",
  42256=>"000000000",
  42257=>"001111101",
  42258=>"000000101",
  42259=>"111111111",
  42260=>"001001111",
  42261=>"111111110",
  42262=>"100100100",
  42263=>"000000000",
  42264=>"000000111",
  42265=>"111001111",
  42266=>"111111111",
  42267=>"000000000",
  42268=>"010011001",
  42269=>"110110000",
  42270=>"111000000",
  42271=>"100110110",
  42272=>"111111000",
  42273=>"011011111",
  42274=>"111011000",
  42275=>"000100101",
  42276=>"000000000",
  42277=>"110111111",
  42278=>"000100111",
  42279=>"101111000",
  42280=>"000000100",
  42281=>"100000111",
  42282=>"111111011",
  42283=>"000000000",
  42284=>"111011000",
  42285=>"000001001",
  42286=>"011011000",
  42287=>"111001000",
  42288=>"110111111",
  42289=>"111100000",
  42290=>"000000010",
  42291=>"000000000",
  42292=>"000100000",
  42293=>"000110011",
  42294=>"111000010",
  42295=>"000000001",
  42296=>"010110010",
  42297=>"001011011",
  42298=>"000001111",
  42299=>"111111111",
  42300=>"100100000",
  42301=>"111111111",
  42302=>"111000000",
  42303=>"111101000",
  42304=>"000111111",
  42305=>"100111000",
  42306=>"000000101",
  42307=>"001001111",
  42308=>"111111011",
  42309=>"110100110",
  42310=>"111111000",
  42311=>"000110010",
  42312=>"000000000",
  42313=>"000000000",
  42314=>"011111111",
  42315=>"011111111",
  42316=>"011100100",
  42317=>"111111011",
  42318=>"000100001",
  42319=>"011011111",
  42320=>"000000110",
  42321=>"001111111",
  42322=>"000010111",
  42323=>"001000001",
  42324=>"110011010",
  42325=>"011111001",
  42326=>"001000000",
  42327=>"100110111",
  42328=>"001000001",
  42329=>"000010000",
  42330=>"000100100",
  42331=>"000000101",
  42332=>"000000000",
  42333=>"001000100",
  42334=>"000000101",
  42335=>"000000000",
  42336=>"111111100",
  42337=>"000001111",
  42338=>"011011000",
  42339=>"000111111",
  42340=>"001000010",
  42341=>"000000000",
  42342=>"000111111",
  42343=>"100000010",
  42344=>"111110110",
  42345=>"000111111",
  42346=>"000000011",
  42347=>"000000000",
  42348=>"111110100",
  42349=>"000000110",
  42350=>"111100110",
  42351=>"000001001",
  42352=>"111000000",
  42353=>"011000000",
  42354=>"111111111",
  42355=>"101111101",
  42356=>"110000110",
  42357=>"000000111",
  42358=>"000000000",
  42359=>"111111110",
  42360=>"000011111",
  42361=>"000000101",
  42362=>"001000111",
  42363=>"111111111",
  42364=>"011111100",
  42365=>"110111111",
  42366=>"001000000",
  42367=>"001000010",
  42368=>"110110110",
  42369=>"111111000",
  42370=>"111111111",
  42371=>"000111111",
  42372=>"001000111",
  42373=>"111111001",
  42374=>"010111101",
  42375=>"101100000",
  42376=>"001111111",
  42377=>"111111111",
  42378=>"000000000",
  42379=>"010111111",
  42380=>"001011011",
  42381=>"110111111",
  42382=>"000000001",
  42383=>"000000110",
  42384=>"000000000",
  42385=>"001001001",
  42386=>"111111000",
  42387=>"001000000",
  42388=>"111111111",
  42389=>"110110110",
  42390=>"111101000",
  42391=>"000000000",
  42392=>"111000000",
  42393=>"011111111",
  42394=>"001100111",
  42395=>"111111000",
  42396=>"001001101",
  42397=>"000111000",
  42398=>"001101011",
  42399=>"000000000",
  42400=>"111000100",
  42401=>"110000011",
  42402=>"100000000",
  42403=>"001001001",
  42404=>"111111110",
  42405=>"110110010",
  42406=>"100100000",
  42407=>"100111111",
  42408=>"011000010",
  42409=>"000000001",
  42410=>"110111111",
  42411=>"000010111",
  42412=>"000000000",
  42413=>"101101111",
  42414=>"111111111",
  42415=>"000110111",
  42416=>"011111011",
  42417=>"111111100",
  42418=>"111111111",
  42419=>"000000000",
  42420=>"000000000",
  42421=>"110110011",
  42422=>"000000101",
  42423=>"001101111",
  42424=>"000000000",
  42425=>"000001100",
  42426=>"000000101",
  42427=>"111111111",
  42428=>"000000000",
  42429=>"111001000",
  42430=>"111001001",
  42431=>"001001001",
  42432=>"000000111",
  42433=>"000000000",
  42434=>"000010000",
  42435=>"000000000",
  42436=>"001000011",
  42437=>"001011011",
  42438=>"011111111",
  42439=>"111111000",
  42440=>"000000000",
  42441=>"000000000",
  42442=>"001001001",
  42443=>"111111111",
  42444=>"010010000",
  42445=>"000000100",
  42446=>"110110100",
  42447=>"000010110",
  42448=>"011001000",
  42449=>"000100101",
  42450=>"000001111",
  42451=>"010000111",
  42452=>"100111111",
  42453=>"000000000",
  42454=>"001011011",
  42455=>"110100100",
  42456=>"000101111",
  42457=>"000000100",
  42458=>"000101100",
  42459=>"111011000",
  42460=>"111001001",
  42461=>"111111010",
  42462=>"011110100",
  42463=>"100100001",
  42464=>"000000000",
  42465=>"111111111",
  42466=>"000000000",
  42467=>"110111011",
  42468=>"011000000",
  42469=>"000000000",
  42470=>"111111111",
  42471=>"011000000",
  42472=>"100111000",
  42473=>"111111111",
  42474=>"001111111",
  42475=>"000011111",
  42476=>"101101111",
  42477=>"010000000",
  42478=>"000000011",
  42479=>"000000000",
  42480=>"001011111",
  42481=>"000000001",
  42482=>"000000101",
  42483=>"011111000",
  42484=>"000000111",
  42485=>"000000000",
  42486=>"011111111",
  42487=>"000011011",
  42488=>"000001011",
  42489=>"000001001",
  42490=>"001000000",
  42491=>"001000000",
  42492=>"000001111",
  42493=>"001001001",
  42494=>"000000111",
  42495=>"000111111",
  42496=>"000000000",
  42497=>"100000000",
  42498=>"000000000",
  42499=>"111111111",
  42500=>"111111111",
  42501=>"100000000",
  42502=>"010010111",
  42503=>"000100101",
  42504=>"111111100",
  42505=>"000000111",
  42506=>"000000010",
  42507=>"111111001",
  42508=>"010110110",
  42509=>"001011100",
  42510=>"111111011",
  42511=>"000011000",
  42512=>"110111111",
  42513=>"111000000",
  42514=>"111000000",
  42515=>"000000000",
  42516=>"110111111",
  42517=>"111111111",
  42518=>"010100111",
  42519=>"100100000",
  42520=>"000101001",
  42521=>"100111111",
  42522=>"111111101",
  42523=>"000011000",
  42524=>"001001001",
  42525=>"110111111",
  42526=>"011011011",
  42527=>"110100111",
  42528=>"011111000",
  42529=>"000000111",
  42530=>"000000000",
  42531=>"001111111",
  42532=>"111000101",
  42533=>"001000000",
  42534=>"011001111",
  42535=>"100100000",
  42536=>"111001001",
  42537=>"001001111",
  42538=>"111111111",
  42539=>"000001000",
  42540=>"110100100",
  42541=>"011001000",
  42542=>"111100100",
  42543=>"000000000",
  42544=>"000011011",
  42545=>"011010110",
  42546=>"111111111",
  42547=>"100110000",
  42548=>"111010000",
  42549=>"110000111",
  42550=>"000011111",
  42551=>"110110111",
  42552=>"110101000",
  42553=>"000000000",
  42554=>"000000100",
  42555=>"000000000",
  42556=>"111111111",
  42557=>"000011111",
  42558=>"110110100",
  42559=>"000000000",
  42560=>"100011111",
  42561=>"001001000",
  42562=>"011010010",
  42563=>"000110110",
  42564=>"000110000",
  42565=>"011011011",
  42566=>"000011000",
  42567=>"000000000",
  42568=>"100110111",
  42569=>"000000000",
  42570=>"010011001",
  42571=>"000100101",
  42572=>"000000000",
  42573=>"111010000",
  42574=>"011000000",
  42575=>"000111111",
  42576=>"000111110",
  42577=>"001111101",
  42578=>"000110110",
  42579=>"000000000",
  42580=>"000000000",
  42581=>"011000010",
  42582=>"000111101",
  42583=>"000000000",
  42584=>"010010001",
  42585=>"000000100",
  42586=>"000111000",
  42587=>"111111100",
  42588=>"111111111",
  42589=>"111101100",
  42590=>"100101101",
  42591=>"000101000",
  42592=>"001111111",
  42593=>"010111111",
  42594=>"010110110",
  42595=>"001000000",
  42596=>"111101000",
  42597=>"000000100",
  42598=>"110000000",
  42599=>"111100001",
  42600=>"000000000",
  42601=>"000000001",
  42602=>"000000001",
  42603=>"010010000",
  42604=>"011111111",
  42605=>"000000000",
  42606=>"111111111",
  42607=>"001100111",
  42608=>"001100100",
  42609=>"100110000",
  42610=>"001000001",
  42611=>"100100101",
  42612=>"000000000",
  42613=>"000000000",
  42614=>"000000000",
  42615=>"000000110",
  42616=>"111011000",
  42617=>"000001001",
  42618=>"111001111",
  42619=>"000111100",
  42620=>"011011011",
  42621=>"000010110",
  42622=>"111111111",
  42623=>"011000000",
  42624=>"111100111",
  42625=>"000111101",
  42626=>"100100000",
  42627=>"000111111",
  42628=>"111111111",
  42629=>"001001000",
  42630=>"111111111",
  42631=>"100000000",
  42632=>"110110000",
  42633=>"111111000",
  42634=>"000000000",
  42635=>"001001100",
  42636=>"011010000",
  42637=>"000110100",
  42638=>"100000000",
  42639=>"000000000",
  42640=>"111110111",
  42641=>"111111000",
  42642=>"100111100",
  42643=>"111000000",
  42644=>"001011011",
  42645=>"111110100",
  42646=>"111111000",
  42647=>"000111111",
  42648=>"000111000",
  42649=>"111111110",
  42650=>"000001011",
  42651=>"111111000",
  42652=>"000111101",
  42653=>"110110010",
  42654=>"000011000",
  42655=>"000000000",
  42656=>"000001011",
  42657=>"000000000",
  42658=>"111000000",
  42659=>"111101101",
  42660=>"011011111",
  42661=>"000011001",
  42662=>"011001000",
  42663=>"001000111",
  42664=>"000011100",
  42665=>"000000000",
  42666=>"000000000",
  42667=>"000110111",
  42668=>"000011111",
  42669=>"001001001",
  42670=>"010000000",
  42671=>"111111111",
  42672=>"000000000",
  42673=>"000000000",
  42674=>"111111111",
  42675=>"000000000",
  42676=>"111011011",
  42677=>"000010110",
  42678=>"111110000",
  42679=>"000000000",
  42680=>"110111111",
  42681=>"111111111",
  42682=>"111001111",
  42683=>"010110000",
  42684=>"111011000",
  42685=>"111100000",
  42686=>"001111000",
  42687=>"111011011",
  42688=>"111111110",
  42689=>"010000100",
  42690=>"011111001",
  42691=>"000000000",
  42692=>"111111111",
  42693=>"000000000",
  42694=>"100000111",
  42695=>"000101101",
  42696=>"110100000",
  42697=>"100110100",
  42698=>"001000100",
  42699=>"111000010",
  42700=>"000010100",
  42701=>"110000110",
  42702=>"000011000",
  42703=>"011000111",
  42704=>"100000000",
  42705=>"111111001",
  42706=>"110000000",
  42707=>"111111111",
  42708=>"100000111",
  42709=>"000100100",
  42710=>"001000000",
  42711=>"000000001",
  42712=>"000000000",
  42713=>"010111000",
  42714=>"111111110",
  42715=>"111111111",
  42716=>"000111110",
  42717=>"110111111",
  42718=>"000000000",
  42719=>"000111111",
  42720=>"000000000",
  42721=>"000001000",
  42722=>"111000000",
  42723=>"110111100",
  42724=>"111001011",
  42725=>"111111001",
  42726=>"000001000",
  42727=>"111111100",
  42728=>"000000000",
  42729=>"111000000",
  42730=>"111111111",
  42731=>"000000001",
  42732=>"010110011",
  42733=>"111111111",
  42734=>"111000000",
  42735=>"011011000",
  42736=>"111111111",
  42737=>"001101100",
  42738=>"000000000",
  42739=>"000000000",
  42740=>"000000111",
  42741=>"100111100",
  42742=>"111111100",
  42743=>"010011100",
  42744=>"000000000",
  42745=>"111111111",
  42746=>"000111001",
  42747=>"111111111",
  42748=>"101001111",
  42749=>"000101111",
  42750=>"010110111",
  42751=>"110101100",
  42752=>"000000000",
  42753=>"111111111",
  42754=>"111001001",
  42755=>"000101000",
  42756=>"000110110",
  42757=>"000001001",
  42758=>"000000001",
  42759=>"000000111",
  42760=>"100111111",
  42761=>"111101101",
  42762=>"000110000",
  42763=>"001111110",
  42764=>"111111111",
  42765=>"001111110",
  42766=>"011101101",
  42767=>"000000000",
  42768=>"110111111",
  42769=>"111110111",
  42770=>"111110000",
  42771=>"111111111",
  42772=>"111111000",
  42773=>"010111111",
  42774=>"011011001",
  42775=>"111111111",
  42776=>"010010111",
  42777=>"101100100",
  42778=>"000000000",
  42779=>"000000000",
  42780=>"101111111",
  42781=>"111111100",
  42782=>"000000000",
  42783=>"101111000",
  42784=>"111111111",
  42785=>"100111111",
  42786=>"000000000",
  42787=>"000000000",
  42788=>"111111100",
  42789=>"111100011",
  42790=>"001011011",
  42791=>"000001101",
  42792=>"111100101",
  42793=>"111111111",
  42794=>"000001000",
  42795=>"000000000",
  42796=>"011111111",
  42797=>"111000101",
  42798=>"000000000",
  42799=>"011111111",
  42800=>"000001001",
  42801=>"000000111",
  42802=>"000011111",
  42803=>"001111001",
  42804=>"000000000",
  42805=>"111111000",
  42806=>"000100100",
  42807=>"111111111",
  42808=>"110111111",
  42809=>"111111000",
  42810=>"111110110",
  42811=>"000000000",
  42812=>"000000011",
  42813=>"000000001",
  42814=>"111111111",
  42815=>"011111011",
  42816=>"000000101",
  42817=>"000110111",
  42818=>"110111111",
  42819=>"111100100",
  42820=>"111111111",
  42821=>"000111110",
  42822=>"001000000",
  42823=>"111000000",
  42824=>"000000001",
  42825=>"111000000",
  42826=>"000000000",
  42827=>"100000001",
  42828=>"111111100",
  42829=>"111011111",
  42830=>"000111100",
  42831=>"001001101",
  42832=>"110110110",
  42833=>"111111110",
  42834=>"000000011",
  42835=>"000000010",
  42836=>"111111111",
  42837=>"111000111",
  42838=>"111111111",
  42839=>"010011000",
  42840=>"000010110",
  42841=>"111100000",
  42842=>"101111111",
  42843=>"000110110",
  42844=>"000000110",
  42845=>"111111100",
  42846=>"111111000",
  42847=>"110111111",
  42848=>"100101001",
  42849=>"000000000",
  42850=>"110111101",
  42851=>"000000000",
  42852=>"010111111",
  42853=>"000000000",
  42854=>"100111000",
  42855=>"111111000",
  42856=>"000011111",
  42857=>"101111100",
  42858=>"111000000",
  42859=>"111110110",
  42860=>"010110111",
  42861=>"000000110",
  42862=>"011000100",
  42863=>"101111001",
  42864=>"111111101",
  42865=>"111111111",
  42866=>"000100000",
  42867=>"111111111",
  42868=>"000010010",
  42869=>"011001000",
  42870=>"000110000",
  42871=>"111101111",
  42872=>"000000000",
  42873=>"101110000",
  42874=>"111000000",
  42875=>"110111111",
  42876=>"001001000",
  42877=>"000111111",
  42878=>"000111000",
  42879=>"111000000",
  42880=>"110110010",
  42881=>"111111001",
  42882=>"110100101",
  42883=>"000001000",
  42884=>"111111111",
  42885=>"101101101",
  42886=>"000100001",
  42887=>"010111110",
  42888=>"111011111",
  42889=>"000000111",
  42890=>"101111111",
  42891=>"000000000",
  42892=>"111111101",
  42893=>"100000111",
  42894=>"000000100",
  42895=>"011111011",
  42896=>"101011001",
  42897=>"100111000",
  42898=>"111111100",
  42899=>"110100000",
  42900=>"111111111",
  42901=>"001000000",
  42902=>"010000000",
  42903=>"100111111",
  42904=>"111111100",
  42905=>"011010010",
  42906=>"000000000",
  42907=>"000000101",
  42908=>"000000101",
  42909=>"000000000",
  42910=>"111110111",
  42911=>"111111011",
  42912=>"111111111",
  42913=>"111110101",
  42914=>"000110111",
  42915=>"100111111",
  42916=>"000001100",
  42917=>"000000000",
  42918=>"000000100",
  42919=>"111110000",
  42920=>"000100000",
  42921=>"011111111",
  42922=>"000000000",
  42923=>"111011111",
  42924=>"001000001",
  42925=>"000100000",
  42926=>"000111111",
  42927=>"111111111",
  42928=>"000000111",
  42929=>"111001111",
  42930=>"000000000",
  42931=>"000110110",
  42932=>"111110110",
  42933=>"111111111",
  42934=>"111111111",
  42935=>"000000011",
  42936=>"000111111",
  42937=>"000000000",
  42938=>"100100100",
  42939=>"000111110",
  42940=>"000010111",
  42941=>"000111000",
  42942=>"111010000",
  42943=>"001001000",
  42944=>"000000000",
  42945=>"010000000",
  42946=>"000000000",
  42947=>"001000000",
  42948=>"000110000",
  42949=>"001001001",
  42950=>"000111111",
  42951=>"001000001",
  42952=>"000110111",
  42953=>"000000100",
  42954=>"000001000",
  42955=>"000000111",
  42956=>"000000111",
  42957=>"111111100",
  42958=>"000101000",
  42959=>"111111111",
  42960=>"100100100",
  42961=>"011111110",
  42962=>"000000000",
  42963=>"000000101",
  42964=>"111011001",
  42965=>"000111011",
  42966=>"111111111",
  42967=>"000000000",
  42968=>"000110111",
  42969=>"000000010",
  42970=>"000000000",
  42971=>"111111111",
  42972=>"111011111",
  42973=>"000010000",
  42974=>"100100000",
  42975=>"111001011",
  42976=>"011111111",
  42977=>"111100101",
  42978=>"010000000",
  42979=>"000010110",
  42980=>"000000000",
  42981=>"000000000",
  42982=>"001110110",
  42983=>"000100110",
  42984=>"111111000",
  42985=>"100000000",
  42986=>"000000111",
  42987=>"000000001",
  42988=>"110110000",
  42989=>"000100000",
  42990=>"111111111",
  42991=>"111111000",
  42992=>"111111111",
  42993=>"000000000",
  42994=>"000010111",
  42995=>"100110001",
  42996=>"000000100",
  42997=>"001111111",
  42998=>"111111100",
  42999=>"111111000",
  43000=>"101000011",
  43001=>"110100101",
  43002=>"000000000",
  43003=>"001000100",
  43004=>"000011111",
  43005=>"000001001",
  43006=>"111111111",
  43007=>"111110111",
  43008=>"111111001",
  43009=>"110111111",
  43010=>"111000000",
  43011=>"111111001",
  43012=>"000000000",
  43013=>"000000011",
  43014=>"110000000",
  43015=>"000001111",
  43016=>"000001011",
  43017=>"000000000",
  43018=>"000000100",
  43019=>"111001101",
  43020=>"111011111",
  43021=>"111111111",
  43022=>"100100100",
  43023=>"111111111",
  43024=>"110110111",
  43025=>"111111100",
  43026=>"111011011",
  43027=>"000000000",
  43028=>"111001001",
  43029=>"000000001",
  43030=>"000000000",
  43031=>"001101110",
  43032=>"001001001",
  43033=>"101001001",
  43034=>"001000000",
  43035=>"011010110",
  43036=>"111001000",
  43037=>"000000001",
  43038=>"011011111",
  43039=>"100000111",
  43040=>"111111111",
  43041=>"111000100",
  43042=>"100111111",
  43043=>"111111111",
  43044=>"110111000",
  43045=>"110110000",
  43046=>"011000000",
  43047=>"001001000",
  43048=>"000010001",
  43049=>"011111011",
  43050=>"101000000",
  43051=>"000000101",
  43052=>"000000000",
  43053=>"011111111",
  43054=>"111000101",
  43055=>"100000000",
  43056=>"000000000",
  43057=>"111011000",
  43058=>"111110000",
  43059=>"000000000",
  43060=>"001111111",
  43061=>"011011011",
  43062=>"000011011",
  43063=>"111111111",
  43064=>"000000011",
  43065=>"000101111",
  43066=>"111111111",
  43067=>"111111111",
  43068=>"000001001",
  43069=>"000000011",
  43070=>"000110111",
  43071=>"000000000",
  43072=>"000001011",
  43073=>"011011011",
  43074=>"010000001",
  43075=>"000000011",
  43076=>"100100101",
  43077=>"111100100",
  43078=>"011001000",
  43079=>"000001000",
  43080=>"100100100",
  43081=>"000000101",
  43082=>"000000111",
  43083=>"000000000",
  43084=>"000000111",
  43085=>"111111111",
  43086=>"001000000",
  43087=>"100111111",
  43088=>"000000000",
  43089=>"001001001",
  43090=>"000001000",
  43091=>"111111011",
  43092=>"111111111",
  43093=>"000110111",
  43094=>"011011011",
  43095=>"000000000",
  43096=>"011000000",
  43097=>"000000000",
  43098=>"000111111",
  43099=>"101001100",
  43100=>"000000000",
  43101=>"101111111",
  43102=>"111011011",
  43103=>"110011111",
  43104=>"111111111",
  43105=>"011010000",
  43106=>"000000111",
  43107=>"101000000",
  43108=>"111111010",
  43109=>"111111100",
  43110=>"000000000",
  43111=>"000000000",
  43112=>"011000000",
  43113=>"111101101",
  43114=>"000000000",
  43115=>"111110110",
  43116=>"000111100",
  43117=>"011111111",
  43118=>"000000111",
  43119=>"000000000",
  43120=>"111111111",
  43121=>"100100000",
  43122=>"001001101",
  43123=>"000111111",
  43124=>"111111111",
  43125=>"100101111",
  43126=>"000000001",
  43127=>"000000000",
  43128=>"000000000",
  43129=>"111111111",
  43130=>"000000000",
  43131=>"111111110",
  43132=>"100111111",
  43133=>"111011000",
  43134=>"000001111",
  43135=>"011011001",
  43136=>"001000000",
  43137=>"000000001",
  43138=>"000010111",
  43139=>"110110100",
  43140=>"100000000",
  43141=>"000000000",
  43142=>"111111011",
  43143=>"111111111",
  43144=>"001000000",
  43145=>"111100000",
  43146=>"000001000",
  43147=>"111111111",
  43148=>"001001101",
  43149=>"100111100",
  43150=>"111111001",
  43151=>"111000011",
  43152=>"000000000",
  43153=>"001001000",
  43154=>"000000000",
  43155=>"111011000",
  43156=>"000000000",
  43157=>"101001111",
  43158=>"000001111",
  43159=>"000000000",
  43160=>"110000011",
  43161=>"111111111",
  43162=>"111111111",
  43163=>"111001101",
  43164=>"111111111",
  43165=>"111111111",
  43166=>"000000100",
  43167=>"000000100",
  43168=>"000000000",
  43169=>"111111111",
  43170=>"001011111",
  43171=>"101111111",
  43172=>"011111101",
  43173=>"111101000",
  43174=>"111111000",
  43175=>"100100110",
  43176=>"110111111",
  43177=>"111111111",
  43178=>"110111111",
  43179=>"111111111",
  43180=>"000000100",
  43181=>"000000000",
  43182=>"111111111",
  43183=>"000101111",
  43184=>"000000000",
  43185=>"100000011",
  43186=>"101111111",
  43187=>"000000000",
  43188=>"111110100",
  43189=>"111111000",
  43190=>"000000110",
  43191=>"111110000",
  43192=>"000011111",
  43193=>"000000011",
  43194=>"001000100",
  43195=>"000001001",
  43196=>"111111100",
  43197=>"000111111",
  43198=>"011001011",
  43199=>"011011011",
  43200=>"011001001",
  43201=>"000000110",
  43202=>"000001011",
  43203=>"011111111",
  43204=>"000100101",
  43205=>"111111000",
  43206=>"111111111",
  43207=>"001000111",
  43208=>"000000000",
  43209=>"001011111",
  43210=>"001001101",
  43211=>"000000000",
  43212=>"001000100",
  43213=>"111111111",
  43214=>"000000000",
  43215=>"000000100",
  43216=>"000000000",
  43217=>"000000000",
  43218=>"101111111",
  43219=>"000010111",
  43220=>"000000000",
  43221=>"110111111",
  43222=>"000111000",
  43223=>"110011010",
  43224=>"000000001",
  43225=>"000000111",
  43226=>"000000000",
  43227=>"000000111",
  43228=>"000000000",
  43229=>"101001000",
  43230=>"111101001",
  43231=>"000000000",
  43232=>"000111111",
  43233=>"111111011",
  43234=>"000000000",
  43235=>"000100010",
  43236=>"110000000",
  43237=>"111000100",
  43238=>"001111000",
  43239=>"100000001",
  43240=>"000111111",
  43241=>"011001111",
  43242=>"011111100",
  43243=>"011111111",
  43244=>"111000000",
  43245=>"000000001",
  43246=>"000111111",
  43247=>"000100000",
  43248=>"111111011",
  43249=>"111111011",
  43250=>"000011111",
  43251=>"001011111",
  43252=>"111111111",
  43253=>"111111111",
  43254=>"000000000",
  43255=>"011001111",
  43256=>"000111111",
  43257=>"000000001",
  43258=>"110111111",
  43259=>"001001000",
  43260=>"000010001",
  43261=>"000111111",
  43262=>"000000000",
  43263=>"011111111",
  43264=>"110111111",
  43265=>"100100101",
  43266=>"000000000",
  43267=>"111111111",
  43268=>"000001111",
  43269=>"000011010",
  43270=>"000101111",
  43271=>"000000111",
  43272=>"010010011",
  43273=>"000000000",
  43274=>"111100101",
  43275=>"111111111",
  43276=>"111111011",
  43277=>"000000000",
  43278=>"110100111",
  43279=>"101111101",
  43280=>"111100111",
  43281=>"110100000",
  43282=>"000000000",
  43283=>"001001000",
  43284=>"000001000",
  43285=>"111111111",
  43286=>"101001001",
  43287=>"111111111",
  43288=>"111011011",
  43289=>"000000010",
  43290=>"111111100",
  43291=>"111111111",
  43292=>"111111111",
  43293=>"000000010",
  43294=>"000000000",
  43295=>"000000111",
  43296=>"001100000",
  43297=>"110000000",
  43298=>"010000000",
  43299=>"000000000",
  43300=>"001011000",
  43301=>"111111111",
  43302=>"100110111",
  43303=>"001000100",
  43304=>"101111111",
  43305=>"111101101",
  43306=>"011111100",
  43307=>"110000000",
  43308=>"101000000",
  43309=>"010000000",
  43310=>"100000000",
  43311=>"110110111",
  43312=>"011000111",
  43313=>"100100000",
  43314=>"011000000",
  43315=>"000000011",
  43316=>"111101000",
  43317=>"000011111",
  43318=>"001001001",
  43319=>"000000101",
  43320=>"000000011",
  43321=>"000000111",
  43322=>"111111100",
  43323=>"000000000",
  43324=>"011111000",
  43325=>"001111111",
  43326=>"010110100",
  43327=>"111110000",
  43328=>"000111000",
  43329=>"111111110",
  43330=>"111111111",
  43331=>"111101111",
  43332=>"001000000",
  43333=>"101000001",
  43334=>"000000000",
  43335=>"101000000",
  43336=>"000000000",
  43337=>"000000000",
  43338=>"000000000",
  43339=>"000000001",
  43340=>"111111111",
  43341=>"000100111",
  43342=>"111111010",
  43343=>"001011111",
  43344=>"011011111",
  43345=>"110111011",
  43346=>"001000001",
  43347=>"011000111",
  43348=>"000111001",
  43349=>"111111111",
  43350=>"000000000",
  43351=>"100111111",
  43352=>"000010111",
  43353=>"000000000",
  43354=>"111111111",
  43355=>"101011011",
  43356=>"000000000",
  43357=>"000000000",
  43358=>"110111011",
  43359=>"101111111",
  43360=>"000000000",
  43361=>"111111111",
  43362=>"001111111",
  43363=>"111111111",
  43364=>"000010011",
  43365=>"111111111",
  43366=>"001000111",
  43367=>"110111111",
  43368=>"001000000",
  43369=>"000000000",
  43370=>"111111111",
  43371=>"101001011",
  43372=>"111111001",
  43373=>"011011111",
  43374=>"000000111",
  43375=>"000000000",
  43376=>"100000000",
  43377=>"000010000",
  43378=>"010000000",
  43379=>"000100100",
  43380=>"110111001",
  43381=>"000000000",
  43382=>"100111001",
  43383=>"111111111",
  43384=>"000111111",
  43385=>"010111111",
  43386=>"000000000",
  43387=>"000101111",
  43388=>"000000110",
  43389=>"111111111",
  43390=>"000000111",
  43391=>"000000111",
  43392=>"110110111",
  43393=>"011011111",
  43394=>"101000001",
  43395=>"111111111",
  43396=>"011101000",
  43397=>"010111111",
  43398=>"101000000",
  43399=>"001110110",
  43400=>"000000000",
  43401=>"000000000",
  43402=>"000001011",
  43403=>"111111111",
  43404=>"000000000",
  43405=>"101101111",
  43406=>"000000101",
  43407=>"000110010",
  43408=>"000001011",
  43409=>"000000111",
  43410=>"000000000",
  43411=>"100111100",
  43412=>"000011111",
  43413=>"010010010",
  43414=>"111001000",
  43415=>"000011011",
  43416=>"111111111",
  43417=>"111001001",
  43418=>"111111111",
  43419=>"111111111",
  43420=>"101100111",
  43421=>"111111011",
  43422=>"111101000",
  43423=>"000000000",
  43424=>"000000000",
  43425=>"110100000",
  43426=>"100000000",
  43427=>"000111000",
  43428=>"110111111",
  43429=>"000011111",
  43430=>"001000000",
  43431=>"011111111",
  43432=>"100110000",
  43433=>"111111110",
  43434=>"000000101",
  43435=>"011001111",
  43436=>"000000000",
  43437=>"000011110",
  43438=>"101111110",
  43439=>"011111111",
  43440=>"111111000",
  43441=>"001000000",
  43442=>"000000000",
  43443=>"000000000",
  43444=>"000000000",
  43445=>"111111111",
  43446=>"000000000",
  43447=>"000000111",
  43448=>"000111111",
  43449=>"000001101",
  43450=>"100100100",
  43451=>"111000000",
  43452=>"000001111",
  43453=>"000110111",
  43454=>"111011011",
  43455=>"101101101",
  43456=>"000011110",
  43457=>"111111111",
  43458=>"000000000",
  43459=>"000000000",
  43460=>"000000100",
  43461=>"111110001",
  43462=>"111111111",
  43463=>"000110111",
  43464=>"000000001",
  43465=>"010110110",
  43466=>"000000011",
  43467=>"011010111",
  43468=>"111111001",
  43469=>"000000101",
  43470=>"111111001",
  43471=>"011111011",
  43472=>"111010000",
  43473=>"111100001",
  43474=>"011100100",
  43475=>"001000001",
  43476=>"001111001",
  43477=>"000000000",
  43478=>"111111010",
  43479=>"000000010",
  43480=>"000001000",
  43481=>"000000000",
  43482=>"111111111",
  43483=>"001101111",
  43484=>"111101111",
  43485=>"111111000",
  43486=>"110000000",
  43487=>"101100101",
  43488=>"101011000",
  43489=>"010000010",
  43490=>"001000000",
  43491=>"111111111",
  43492=>"100001000",
  43493=>"110110110",
  43494=>"011011011",
  43495=>"000000000",
  43496=>"000000001",
  43497=>"111111111",
  43498=>"000011111",
  43499=>"111111110",
  43500=>"111111111",
  43501=>"000100011",
  43502=>"000000000",
  43503=>"000111111",
  43504=>"000000000",
  43505=>"111111111",
  43506=>"111110100",
  43507=>"110010000",
  43508=>"110111111",
  43509=>"100100100",
  43510=>"111111111",
  43511=>"110100000",
  43512=>"111111111",
  43513=>"011011011",
  43514=>"000000001",
  43515=>"111000000",
  43516=>"111011111",
  43517=>"111111111",
  43518=>"101111111",
  43519=>"000000000",
  43520=>"110110110",
  43521=>"000000000",
  43522=>"000000000",
  43523=>"111011111",
  43524=>"011111111",
  43525=>"010000000",
  43526=>"000000000",
  43527=>"000000000",
  43528=>"100000000",
  43529=>"000001011",
  43530=>"011000000",
  43531=>"111111101",
  43532=>"110110110",
  43533=>"100000000",
  43534=>"000100101",
  43535=>"111111111",
  43536=>"000101111",
  43537=>"000111111",
  43538=>"111111111",
  43539=>"001001111",
  43540=>"000000000",
  43541=>"010000111",
  43542=>"111111111",
  43543=>"001110111",
  43544=>"111111110",
  43545=>"100000000",
  43546=>"111101000",
  43547=>"011011111",
  43548=>"011011111",
  43549=>"111111111",
  43550=>"111111111",
  43551=>"000000000",
  43552=>"111000101",
  43553=>"000000111",
  43554=>"111111000",
  43555=>"111111111",
  43556=>"000011101",
  43557=>"000001011",
  43558=>"111111111",
  43559=>"001001000",
  43560=>"111111111",
  43561=>"000100000",
  43562=>"111111000",
  43563=>"000000000",
  43564=>"000000000",
  43565=>"111111110",
  43566=>"111100000",
  43567=>"110111000",
  43568=>"111001010",
  43569=>"000110010",
  43570=>"001000001",
  43571=>"010000100",
  43572=>"110111111",
  43573=>"100110010",
  43574=>"000000001",
  43575=>"100111111",
  43576=>"100000000",
  43577=>"111111111",
  43578=>"000000011",
  43579=>"000000111",
  43580=>"000000001",
  43581=>"010010001",
  43582=>"001111111",
  43583=>"000000001",
  43584=>"010000001",
  43585=>"111110111",
  43586=>"101101000",
  43587=>"000000111",
  43588=>"100100000",
  43589=>"110111010",
  43590=>"111111111",
  43591=>"111111111",
  43592=>"111000111",
  43593=>"001000000",
  43594=>"000100001",
  43595=>"111111111",
  43596=>"000000001",
  43597=>"100001000",
  43598=>"111000000",
  43599=>"111011001",
  43600=>"111111111",
  43601=>"000000111",
  43602=>"110111111",
  43603=>"100100110",
  43604=>"000000000",
  43605=>"000001000",
  43606=>"111111111",
  43607=>"011001011",
  43608=>"000000111",
  43609=>"100100001",
  43610=>"100110111",
  43611=>"011111111",
  43612=>"000111111",
  43613=>"000000000",
  43614=>"111111111",
  43615=>"100000000",
  43616=>"111110110",
  43617=>"110110110",
  43618=>"110111111",
  43619=>"111110010",
  43620=>"011011111",
  43621=>"111011111",
  43622=>"011111001",
  43623=>"000000000",
  43624=>"000000000",
  43625=>"111111111",
  43626=>"111111001",
  43627=>"011110110",
  43628=>"000100100",
  43629=>"000000010",
  43630=>"111000000",
  43631=>"001011011",
  43632=>"110111111",
  43633=>"000101100",
  43634=>"111111111",
  43635=>"000001111",
  43636=>"111111111",
  43637=>"000110111",
  43638=>"000000000",
  43639=>"000111111",
  43640=>"011001000",
  43641=>"000000100",
  43642=>"000110111",
  43643=>"000000000",
  43644=>"100000000",
  43645=>"001000000",
  43646=>"101111111",
  43647=>"110111100",
  43648=>"111111111",
  43649=>"111111111",
  43650=>"111000000",
  43651=>"000100111",
  43652=>"111111100",
  43653=>"000000000",
  43654=>"111111111",
  43655=>"000100110",
  43656=>"111110010",
  43657=>"000000000",
  43658=>"000000010",
  43659=>"000001011",
  43660=>"111111111",
  43661=>"000000000",
  43662=>"111111111",
  43663=>"000000000",
  43664=>"000000000",
  43665=>"000100100",
  43666=>"011000111",
  43667=>"000111011",
  43668=>"000000110",
  43669=>"110110010",
  43670=>"000000000",
  43671=>"001000000",
  43672=>"111111111",
  43673=>"101001011",
  43674=>"011000000",
  43675=>"111001101",
  43676=>"110000000",
  43677=>"000000000",
  43678=>"111001000",
  43679=>"111111111",
  43680=>"111110100",
  43681=>"111000000",
  43682=>"000000000",
  43683=>"000000000",
  43684=>"000111111",
  43685=>"110110111",
  43686=>"111101000",
  43687=>"111100000",
  43688=>"111001111",
  43689=>"101100100",
  43690=>"111111111",
  43691=>"111101111",
  43692=>"000000011",
  43693=>"111110100",
  43694=>"011001111",
  43695=>"000000011",
  43696=>"100000000",
  43697=>"111100100",
  43698=>"111111111",
  43699=>"111111000",
  43700=>"110010000",
  43701=>"000000000",
  43702=>"101111111",
  43703=>"000000100",
  43704=>"100000111",
  43705=>"111111111",
  43706=>"000111111",
  43707=>"110110000",
  43708=>"011000000",
  43709=>"111011011",
  43710=>"111111011",
  43711=>"000000001",
  43712=>"111111111",
  43713=>"000000100",
  43714=>"000000000",
  43715=>"101111111",
  43716=>"100101111",
  43717=>"111110111",
  43718=>"000110111",
  43719=>"111111111",
  43720=>"111111111",
  43721=>"000000000",
  43722=>"111111010",
  43723=>"000100000",
  43724=>"000101111",
  43725=>"100100111",
  43726=>"110110000",
  43727=>"110000100",
  43728=>"000000000",
  43729=>"000111111",
  43730=>"000000000",
  43731=>"000000000",
  43732=>"001000000",
  43733=>"100000110",
  43734=>"000000010",
  43735=>"000000000",
  43736=>"011111111",
  43737=>"000000000",
  43738=>"111111111",
  43739=>"010000111",
  43740=>"111110100",
  43741=>"110000000",
  43742=>"110111111",
  43743=>"111111001",
  43744=>"000000000",
  43745=>"010110110",
  43746=>"110000000",
  43747=>"111111111",
  43748=>"011111111",
  43749=>"111110110",
  43750=>"010000000",
  43751=>"111111111",
  43752=>"000000000",
  43753=>"111111111",
  43754=>"100000000",
  43755=>"110100100",
  43756=>"000000101",
  43757=>"000000000",
  43758=>"110100010",
  43759=>"010000000",
  43760=>"110111111",
  43761=>"111111111",
  43762=>"000000000",
  43763=>"000000110",
  43764=>"111111110",
  43765=>"011000000",
  43766=>"111111111",
  43767=>"000000000",
  43768=>"000111000",
  43769=>"111110110",
  43770=>"000000000",
  43771=>"000000000",
  43772=>"110111011",
  43773=>"011001000",
  43774=>"011000000",
  43775=>"000000001",
  43776=>"010011111",
  43777=>"111100000",
  43778=>"000000000",
  43779=>"000000010",
  43780=>"000000000",
  43781=>"000110000",
  43782=>"111111110",
  43783=>"000000111",
  43784=>"000000000",
  43785=>"111100000",
  43786=>"110000000",
  43787=>"111100100",
  43788=>"011011111",
  43789=>"000000000",
  43790=>"111111111",
  43791=>"000110101",
  43792=>"111011100",
  43793=>"000000000",
  43794=>"001000000",
  43795=>"000001001",
  43796=>"000000000",
  43797=>"010111010",
  43798=>"001000000",
  43799=>"000000000",
  43800=>"000000010",
  43801=>"100000000",
  43802=>"111111111",
  43803=>"111110000",
  43804=>"110110100",
  43805=>"011111110",
  43806=>"000000000",
  43807=>"000001111",
  43808=>"111111001",
  43809=>"100000000",
  43810=>"111110000",
  43811=>"101111111",
  43812=>"111100000",
  43813=>"111111110",
  43814=>"111111111",
  43815=>"000101111",
  43816=>"111111110",
  43817=>"000001001",
  43818=>"000011111",
  43819=>"000000000",
  43820=>"010110000",
  43821=>"000000101",
  43822=>"000000000",
  43823=>"000100111",
  43824=>"110100000",
  43825=>"010010001",
  43826=>"011011000",
  43827=>"000000000",
  43828=>"110000000",
  43829=>"111111101",
  43830=>"010000000",
  43831=>"000000111",
  43832=>"000000000",
  43833=>"000000000",
  43834=>"000000000",
  43835=>"000001000",
  43836=>"111111110",
  43837=>"111001010",
  43838=>"000000000",
  43839=>"110100000",
  43840=>"000000000",
  43841=>"000000000",
  43842=>"111111111",
  43843=>"111011011",
  43844=>"111111111",
  43845=>"000000000",
  43846=>"000000000",
  43847=>"011111000",
  43848=>"000000000",
  43849=>"000000000",
  43850=>"111111110",
  43851=>"000000000",
  43852=>"000001011",
  43853=>"111011000",
  43854=>"111100111",
  43855=>"111111111",
  43856=>"110100100",
  43857=>"101101000",
  43858=>"110110000",
  43859=>"111110100",
  43860=>"111111000",
  43861=>"000010001",
  43862=>"111000011",
  43863=>"100111111",
  43864=>"111011000",
  43865=>"100000000",
  43866=>"111111111",
  43867=>"001000111",
  43868=>"000111100",
  43869=>"000000101",
  43870=>"111111110",
  43871=>"001011001",
  43872=>"000000100",
  43873=>"001000010",
  43874=>"110110111",
  43875=>"111111111",
  43876=>"000000000",
  43877=>"001000000",
  43878=>"111001111",
  43879=>"110000000",
  43880=>"110110110",
  43881=>"000010111",
  43882=>"010111111",
  43883=>"111111100",
  43884=>"110110100",
  43885=>"000000000",
  43886=>"010011000",
  43887=>"111111111",
  43888=>"111111011",
  43889=>"100000000",
  43890=>"111111110",
  43891=>"100000101",
  43892=>"010000001",
  43893=>"000000000",
  43894=>"111000000",
  43895=>"010100100",
  43896=>"000001101",
  43897=>"111111000",
  43898=>"111111000",
  43899=>"111111111",
  43900=>"001101111",
  43901=>"000000000",
  43902=>"111001000",
  43903=>"000100000",
  43904=>"111111111",
  43905=>"000000101",
  43906=>"000000000",
  43907=>"000000000",
  43908=>"000010011",
  43909=>"001000111",
  43910=>"000000100",
  43911=>"111000100",
  43912=>"111110100",
  43913=>"110000000",
  43914=>"100000000",
  43915=>"001111111",
  43916=>"111111111",
  43917=>"011001111",
  43918=>"000000111",
  43919=>"111111111",
  43920=>"000000000",
  43921=>"001111111",
  43922=>"001111111",
  43923=>"111111111",
  43924=>"000000000",
  43925=>"000100100",
  43926=>"001001001",
  43927=>"111111010",
  43928=>"111111111",
  43929=>"111111111",
  43930=>"111111101",
  43931=>"111111000",
  43932=>"111000000",
  43933=>"000111111",
  43934=>"010011001",
  43935=>"000000000",
  43936=>"000000000",
  43937=>"111010000",
  43938=>"000000101",
  43939=>"000000011",
  43940=>"111111111",
  43941=>"101111111",
  43942=>"101000000",
  43943=>"111111001",
  43944=>"111110000",
  43945=>"110100000",
  43946=>"111111011",
  43947=>"000000000",
  43948=>"111101101",
  43949=>"111000001",
  43950=>"110010111",
  43951=>"000000010",
  43952=>"000000011",
  43953=>"111110010",
  43954=>"111000111",
  43955=>"011011111",
  43956=>"111111000",
  43957=>"000000100",
  43958=>"000000000",
  43959=>"011111111",
  43960=>"000000000",
  43961=>"111011001",
  43962=>"010111011",
  43963=>"111111011",
  43964=>"000000100",
  43965=>"111111111",
  43966=>"110000000",
  43967=>"011011110",
  43968=>"001001001",
  43969=>"111111101",
  43970=>"011001000",
  43971=>"110111000",
  43972=>"001101111",
  43973=>"111100000",
  43974=>"010000000",
  43975=>"010010000",
  43976=>"111110111",
  43977=>"111111111",
  43978=>"100000100",
  43979=>"000000000",
  43980=>"000000000",
  43981=>"111111111",
  43982=>"011001000",
  43983=>"111111011",
  43984=>"111111000",
  43985=>"111000000",
  43986=>"000001011",
  43987=>"000010000",
  43988=>"011011111",
  43989=>"011000000",
  43990=>"110000001",
  43991=>"001011111",
  43992=>"000100110",
  43993=>"111000000",
  43994=>"011010000",
  43995=>"011000001",
  43996=>"100110111",
  43997=>"101000101",
  43998=>"000000111",
  43999=>"111111110",
  44000=>"111111111",
  44001=>"110111110",
  44002=>"011111011",
  44003=>"001000000",
  44004=>"111011110",
  44005=>"110111011",
  44006=>"000100101",
  44007=>"000000111",
  44008=>"001111101",
  44009=>"000000100",
  44010=>"010011000",
  44011=>"000000001",
  44012=>"000000000",
  44013=>"000000101",
  44014=>"100111111",
  44015=>"000100100",
  44016=>"000000000",
  44017=>"111111011",
  44018=>"000000011",
  44019=>"000100111",
  44020=>"111000111",
  44021=>"111101101",
  44022=>"110000000",
  44023=>"110010110",
  44024=>"001001001",
  44025=>"100100011",
  44026=>"000010110",
  44027=>"111111011",
  44028=>"001000000",
  44029=>"101001011",
  44030=>"110010111",
  44031=>"111111111",
  44032=>"111111111",
  44033=>"111100000",
  44034=>"000100110",
  44035=>"000001111",
  44036=>"000000000",
  44037=>"001001001",
  44038=>"000000000",
  44039=>"100111111",
  44040=>"000000101",
  44041=>"100000100",
  44042=>"111111111",
  44043=>"000000011",
  44044=>"001000000",
  44045=>"110111111",
  44046=>"000100111",
  44047=>"000000000",
  44048=>"010111110",
  44049=>"010000000",
  44050=>"001001111",
  44051=>"101000000",
  44052=>"111011001",
  44053=>"111000000",
  44054=>"111111111",
  44055=>"111111111",
  44056=>"000000000",
  44057=>"001001001",
  44058=>"000111111",
  44059=>"011001111",
  44060=>"001001000",
  44061=>"000000001",
  44062=>"000110101",
  44063=>"000111111",
  44064=>"111111000",
  44065=>"010100000",
  44066=>"001100000",
  44067=>"111111111",
  44068=>"111000000",
  44069=>"000000000",
  44070=>"111011000",
  44071=>"000000000",
  44072=>"001101111",
  44073=>"101101000",
  44074=>"111001101",
  44075=>"010011011",
  44076=>"100111111",
  44077=>"111111110",
  44078=>"111111110",
  44079=>"000000000",
  44080=>"111111111",
  44081=>"001110111",
  44082=>"100100100",
  44083=>"111111001",
  44084=>"111111111",
  44085=>"111011011",
  44086=>"000101111",
  44087=>"001111110",
  44088=>"111111100",
  44089=>"110000011",
  44090=>"111111110",
  44091=>"101000111",
  44092=>"111111111",
  44093=>"101111111",
  44094=>"011011110",
  44095=>"101000101",
  44096=>"111011011",
  44097=>"001001000",
  44098=>"111010111",
  44099=>"111111010",
  44100=>"000011011",
  44101=>"001010010",
  44102=>"101101111",
  44103=>"111100100",
  44104=>"111111111",
  44105=>"101000001",
  44106=>"111111111",
  44107=>"010111111",
  44108=>"111111111",
  44109=>"111111110",
  44110=>"001000100",
  44111=>"011011111",
  44112=>"101111111",
  44113=>"111111101",
  44114=>"000000001",
  44115=>"000000000",
  44116=>"000000000",
  44117=>"100000000",
  44118=>"111000100",
  44119=>"010000000",
  44120=>"000111111",
  44121=>"101000000",
  44122=>"001000000",
  44123=>"110110110",
  44124=>"000000101",
  44125=>"010000000",
  44126=>"001000011",
  44127=>"010111011",
  44128=>"000000000",
  44129=>"000001111",
  44130=>"111111001",
  44131=>"100101111",
  44132=>"111011001",
  44133=>"011111011",
  44134=>"111111111",
  44135=>"010111011",
  44136=>"111111111",
  44137=>"010000000",
  44138=>"000001111",
  44139=>"001111111",
  44140=>"000000100",
  44141=>"111111111",
  44142=>"001001001",
  44143=>"000101011",
  44144=>"011110111",
  44145=>"000111111",
  44146=>"001001111",
  44147=>"001000100",
  44148=>"000000011",
  44149=>"111011001",
  44150=>"111111101",
  44151=>"111001000",
  44152=>"110000000",
  44153=>"111111000",
  44154=>"000100100",
  44155=>"000000000",
  44156=>"100100000",
  44157=>"001100111",
  44158=>"000100100",
  44159=>"110000000",
  44160=>"000000000",
  44161=>"000001111",
  44162=>"111000000",
  44163=>"001001011",
  44164=>"111111011",
  44165=>"000000000",
  44166=>"111111110",
  44167=>"111111011",
  44168=>"000000000",
  44169=>"111101111",
  44170=>"111101111",
  44171=>"111111110",
  44172=>"100000000",
  44173=>"000000000",
  44174=>"000000000",
  44175=>"000000000",
  44176=>"101101111",
  44177=>"101100101",
  44178=>"000000000",
  44179=>"101101101",
  44180=>"100011111",
  44181=>"000000000",
  44182=>"111111100",
  44183=>"100000000",
  44184=>"001101111",
  44185=>"111111110",
  44186=>"000000011",
  44187=>"010110000",
  44188=>"000011001",
  44189=>"111000000",
  44190=>"101000111",
  44191=>"111111000",
  44192=>"000000110",
  44193=>"111111111",
  44194=>"000000010",
  44195=>"000000000",
  44196=>"111111111",
  44197=>"110110111",
  44198=>"010111111",
  44199=>"011111110",
  44200=>"000001000",
  44201=>"110010000",
  44202=>"000010000",
  44203=>"111111111",
  44204=>"000000000",
  44205=>"111111100",
  44206=>"110101111",
  44207=>"001001000",
  44208=>"111010000",
  44209=>"010000000",
  44210=>"011111111",
  44211=>"111111111",
  44212=>"110110111",
  44213=>"101101000",
  44214=>"000000100",
  44215=>"100000000",
  44216=>"110101111",
  44217=>"001101000",
  44218=>"100001111",
  44219=>"110110110",
  44220=>"000000000",
  44221=>"000010000",
  44222=>"111111111",
  44223=>"001000100",
  44224=>"111111011",
  44225=>"100000000",
  44226=>"111111101",
  44227=>"111111111",
  44228=>"011111111",
  44229=>"111111010",
  44230=>"000000000",
  44231=>"000111111",
  44232=>"110111111",
  44233=>"111111010",
  44234=>"111000111",
  44235=>"100100101",
  44236=>"110000000",
  44237=>"011111011",
  44238=>"010000010",
  44239=>"001000000",
  44240=>"111111001",
  44241=>"011001010",
  44242=>"000111111",
  44243=>"000000111",
  44244=>"111101000",
  44245=>"000000111",
  44246=>"000000000",
  44247=>"111000100",
  44248=>"011111111",
  44249=>"100110000",
  44250=>"000000000",
  44251=>"111111111",
  44252=>"110000000",
  44253=>"111011111",
  44254=>"111111111",
  44255=>"001001000",
  44256=>"111111111",
  44257=>"101111000",
  44258=>"000000000",
  44259=>"011000110",
  44260=>"001001000",
  44261=>"111111011",
  44262=>"111111111",
  44263=>"111110000",
  44264=>"111111111",
  44265=>"001001111",
  44266=>"000000000",
  44267=>"000000000",
  44268=>"111101101",
  44269=>"000000000",
  44270=>"111111111",
  44271=>"111111111",
  44272=>"000000000",
  44273=>"101010111",
  44274=>"111000000",
  44275=>"001001001",
  44276=>"000001111",
  44277=>"010011010",
  44278=>"111111111",
  44279=>"000000001",
  44280=>"001000000",
  44281=>"011111010",
  44282=>"000000000",
  44283=>"101101101",
  44284=>"000100100",
  44285=>"110110000",
  44286=>"111001110",
  44287=>"000001111",
  44288=>"010111100",
  44289=>"010011011",
  44290=>"111111111",
  44291=>"000000000",
  44292=>"011111100",
  44293=>"111111111",
  44294=>"101000000",
  44295=>"101000111",
  44296=>"001000000",
  44297=>"010000011",
  44298=>"000000111",
  44299=>"000000000",
  44300=>"000000011",
  44301=>"110101111",
  44302=>"111111100",
  44303=>"111111011",
  44304=>"000000010",
  44305=>"100001111",
  44306=>"101000001",
  44307=>"110110110",
  44308=>"001111111",
  44309=>"001111111",
  44310=>"110110110",
  44311=>"100111111",
  44312=>"000001111",
  44313=>"111000000",
  44314=>"111001001",
  44315=>"111111111",
  44316=>"000000000",
  44317=>"000010111",
  44318=>"111111111",
  44319=>"000000000",
  44320=>"111111111",
  44321=>"101101101",
  44322=>"000000111",
  44323=>"111111000",
  44324=>"000000010",
  44325=>"101000001",
  44326=>"111000100",
  44327=>"111010110",
  44328=>"000000010",
  44329=>"000001001",
  44330=>"011011010",
  44331=>"101001001",
  44332=>"110110110",
  44333=>"000001001",
  44334=>"111000110",
  44335=>"000000111",
  44336=>"000000110",
  44337=>"000000000",
  44338=>"111111111",
  44339=>"010111111",
  44340=>"000000000",
  44341=>"001001111",
  44342=>"000000000",
  44343=>"000000011",
  44344=>"000100100",
  44345=>"111110001",
  44346=>"111111111",
  44347=>"110110000",
  44348=>"111001001",
  44349=>"000000000",
  44350=>"000000000",
  44351=>"111000111",
  44352=>"111100100",
  44353=>"111101111",
  44354=>"111111111",
  44355=>"000000000",
  44356=>"000000000",
  44357=>"111111111",
  44358=>"000000000",
  44359=>"111100110",
  44360=>"111111111",
  44361=>"010111111",
  44362=>"111111011",
  44363=>"011000110",
  44364=>"111101111",
  44365=>"000000111",
  44366=>"111110110",
  44367=>"110011010",
  44368=>"011111011",
  44369=>"111000000",
  44370=>"111010011",
  44371=>"010011111",
  44372=>"000000000",
  44373=>"011011001",
  44374=>"111111111",
  44375=>"111111111",
  44376=>"000001011",
  44377=>"000000000",
  44378=>"111000000",
  44379=>"001000100",
  44380=>"110110000",
  44381=>"000000001",
  44382=>"001000000",
  44383=>"000000101",
  44384=>"100000101",
  44385=>"000000001",
  44386=>"100101101",
  44387=>"111111111",
  44388=>"111111111",
  44389=>"000000000",
  44390=>"000000000",
  44391=>"111000000",
  44392=>"100110110",
  44393=>"100000000",
  44394=>"000111111",
  44395=>"100000111",
  44396=>"111111011",
  44397=>"111111101",
  44398=>"111111111",
  44399=>"111001000",
  44400=>"010111111",
  44401=>"111110000",
  44402=>"111111111",
  44403=>"111111000",
  44404=>"000000000",
  44405=>"000000100",
  44406=>"000000110",
  44407=>"111000000",
  44408=>"111111011",
  44409=>"110111111",
  44410=>"011001011",
  44411=>"000010001",
  44412=>"111001000",
  44413=>"000001111",
  44414=>"100000001",
  44415=>"111100111",
  44416=>"000100110",
  44417=>"000000000",
  44418=>"110110000",
  44419=>"000000000",
  44420=>"111111000",
  44421=>"000000000",
  44422=>"000000011",
  44423=>"000000010",
  44424=>"111101111",
  44425=>"111111111",
  44426=>"111111111",
  44427=>"100000100",
  44428=>"111111111",
  44429=>"011111110",
  44430=>"011111100",
  44431=>"000000000",
  44432=>"110111000",
  44433=>"111111110",
  44434=>"000011000",
  44435=>"111011000",
  44436=>"000001101",
  44437=>"010110000",
  44438=>"111111010",
  44439=>"000000000",
  44440=>"101000000",
  44441=>"000000000",
  44442=>"000010000",
  44443=>"111111111",
  44444=>"001000111",
  44445=>"001000000",
  44446=>"000000000",
  44447=>"000000001",
  44448=>"000000000",
  44449=>"110110110",
  44450=>"000000101",
  44451=>"000000000",
  44452=>"000000000",
  44453=>"111111111",
  44454=>"111101111",
  44455=>"000000000",
  44456=>"000000000",
  44457=>"011001000",
  44458=>"111100100",
  44459=>"001000001",
  44460=>"000000000",
  44461=>"110111011",
  44462=>"111010000",
  44463=>"000001000",
  44464=>"111000110",
  44465=>"000000000",
  44466=>"000000000",
  44467=>"111111100",
  44468=>"101101101",
  44469=>"100001101",
  44470=>"000000111",
  44471=>"101111111",
  44472=>"111111111",
  44473=>"111111010",
  44474=>"000000110",
  44475=>"111011011",
  44476=>"000011111",
  44477=>"110111111",
  44478=>"000101000",
  44479=>"010011011",
  44480=>"000011111",
  44481=>"111111111",
  44482=>"111001101",
  44483=>"000000001",
  44484=>"000000000",
  44485=>"111011000",
  44486=>"110111101",
  44487=>"110000000",
  44488=>"001101001",
  44489=>"011010011",
  44490=>"000000000",
  44491=>"000010111",
  44492=>"111000000",
  44493=>"110111111",
  44494=>"111000000",
  44495=>"000100111",
  44496=>"101111111",
  44497=>"011111111",
  44498=>"111111111",
  44499=>"000011011",
  44500=>"000000001",
  44501=>"110100000",
  44502=>"000000000",
  44503=>"000001001",
  44504=>"101000111",
  44505=>"111000000",
  44506=>"000000010",
  44507=>"000000001",
  44508=>"111000000",
  44509=>"011100100",
  44510=>"000000010",
  44511=>"110111111",
  44512=>"111111111",
  44513=>"001001101",
  44514=>"001001111",
  44515=>"001011011",
  44516=>"100000111",
  44517=>"000100001",
  44518=>"111111101",
  44519=>"000000000",
  44520=>"111110011",
  44521=>"000000000",
  44522=>"100111111",
  44523=>"111111101",
  44524=>"000000000",
  44525=>"101100110",
  44526=>"101000101",
  44527=>"011011001",
  44528=>"000000100",
  44529=>"000101000",
  44530=>"101000000",
  44531=>"000100110",
  44532=>"000000000",
  44533=>"000111000",
  44534=>"000000000",
  44535=>"110110010",
  44536=>"101001000",
  44537=>"111111011",
  44538=>"001111111",
  44539=>"011001001",
  44540=>"111011000",
  44541=>"110111110",
  44542=>"111111000",
  44543=>"000000000",
  44544=>"010111111",
  44545=>"000000000",
  44546=>"000000111",
  44547=>"110111111",
  44548=>"110111101",
  44549=>"000000101",
  44550=>"111111111",
  44551=>"000000000",
  44552=>"000010100",
  44553=>"011111110",
  44554=>"111111000",
  44555=>"011001111",
  44556=>"110110110",
  44557=>"111111110",
  44558=>"000100111",
  44559=>"001000000",
  44560=>"000100101",
  44561=>"000000000",
  44562=>"000000000",
  44563=>"000000000",
  44564=>"111111111",
  44565=>"000011111",
  44566=>"000111110",
  44567=>"110100110",
  44568=>"100100100",
  44569=>"000000100",
  44570=>"000000111",
  44571=>"000001111",
  44572=>"100100100",
  44573=>"111111101",
  44574=>"111111111",
  44575=>"000000000",
  44576=>"111111110",
  44577=>"000000000",
  44578=>"000001001",
  44579=>"001001001",
  44580=>"110111111",
  44581=>"101100100",
  44582=>"111101100",
  44583=>"000000000",
  44584=>"001000011",
  44585=>"111111111",
  44586=>"000000000",
  44587=>"011001011",
  44588=>"011001000",
  44589=>"011001001",
  44590=>"000000000",
  44591=>"111111100",
  44592=>"000100000",
  44593=>"000000000",
  44594=>"111001000",
  44595=>"001000000",
  44596=>"011001001",
  44597=>"110111111",
  44598=>"000110111",
  44599=>"010111111",
  44600=>"111000000",
  44601=>"000000111",
  44602=>"000010010",
  44603=>"000000000",
  44604=>"000000000",
  44605=>"101000000",
  44606=>"000001111",
  44607=>"101000001",
  44608=>"111011001",
  44609=>"000000101",
  44610=>"010111111",
  44611=>"001100110",
  44612=>"000000000",
  44613=>"110110000",
  44614=>"000000100",
  44615=>"000000111",
  44616=>"011111111",
  44617=>"111111000",
  44618=>"101000000",
  44619=>"111111101",
  44620=>"111111100",
  44621=>"101000000",
  44622=>"000010011",
  44623=>"000100100",
  44624=>"001011011",
  44625=>"000100000",
  44626=>"000000000",
  44627=>"111111111",
  44628=>"000100111",
  44629=>"111001100",
  44630=>"111111111",
  44631=>"110110110",
  44632=>"111011000",
  44633=>"111000000",
  44634=>"110000000",
  44635=>"000001011",
  44636=>"000000000",
  44637=>"000100100",
  44638=>"111111101",
  44639=>"000011011",
  44640=>"111000000",
  44641=>"000010011",
  44642=>"101001101",
  44643=>"000001000",
  44644=>"110111000",
  44645=>"010000000",
  44646=>"110111111",
  44647=>"000000100",
  44648=>"111111111",
  44649=>"111100000",
  44650=>"111111111",
  44651=>"111111111",
  44652=>"000011111",
  44653=>"000000001",
  44654=>"000000100",
  44655=>"000000001",
  44656=>"011010110",
  44657=>"001000000",
  44658=>"011011111",
  44659=>"000000001",
  44660=>"111111111",
  44661=>"000000100",
  44662=>"100000100",
  44663=>"000000011",
  44664=>"000000110",
  44665=>"111001000",
  44666=>"000000000",
  44667=>"100000000",
  44668=>"000000000",
  44669=>"111111111",
  44670=>"000000000",
  44671=>"101001101",
  44672=>"000000000",
  44673=>"001000111",
  44674=>"110000000",
  44675=>"000000011",
  44676=>"000011011",
  44677=>"000010010",
  44678=>"111011011",
  44679=>"111111111",
  44680=>"110010111",
  44681=>"010000001",
  44682=>"010011000",
  44683=>"111111111",
  44684=>"000101111",
  44685=>"110111111",
  44686=>"011111111",
  44687=>"010000000",
  44688=>"101000000",
  44689=>"001111100",
  44690=>"011011011",
  44691=>"001001001",
  44692=>"111111111",
  44693=>"000110110",
  44694=>"000010010",
  44695=>"001000001",
  44696=>"111000000",
  44697=>"111111111",
  44698=>"111011011",
  44699=>"110110100",
  44700=>"110111111",
  44701=>"111111111",
  44702=>"111111111",
  44703=>"000000000",
  44704=>"110000000",
  44705=>"010011011",
  44706=>"000110111",
  44707=>"111111111",
  44708=>"000000000",
  44709=>"000100111",
  44710=>"101100101",
  44711=>"000101111",
  44712=>"111111111",
  44713=>"011000001",
  44714=>"111000000",
  44715=>"111111111",
  44716=>"000000100",
  44717=>"000001001",
  44718=>"111000000",
  44719=>"001000001",
  44720=>"000000000",
  44721=>"000000001",
  44722=>"111100000",
  44723=>"111000001",
  44724=>"000011001",
  44725=>"101001101",
  44726=>"010111011",
  44727=>"111001000",
  44728=>"000000000",
  44729=>"011110110",
  44730=>"101000000",
  44731=>"011000100",
  44732=>"111110000",
  44733=>"111111111",
  44734=>"000000110",
  44735=>"011111011",
  44736=>"110111111",
  44737=>"000000000",
  44738=>"111111111",
  44739=>"000000001",
  44740=>"000001001",
  44741=>"111000000",
  44742=>"001100101",
  44743=>"101110100",
  44744=>"100111111",
  44745=>"110100100",
  44746=>"000000110",
  44747=>"100100000",
  44748=>"011011111",
  44749=>"000000000",
  44750=>"011111111",
  44751=>"100000101",
  44752=>"111111110",
  44753=>"100100000",
  44754=>"100110000",
  44755=>"110111110",
  44756=>"110111111",
  44757=>"111111100",
  44758=>"000000000",
  44759=>"000111111",
  44760=>"000000111",
  44761=>"100000000",
  44762=>"011111111",
  44763=>"010010000",
  44764=>"110010000",
  44765=>"000000001",
  44766=>"111100000",
  44767=>"110000000",
  44768=>"110100100",
  44769=>"000000010",
  44770=>"010010111",
  44771=>"111111011",
  44772=>"000000100",
  44773=>"000000000",
  44774=>"000000111",
  44775=>"111000000",
  44776=>"010000000",
  44777=>"010000100",
  44778=>"001000000",
  44779=>"010010010",
  44780=>"111101000",
  44781=>"111000000",
  44782=>"100100001",
  44783=>"010110110",
  44784=>"111101101",
  44785=>"111111111",
  44786=>"110111111",
  44787=>"011100000",
  44788=>"000000000",
  44789=>"000011111",
  44790=>"011111111",
  44791=>"111111111",
  44792=>"111111111",
  44793=>"111111111",
  44794=>"001001000",
  44795=>"111100000",
  44796=>"110111111",
  44797=>"001001000",
  44798=>"110010000",
  44799=>"000111011",
  44800=>"000000000",
  44801=>"000101101",
  44802=>"111111111",
  44803=>"000111100",
  44804=>"001001101",
  44805=>"010111011",
  44806=>"111001000",
  44807=>"111111000",
  44808=>"000000000",
  44809=>"110000100",
  44810=>"000011011",
  44811=>"000000110",
  44812=>"110000100",
  44813=>"111111001",
  44814=>"000000000",
  44815=>"000000000",
  44816=>"000000111",
  44817=>"010111101",
  44818=>"110110111",
  44819=>"000000000",
  44820=>"000000000",
  44821=>"000000000",
  44822=>"001111001",
  44823=>"110111110",
  44824=>"001111111",
  44825=>"111111010",
  44826=>"110111100",
  44827=>"000100001",
  44828=>"110110110",
  44829=>"111111110",
  44830=>"000000000",
  44831=>"111000001",
  44832=>"001000010",
  44833=>"111111000",
  44834=>"111000000",
  44835=>"001011111",
  44836=>"000100100",
  44837=>"000000111",
  44838=>"011001000",
  44839=>"111111000",
  44840=>"011001011",
  44841=>"111111110",
  44842=>"000000000",
  44843=>"111101111",
  44844=>"000000111",
  44845=>"001001101",
  44846=>"000100000",
  44847=>"000000110",
  44848=>"011111111",
  44849=>"111100111",
  44850=>"000000000",
  44851=>"111000000",
  44852=>"111001111",
  44853=>"011011011",
  44854=>"000000000",
  44855=>"011000000",
  44856=>"001000000",
  44857=>"001000101",
  44858=>"100000000",
  44859=>"111001101",
  44860=>"100000000",
  44861=>"000000000",
  44862=>"000100100",
  44863=>"000000111",
  44864=>"111111100",
  44865=>"111111110",
  44866=>"111111111",
  44867=>"110110111",
  44868=>"001011011",
  44869=>"110110010",
  44870=>"100111111",
  44871=>"000001101",
  44872=>"000000000",
  44873=>"111111000",
  44874=>"111111001",
  44875=>"111111111",
  44876=>"111111111",
  44877=>"111110000",
  44878=>"000010001",
  44879=>"100110110",
  44880=>"111011001",
  44881=>"000000000",
  44882=>"111111010",
  44883=>"111100100",
  44884=>"100010011",
  44885=>"001001001",
  44886=>"111001000",
  44887=>"000000000",
  44888=>"000000000",
  44889=>"000000011",
  44890=>"000001101",
  44891=>"111001000",
  44892=>"111111000",
  44893=>"000000000",
  44894=>"010110011",
  44895=>"111001101",
  44896=>"011000010",
  44897=>"100100000",
  44898=>"011001000",
  44899=>"000000111",
  44900=>"110110111",
  44901=>"111111110",
  44902=>"111000000",
  44903=>"000110100",
  44904=>"011001110",
  44905=>"000000010",
  44906=>"110111000",
  44907=>"110111111",
  44908=>"000000010",
  44909=>"101000101",
  44910=>"111111111",
  44911=>"000000101",
  44912=>"000000000",
  44913=>"000000111",
  44914=>"111111011",
  44915=>"111101111",
  44916=>"110000100",
  44917=>"001111000",
  44918=>"111111011",
  44919=>"000000000",
  44920=>"000000000",
  44921=>"100100100",
  44922=>"110010111",
  44923=>"100000000",
  44924=>"000000110",
  44925=>"001001111",
  44926=>"110110110",
  44927=>"000010111",
  44928=>"001000100",
  44929=>"011000010",
  44930=>"110111111",
  44931=>"100110111",
  44932=>"110110110",
  44933=>"000000011",
  44934=>"000000111",
  44935=>"011011011",
  44936=>"110010111",
  44937=>"000110011",
  44938=>"100100100",
  44939=>"011011111",
  44940=>"111011111",
  44941=>"000000000",
  44942=>"001000110",
  44943=>"000001111",
  44944=>"100100111",
  44945=>"001111111",
  44946=>"111110111",
  44947=>"100101111",
  44948=>"100101111",
  44949=>"000000000",
  44950=>"111011000",
  44951=>"001001001",
  44952=>"111111111",
  44953=>"000100111",
  44954=>"111000101",
  44955=>"001000100",
  44956=>"110111110",
  44957=>"111111011",
  44958=>"000001111",
  44959=>"110000000",
  44960=>"000000000",
  44961=>"100000000",
  44962=>"000000000",
  44963=>"111111111",
  44964=>"000000111",
  44965=>"111101001",
  44966=>"101101000",
  44967=>"100110000",
  44968=>"110100000",
  44969=>"001001111",
  44970=>"000000000",
  44971=>"111101011",
  44972=>"000000101",
  44973=>"010011000",
  44974=>"000000000",
  44975=>"110100110",
  44976=>"000000011",
  44977=>"100000000",
  44978=>"010001000",
  44979=>"111111000",
  44980=>"001000001",
  44981=>"001001001",
  44982=>"011000000",
  44983=>"000000000",
  44984=>"111100100",
  44985=>"001000000",
  44986=>"010000000",
  44987=>"000000000",
  44988=>"111101101",
  44989=>"000111111",
  44990=>"001001111",
  44991=>"001001101",
  44992=>"011111000",
  44993=>"000000000",
  44994=>"111111000",
  44995=>"000000000",
  44996=>"111101001",
  44997=>"111111100",
  44998=>"011111111",
  44999=>"111101001",
  45000=>"000000000",
  45001=>"111001000",
  45002=>"111000101",
  45003=>"111111001",
  45004=>"000000000",
  45005=>"000000000",
  45006=>"111001000",
  45007=>"110111110",
  45008=>"011011000",
  45009=>"011111111",
  45010=>"101011001",
  45011=>"000000100",
  45012=>"100100001",
  45013=>"000000100",
  45014=>"100000000",
  45015=>"001001011",
  45016=>"000000101",
  45017=>"010000100",
  45018=>"111111000",
  45019=>"101000100",
  45020=>"111111111",
  45021=>"011000000",
  45022=>"100100100",
  45023=>"000111111",
  45024=>"011111110",
  45025=>"000110110",
  45026=>"111000110",
  45027=>"000000011",
  45028=>"101100000",
  45029=>"111111111",
  45030=>"000000000",
  45031=>"110111111",
  45032=>"001000000",
  45033=>"100001000",
  45034=>"110010010",
  45035=>"111111101",
  45036=>"100000000",
  45037=>"101100111",
  45038=>"111111111",
  45039=>"111110011",
  45040=>"100100100",
  45041=>"110000111",
  45042=>"010011011",
  45043=>"111100100",
  45044=>"000000001",
  45045=>"110000000",
  45046=>"000000101",
  45047=>"011010000",
  45048=>"010001011",
  45049=>"110000000",
  45050=>"000000000",
  45051=>"111000000",
  45052=>"111100110",
  45053=>"000000000",
  45054=>"001000000",
  45055=>"111001111",
  45056=>"110000000",
  45057=>"000000111",
  45058=>"111111111",
  45059=>"110000001",
  45060=>"111111111",
  45061=>"000000111",
  45062=>"000011111",
  45063=>"001111111",
  45064=>"101111000",
  45065=>"001011000",
  45066=>"001001000",
  45067=>"000000000",
  45068=>"000000010",
  45069=>"101000000",
  45070=>"000000100",
  45071=>"001011000",
  45072=>"110001011",
  45073=>"000111111",
  45074=>"000110100",
  45075=>"000010000",
  45076=>"100000000",
  45077=>"000000111",
  45078=>"100110111",
  45079=>"000100110",
  45080=>"111111111",
  45081=>"010010000",
  45082=>"000000000",
  45083=>"011011011",
  45084=>"000000000",
  45085=>"110000000",
  45086=>"001001001",
  45087=>"111111111",
  45088=>"000000000",
  45089=>"000000001",
  45090=>"000000000",
  45091=>"000000000",
  45092=>"111111001",
  45093=>"000000000",
  45094=>"000100111",
  45095=>"011000000",
  45096=>"111100000",
  45097=>"000000011",
  45098=>"000000000",
  45099=>"100111111",
  45100=>"001101111",
  45101=>"000101111",
  45102=>"111111111",
  45103=>"000010000",
  45104=>"000000001",
  45105=>"000000000",
  45106=>"011000100",
  45107=>"100000111",
  45108=>"111111111",
  45109=>"000000100",
  45110=>"001000100",
  45111=>"000111111",
  45112=>"111111000",
  45113=>"000000000",
  45114=>"000000000",
  45115=>"000000111",
  45116=>"111001001",
  45117=>"111111111",
  45118=>"111101111",
  45119=>"000000000",
  45120=>"011111000",
  45121=>"111111111",
  45122=>"111111111",
  45123=>"111111111",
  45124=>"000000000",
  45125=>"110100000",
  45126=>"000000000",
  45127=>"111111111",
  45128=>"011001001",
  45129=>"010000000",
  45130=>"001111111",
  45131=>"111111000",
  45132=>"000000000",
  45133=>"000010111",
  45134=>"011000000",
  45135=>"111000111",
  45136=>"000111110",
  45137=>"000000001",
  45138=>"011111000",
  45139=>"000000011",
  45140=>"000000000",
  45141=>"111101000",
  45142=>"111011111",
  45143=>"111000111",
  45144=>"111000100",
  45145=>"000000010",
  45146=>"111001000",
  45147=>"111000000",
  45148=>"000000000",
  45149=>"000000111",
  45150=>"111111111",
  45151=>"100100000",
  45152=>"000000000",
  45153=>"111111000",
  45154=>"110000000",
  45155=>"000000111",
  45156=>"001111111",
  45157=>"000000000",
  45158=>"100111111",
  45159=>"000100110",
  45160=>"000011000",
  45161=>"111111111",
  45162=>"000000000",
  45163=>"111110000",
  45164=>"111111110",
  45165=>"000111101",
  45166=>"111110100",
  45167=>"111111111",
  45168=>"010110111",
  45169=>"000001011",
  45170=>"111101000",
  45171=>"110110001",
  45172=>"000000000",
  45173=>"111110100",
  45174=>"111111111",
  45175=>"000000000",
  45176=>"110110100",
  45177=>"000000110",
  45178=>"000000000",
  45179=>"000000000",
  45180=>"110111111",
  45181=>"111000000",
  45182=>"000000000",
  45183=>"000010111",
  45184=>"001101111",
  45185=>"110000000",
  45186=>"111000000",
  45187=>"000000100",
  45188=>"000110110",
  45189=>"111000000",
  45190=>"000000000",
  45191=>"110000110",
  45192=>"110100000",
  45193=>"111000000",
  45194=>"011000000",
  45195=>"000001001",
  45196=>"000110111",
  45197=>"000000000",
  45198=>"110111111",
  45199=>"111111001",
  45200=>"111111111",
  45201=>"111011111",
  45202=>"011010000",
  45203=>"000000000",
  45204=>"000000111",
  45205=>"000000001",
  45206=>"111111111",
  45207=>"111111111",
  45208=>"000000000",
  45209=>"111111101",
  45210=>"111000101",
  45211=>"000011001",
  45212=>"000000000",
  45213=>"000000100",
  45214=>"000000000",
  45215=>"000000000",
  45216=>"111111000",
  45217=>"001011001",
  45218=>"110111110",
  45219=>"000000000",
  45220=>"000000000",
  45221=>"000011111",
  45222=>"111111111",
  45223=>"111111111",
  45224=>"111001011",
  45225=>"000000000",
  45226=>"111111111",
  45227=>"110010000",
  45228=>"111111111",
  45229=>"000000000",
  45230=>"000000000",
  45231=>"111100000",
  45232=>"000010000",
  45233=>"111111111",
  45234=>"110110110",
  45235=>"111111111",
  45236=>"000000001",
  45237=>"111111111",
  45238=>"111001101",
  45239=>"111111000",
  45240=>"111100001",
  45241=>"000000111",
  45242=>"000000000",
  45243=>"111111111",
  45244=>"000100101",
  45245=>"111111111",
  45246=>"000000000",
  45247=>"011011000",
  45248=>"111111111",
  45249=>"000000000",
  45250=>"000000000",
  45251=>"000000111",
  45252=>"000000110",
  45253=>"000000000",
  45254=>"111111010",
  45255=>"000011000",
  45256=>"000111101",
  45257=>"000011111",
  45258=>"111111010",
  45259=>"010000110",
  45260=>"111111000",
  45261=>"111111111",
  45262=>"000000101",
  45263=>"000000000",
  45264=>"111111000",
  45265=>"000110000",
  45266=>"111111111",
  45267=>"000010111",
  45268=>"001000111",
  45269=>"000111111",
  45270=>"000000000",
  45271=>"111111110",
  45272=>"000000000",
  45273=>"111111111",
  45274=>"111100000",
  45275=>"110111111",
  45276=>"001000000",
  45277=>"100110111",
  45278=>"001111111",
  45279=>"000000000",
  45280=>"000000010",
  45281=>"000011111",
  45282=>"101101000",
  45283=>"111001000",
  45284=>"111111111",
  45285=>"110110000",
  45286=>"000000000",
  45287=>"111100101",
  45288=>"001001001",
  45289=>"001110111",
  45290=>"001000000",
  45291=>"001111111",
  45292=>"111111000",
  45293=>"111110111",
  45294=>"110010000",
  45295=>"000111111",
  45296=>"111100111",
  45297=>"000010000",
  45298=>"000111101",
  45299=>"000000001",
  45300=>"000000011",
  45301=>"111000000",
  45302=>"110111000",
  45303=>"000100100",
  45304=>"000000000",
  45305=>"111111000",
  45306=>"111001000",
  45307=>"011011000",
  45308=>"001001111",
  45309=>"000110110",
  45310=>"000110110",
  45311=>"111111101",
  45312=>"000000000",
  45313=>"111111011",
  45314=>"000000011",
  45315=>"110111000",
  45316=>"110110000",
  45317=>"111110110",
  45318=>"000111111",
  45319=>"111101000",
  45320=>"110100000",
  45321=>"000000111",
  45322=>"111100000",
  45323=>"000000111",
  45324=>"110000000",
  45325=>"111001111",
  45326=>"000000111",
  45327=>"111011000",
  45328=>"111111000",
  45329=>"111001001",
  45330=>"000000000",
  45331=>"111100111",
  45332=>"000000000",
  45333=>"000000111",
  45334=>"110110111",
  45335=>"011011111",
  45336=>"100111111",
  45337=>"000000000",
  45338=>"111011111",
  45339=>"100100111",
  45340=>"111000000",
  45341=>"111101111",
  45342=>"001000000",
  45343=>"111111111",
  45344=>"111111111",
  45345=>"010000000",
  45346=>"011010000",
  45347=>"111100000",
  45348=>"010000000",
  45349=>"000111101",
  45350=>"000001011",
  45351=>"100100001",
  45352=>"000000111",
  45353=>"001111000",
  45354=>"000000000",
  45355=>"000000000",
  45356=>"111100110",
  45357=>"111000001",
  45358=>"000000000",
  45359=>"010000000",
  45360=>"000000000",
  45361=>"000000000",
  45362=>"111101111",
  45363=>"110111111",
  45364=>"111111111",
  45365=>"111111100",
  45366=>"011000011",
  45367=>"011111111",
  45368=>"110110000",
  45369=>"000000000",
  45370=>"000111111",
  45371=>"000000000",
  45372=>"111001111",
  45373=>"001001000",
  45374=>"111111111",
  45375=>"000111111",
  45376=>"000000000",
  45377=>"000000000",
  45378=>"000000000",
  45379=>"111111111",
  45380=>"111111111",
  45381=>"111111110",
  45382=>"111111111",
  45383=>"111111100",
  45384=>"000000011",
  45385=>"111111000",
  45386=>"000000000",
  45387=>"100100000",
  45388=>"000000111",
  45389=>"100000111",
  45390=>"111101111",
  45391=>"111111100",
  45392=>"110110100",
  45393=>"000000111",
  45394=>"101000000",
  45395=>"111111011",
  45396=>"000000000",
  45397=>"001001001",
  45398=>"100000000",
  45399=>"111011000",
  45400=>"110100000",
  45401=>"000000000",
  45402=>"101100000",
  45403=>"011000001",
  45404=>"000000001",
  45405=>"101001100",
  45406=>"000000000",
  45407=>"011011111",
  45408=>"000000001",
  45409=>"111111111",
  45410=>"011111111",
  45411=>"111111011",
  45412=>"111111111",
  45413=>"111111111",
  45414=>"000000000",
  45415=>"111111111",
  45416=>"011011001",
  45417=>"010110000",
  45418=>"000000000",
  45419=>"000000011",
  45420=>"100100110",
  45421=>"111111100",
  45422=>"000000000",
  45423=>"011011111",
  45424=>"111111111",
  45425=>"000000000",
  45426=>"111001000",
  45427=>"000011011",
  45428=>"111111011",
  45429=>"110111111",
  45430=>"010010010",
  45431=>"111011011",
  45432=>"000000000",
  45433=>"111010111",
  45434=>"111111000",
  45435=>"010010010",
  45436=>"000000000",
  45437=>"110001000",
  45438=>"111111000",
  45439=>"111111110",
  45440=>"001001111",
  45441=>"101000000",
  45442=>"111000000",
  45443=>"000011000",
  45444=>"000000111",
  45445=>"111111111",
  45446=>"000111001",
  45447=>"111111000",
  45448=>"011001000",
  45449=>"000001111",
  45450=>"000100001",
  45451=>"111111000",
  45452=>"111111111",
  45453=>"000010000",
  45454=>"100000000",
  45455=>"000000000",
  45456=>"111111111",
  45457=>"111111111",
  45458=>"111111011",
  45459=>"111111111",
  45460=>"111111111",
  45461=>"000000000",
  45462=>"000000100",
  45463=>"000000100",
  45464=>"001011111",
  45465=>"110000000",
  45466=>"111111111",
  45467=>"000000000",
  45468=>"110100000",
  45469=>"000110111",
  45470=>"000000000",
  45471=>"000000000",
  45472=>"111111100",
  45473=>"001100000",
  45474=>"000000001",
  45475=>"111111111",
  45476=>"001111111",
  45477=>"000000000",
  45478=>"000000000",
  45479=>"110010010",
  45480=>"111000000",
  45481=>"111111011",
  45482=>"111111111",
  45483=>"000000111",
  45484=>"000000000",
  45485=>"011001001",
  45486=>"000000010",
  45487=>"000000111",
  45488=>"010111111",
  45489=>"111111010",
  45490=>"000100100",
  45491=>"000001000",
  45492=>"010111111",
  45493=>"000000100",
  45494=>"111111111",
  45495=>"000000000",
  45496=>"000010000",
  45497=>"000110101",
  45498=>"000000111",
  45499=>"111011111",
  45500=>"011111111",
  45501=>"110100111",
  45502=>"010010111",
  45503=>"011011010",
  45504=>"000000000",
  45505=>"000010111",
  45506=>"000000011",
  45507=>"000000000",
  45508=>"001000100",
  45509=>"101111100",
  45510=>"101001111",
  45511=>"000111111",
  45512=>"000110000",
  45513=>"111100000",
  45514=>"000000000",
  45515=>"111111111",
  45516=>"011011111",
  45517=>"111111111",
  45518=>"000000000",
  45519=>"011111111",
  45520=>"011000000",
  45521=>"110111111",
  45522=>"000111111",
  45523=>"000000000",
  45524=>"111111111",
  45525=>"111101111",
  45526=>"000000000",
  45527=>"010000100",
  45528=>"000000000",
  45529=>"010000000",
  45530=>"110111111",
  45531=>"111001011",
  45532=>"000000011",
  45533=>"000101001",
  45534=>"111111111",
  45535=>"001001011",
  45536=>"111011111",
  45537=>"000111111",
  45538=>"000000111",
  45539=>"000000000",
  45540=>"111111111",
  45541=>"111101111",
  45542=>"111000000",
  45543=>"100100111",
  45544=>"100101111",
  45545=>"000000010",
  45546=>"110000000",
  45547=>"000011011",
  45548=>"000000111",
  45549=>"111010010",
  45550=>"000000000",
  45551=>"000000111",
  45552=>"000000000",
  45553=>"000000000",
  45554=>"001100100",
  45555=>"111110000",
  45556=>"000000000",
  45557=>"110111111",
  45558=>"000011011",
  45559=>"110010000",
  45560=>"000000111",
  45561=>"110110100",
  45562=>"000000000",
  45563=>"111111111",
  45564=>"000000000",
  45565=>"111111111",
  45566=>"010000111",
  45567=>"100110110",
  45568=>"000000000",
  45569=>"011111111",
  45570=>"000000011",
  45571=>"111110000",
  45572=>"000000000",
  45573=>"011001100",
  45574=>"100100000",
  45575=>"100000100",
  45576=>"111111010",
  45577=>"111111000",
  45578=>"000000110",
  45579=>"111111111",
  45580=>"000100100",
  45581=>"111111110",
  45582=>"000000000",
  45583=>"100110111",
  45584=>"110001001",
  45585=>"000111111",
  45586=>"100100100",
  45587=>"111011111",
  45588=>"000000011",
  45589=>"111101111",
  45590=>"000000000",
  45591=>"111111111",
  45592=>"111100100",
  45593=>"110111111",
  45594=>"001101001",
  45595=>"000100111",
  45596=>"111111111",
  45597=>"100100111",
  45598=>"001011111",
  45599=>"000100111",
  45600=>"100100111",
  45601=>"111111111",
  45602=>"111011001",
  45603=>"110000111",
  45604=>"111110000",
  45605=>"111111111",
  45606=>"100000111",
  45607=>"111111010",
  45608=>"001011111",
  45609=>"001111000",
  45610=>"111111110",
  45611=>"101000000",
  45612=>"111000000",
  45613=>"100000100",
  45614=>"000111110",
  45615=>"000000000",
  45616=>"111101000",
  45617=>"000000110",
  45618=>"111111001",
  45619=>"000000000",
  45620=>"000100000",
  45621=>"000000111",
  45622=>"000000000",
  45623=>"101100111",
  45624=>"111111000",
  45625=>"100000111",
  45626=>"110010000",
  45627=>"011001000",
  45628=>"000000110",
  45629=>"111111111",
  45630=>"000000001",
  45631=>"111111000",
  45632=>"100000000",
  45633=>"000000000",
  45634=>"000110111",
  45635=>"011000111",
  45636=>"001000000",
  45637=>"011111110",
  45638=>"111000000",
  45639=>"111000000",
  45640=>"011111011",
  45641=>"101000111",
  45642=>"111100111",
  45643=>"000000001",
  45644=>"111111000",
  45645=>"000000111",
  45646=>"001000010",
  45647=>"111000100",
  45648=>"000000000",
  45649=>"001001001",
  45650=>"000000111",
  45651=>"011000001",
  45652=>"000000000",
  45653=>"010000000",
  45654=>"111111000",
  45655=>"111111000",
  45656=>"011111111",
  45657=>"111000111",
  45658=>"111111000",
  45659=>"000000100",
  45660=>"000000000",
  45661=>"000000111",
  45662=>"110000000",
  45663=>"000011000",
  45664=>"000000111",
  45665=>"111111011",
  45666=>"001001001",
  45667=>"000001110",
  45668=>"111110000",
  45669=>"100100000",
  45670=>"001001111",
  45671=>"110001000",
  45672=>"011011111",
  45673=>"000000000",
  45674=>"100000110",
  45675=>"000001111",
  45676=>"011000100",
  45677=>"000000111",
  45678=>"111011001",
  45679=>"111111111",
  45680=>"111111110",
  45681=>"000000001",
  45682=>"100100000",
  45683=>"001001111",
  45684=>"000000000",
  45685=>"000100111",
  45686=>"000010111",
  45687=>"000000110",
  45688=>"000000000",
  45689=>"000000001",
  45690=>"001001111",
  45691=>"000000111",
  45692=>"100100100",
  45693=>"100100110",
  45694=>"000000000",
  45695=>"000000000",
  45696=>"110111111",
  45697=>"110111111",
  45698=>"011011000",
  45699=>"111100110",
  45700=>"000100100",
  45701=>"000000000",
  45702=>"110011000",
  45703=>"000011111",
  45704=>"111111000",
  45705=>"001000000",
  45706=>"111010000",
  45707=>"111111111",
  45708=>"000000101",
  45709=>"101001100",
  45710=>"110100000",
  45711=>"000010010",
  45712=>"000000000",
  45713=>"000000000",
  45714=>"111111000",
  45715=>"000000111",
  45716=>"111111001",
  45717=>"111011110",
  45718=>"001101011",
  45719=>"111111000",
  45720=>"100000000",
  45721=>"111111000",
  45722=>"000000000",
  45723=>"000000111",
  45724=>"110110000",
  45725=>"000000000",
  45726=>"111111111",
  45727=>"111111000",
  45728=>"111111111",
  45729=>"000111111",
  45730=>"010011110",
  45731=>"111111111",
  45732=>"000000000",
  45733=>"110000000",
  45734=>"111101111",
  45735=>"100100110",
  45736=>"000000010",
  45737=>"001111111",
  45738=>"111000000",
  45739=>"000000111",
  45740=>"001000001",
  45741=>"111111111",
  45742=>"110111111",
  45743=>"101110110",
  45744=>"111110000",
  45745=>"000101110",
  45746=>"110111011",
  45747=>"000001000",
  45748=>"000000000",
  45749=>"110000000",
  45750=>"000000000",
  45751=>"000100000",
  45752=>"100000000",
  45753=>"111001111",
  45754=>"000000000",
  45755=>"110100100",
  45756=>"001000000",
  45757=>"000000111",
  45758=>"000101011",
  45759=>"111110111",
  45760=>"111111001",
  45761=>"111111000",
  45762=>"111000000",
  45763=>"111111111",
  45764=>"111111110",
  45765=>"000000000",
  45766=>"000011111",
  45767=>"111000100",
  45768=>"011111110",
  45769=>"011001000",
  45770=>"111100000",
  45771=>"010111111",
  45772=>"101001011",
  45773=>"000111111",
  45774=>"111111010",
  45775=>"111111000",
  45776=>"111111100",
  45777=>"011111000",
  45778=>"001000000",
  45779=>"111101111",
  45780=>"111111111",
  45781=>"000000000",
  45782=>"001000000",
  45783=>"011010001",
  45784=>"000000010",
  45785=>"000000111",
  45786=>"111111101",
  45787=>"010010110",
  45788=>"111111010",
  45789=>"111111000",
  45790=>"000001111",
  45791=>"000000111",
  45792=>"111000000",
  45793=>"011011111",
  45794=>"111000000",
  45795=>"100000000",
  45796=>"000000000",
  45797=>"000110111",
  45798=>"100000000",
  45799=>"000000001",
  45800=>"111111000",
  45801=>"000000011",
  45802=>"000000000",
  45803=>"001001111",
  45804=>"000111111",
  45805=>"000000011",
  45806=>"111111011",
  45807=>"111001000",
  45808=>"110110000",
  45809=>"001000000",
  45810=>"000000111",
  45811=>"000000001",
  45812=>"110111111",
  45813=>"000100101",
  45814=>"000100011",
  45815=>"111000010",
  45816=>"000000100",
  45817=>"000001111",
  45818=>"000000000",
  45819=>"000100110",
  45820=>"000000000",
  45821=>"011100000",
  45822=>"000010000",
  45823=>"100000000",
  45824=>"100000100",
  45825=>"001001000",
  45826=>"111111111",
  45827=>"111000000",
  45828=>"011011011",
  45829=>"111111111",
  45830=>"000000000",
  45831=>"111000000",
  45832=>"110011010",
  45833=>"000000000",
  45834=>"000000000",
  45835=>"000000000",
  45836=>"111111101",
  45837=>"000000000",
  45838=>"000000111",
  45839=>"111101100",
  45840=>"000001001",
  45841=>"000110111",
  45842=>"001000111",
  45843=>"000000100",
  45844=>"011001000",
  45845=>"000000001",
  45846=>"100111111",
  45847=>"000000111",
  45848=>"001001111",
  45849=>"111110000",
  45850=>"000000000",
  45851=>"111110110",
  45852=>"110110000",
  45853=>"000000000",
  45854=>"000000000",
  45855=>"111011111",
  45856=>"000001000",
  45857=>"111111110",
  45858=>"111111111",
  45859=>"001000000",
  45860=>"011011000",
  45861=>"000100110",
  45862=>"111111111",
  45863=>"000000000",
  45864=>"111011000",
  45865=>"000001000",
  45866=>"001000111",
  45867=>"101001111",
  45868=>"000001111",
  45869=>"000000000",
  45870=>"111000000",
  45871=>"000000111",
  45872=>"110111000",
  45873=>"110010000",
  45874=>"110111110",
  45875=>"001001011",
  45876=>"000010000",
  45877=>"001000000",
  45878=>"001000000",
  45879=>"001000000",
  45880=>"000000000",
  45881=>"000000111",
  45882=>"111000000",
  45883=>"000000000",
  45884=>"100000000",
  45885=>"000000000",
  45886=>"000000000",
  45887=>"111111000",
  45888=>"000000000",
  45889=>"111111111",
  45890=>"100100000",
  45891=>"001011000",
  45892=>"000011111",
  45893=>"011000000",
  45894=>"010011000",
  45895=>"101000000",
  45896=>"000000100",
  45897=>"000111111",
  45898=>"001000000",
  45899=>"000000000",
  45900=>"111111111",
  45901=>"111111110",
  45902=>"111111111",
  45903=>"111111011",
  45904=>"000101001",
  45905=>"110000000",
  45906=>"111110011",
  45907=>"111111111",
  45908=>"111000000",
  45909=>"001001001",
  45910=>"111011000",
  45911=>"000000011",
  45912=>"111100111",
  45913=>"111000000",
  45914=>"111111111",
  45915=>"110110110",
  45916=>"001101001",
  45917=>"000111111",
  45918=>"111000000",
  45919=>"000000000",
  45920=>"000110111",
  45921=>"001000111",
  45922=>"100110000",
  45923=>"101100100",
  45924=>"001001000",
  45925=>"000000110",
  45926=>"000000000",
  45927=>"111111111",
  45928=>"111111110",
  45929=>"000000000",
  45930=>"001111001",
  45931=>"111010000",
  45932=>"110111000",
  45933=>"000100000",
  45934=>"111100100",
  45935=>"001000000",
  45936=>"000011000",
  45937=>"000000000",
  45938=>"111111111",
  45939=>"111111110",
  45940=>"000111111",
  45941=>"010000010",
  45942=>"100000010",
  45943=>"000001001",
  45944=>"000110111",
  45945=>"111011000",
  45946=>"000000001",
  45947=>"111111111",
  45948=>"111111111",
  45949=>"111110110",
  45950=>"100000000",
  45951=>"000000111",
  45952=>"011111001",
  45953=>"111111111",
  45954=>"001011001",
  45955=>"000000000",
  45956=>"000000000",
  45957=>"000111000",
  45958=>"111000111",
  45959=>"011000011",
  45960=>"111000000",
  45961=>"111101001",
  45962=>"111101101",
  45963=>"000000011",
  45964=>"011011011",
  45965=>"100111000",
  45966=>"111111111",
  45967=>"000000111",
  45968=>"000000000",
  45969=>"000000000",
  45970=>"000100110",
  45971=>"000000000",
  45972=>"111110000",
  45973=>"000110110",
  45974=>"111110000",
  45975=>"000111000",
  45976=>"000000111",
  45977=>"000011010",
  45978=>"111111010",
  45979=>"000000010",
  45980=>"000000111",
  45981=>"111010000",
  45982=>"000000010",
  45983=>"111111111",
  45984=>"111111111",
  45985=>"010010000",
  45986=>"101000000",
  45987=>"000000111",
  45988=>"101111000",
  45989=>"011011000",
  45990=>"001000000",
  45991=>"010000000",
  45992=>"000010000",
  45993=>"000011001",
  45994=>"110000000",
  45995=>"000010000",
  45996=>"111111111",
  45997=>"011110111",
  45998=>"000101111",
  45999=>"001111000",
  46000=>"111001001",
  46001=>"000110100",
  46002=>"000000000",
  46003=>"000000000",
  46004=>"000111011",
  46005=>"001000000",
  46006=>"000000000",
  46007=>"110110000",
  46008=>"111110000",
  46009=>"011000000",
  46010=>"000000000",
  46011=>"111110000",
  46012=>"000110100",
  46013=>"110111010",
  46014=>"001001001",
  46015=>"111111100",
  46016=>"111011000",
  46017=>"101111111",
  46018=>"000000111",
  46019=>"000100000",
  46020=>"101110010",
  46021=>"000000000",
  46022=>"110111100",
  46023=>"111111101",
  46024=>"111111111",
  46025=>"000000000",
  46026=>"000000000",
  46027=>"111111111",
  46028=>"000000000",
  46029=>"001111111",
  46030=>"101000000",
  46031=>"000110011",
  46032=>"000010000",
  46033=>"000001001",
  46034=>"111000000",
  46035=>"011000000",
  46036=>"100000000",
  46037=>"101101000",
  46038=>"111000100",
  46039=>"000000100",
  46040=>"000000111",
  46041=>"110111111",
  46042=>"000000000",
  46043=>"011000000",
  46044=>"000000000",
  46045=>"111111011",
  46046=>"111111000",
  46047=>"110110100",
  46048=>"111011001",
  46049=>"111111111",
  46050=>"111111111",
  46051=>"111111001",
  46052=>"111111111",
  46053=>"000111111",
  46054=>"000011111",
  46055=>"111111111",
  46056=>"010000000",
  46057=>"111111111",
  46058=>"111111010",
  46059=>"010111111",
  46060=>"000001001",
  46061=>"111111110",
  46062=>"000000000",
  46063=>"000100110",
  46064=>"100000100",
  46065=>"111111111",
  46066=>"001001011",
  46067=>"000000000",
  46068=>"111111111",
  46069=>"000000000",
  46070=>"001011010",
  46071=>"000001111",
  46072=>"000010000",
  46073=>"111111110",
  46074=>"011001000",
  46075=>"111101111",
  46076=>"000011000",
  46077=>"000000000",
  46078=>"000000110",
  46079=>"000011111",
  46080=>"110110110",
  46081=>"111110000",
  46082=>"101000000",
  46083=>"000000000",
  46084=>"000000000",
  46085=>"000000000",
  46086=>"000000000",
  46087=>"111111101",
  46088=>"110111111",
  46089=>"000000001",
  46090=>"010000000",
  46091=>"000000110",
  46092=>"000000000",
  46093=>"111011000",
  46094=>"000000000",
  46095=>"000000110",
  46096=>"111000000",
  46097=>"000100000",
  46098=>"110110000",
  46099=>"000000000",
  46100=>"000010000",
  46101=>"000000000",
  46102=>"000100111",
  46103=>"100000000",
  46104=>"000000000",
  46105=>"101001101",
  46106=>"111111111",
  46107=>"001011011",
  46108=>"111111111",
  46109=>"000110000",
  46110=>"111111111",
  46111=>"001011111",
  46112=>"000010111",
  46113=>"111111111",
  46114=>"000000000",
  46115=>"011011111",
  46116=>"000110111",
  46117=>"100000000",
  46118=>"000110111",
  46119=>"000000111",
  46120=>"100010001",
  46121=>"000111111",
  46122=>"001000000",
  46123=>"001000000",
  46124=>"000000110",
  46125=>"000000000",
  46126=>"111111111",
  46127=>"111111111",
  46128=>"111111000",
  46129=>"000000000",
  46130=>"100000001",
  46131=>"111111111",
  46132=>"111101111",
  46133=>"000100110",
  46134=>"110011111",
  46135=>"000000100",
  46136=>"111111111",
  46137=>"011011001",
  46138=>"000000000",
  46139=>"111111111",
  46140=>"000000111",
  46141=>"000000000",
  46142=>"000010101",
  46143=>"000000000",
  46144=>"011111011",
  46145=>"111111111",
  46146=>"111110110",
  46147=>"000011111",
  46148=>"110111110",
  46149=>"111110110",
  46150=>"111111000",
  46151=>"111000000",
  46152=>"111111111",
  46153=>"111000000",
  46154=>"010000100",
  46155=>"110111110",
  46156=>"111111111",
  46157=>"000000000",
  46158=>"001000000",
  46159=>"011000000",
  46160=>"011011111",
  46161=>"000000000",
  46162=>"000100111",
  46163=>"111111111",
  46164=>"000000110",
  46165=>"100000000",
  46166=>"001001111",
  46167=>"010111111",
  46168=>"000000000",
  46169=>"111111111",
  46170=>"000000111",
  46171=>"000000000",
  46172=>"000000101",
  46173=>"000000000",
  46174=>"011111000",
  46175=>"110110111",
  46176=>"100110110",
  46177=>"000000000",
  46178=>"111111111",
  46179=>"000000000",
  46180=>"000000000",
  46181=>"000000010",
  46182=>"000000000",
  46183=>"101100101",
  46184=>"000000000",
  46185=>"001001000",
  46186=>"111111111",
  46187=>"111111000",
  46188=>"000000100",
  46189=>"111111111",
  46190=>"111111011",
  46191=>"000000000",
  46192=>"010110110",
  46193=>"000011111",
  46194=>"100111111",
  46195=>"000000000",
  46196=>"100000000",
  46197=>"000000100",
  46198=>"000000000",
  46199=>"100111110",
  46200=>"000000000",
  46201=>"000001000",
  46202=>"100110111",
  46203=>"000000000",
  46204=>"001001000",
  46205=>"111111111",
  46206=>"100000000",
  46207=>"000000000",
  46208=>"111111111",
  46209=>"010111111",
  46210=>"110110111",
  46211=>"010110110",
  46212=>"111111111",
  46213=>"001001111",
  46214=>"111111111",
  46215=>"000010010",
  46216=>"111111110",
  46217=>"011000000",
  46218=>"000010110",
  46219=>"000000001",
  46220=>"000010110",
  46221=>"111111111",
  46222=>"100111111",
  46223=>"111111111",
  46224=>"011111110",
  46225=>"100110110",
  46226=>"111111111",
  46227=>"111111110",
  46228=>"000100110",
  46229=>"000000000",
  46230=>"111111111",
  46231=>"000111111",
  46232=>"000110111",
  46233=>"111101111",
  46234=>"000000101",
  46235=>"101111110",
  46236=>"000000011",
  46237=>"010010010",
  46238=>"100000111",
  46239=>"111111111",
  46240=>"111111111",
  46241=>"110111011",
  46242=>"101000000",
  46243=>"111111111",
  46244=>"000000110",
  46245=>"111000000",
  46246=>"000000000",
  46247=>"100111111",
  46248=>"111111111",
  46249=>"110111111",
  46250=>"011000000",
  46251=>"000000000",
  46252=>"000000001",
  46253=>"111111111",
  46254=>"001000101",
  46255=>"110110110",
  46256=>"000000111",
  46257=>"110110110",
  46258=>"111111111",
  46259=>"000000000",
  46260=>"111100000",
  46261=>"000010000",
  46262=>"000110111",
  46263=>"111111111",
  46264=>"111111111",
  46265=>"000110000",
  46266=>"000000100",
  46267=>"000010111",
  46268=>"111001001",
  46269=>"111111111",
  46270=>"000000000",
  46271=>"000010110",
  46272=>"000000000",
  46273=>"000000111",
  46274=>"000110100",
  46275=>"110110010",
  46276=>"111111111",
  46277=>"011000000",
  46278=>"011110111",
  46279=>"000000000",
  46280=>"110110111",
  46281=>"110000000",
  46282=>"110010000",
  46283=>"000000000",
  46284=>"100000000",
  46285=>"000000000",
  46286=>"110000000",
  46287=>"110111001",
  46288=>"111111111",
  46289=>"101000000",
  46290=>"000110000",
  46291=>"000010000",
  46292=>"100000000",
  46293=>"001011011",
  46294=>"010000000",
  46295=>"010000000",
  46296=>"000000000",
  46297=>"110111001",
  46298=>"000001001",
  46299=>"000000000",
  46300=>"111111111",
  46301=>"000000000",
  46302=>"000000000",
  46303=>"110011011",
  46304=>"000000000",
  46305=>"001111000",
  46306=>"100000111",
  46307=>"000000000",
  46308=>"100000000",
  46309=>"100100100",
  46310=>"000000001",
  46311=>"000111111",
  46312=>"111111111",
  46313=>"100100111",
  46314=>"000110111",
  46315=>"110010000",
  46316=>"000000000",
  46317=>"111111111",
  46318=>"010010011",
  46319=>"111111110",
  46320=>"111111111",
  46321=>"111111111",
  46322=>"110110111",
  46323=>"000000110",
  46324=>"111111111",
  46325=>"111111111",
  46326=>"111011111",
  46327=>"111100111",
  46328=>"010000000",
  46329=>"100000000",
  46330=>"000000000",
  46331=>"000000000",
  46332=>"111100110",
  46333=>"111000110",
  46334=>"000001111",
  46335=>"100100100",
  46336=>"110111111",
  46337=>"000100100",
  46338=>"111111111",
  46339=>"001011001",
  46340=>"111111111",
  46341=>"000000100",
  46342=>"111111100",
  46343=>"011011100",
  46344=>"000000000",
  46345=>"111000000",
  46346=>"111110111",
  46347=>"000001000",
  46348=>"111111111",
  46349=>"100110111",
  46350=>"000000000",
  46351=>"101110111",
  46352=>"111111000",
  46353=>"110111000",
  46354=>"000000000",
  46355=>"000000111",
  46356=>"111111010",
  46357=>"000000011",
  46358=>"101101101",
  46359=>"110111000",
  46360=>"110111111",
  46361=>"111111111",
  46362=>"111011000",
  46363=>"110110100",
  46364=>"001001111",
  46365=>"111111000",
  46366=>"111111111",
  46367=>"110110000",
  46368=>"111011001",
  46369=>"100000000",
  46370=>"001011011",
  46371=>"000000001",
  46372=>"011011001",
  46373=>"111111111",
  46374=>"111111100",
  46375=>"111111111",
  46376=>"111111111",
  46377=>"111111111",
  46378=>"000110011",
  46379=>"001111111",
  46380=>"000000000",
  46381=>"110111111",
  46382=>"000000000",
  46383=>"000000100",
  46384=>"000000000",
  46385=>"110110111",
  46386=>"111111011",
  46387=>"111111111",
  46388=>"000000000",
  46389=>"000000111",
  46390=>"000000000",
  46391=>"010110110",
  46392=>"000000000",
  46393=>"000100000",
  46394=>"000000100",
  46395=>"111111111",
  46396=>"111000100",
  46397=>"000000010",
  46398=>"111111111",
  46399=>"000010110",
  46400=>"000000110",
  46401=>"111110110",
  46402=>"001111111",
  46403=>"000000001",
  46404=>"001000000",
  46405=>"010011000",
  46406=>"111111000",
  46407=>"110110100",
  46408=>"000001001",
  46409=>"100111010",
  46410=>"100111011",
  46411=>"000110110",
  46412=>"111111111",
  46413=>"100111111",
  46414=>"010011000",
  46415=>"111111111",
  46416=>"100111111",
  46417=>"111111101",
  46418=>"111110110",
  46419=>"000000000",
  46420=>"000000000",
  46421=>"001000000",
  46422=>"000000000",
  46423=>"100110111",
  46424=>"000000000",
  46425=>"000000000",
  46426=>"111111011",
  46427=>"111111111",
  46428=>"011111110",
  46429=>"111111000",
  46430=>"111011111",
  46431=>"000111111",
  46432=>"100000000",
  46433=>"000000000",
  46434=>"100101100",
  46435=>"000000000",
  46436=>"110110100",
  46437=>"000111000",
  46438=>"000000001",
  46439=>"100000111",
  46440=>"000100110",
  46441=>"100101111",
  46442=>"111111010",
  46443=>"110100000",
  46444=>"000100000",
  46445=>"000011111",
  46446=>"000110010",
  46447=>"011001000",
  46448=>"011000000",
  46449=>"100100111",
  46450=>"000000110",
  46451=>"001001001",
  46452=>"100110110",
  46453=>"111111111",
  46454=>"000000111",
  46455=>"000000000",
  46456=>"111111110",
  46457=>"000000000",
  46458=>"000000000",
  46459=>"111110110",
  46460=>"011111111",
  46461=>"011000000",
  46462=>"000000011",
  46463=>"111111101",
  46464=>"000111111",
  46465=>"110100100",
  46466=>"100000000",
  46467=>"000000000",
  46468=>"000000000",
  46469=>"111111111",
  46470=>"111011100",
  46471=>"111111111",
  46472=>"010010010",
  46473=>"000000000",
  46474=>"111111111",
  46475=>"011001001",
  46476=>"000000000",
  46477=>"001101111",
  46478=>"100000001",
  46479=>"110000000",
  46480=>"010000000",
  46481=>"000000000",
  46482=>"000111111",
  46483=>"000000001",
  46484=>"000000000",
  46485=>"000000000",
  46486=>"111001000",
  46487=>"000000000",
  46488=>"000000000",
  46489=>"111010010",
  46490=>"101001001",
  46491=>"111111001",
  46492=>"111110100",
  46493=>"000000110",
  46494=>"011000000",
  46495=>"000000000",
  46496=>"110110000",
  46497=>"101111110",
  46498=>"000100101",
  46499=>"111111111",
  46500=>"111111111",
  46501=>"000011000",
  46502=>"000000100",
  46503=>"111000000",
  46504=>"100100000",
  46505=>"010111111",
  46506=>"111111111",
  46507=>"000000000",
  46508=>"000000000",
  46509=>"111111011",
  46510=>"110111111",
  46511=>"111101000",
  46512=>"111111000",
  46513=>"000000000",
  46514=>"000101000",
  46515=>"100000000",
  46516=>"111111111",
  46517=>"011110111",
  46518=>"011111111",
  46519=>"111110111",
  46520=>"111111111",
  46521=>"111111011",
  46522=>"111111111",
  46523=>"000000001",
  46524=>"000000000",
  46525=>"111111111",
  46526=>"000000000",
  46527=>"100111111",
  46528=>"000001000",
  46529=>"111111000",
  46530=>"000000000",
  46531=>"111111111",
  46532=>"000000000",
  46533=>"000100100",
  46534=>"000000000",
  46535=>"000000000",
  46536=>"000010111",
  46537=>"111111111",
  46538=>"000000100",
  46539=>"110110111",
  46540=>"111111100",
  46541=>"001000000",
  46542=>"111001100",
  46543=>"111011001",
  46544=>"001011111",
  46545=>"111111111",
  46546=>"000000000",
  46547=>"000000000",
  46548=>"111100100",
  46549=>"100000000",
  46550=>"001111000",
  46551=>"001001001",
  46552=>"000000100",
  46553=>"000100101",
  46554=>"000000110",
  46555=>"111011111",
  46556=>"000000000",
  46557=>"000000000",
  46558=>"000000000",
  46559=>"111111111",
  46560=>"110111111",
  46561=>"000000100",
  46562=>"111111111",
  46563=>"000000000",
  46564=>"011011110",
  46565=>"111101111",
  46566=>"011011010",
  46567=>"000000000",
  46568=>"000000000",
  46569=>"100110110",
  46570=>"000000000",
  46571=>"111111111",
  46572=>"000000000",
  46573=>"111111111",
  46574=>"111111111",
  46575=>"001011111",
  46576=>"110111111",
  46577=>"110000100",
  46578=>"000000111",
  46579=>"000011011",
  46580=>"000000000",
  46581=>"100000000",
  46582=>"111111111",
  46583=>"011011000",
  46584=>"111111111",
  46585=>"100000000",
  46586=>"000110110",
  46587=>"000010000",
  46588=>"000000000",
  46589=>"111111111",
  46590=>"000000000",
  46591=>"000000000",
  46592=>"111101111",
  46593=>"000000000",
  46594=>"100100101",
  46595=>"101000110",
  46596=>"000011111",
  46597=>"110110110",
  46598=>"001101111",
  46599=>"111111111",
  46600=>"111101101",
  46601=>"000011111",
  46602=>"010110110",
  46603=>"110110110",
  46604=>"001000110",
  46605=>"100111111",
  46606=>"110001001",
  46607=>"001001001",
  46608=>"111111111",
  46609=>"000000111",
  46610=>"111111101",
  46611=>"110110010",
  46612=>"111011101",
  46613=>"111000001",
  46614=>"000000000",
  46615=>"010011011",
  46616=>"000000000",
  46617=>"100011110",
  46618=>"000001000",
  46619=>"010110111",
  46620=>"110110000",
  46621=>"111000000",
  46622=>"011011011",
  46623=>"111111110",
  46624=>"100000000",
  46625=>"000000110",
  46626=>"000110111",
  46627=>"001111001",
  46628=>"101000000",
  46629=>"111001011",
  46630=>"000000001",
  46631=>"110000000",
  46632=>"001000001",
  46633=>"001111111",
  46634=>"000000000",
  46635=>"011011010",
  46636=>"010111011",
  46637=>"000001110",
  46638=>"000110100",
  46639=>"101000000",
  46640=>"010111111",
  46641=>"111111111",
  46642=>"000001000",
  46643=>"011010010",
  46644=>"000000001",
  46645=>"001001001",
  46646=>"111001011",
  46647=>"000000000",
  46648=>"110110000",
  46649=>"011001101",
  46650=>"011111011",
  46651=>"010000000",
  46652=>"111110110",
  46653=>"000000111",
  46654=>"011001101",
  46655=>"110000000",
  46656=>"111110110",
  46657=>"000000000",
  46658=>"110110111",
  46659=>"000000000",
  46660=>"000000000",
  46661=>"000000001",
  46662=>"000000000",
  46663=>"100000111",
  46664=>"011011000",
  46665=>"111101101",
  46666=>"101111111",
  46667=>"000001001",
  46668=>"110110010",
  46669=>"111011111",
  46670=>"011010010",
  46671=>"011111110",
  46672=>"000000000",
  46673=>"111111000",
  46674=>"111111001",
  46675=>"000000100",
  46676=>"110000000",
  46677=>"001001001",
  46678=>"100000001",
  46679=>"101101101",
  46680=>"001001001",
  46681=>"101100101",
  46682=>"111111111",
  46683=>"100100110",
  46684=>"000000001",
  46685=>"001011111",
  46686=>"111111111",
  46687=>"111001000",
  46688=>"101101101",
  46689=>"010010010",
  46690=>"111111101",
  46691=>"000000000",
  46692=>"110110110",
  46693=>"101001111",
  46694=>"110100000",
  46695=>"111111111",
  46696=>"111111111",
  46697=>"111000000",
  46698=>"001000000",
  46699=>"011111111",
  46700=>"100101101",
  46701=>"000000000",
  46702=>"001010000",
  46703=>"001101111",
  46704=>"110011111",
  46705=>"100001111",
  46706=>"010110111",
  46707=>"111010000",
  46708=>"110000000",
  46709=>"011010010",
  46710=>"000000000",
  46711=>"001111111",
  46712=>"111101101",
  46713=>"100000000",
  46714=>"000000000",
  46715=>"010010000",
  46716=>"100110110",
  46717=>"000110111",
  46718=>"000000110",
  46719=>"000001000",
  46720=>"000000101",
  46721=>"111111111",
  46722=>"111111111",
  46723=>"100101101",
  46724=>"100111111",
  46725=>"111111111",
  46726=>"100000010",
  46727=>"010010010",
  46728=>"110000000",
  46729=>"000000010",
  46730=>"110111010",
  46731=>"100000100",
  46732=>"110111111",
  46733=>"000110110",
  46734=>"000000000",
  46735=>"111001001",
  46736=>"001101001",
  46737=>"000000001",
  46738=>"000000000",
  46739=>"000100100",
  46740=>"111111111",
  46741=>"001000000",
  46742=>"111111111",
  46743=>"111111111",
  46744=>"000001001",
  46745=>"101000000",
  46746=>"111111111",
  46747=>"000000011",
  46748=>"000000000",
  46749=>"000000000",
  46750=>"110111111",
  46751=>"000000000",
  46752=>"111101101",
  46753=>"000000000",
  46754=>"101101111",
  46755=>"111111111",
  46756=>"001001000",
  46757=>"101011100",
  46758=>"001000000",
  46759=>"011011111",
  46760=>"101101101",
  46761=>"000000000",
  46762=>"101000101",
  46763=>"110110000",
  46764=>"000000000",
  46765=>"001000100",
  46766=>"001001111",
  46767=>"000000000",
  46768=>"010010000",
  46769=>"011011011",
  46770=>"001111011",
  46771=>"111000000",
  46772=>"111001000",
  46773=>"000110111",
  46774=>"001001111",
  46775=>"000000000",
  46776=>"000001001",
  46777=>"011001001",
  46778=>"001001101",
  46779=>"001001111",
  46780=>"111011001",
  46781=>"011000000",
  46782=>"000001111",
  46783=>"001001001",
  46784=>"010000000",
  46785=>"100110100",
  46786=>"110110100",
  46787=>"000010110",
  46788=>"111111101",
  46789=>"000000000",
  46790=>"111110000",
  46791=>"101111001",
  46792=>"111111111",
  46793=>"110110010",
  46794=>"010110010",
  46795=>"101111111",
  46796=>"111000000",
  46797=>"000001111",
  46798=>"101000000",
  46799=>"001000011",
  46800=>"000000110",
  46801=>"000000111",
  46802=>"000000000",
  46803=>"000000000",
  46804=>"001000101",
  46805=>"000000000",
  46806=>"111111111",
  46807=>"001101111",
  46808=>"111111111",
  46809=>"010100000",
  46810=>"001000000",
  46811=>"011010010",
  46812=>"010110100",
  46813=>"000000000",
  46814=>"000111111",
  46815=>"000000000",
  46816=>"111101000",
  46817=>"011111111",
  46818=>"111101110",
  46819=>"001000001",
  46820=>"110110010",
  46821=>"001001000",
  46822=>"011010110",
  46823=>"000000001",
  46824=>"011111110",
  46825=>"011001001",
  46826=>"011011101",
  46827=>"111111000",
  46828=>"100100001",
  46829=>"111101101",
  46830=>"000010110",
  46831=>"000000000",
  46832=>"111100111",
  46833=>"000000100",
  46834=>"111111011",
  46835=>"101101111",
  46836=>"000000110",
  46837=>"111001000",
  46838=>"001001011",
  46839=>"010111011",
  46840=>"111111110",
  46841=>"100101000",
  46842=>"111110111",
  46843=>"000010110",
  46844=>"100110111",
  46845=>"110110110",
  46846=>"111001011",
  46847=>"001011011",
  46848=>"000000000",
  46849=>"001000001",
  46850=>"111111101",
  46851=>"010110010",
  46852=>"111111011",
  46853=>"000000000",
  46854=>"000000000",
  46855=>"101001101",
  46856=>"000000011",
  46857=>"100000000",
  46858=>"000111110",
  46859=>"001011001",
  46860=>"011000000",
  46861=>"110000101",
  46862=>"001111111",
  46863=>"110110000",
  46864=>"111111001",
  46865=>"000000001",
  46866=>"110000000",
  46867=>"010110110",
  46868=>"111001000",
  46869=>"101001000",
  46870=>"000000000",
  46871=>"000001001",
  46872=>"000000000",
  46873=>"000000100",
  46874=>"001001001",
  46875=>"000000110",
  46876=>"000000000",
  46877=>"111010011",
  46878=>"000000000",
  46879=>"000000000",
  46880=>"010010010",
  46881=>"001001101",
  46882=>"011011010",
  46883=>"101111111",
  46884=>"001100000",
  46885=>"011111111",
  46886=>"100100101",
  46887=>"110111111",
  46888=>"001001001",
  46889=>"111111111",
  46890=>"111010001",
  46891=>"001000000",
  46892=>"110100000",
  46893=>"110110111",
  46894=>"000110010",
  46895=>"001000000",
  46896=>"110110110",
  46897=>"010000000",
  46898=>"011000000",
  46899=>"110110100",
  46900=>"111111111",
  46901=>"100111111",
  46902=>"101101001",
  46903=>"111111111",
  46904=>"101101100",
  46905=>"001000000",
  46906=>"000000000",
  46907=>"111001001",
  46908=>"000001001",
  46909=>"000110110",
  46910=>"000000001",
  46911=>"111100100",
  46912=>"000111111",
  46913=>"111000000",
  46914=>"000000000",
  46915=>"101101101",
  46916=>"111001000",
  46917=>"111111111",
  46918=>"101111111",
  46919=>"001001001",
  46920=>"001000010",
  46921=>"000000010",
  46922=>"101001001",
  46923=>"101100100",
  46924=>"000010010",
  46925=>"001101110",
  46926=>"111011010",
  46927=>"110111111",
  46928=>"100110110",
  46929=>"101001111",
  46930=>"100110000",
  46931=>"001001101",
  46932=>"001001000",
  46933=>"001001001",
  46934=>"111111111",
  46935=>"100000111",
  46936=>"101001011",
  46937=>"000000000",
  46938=>"100111011",
  46939=>"000000000",
  46940=>"011001000",
  46941=>"000100111",
  46942=>"111111110",
  46943=>"111111011",
  46944=>"100000001",
  46945=>"111111100",
  46946=>"100100000",
  46947=>"101100111",
  46948=>"001001001",
  46949=>"011111111",
  46950=>"000001111",
  46951=>"101000001",
  46952=>"001001001",
  46953=>"111101101",
  46954=>"000000000",
  46955=>"110110110",
  46956=>"100100100",
  46957=>"000000000",
  46958=>"000001000",
  46959=>"111110010",
  46960=>"000001101",
  46961=>"000000010",
  46962=>"111001011",
  46963=>"101111111",
  46964=>"000000000",
  46965=>"000001000",
  46966=>"111111011",
  46967=>"000000111",
  46968=>"101101101",
  46969=>"010010010",
  46970=>"111100100",
  46971=>"011001001",
  46972=>"010110000",
  46973=>"001001001",
  46974=>"000001000",
  46975=>"000000000",
  46976=>"001001000",
  46977=>"001001001",
  46978=>"100000100",
  46979=>"000111011",
  46980=>"101101111",
  46981=>"010010010",
  46982=>"100000001",
  46983=>"100111111",
  46984=>"000000100",
  46985=>"110110101",
  46986=>"111110010",
  46987=>"010110110",
  46988=>"000001111",
  46989=>"111111110",
  46990=>"010111011",
  46991=>"111111111",
  46992=>"000000000",
  46993=>"011111111",
  46994=>"101000111",
  46995=>"001000000",
  46996=>"000010010",
  46997=>"010000000",
  46998=>"001001001",
  46999=>"101111111",
  47000=>"011011111",
  47001=>"000000100",
  47002=>"000010010",
  47003=>"000010110",
  47004=>"101101111",
  47005=>"000010010",
  47006=>"111001101",
  47007=>"000000000",
  47008=>"111100111",
  47009=>"111111110",
  47010=>"111101101",
  47011=>"101101001",
  47012=>"000001111",
  47013=>"110101000",
  47014=>"101001000",
  47015=>"110110110",
  47016=>"001000000",
  47017=>"111011011",
  47018=>"111011000",
  47019=>"111101111",
  47020=>"000000001",
  47021=>"111101001",
  47022=>"001000000",
  47023=>"000011011",
  47024=>"000000000",
  47025=>"000000000",
  47026=>"111111101",
  47027=>"111111101",
  47028=>"001111111",
  47029=>"110110110",
  47030=>"111111110",
  47031=>"010110110",
  47032=>"110000010",
  47033=>"010010110",
  47034=>"011000000",
  47035=>"101101111",
  47036=>"000100100",
  47037=>"000001010",
  47038=>"101000110",
  47039=>"111111110",
  47040=>"010110010",
  47041=>"000000000",
  47042=>"111010010",
  47043=>"001111111",
  47044=>"110110010",
  47045=>"011000000",
  47046=>"101001001",
  47047=>"000001111",
  47048=>"001101101",
  47049=>"110110000",
  47050=>"000000000",
  47051=>"111111011",
  47052=>"010111111",
  47053=>"000000000",
  47054=>"000001000",
  47055=>"101011000",
  47056=>"111000101",
  47057=>"101100101",
  47058=>"011111111",
  47059=>"011011011",
  47060=>"111101000",
  47061=>"111111000",
  47062=>"111011010",
  47063=>"100100111",
  47064=>"111111011",
  47065=>"110110000",
  47066=>"000011001",
  47067=>"001100101",
  47068=>"111111111",
  47069=>"001001001",
  47070=>"100001101",
  47071=>"000001001",
  47072=>"111011011",
  47073=>"000000000",
  47074=>"000000100",
  47075=>"100101111",
  47076=>"001111111",
  47077=>"111011011",
  47078=>"110110010",
  47079=>"101101101",
  47080=>"110110110",
  47081=>"000000011",
  47082=>"000000111",
  47083=>"110110111",
  47084=>"001000001",
  47085=>"010110110",
  47086=>"000111111",
  47087=>"111000000",
  47088=>"000000101",
  47089=>"111101101",
  47090=>"010111011",
  47091=>"001001001",
  47092=>"001001011",
  47093=>"000000100",
  47094=>"111110001",
  47095=>"011011001",
  47096=>"010010000",
  47097=>"000000010",
  47098=>"000010110",
  47099=>"101101000",
  47100=>"110110000",
  47101=>"111001111",
  47102=>"011000000",
  47103=>"000000111",
  47104=>"111111000",
  47105=>"000000110",
  47106=>"001000001",
  47107=>"000011011",
  47108=>"111111011",
  47109=>"111000000",
  47110=>"111111111",
  47111=>"101111111",
  47112=>"011010111",
  47113=>"000000100",
  47114=>"100000001",
  47115=>"100000000",
  47116=>"111110110",
  47117=>"111000000",
  47118=>"111101011",
  47119=>"111000000",
  47120=>"001000000",
  47121=>"111111111",
  47122=>"111111111",
  47123=>"000000000",
  47124=>"000000100",
  47125=>"000111111",
  47126=>"100000000",
  47127=>"110110000",
  47128=>"111000100",
  47129=>"110100000",
  47130=>"111111111",
  47131=>"011100100",
  47132=>"111101111",
  47133=>"000110111",
  47134=>"101101000",
  47135=>"000100111",
  47136=>"000110110",
  47137=>"111101000",
  47138=>"110111110",
  47139=>"111111011",
  47140=>"000000000",
  47141=>"000000111",
  47142=>"111111111",
  47143=>"000111111",
  47144=>"001000111",
  47145=>"111111101",
  47146=>"111111111",
  47147=>"111110100",
  47148=>"100100000",
  47149=>"000110111",
  47150=>"111100001",
  47151=>"110000001",
  47152=>"100110111",
  47153=>"111111000",
  47154=>"001001000",
  47155=>"011000000",
  47156=>"010110010",
  47157=>"100100100",
  47158=>"111000001",
  47159=>"001000000",
  47160=>"000000001",
  47161=>"110000001",
  47162=>"010011000",
  47163=>"111111111",
  47164=>"100100100",
  47165=>"111111010",
  47166=>"111001000",
  47167=>"111111111",
  47168=>"011000000",
  47169=>"011010010",
  47170=>"111000000",
  47171=>"111111111",
  47172=>"100110111",
  47173=>"111111111",
  47174=>"000000111",
  47175=>"111111111",
  47176=>"000110000",
  47177=>"010111111",
  47178=>"000000000",
  47179=>"111111011",
  47180=>"000000111",
  47181=>"001001000",
  47182=>"100100100",
  47183=>"000110110",
  47184=>"111111111",
  47185=>"000000000",
  47186=>"110111111",
  47187=>"000000110",
  47188=>"000000000",
  47189=>"001111111",
  47190=>"000011111",
  47191=>"000000000",
  47192=>"000000000",
  47193=>"000000101",
  47194=>"000010111",
  47195=>"111010000",
  47196=>"111111111",
  47197=>"000000000",
  47198=>"111111100",
  47199=>"111000011",
  47200=>"000000001",
  47201=>"000110110",
  47202=>"011000000",
  47203=>"111011110",
  47204=>"111000000",
  47205=>"100000100",
  47206=>"110110110",
  47207=>"111000000",
  47208=>"001011111",
  47209=>"001001001",
  47210=>"111111010",
  47211=>"111111111",
  47212=>"011010000",
  47213=>"111111111",
  47214=>"001101111",
  47215=>"111110110",
  47216=>"111111111",
  47217=>"001011011",
  47218=>"100000000",
  47219=>"101100110",
  47220=>"111111011",
  47221=>"111111110",
  47222=>"001011111",
  47223=>"110111010",
  47224=>"000000000",
  47225=>"001001111",
  47226=>"001000000",
  47227=>"111111111",
  47228=>"100100101",
  47229=>"100100011",
  47230=>"011001100",
  47231=>"000011111",
  47232=>"101000000",
  47233=>"100111000",
  47234=>"111111111",
  47235=>"010011101",
  47236=>"001001000",
  47237=>"111101111",
  47238=>"011101111",
  47239=>"001111100",
  47240=>"000110111",
  47241=>"010110101",
  47242=>"011111111",
  47243=>"000000011",
  47244=>"111011111",
  47245=>"000000000",
  47246=>"001001001",
  47247=>"111111111",
  47248=>"101100101",
  47249=>"010110111",
  47250=>"111100000",
  47251=>"111001111",
  47252=>"111001000",
  47253=>"100110110",
  47254=>"111111000",
  47255=>"000000000",
  47256=>"000000000",
  47257=>"100010001",
  47258=>"000000000",
  47259=>"000000101",
  47260=>"101000000",
  47261=>"001000000",
  47262=>"100000001",
  47263=>"010010000",
  47264=>"111111111",
  47265=>"111011111",
  47266=>"111111111",
  47267=>"100111111",
  47268=>"101111001",
  47269=>"111110110",
  47270=>"001000000",
  47271=>"111110100",
  47272=>"000000000",
  47273=>"000000000",
  47274=>"001000000",
  47275=>"100100100",
  47276=>"001001001",
  47277=>"000000000",
  47278=>"000000001",
  47279=>"000000000",
  47280=>"110111111",
  47281=>"111110100",
  47282=>"010111000",
  47283=>"001111000",
  47284=>"111110000",
  47285=>"111111011",
  47286=>"100001000",
  47287=>"000000000",
  47288=>"110101011",
  47289=>"111111010",
  47290=>"000000000",
  47291=>"111110000",
  47292=>"000100110",
  47293=>"000000000",
  47294=>"111111111",
  47295=>"101111110",
  47296=>"101001000",
  47297=>"111111111",
  47298=>"100000000",
  47299=>"111111010",
  47300=>"000000000",
  47301=>"000111111",
  47302=>"000000000",
  47303=>"111111011",
  47304=>"000000000",
  47305=>"000110111",
  47306=>"001001101",
  47307=>"111111111",
  47308=>"000000110",
  47309=>"100100100",
  47310=>"111100000",
  47311=>"010100100",
  47312=>"111111111",
  47313=>"111001111",
  47314=>"100000100",
  47315=>"001000000",
  47316=>"110111000",
  47317=>"000000000",
  47318=>"000000000",
  47319=>"111010000",
  47320=>"111111100",
  47321=>"111111010",
  47322=>"111111111",
  47323=>"100110010",
  47324=>"000000000",
  47325=>"100101111",
  47326=>"000000000",
  47327=>"111111000",
  47328=>"001001011",
  47329=>"000000000",
  47330=>"000110110",
  47331=>"110010000",
  47332=>"101111111",
  47333=>"100000000",
  47334=>"110010010",
  47335=>"000000011",
  47336=>"000000111",
  47337=>"111111111",
  47338=>"111111111",
  47339=>"111110111",
  47340=>"000000111",
  47341=>"100111011",
  47342=>"111111101",
  47343=>"000111111",
  47344=>"111001000",
  47345=>"110110100",
  47346=>"001000000",
  47347=>"000000000",
  47348=>"001000001",
  47349=>"111111100",
  47350=>"100100100",
  47351=>"110000111",
  47352=>"000010111",
  47353=>"000000000",
  47354=>"000110000",
  47355=>"111000000",
  47356=>"111110011",
  47357=>"001000000",
  47358=>"111010000",
  47359=>"111110010",
  47360=>"011111010",
  47361=>"100000000",
  47362=>"010010111",
  47363=>"111111110",
  47364=>"000000000",
  47365=>"000000000",
  47366=>"011011011",
  47367=>"000001001",
  47368=>"010000000",
  47369=>"100110111",
  47370=>"101101101",
  47371=>"111111010",
  47372=>"100000100",
  47373=>"000111111",
  47374=>"111111111",
  47375=>"010110000",
  47376=>"000000000",
  47377=>"111100111",
  47378=>"000000000",
  47379=>"001011001",
  47380=>"001000111",
  47381=>"111100111",
  47382=>"111111111",
  47383=>"011111110",
  47384=>"111111111",
  47385=>"111111001",
  47386=>"000000100",
  47387=>"111111010",
  47388=>"110100100",
  47389=>"000000110",
  47390=>"111101000",
  47391=>"011011111",
  47392=>"101101111",
  47393=>"110111011",
  47394=>"010010000",
  47395=>"000000110",
  47396=>"001001111",
  47397=>"111100111",
  47398=>"000111111",
  47399=>"110000011",
  47400=>"110111111",
  47401=>"110100000",
  47402=>"000000000",
  47403=>"000000000",
  47404=>"000000000",
  47405=>"111110000",
  47406=>"111100111",
  47407=>"000000110",
  47408=>"001101000",
  47409=>"000000000",
  47410=>"111111111",
  47411=>"111111000",
  47412=>"110000000",
  47413=>"110111111",
  47414=>"001101100",
  47415=>"001000000",
  47416=>"000110000",
  47417=>"001000001",
  47418=>"111111111",
  47419=>"110110000",
  47420=>"001001001",
  47421=>"000000110",
  47422=>"111111111",
  47423=>"111110111",
  47424=>"111001001",
  47425=>"000110110",
  47426=>"000001001",
  47427=>"000000110",
  47428=>"000000110",
  47429=>"000100100",
  47430=>"101001000",
  47431=>"000000000",
  47432=>"000000000",
  47433=>"001000000",
  47434=>"011011111",
  47435=>"101111111",
  47436=>"111000101",
  47437=>"000011011",
  47438=>"100000100",
  47439=>"000010110",
  47440=>"000000011",
  47441=>"000111111",
  47442=>"111111111",
  47443=>"000000000",
  47444=>"000111111",
  47445=>"011011011",
  47446=>"100000000",
  47447=>"111110100",
  47448=>"111111111",
  47449=>"000000111",
  47450=>"000000000",
  47451=>"000000001",
  47452=>"100000001",
  47453=>"010111011",
  47454=>"000110111",
  47455=>"000000000",
  47456=>"100001111",
  47457=>"111100000",
  47458=>"001000001",
  47459=>"100000101",
  47460=>"011000000",
  47461=>"000000000",
  47462=>"000000000",
  47463=>"000111110",
  47464=>"001001001",
  47465=>"110100101",
  47466=>"111000111",
  47467=>"000000011",
  47468=>"000000000",
  47469=>"111110000",
  47470=>"111110000",
  47471=>"111000111",
  47472=>"100100111",
  47473=>"111111110",
  47474=>"000000000",
  47475=>"111111111",
  47476=>"001011000",
  47477=>"111111111",
  47478=>"000000000",
  47479=>"000000100",
  47480=>"111000001",
  47481=>"001100111",
  47482=>"000000000",
  47483=>"100100100",
  47484=>"001000011",
  47485=>"100110100",
  47486=>"111100000",
  47487=>"000001101",
  47488=>"000100110",
  47489=>"111111111",
  47490=>"111111110",
  47491=>"000000010",
  47492=>"000000111",
  47493=>"000110111",
  47494=>"111011111",
  47495=>"111000000",
  47496=>"000000111",
  47497=>"000000110",
  47498=>"000000111",
  47499=>"000011011",
  47500=>"000100111",
  47501=>"000110110",
  47502=>"000000000",
  47503=>"100111011",
  47504=>"100100101",
  47505=>"000000100",
  47506=>"100000000",
  47507=>"000010011",
  47508=>"111111111",
  47509=>"000000000",
  47510=>"001001001",
  47511=>"110110000",
  47512=>"111111111",
  47513=>"111111111",
  47514=>"101000000",
  47515=>"000000101",
  47516=>"000110100",
  47517=>"111111110",
  47518=>"100000000",
  47519=>"110111110",
  47520=>"111101010",
  47521=>"100110111",
  47522=>"010110010",
  47523=>"001111101",
  47524=>"000000101",
  47525=>"110111111",
  47526=>"100000101",
  47527=>"000000000",
  47528=>"000011011",
  47529=>"000000000",
  47530=>"011000111",
  47531=>"000010011",
  47532=>"100110111",
  47533=>"111000000",
  47534=>"000111111",
  47535=>"111001111",
  47536=>"111101111",
  47537=>"110100100",
  47538=>"110000000",
  47539=>"111111111",
  47540=>"111111111",
  47541=>"110000000",
  47542=>"111111111",
  47543=>"111111110",
  47544=>"101001001",
  47545=>"111111000",
  47546=>"110000000",
  47547=>"100000111",
  47548=>"001000000",
  47549=>"001100000",
  47550=>"101100010",
  47551=>"101100100",
  47552=>"011111110",
  47553=>"000011111",
  47554=>"111111000",
  47555=>"000011111",
  47556=>"010111111",
  47557=>"000000100",
  47558=>"000000000",
  47559=>"111111111",
  47560=>"001000000",
  47561=>"110110010",
  47562=>"000000000",
  47563=>"000000000",
  47564=>"111111110",
  47565=>"111000000",
  47566=>"110000101",
  47567=>"110100111",
  47568=>"111111111",
  47569=>"000100100",
  47570=>"010110111",
  47571=>"000000111",
  47572=>"101100100",
  47573=>"011011001",
  47574=>"000000110",
  47575=>"010010000",
  47576=>"110000000",
  47577=>"000000000",
  47578=>"111100111",
  47579=>"001110000",
  47580=>"111111111",
  47581=>"110110110",
  47582=>"000000111",
  47583=>"111100111",
  47584=>"111111110",
  47585=>"111110110",
  47586=>"111111011",
  47587=>"000001001",
  47588=>"111011000",
  47589=>"101011001",
  47590=>"000000000",
  47591=>"101001101",
  47592=>"010010000",
  47593=>"111111111",
  47594=>"111111000",
  47595=>"111100100",
  47596=>"010110111",
  47597=>"011011010",
  47598=>"010110110",
  47599=>"100000000",
  47600=>"111111110",
  47601=>"111000100",
  47602=>"111111111",
  47603=>"000000000",
  47604=>"101101111",
  47605=>"100110111",
  47606=>"111000000",
  47607=>"001100000",
  47608=>"111001000",
  47609=>"100110010",
  47610=>"111111001",
  47611=>"000000000",
  47612=>"111110111",
  47613=>"111111111",
  47614=>"111111110",
  47615=>"111101111",
  47616=>"111111111",
  47617=>"111000000",
  47618=>"111111111",
  47619=>"110000010",
  47620=>"000000000",
  47621=>"001001011",
  47622=>"001000101",
  47623=>"111111111",
  47624=>"000000000",
  47625=>"100100110",
  47626=>"101001001",
  47627=>"000010110",
  47628=>"000000000",
  47629=>"000000001",
  47630=>"000000000",
  47631=>"000110100",
  47632=>"000000111",
  47633=>"000110111",
  47634=>"111001101",
  47635=>"001000111",
  47636=>"000000000",
  47637=>"000101111",
  47638=>"011000000",
  47639=>"010110110",
  47640=>"111111111",
  47641=>"111111111",
  47642=>"001001101",
  47643=>"010111011",
  47644=>"111001000",
  47645=>"110000000",
  47646=>"000001101",
  47647=>"000101111",
  47648=>"111000000",
  47649=>"111010000",
  47650=>"000000000",
  47651=>"111000000",
  47652=>"110111000",
  47653=>"101000110",
  47654=>"111101111",
  47655=>"111111000",
  47656=>"000001111",
  47657=>"001001101",
  47658=>"001000000",
  47659=>"000000000",
  47660=>"101101111",
  47661=>"111111111",
  47662=>"001001001",
  47663=>"101000000",
  47664=>"000000000",
  47665=>"000000100",
  47666=>"000000000",
  47667=>"000000000",
  47668=>"001100100",
  47669=>"110111111",
  47670=>"111111110",
  47671=>"111111111",
  47672=>"110111111",
  47673=>"001001111",
  47674=>"111111111",
  47675=>"111101111",
  47676=>"010000111",
  47677=>"111000000",
  47678=>"011111011",
  47679=>"000000000",
  47680=>"011010000",
  47681=>"001001000",
  47682=>"000000000",
  47683=>"000000001",
  47684=>"110110110",
  47685=>"111011110",
  47686=>"001110110",
  47687=>"111111111",
  47688=>"111111000",
  47689=>"100000000",
  47690=>"111110110",
  47691=>"011010000",
  47692=>"110110000",
  47693=>"010010010",
  47694=>"111110010",
  47695=>"000000000",
  47696=>"000111011",
  47697=>"001000000",
  47698=>"100001000",
  47699=>"001001011",
  47700=>"000111100",
  47701=>"000000000",
  47702=>"001000111",
  47703=>"110110010",
  47704=>"001000000",
  47705=>"111101111",
  47706=>"111011000",
  47707=>"000001111",
  47708=>"000000011",
  47709=>"011110111",
  47710=>"101000101",
  47711=>"000000000",
  47712=>"100000100",
  47713=>"111101111",
  47714=>"000000000",
  47715=>"000001101",
  47716=>"110110111",
  47717=>"000000000",
  47718=>"110110010",
  47719=>"000000110",
  47720=>"001011111",
  47721=>"101011111",
  47722=>"001000000",
  47723=>"001001100",
  47724=>"011110000",
  47725=>"111000000",
  47726=>"000110110",
  47727=>"111110110",
  47728=>"100101111",
  47729=>"111111111",
  47730=>"100000000",
  47731=>"000010010",
  47732=>"000001001",
  47733=>"001000000",
  47734=>"000000010",
  47735=>"001001001",
  47736=>"111010111",
  47737=>"100000000",
  47738=>"001100101",
  47739=>"000000010",
  47740=>"110110100",
  47741=>"000000000",
  47742=>"000000000",
  47743=>"000000000",
  47744=>"110000000",
  47745=>"111100111",
  47746=>"000000000",
  47747=>"100110111",
  47748=>"000000000",
  47749=>"000000000",
  47750=>"110110000",
  47751=>"010111111",
  47752=>"001000101",
  47753=>"000000000",
  47754=>"000000000",
  47755=>"000000000",
  47756=>"000001001",
  47757=>"110111011",
  47758=>"000000111",
  47759=>"000111000",
  47760=>"010111111",
  47761=>"000001011",
  47762=>"111111111",
  47763=>"001111111",
  47764=>"001001000",
  47765=>"000000111",
  47766=>"000000000",
  47767=>"011000001",
  47768=>"001001100",
  47769=>"111111011",
  47770=>"000000000",
  47771=>"000000111",
  47772=>"011000111",
  47773=>"110000000",
  47774=>"111111010",
  47775=>"101111011",
  47776=>"001001001",
  47777=>"110111111",
  47778=>"111111111",
  47779=>"111010000",
  47780=>"111001001",
  47781=>"000000000",
  47782=>"111111011",
  47783=>"010111011",
  47784=>"000000000",
  47785=>"000000000",
  47786=>"100100101",
  47787=>"110111111",
  47788=>"011000000",
  47789=>"100110111",
  47790=>"000000000",
  47791=>"000101100",
  47792=>"111000000",
  47793=>"001000000",
  47794=>"111111000",
  47795=>"010011000",
  47796=>"001111111",
  47797=>"111111111",
  47798=>"111111110",
  47799=>"111111000",
  47800=>"111111000",
  47801=>"010000001",
  47802=>"111111111",
  47803=>"100111111",
  47804=>"101000111",
  47805=>"000010111",
  47806=>"000000000",
  47807=>"111011011",
  47808=>"100000000",
  47809=>"111110000",
  47810=>"110100001",
  47811=>"000011001",
  47812=>"110000000",
  47813=>"000000000",
  47814=>"000000001",
  47815=>"010011000",
  47816=>"011010010",
  47817=>"110111111",
  47818=>"001011100",
  47819=>"111111110",
  47820=>"111111111",
  47821=>"110111111",
  47822=>"000001001",
  47823=>"111100000",
  47824=>"001000000",
  47825=>"000000010",
  47826=>"110111111",
  47827=>"000000101",
  47828=>"110110110",
  47829=>"000000000",
  47830=>"000000010",
  47831=>"011011100",
  47832=>"111111111",
  47833=>"000000111",
  47834=>"111101111",
  47835=>"110110110",
  47836=>"111111111",
  47837=>"000001001",
  47838=>"000011011",
  47839=>"111001001",
  47840=>"000000001",
  47841=>"011111111",
  47842=>"111000000",
  47843=>"101001001",
  47844=>"000010110",
  47845=>"101101101",
  47846=>"111111111",
  47847=>"000000000",
  47848=>"000000000",
  47849=>"000000101",
  47850=>"000000000",
  47851=>"000000001",
  47852=>"111111111",
  47853=>"000000010",
  47854=>"000000000",
  47855=>"111000000",
  47856=>"101111111",
  47857=>"011011111",
  47858=>"000001011",
  47859=>"011101000",
  47860=>"000000111",
  47861=>"111000000",
  47862=>"011111011",
  47863=>"110110000",
  47864=>"111110000",
  47865=>"000111111",
  47866=>"001011000",
  47867=>"000011011",
  47868=>"000001001",
  47869=>"001001001",
  47870=>"110100111",
  47871=>"000000000",
  47872=>"001001101",
  47873=>"001011011",
  47874=>"111111111",
  47875=>"111110111",
  47876=>"000000000",
  47877=>"000000000",
  47878=>"111100000",
  47879=>"111111000",
  47880=>"000000000",
  47881=>"101000000",
  47882=>"000000000",
  47883=>"001001111",
  47884=>"001001001",
  47885=>"111111111",
  47886=>"000000000",
  47887=>"111011000",
  47888=>"000000000",
  47889=>"000100111",
  47890=>"101111111",
  47891=>"010100000",
  47892=>"000000000",
  47893=>"001000000",
  47894=>"001011011",
  47895=>"000000001",
  47896=>"000000101",
  47897=>"000000000",
  47898=>"111111110",
  47899=>"111001111",
  47900=>"011011000",
  47901=>"000111111",
  47902=>"101000000",
  47903=>"110100010",
  47904=>"110111001",
  47905=>"000000000",
  47906=>"011010000",
  47907=>"000100000",
  47908=>"000000000",
  47909=>"111111111",
  47910=>"100100111",
  47911=>"111111100",
  47912=>"000011111",
  47913=>"111111110",
  47914=>"000000001",
  47915=>"011000000",
  47916=>"100000111",
  47917=>"000000001",
  47918=>"001000000",
  47919=>"000000111",
  47920=>"100110100",
  47921=>"000000000",
  47922=>"111111000",
  47923=>"000001001",
  47924=>"000000011",
  47925=>"000011111",
  47926=>"001001000",
  47927=>"111001111",
  47928=>"001111000",
  47929=>"001001101",
  47930=>"000000000",
  47931=>"000010010",
  47932=>"000000010",
  47933=>"110110000",
  47934=>"000010010",
  47935=>"111111000",
  47936=>"000000011",
  47937=>"111111110",
  47938=>"011001011",
  47939=>"000001000",
  47940=>"000001000",
  47941=>"111111111",
  47942=>"000111111",
  47943=>"111000000",
  47944=>"000000000",
  47945=>"010011011",
  47946=>"000000001",
  47947=>"111000000",
  47948=>"001010111",
  47949=>"000000011",
  47950=>"111100001",
  47951=>"011001011",
  47952=>"000000000",
  47953=>"111011111",
  47954=>"000000100",
  47955=>"000000100",
  47956=>"000000000",
  47957=>"011011011",
  47958=>"011001001",
  47959=>"110110010",
  47960=>"001001001",
  47961=>"001000000",
  47962=>"000111011",
  47963=>"101101111",
  47964=>"001011011",
  47965=>"010010010",
  47966=>"001000000",
  47967=>"110110110",
  47968=>"111000001",
  47969=>"111100011",
  47970=>"011001011",
  47971=>"101101111",
  47972=>"101111111",
  47973=>"000000111",
  47974=>"111001000",
  47975=>"001000000",
  47976=>"001001000",
  47977=>"000010000",
  47978=>"111111111",
  47979=>"000110110",
  47980=>"111110100",
  47981=>"010011111",
  47982=>"101111111",
  47983=>"000011011",
  47984=>"000000011",
  47985=>"000011011",
  47986=>"111111111",
  47987=>"000111001",
  47988=>"111011000",
  47989=>"100110110",
  47990=>"011011000",
  47991=>"111011001",
  47992=>"001000111",
  47993=>"111111111",
  47994=>"000000000",
  47995=>"000000000",
  47996=>"000000000",
  47997=>"000000000",
  47998=>"000000001",
  47999=>"101101000",
  48000=>"000000111",
  48001=>"000000010",
  48002=>"111111001",
  48003=>"000000011",
  48004=>"111111111",
  48005=>"000000000",
  48006=>"111000100",
  48007=>"111111111",
  48008=>"000001111",
  48009=>"001111111",
  48010=>"000000100",
  48011=>"111111000",
  48012=>"111000000",
  48013=>"100000000",
  48014=>"011110001",
  48015=>"000000000",
  48016=>"100000001",
  48017=>"111111111",
  48018=>"110110000",
  48019=>"001000000",
  48020=>"111111111",
  48021=>"000000010",
  48022=>"011000000",
  48023=>"001001001",
  48024=>"011001000",
  48025=>"110110111",
  48026=>"111111010",
  48027=>"000000000",
  48028=>"100100110",
  48029=>"000000001",
  48030=>"001001001",
  48031=>"111110111",
  48032=>"010111110",
  48033=>"010010010",
  48034=>"111101101",
  48035=>"000000000",
  48036=>"000000000",
  48037=>"001111111",
  48038=>"001001000",
  48039=>"010111110",
  48040=>"111000000",
  48041=>"000000000",
  48042=>"000000000",
  48043=>"001001001",
  48044=>"000010000",
  48045=>"000101000",
  48046=>"000000000",
  48047=>"111001001",
  48048=>"011111111",
  48049=>"110111011",
  48050=>"110111111",
  48051=>"111111111",
  48052=>"000000011",
  48053=>"000000000",
  48054=>"111111010",
  48055=>"110111111",
  48056=>"000011111",
  48057=>"000000000",
  48058=>"000000100",
  48059=>"111111111",
  48060=>"000001001",
  48061=>"111110110",
  48062=>"001011111",
  48063=>"000101101",
  48064=>"000010000",
  48065=>"000010000",
  48066=>"001001001",
  48067=>"000000000",
  48068=>"001000001",
  48069=>"011001001",
  48070=>"001000000",
  48071=>"010111111",
  48072=>"101101111",
  48073=>"000000000",
  48074=>"001001000",
  48075=>"000011000",
  48076=>"000110000",
  48077=>"111101000",
  48078=>"111110010",
  48079=>"000000000",
  48080=>"000000000",
  48081=>"001001011",
  48082=>"111110110",
  48083=>"011011011",
  48084=>"111111001",
  48085=>"000000000",
  48086=>"000000000",
  48087=>"100000000",
  48088=>"000100111",
  48089=>"000000000",
  48090=>"000000000",
  48091=>"111110111",
  48092=>"000001000",
  48093=>"001101101",
  48094=>"001011011",
  48095=>"101000001",
  48096=>"111101111",
  48097=>"110101000",
  48098=>"011011011",
  48099=>"111111010",
  48100=>"111111111",
  48101=>"000000000",
  48102=>"000000000",
  48103=>"111010010",
  48104=>"000000001",
  48105=>"000010010",
  48106=>"111001000",
  48107=>"111111000",
  48108=>"000001101",
  48109=>"000000100",
  48110=>"001000000",
  48111=>"110111111",
  48112=>"000000001",
  48113=>"110111111",
  48114=>"000000010",
  48115=>"001111111",
  48116=>"000010010",
  48117=>"010010111",
  48118=>"000000101",
  48119=>"000000000",
  48120=>"010000000",
  48121=>"001001001",
  48122=>"110111111",
  48123=>"001000100",
  48124=>"111110000",
  48125=>"000000000",
  48126=>"011000000",
  48127=>"111111110",
  48128=>"000111111",
  48129=>"000111010",
  48130=>"000111111",
  48131=>"111110111",
  48132=>"001111011",
  48133=>"000000100",
  48134=>"000011011",
  48135=>"111111111",
  48136=>"101101000",
  48137=>"001000000",
  48138=>"100111111",
  48139=>"000000111",
  48140=>"000100000",
  48141=>"000001111",
  48142=>"011110111",
  48143=>"110110000",
  48144=>"111100000",
  48145=>"111111001",
  48146=>"111111111",
  48147=>"000000001",
  48148=>"000111111",
  48149=>"000000000",
  48150=>"110110000",
  48151=>"011110111",
  48152=>"111111110",
  48153=>"100100000",
  48154=>"000000000",
  48155=>"000000001",
  48156=>"111111111",
  48157=>"111111111",
  48158=>"111111111",
  48159=>"111111100",
  48160=>"001001000",
  48161=>"111111111",
  48162=>"111111100",
  48163=>"000000010",
  48164=>"111100111",
  48165=>"100000100",
  48166=>"000000000",
  48167=>"010111100",
  48168=>"100000000",
  48169=>"000000000",
  48170=>"000000000",
  48171=>"110111110",
  48172=>"011111111",
  48173=>"111111111",
  48174=>"100111111",
  48175=>"000000000",
  48176=>"000000001",
  48177=>"110110000",
  48178=>"001011100",
  48179=>"000000000",
  48180=>"111000000",
  48181=>"001100000",
  48182=>"000000000",
  48183=>"000000000",
  48184=>"010111111",
  48185=>"111000101",
  48186=>"000000000",
  48187=>"011011011",
  48188=>"111111111",
  48189=>"100110100",
  48190=>"100110110",
  48191=>"100000100",
  48192=>"011001101",
  48193=>"011111111",
  48194=>"000000001",
  48195=>"000000000",
  48196=>"001111011",
  48197=>"111111111",
  48198=>"000000000",
  48199=>"100100111",
  48200=>"110000011",
  48201=>"000000000",
  48202=>"111111111",
  48203=>"000111100",
  48204=>"111111111",
  48205=>"000000000",
  48206=>"111111000",
  48207=>"000000000",
  48208=>"111010000",
  48209=>"000000000",
  48210=>"000010000",
  48211=>"011111111",
  48212=>"101000000",
  48213=>"011111111",
  48214=>"000000000",
  48215=>"111001011",
  48216=>"011011000",
  48217=>"000000000",
  48218=>"111111111",
  48219=>"000000001",
  48220=>"111111111",
  48221=>"000000000",
  48222=>"000000000",
  48223=>"001000001",
  48224=>"000000000",
  48225=>"000000000",
  48226=>"000000000",
  48227=>"110110110",
  48228=>"111100100",
  48229=>"000000001",
  48230=>"111111111",
  48231=>"111111111",
  48232=>"111111111",
  48233=>"000100000",
  48234=>"000000000",
  48235=>"000000011",
  48236=>"111110010",
  48237=>"111011011",
  48238=>"000111111",
  48239=>"001000000",
  48240=>"111111111",
  48241=>"110110010",
  48242=>"111011010",
  48243=>"111111111",
  48244=>"101111001",
  48245=>"100000101",
  48246=>"000000000",
  48247=>"001000000",
  48248=>"111111111",
  48249=>"000000001",
  48250=>"111100001",
  48251=>"111111111",
  48252=>"000000000",
  48253=>"101111111",
  48254=>"100000000",
  48255=>"100000000",
  48256=>"011111111",
  48257=>"000000000",
  48258=>"000000000",
  48259=>"111111111",
  48260=>"011111111",
  48261=>"111111111",
  48262=>"011111111",
  48263=>"000000000",
  48264=>"101111111",
  48265=>"110111111",
  48266=>"000000111",
  48267=>"000000000",
  48268=>"000010111",
  48269=>"000000000",
  48270=>"100100000",
  48271=>"101000000",
  48272=>"000000000",
  48273=>"101111111",
  48274=>"000110110",
  48275=>"110110000",
  48276=>"111111111",
  48277=>"111111111",
  48278=>"000000000",
  48279=>"000000000",
  48280=>"111111110",
  48281=>"111111110",
  48282=>"000000000",
  48283=>"100000000",
  48284=>"000000000",
  48285=>"000000000",
  48286=>"000111111",
  48287=>"111111011",
  48288=>"000000000",
  48289=>"000011011",
  48290=>"111111111",
  48291=>"000000000",
  48292=>"000001001",
  48293=>"000110111",
  48294=>"010110111",
  48295=>"100000000",
  48296=>"000000010",
  48297=>"110111110",
  48298=>"111111111",
  48299=>"111111111",
  48300=>"111111111",
  48301=>"011001100",
  48302=>"100000100",
  48303=>"111010110",
  48304=>"000110110",
  48305=>"000100100",
  48306=>"110110000",
  48307=>"111111111",
  48308=>"000000000",
  48309=>"111100100",
  48310=>"000000000",
  48311=>"111111100",
  48312=>"000110110",
  48313=>"000000000",
  48314=>"000000000",
  48315=>"000000110",
  48316=>"001001111",
  48317=>"101101101",
  48318=>"111111111",
  48319=>"000110110",
  48320=>"000010110",
  48321=>"001000000",
  48322=>"111111111",
  48323=>"110111111",
  48324=>"000010000",
  48325=>"011011000",
  48326=>"000000000",
  48327=>"000000010",
  48328=>"111100000",
  48329=>"101100000",
  48330=>"000000000",
  48331=>"111111111",
  48332=>"000010110",
  48333=>"001000000",
  48334=>"100100100",
  48335=>"111101111",
  48336=>"000001001",
  48337=>"001000000",
  48338=>"111111110",
  48339=>"000000000",
  48340=>"001011111",
  48341=>"000100100",
  48342=>"011000000",
  48343=>"000000000",
  48344=>"111111111",
  48345=>"100010111",
  48346=>"000000000",
  48347=>"110010001",
  48348=>"101101111",
  48349=>"111111111",
  48350=>"111111110",
  48351=>"000011111",
  48352=>"000111111",
  48353=>"000000000",
  48354=>"111111111",
  48355=>"000011111",
  48356=>"111101101",
  48357=>"000000100",
  48358=>"110000110",
  48359=>"000000000",
  48360=>"000000001",
  48361=>"111111111",
  48362=>"111111111",
  48363=>"000000000",
  48364=>"000010000",
  48365=>"111111111",
  48366=>"111111000",
  48367=>"100111100",
  48368=>"111111111",
  48369=>"000001000",
  48370=>"011111111",
  48371=>"000000000",
  48372=>"011000000",
  48373=>"100000110",
  48374=>"111111111",
  48375=>"000000000",
  48376=>"110000000",
  48377=>"000010000",
  48378=>"110111111",
  48379=>"011010000",
  48380=>"101100111",
  48381=>"001011011",
  48382=>"111111000",
  48383=>"111111111",
  48384=>"000000000",
  48385=>"011011011",
  48386=>"101111111",
  48387=>"111111111",
  48388=>"001111111",
  48389=>"011011000",
  48390=>"111000000",
  48391=>"001111110",
  48392=>"110110000",
  48393=>"000100101",
  48394=>"111110110",
  48395=>"100111111",
  48396=>"110110110",
  48397=>"111111111",
  48398=>"111111110",
  48399=>"000000100",
  48400=>"110111111",
  48401=>"100000000",
  48402=>"111100001",
  48403=>"000000000",
  48404=>"111111000",
  48405=>"111111001",
  48406=>"110110110",
  48407=>"000000000",
  48408=>"111111111",
  48409=>"000000100",
  48410=>"000000000",
  48411=>"111111100",
  48412=>"000000000",
  48413=>"011101000",
  48414=>"011111011",
  48415=>"000111111",
  48416=>"000110111",
  48417=>"000000000",
  48418=>"100110111",
  48419=>"111110000",
  48420=>"101111110",
  48421=>"111100000",
  48422=>"111111011",
  48423=>"111101000",
  48424=>"111111111",
  48425=>"000000000",
  48426=>"010010001",
  48427=>"111111111",
  48428=>"000000000",
  48429=>"111011011",
  48430=>"111110000",
  48431=>"000000000",
  48432=>"011111111",
  48433=>"111100000",
  48434=>"110111000",
  48435=>"000000100",
  48436=>"110111010",
  48437=>"101011000",
  48438=>"000010000",
  48439=>"000000000",
  48440=>"000000111",
  48441=>"000000000",
  48442=>"101101101",
  48443=>"000100111",
  48444=>"000000011",
  48445=>"000000000",
  48446=>"111011001",
  48447=>"111111111",
  48448=>"010001100",
  48449=>"111111110",
  48450=>"000110110",
  48451=>"000000000",
  48452=>"111111100",
  48453=>"000000000",
  48454=>"111000100",
  48455=>"000000000",
  48456=>"110110100",
  48457=>"000000000",
  48458=>"110111111",
  48459=>"011010000",
  48460=>"001011000",
  48461=>"000011111",
  48462=>"110110100",
  48463=>"111010000",
  48464=>"111010000",
  48465=>"000001001",
  48466=>"011000000",
  48467=>"011011001",
  48468=>"010000000",
  48469=>"000000001",
  48470=>"101000000",
  48471=>"001000000",
  48472=>"010010111",
  48473=>"000110000",
  48474=>"000000000",
  48475=>"111010000",
  48476=>"000000000",
  48477=>"110111110",
  48478=>"000000000",
  48479=>"001011011",
  48480=>"111111111",
  48481=>"111111111",
  48482=>"111110011",
  48483=>"000000000",
  48484=>"111111111",
  48485=>"111111111",
  48486=>"000010000",
  48487=>"111111110",
  48488=>"000000000",
  48489=>"010000000",
  48490=>"111111111",
  48491=>"001011111",
  48492=>"111111111",
  48493=>"001111111",
  48494=>"111111111",
  48495=>"010010000",
  48496=>"000000000",
  48497=>"111110111",
  48498=>"011011000",
  48499=>"100100110",
  48500=>"101111100",
  48501=>"001000001",
  48502=>"000000000",
  48503=>"011000000",
  48504=>"000000011",
  48505=>"000000110",
  48506=>"111111001",
  48507=>"100110100",
  48508=>"000111111",
  48509=>"111111111",
  48510=>"101101111",
  48511=>"000000000",
  48512=>"000000110",
  48513=>"000000000",
  48514=>"111111111",
  48515=>"011111000",
  48516=>"111111000",
  48517=>"111111000",
  48518=>"000000000",
  48519=>"111111111",
  48520=>"001001000",
  48521=>"000001000",
  48522=>"000000111",
  48523=>"111110010",
  48524=>"000111111",
  48525=>"111111111",
  48526=>"110100110",
  48527=>"111111000",
  48528=>"111111011",
  48529=>"000000000",
  48530=>"111111111",
  48531=>"000001101",
  48532=>"111101110",
  48533=>"111101111",
  48534=>"100111011",
  48535=>"001111111",
  48536=>"100100001",
  48537=>"000000000",
  48538=>"100111101",
  48539=>"110100110",
  48540=>"010010000",
  48541=>"000101100",
  48542=>"000000000",
  48543=>"000111111",
  48544=>"111000000",
  48545=>"101001100",
  48546=>"111111111",
  48547=>"000000111",
  48548=>"100110000",
  48549=>"111111111",
  48550=>"111111011",
  48551=>"000000000",
  48552=>"111111000",
  48553=>"000000000",
  48554=>"000111111",
  48555=>"111111100",
  48556=>"111111000",
  48557=>"111001001",
  48558=>"000000110",
  48559=>"000111111",
  48560=>"000000011",
  48561=>"111101000",
  48562=>"100100000",
  48563=>"111111111",
  48564=>"111111010",
  48565=>"100000000",
  48566=>"001101111",
  48567=>"100100000",
  48568=>"111111110",
  48569=>"110111111",
  48570=>"111100111",
  48571=>"101111111",
  48572=>"000100100",
  48573=>"110000000",
  48574=>"000000000",
  48575=>"011011011",
  48576=>"000010000",
  48577=>"111111111",
  48578=>"000010110",
  48579=>"000000001",
  48580=>"000000101",
  48581=>"010000100",
  48582=>"000010000",
  48583=>"000110111",
  48584=>"000001000",
  48585=>"111111100",
  48586=>"000000000",
  48587=>"010010000",
  48588=>"110111000",
  48589=>"110111111",
  48590=>"000000000",
  48591=>"111111101",
  48592=>"000000000",
  48593=>"010111111",
  48594=>"011111111",
  48595=>"111111111",
  48596=>"101100100",
  48597=>"111111111",
  48598=>"000000000",
  48599=>"000000111",
  48600=>"110000000",
  48601=>"111001001",
  48602=>"101101000",
  48603=>"000000000",
  48604=>"010000000",
  48605=>"000000000",
  48606=>"000100000",
  48607=>"110111111",
  48608=>"010110110",
  48609=>"000011011",
  48610=>"000000000",
  48611=>"011110111",
  48612=>"011111011",
  48613=>"101101111",
  48614=>"000001001",
  48615=>"010001111",
  48616=>"000000100",
  48617=>"000000001",
  48618=>"001011011",
  48619=>"110000000",
  48620=>"111111111",
  48621=>"000100100",
  48622=>"100110110",
  48623=>"111111100",
  48624=>"100110111",
  48625=>"000000000",
  48626=>"111111111",
  48627=>"000000000",
  48628=>"000000000",
  48629=>"101101001",
  48630=>"111111111",
  48631=>"100000000",
  48632=>"000000000",
  48633=>"110010110",
  48634=>"001111111",
  48635=>"011001011",
  48636=>"110100100",
  48637=>"000000000",
  48638=>"111111111",
  48639=>"110111111",
  48640=>"001111100",
  48641=>"000000111",
  48642=>"111111000",
  48643=>"000111111",
  48644=>"001001000",
  48645=>"100110100",
  48646=>"111100100",
  48647=>"000000111",
  48648=>"000000000",
  48649=>"001001000",
  48650=>"111111110",
  48651=>"000110000",
  48652=>"011011001",
  48653=>"111111111",
  48654=>"111111011",
  48655=>"101000101",
  48656=>"011000100",
  48657=>"110000000",
  48658=>"111100110",
  48659=>"000000111",
  48660=>"000110000",
  48661=>"111100100",
  48662=>"111001101",
  48663=>"001001111",
  48664=>"010100111",
  48665=>"011011110",
  48666=>"111011000",
  48667=>"000000100",
  48668=>"000000000",
  48669=>"111111111",
  48670=>"110111110",
  48671=>"000011000",
  48672=>"001011000",
  48673=>"000111111",
  48674=>"101100000",
  48675=>"001000000",
  48676=>"000000001",
  48677=>"000000010",
  48678=>"111100111",
  48679=>"000000000",
  48680=>"001011111",
  48681=>"110111111",
  48682=>"110100111",
  48683=>"111111111",
  48684=>"111110111",
  48685=>"000001111",
  48686=>"000000000",
  48687=>"111111111",
  48688=>"000000011",
  48689=>"111101111",
  48690=>"110110110",
  48691=>"111111000",
  48692=>"000000000",
  48693=>"011000000",
  48694=>"101000001",
  48695=>"100111000",
  48696=>"000000000",
  48697=>"111111011",
  48698=>"111111111",
  48699=>"000011111",
  48700=>"011000000",
  48701=>"100111111",
  48702=>"100111111",
  48703=>"000000111",
  48704=>"010101101",
  48705=>"110000000",
  48706=>"111111100",
  48707=>"111111011",
  48708=>"011111011",
  48709=>"010000111",
  48710=>"111111010",
  48711=>"011011011",
  48712=>"000000100",
  48713=>"000000111",
  48714=>"111111111",
  48715=>"000000000",
  48716=>"000000000",
  48717=>"111000111",
  48718=>"100100111",
  48719=>"000111111",
  48720=>"111111111",
  48721=>"000100111",
  48722=>"111000001",
  48723=>"000111110",
  48724=>"111000100",
  48725=>"000000000",
  48726=>"111000001",
  48727=>"111111000",
  48728=>"011001011",
  48729=>"001000111",
  48730=>"111000000",
  48731=>"111110110",
  48732=>"111100000",
  48733=>"000000111",
  48734=>"000100111",
  48735=>"111110000",
  48736=>"000000000",
  48737=>"000100111",
  48738=>"000000000",
  48739=>"111101111",
  48740=>"011111100",
  48741=>"011010111",
  48742=>"111111111",
  48743=>"111000000",
  48744=>"000111111",
  48745=>"111111000",
  48746=>"111001111",
  48747=>"000000111",
  48748=>"110111110",
  48749=>"111111111",
  48750=>"111000000",
  48751=>"000000100",
  48752=>"100100100",
  48753=>"001000000",
  48754=>"111100000",
  48755=>"011111110",
  48756=>"100000100",
  48757=>"000001111",
  48758=>"010000000",
  48759=>"001101111",
  48760=>"010011001",
  48761=>"010010100",
  48762=>"000000000",
  48763=>"000000011",
  48764=>"000011011",
  48765=>"010110110",
  48766=>"111101000",
  48767=>"111111111",
  48768=>"111111111",
  48769=>"000000000",
  48770=>"111011001",
  48771=>"100000000",
  48772=>"111111001",
  48773=>"001001111",
  48774=>"000000110",
  48775=>"110100000",
  48776=>"011111111",
  48777=>"000000000",
  48778=>"000100000",
  48779=>"000000111",
  48780=>"001000000",
  48781=>"000111111",
  48782=>"111110000",
  48783=>"111111010",
  48784=>"111000000",
  48785=>"111111110",
  48786=>"111111110",
  48787=>"111100000",
  48788=>"111101100",
  48789=>"111010000",
  48790=>"111111000",
  48791=>"111111000",
  48792=>"001000101",
  48793=>"000000001",
  48794=>"111000000",
  48795=>"000001000",
  48796=>"000111111",
  48797=>"111000100",
  48798=>"000000111",
  48799=>"110111111",
  48800=>"111111001",
  48801=>"111111111",
  48802=>"111000000",
  48803=>"011000000",
  48804=>"001001111",
  48805=>"001111111",
  48806=>"111101000",
  48807=>"111111100",
  48808=>"000000000",
  48809=>"001000000",
  48810=>"000001011",
  48811=>"000000000",
  48812=>"001111111",
  48813=>"100100000",
  48814=>"001000000",
  48815=>"000000000",
  48816=>"000011011",
  48817=>"100111111",
  48818=>"000111110",
  48819=>"111111001",
  48820=>"111111000",
  48821=>"111111001",
  48822=>"111010111",
  48823=>"000000111",
  48824=>"111101000",
  48825=>"110111111",
  48826=>"100000101",
  48827=>"001011111",
  48828=>"000110000",
  48829=>"111111111",
  48830=>"000100000",
  48831=>"000000100",
  48832=>"101011111",
  48833=>"111111010",
  48834=>"000111111",
  48835=>"000011011",
  48836=>"111111111",
  48837=>"001001000",
  48838=>"000111111",
  48839=>"000011011",
  48840=>"010111111",
  48841=>"000000000",
  48842=>"000010100",
  48843=>"111111111",
  48844=>"000000010",
  48845=>"001000000",
  48846=>"000011111",
  48847=>"000000100",
  48848=>"000100100",
  48849=>"000000010",
  48850=>"000000001",
  48851=>"000000010",
  48852=>"100000101",
  48853=>"000000000",
  48854=>"010111111",
  48855=>"111000000",
  48856=>"111111111",
  48857=>"011111011",
  48858=>"000111111",
  48859=>"000010111",
  48860=>"111111111",
  48861=>"000000000",
  48862=>"111000000",
  48863=>"101111111",
  48864=>"100000000",
  48865=>"000001111",
  48866=>"000000000",
  48867=>"111111111",
  48868=>"000000011",
  48869=>"111111111",
  48870=>"111111111",
  48871=>"001001000",
  48872=>"000000000",
  48873=>"111111000",
  48874=>"010111011",
  48875=>"001111001",
  48876=>"111001000",
  48877=>"000111000",
  48878=>"000000101",
  48879=>"111111111",
  48880=>"100100010",
  48881=>"111111010",
  48882=>"111111111",
  48883=>"111000111",
  48884=>"000000111",
  48885=>"111111111",
  48886=>"100100101",
  48887=>"000010000",
  48888=>"111111111",
  48889=>"111111111",
  48890=>"001111111",
  48891=>"000000111",
  48892=>"100011111",
  48893=>"000111000",
  48894=>"001000000",
  48895=>"111111000",
  48896=>"000000100",
  48897=>"000000000",
  48898=>"111000000",
  48899=>"111111000",
  48900=>"110111010",
  48901=>"001111111",
  48902=>"000000000",
  48903=>"001001000",
  48904=>"000000101",
  48905=>"000000000",
  48906=>"111010000",
  48907=>"110111010",
  48908=>"100000000",
  48909=>"000000111",
  48910=>"011011000",
  48911=>"110110111",
  48912=>"000000000",
  48913=>"000000000",
  48914=>"000000000",
  48915=>"000111111",
  48916=>"001111111",
  48917=>"111111000",
  48918=>"001001011",
  48919=>"111111111",
  48920=>"101000000",
  48921=>"110111111",
  48922=>"000000000",
  48923=>"101111111",
  48924=>"000000000",
  48925=>"111111111",
  48926=>"000000000",
  48927=>"111111110",
  48928=>"111111111",
  48929=>"000000000",
  48930=>"000011111",
  48931=>"000000000",
  48932=>"000011111",
  48933=>"000000000",
  48934=>"100110110",
  48935=>"111110010",
  48936=>"111110111",
  48937=>"111111111",
  48938=>"000111111",
  48939=>"110111111",
  48940=>"110000010",
  48941=>"000111111",
  48942=>"111111111",
  48943=>"100000000",
  48944=>"011011110",
  48945=>"000000111",
  48946=>"111111111",
  48947=>"000000101",
  48948=>"110111000",
  48949=>"111111111",
  48950=>"111111111",
  48951=>"000001000",
  48952=>"111111110",
  48953=>"111100000",
  48954=>"000000000",
  48955=>"111111111",
  48956=>"100000000",
  48957=>"000001111",
  48958=>"000000000",
  48959=>"111111000",
  48960=>"000001011",
  48961=>"110000000",
  48962=>"001011000",
  48963=>"000000000",
  48964=>"111111111",
  48965=>"110110000",
  48966=>"111111001",
  48967=>"111111111",
  48968=>"111000011",
  48969=>"111111001",
  48970=>"000100111",
  48971=>"000111101",
  48972=>"000100111",
  48973=>"000011000",
  48974=>"111111110",
  48975=>"001011111",
  48976=>"000000000",
  48977=>"111111111",
  48978=>"010011000",
  48979=>"000000001",
  48980=>"111111111",
  48981=>"011101111",
  48982=>"110111110",
  48983=>"100111111",
  48984=>"011111111",
  48985=>"111111001",
  48986=>"111000000",
  48987=>"101001100",
  48988=>"010000000",
  48989=>"111111000",
  48990=>"000111011",
  48991=>"111110000",
  48992=>"111101001",
  48993=>"110111111",
  48994=>"101111000",
  48995=>"111000000",
  48996=>"101111111",
  48997=>"111111111",
  48998=>"111101000",
  48999=>"111111110",
  49000=>"100110110",
  49001=>"000111111",
  49002=>"110000100",
  49003=>"000000100",
  49004=>"011011011",
  49005=>"000000101",
  49006=>"110110110",
  49007=>"000000111",
  49008=>"111110000",
  49009=>"000000000",
  49010=>"010000001",
  49011=>"001001011",
  49012=>"111100100",
  49013=>"111111110",
  49014=>"000000000",
  49015=>"010110110",
  49016=>"111111111",
  49017=>"001000000",
  49018=>"111111111",
  49019=>"000000000",
  49020=>"101111111",
  49021=>"000110111",
  49022=>"001000000",
  49023=>"111000000",
  49024=>"000000000",
  49025=>"001111000",
  49026=>"110000110",
  49027=>"000111011",
  49028=>"010010110",
  49029=>"111111111",
  49030=>"100100111",
  49031=>"100000110",
  49032=>"111111111",
  49033=>"000000000",
  49034=>"000100111",
  49035=>"111111001",
  49036=>"000000000",
  49037=>"101001001",
  49038=>"111111010",
  49039=>"000000111",
  49040=>"001001000",
  49041=>"111111111",
  49042=>"001001111",
  49043=>"111001001",
  49044=>"111111111",
  49045=>"111101111",
  49046=>"000000110",
  49047=>"111110000",
  49048=>"001111111",
  49049=>"110110110",
  49050=>"111001111",
  49051=>"111111111",
  49052=>"100110111",
  49053=>"000011111",
  49054=>"111111111",
  49055=>"000000000",
  49056=>"111111111",
  49057=>"111111000",
  49058=>"111111010",
  49059=>"111111011",
  49060=>"000000001",
  49061=>"100000011",
  49062=>"111111111",
  49063=>"111111111",
  49064=>"000001111",
  49065=>"000110111",
  49066=>"111111110",
  49067=>"110100100",
  49068=>"111111110",
  49069=>"101011011",
  49070=>"111011000",
  49071=>"000000000",
  49072=>"110000000",
  49073=>"011000000",
  49074=>"001010010",
  49075=>"111111110",
  49076=>"111111011",
  49077=>"110111111",
  49078=>"001000000",
  49079=>"010110110",
  49080=>"000000111",
  49081=>"000111111",
  49082=>"111000111",
  49083=>"110000000",
  49084=>"111001000",
  49085=>"000000001",
  49086=>"000101111",
  49087=>"000000111",
  49088=>"100111111",
  49089=>"000000100",
  49090=>"000000000",
  49091=>"000000111",
  49092=>"001000000",
  49093=>"000011000",
  49094=>"111010000",
  49095=>"000000000",
  49096=>"101111100",
  49097=>"111101110",
  49098=>"001111000",
  49099=>"111000000",
  49100=>"000101000",
  49101=>"000000000",
  49102=>"000000111",
  49103=>"010111111",
  49104=>"001101001",
  49105=>"101000000",
  49106=>"000000000",
  49107=>"000000111",
  49108=>"111101000",
  49109=>"000000110",
  49110=>"000000111",
  49111=>"110111101",
  49112=>"000000100",
  49113=>"101111111",
  49114=>"111111000",
  49115=>"010010000",
  49116=>"000000000",
  49117=>"111011000",
  49118=>"011000100",
  49119=>"000000111",
  49120=>"100000000",
  49121=>"111101111",
  49122=>"000000001",
  49123=>"000001111",
  49124=>"110000000",
  49125=>"000000000",
  49126=>"000101110",
  49127=>"110111111",
  49128=>"111111110",
  49129=>"111001111",
  49130=>"000011011",
  49131=>"000000100",
  49132=>"100110111",
  49133=>"111111000",
  49134=>"000000000",
  49135=>"000011111",
  49136=>"111000000",
  49137=>"111001001",
  49138=>"101111100",
  49139=>"000000000",
  49140=>"000000111",
  49141=>"001000000",
  49142=>"110111100",
  49143=>"000011010",
  49144=>"000000100",
  49145=>"111011000",
  49146=>"111101100",
  49147=>"111111111",
  49148=>"000100110",
  49149=>"001000000",
  49150=>"111111000",
  49151=>"111110010",
  49152=>"100001001",
  49153=>"000000100",
  49154=>"111111111",
  49155=>"000000000",
  49156=>"111111111",
  49157=>"111100000",
  49158=>"111111111",
  49159=>"111111111",
  49160=>"000000100",
  49161=>"111000000",
  49162=>"111001000",
  49163=>"111001001",
  49164=>"100111001",
  49165=>"010000000",
  49166=>"111100011",
  49167=>"000111111",
  49168=>"000000110",
  49169=>"000111000",
  49170=>"111100001",
  49171=>"111111111",
  49172=>"001111111",
  49173=>"111111000",
  49174=>"011011000",
  49175=>"001000000",
  49176=>"100000101",
  49177=>"111100000",
  49178=>"111111111",
  49179=>"011110000",
  49180=>"111111111",
  49181=>"110100111",
  49182=>"000111111",
  49183=>"001001101",
  49184=>"000001011",
  49185=>"000000000",
  49186=>"111111111",
  49187=>"000000000",
  49188=>"111111111",
  49189=>"000000100",
  49190=>"000000000",
  49191=>"001001000",
  49192=>"011011111",
  49193=>"000000000",
  49194=>"000000100",
  49195=>"111101000",
  49196=>"000110000",
  49197=>"100111111",
  49198=>"100111111",
  49199=>"011001000",
  49200=>"001001001",
  49201=>"001111000",
  49202=>"001111111",
  49203=>"000000000",
  49204=>"100000011",
  49205=>"111111000",
  49206=>"000000000",
  49207=>"111111111",
  49208=>"001001111",
  49209=>"000100101",
  49210=>"011111111",
  49211=>"111110100",
  49212=>"111111111",
  49213=>"111000000",
  49214=>"000000000",
  49215=>"000000100",
  49216=>"011111111",
  49217=>"000000000",
  49218=>"000100000",
  49219=>"001110100",
  49220=>"111111111",
  49221=>"000000000",
  49222=>"111111011",
  49223=>"111111111",
  49224=>"011011111",
  49225=>"000000111",
  49226=>"000000000",
  49227=>"000000000",
  49228=>"000010111",
  49229=>"111111111",
  49230=>"100000110",
  49231=>"000000100",
  49232=>"111110111",
  49233=>"001100100",
  49234=>"001000000",
  49235=>"011001100",
  49236=>"000000000",
  49237=>"000000000",
  49238=>"000001000",
  49239=>"011000000",
  49240=>"100000000",
  49241=>"111111111",
  49242=>"111101101",
  49243=>"000000011",
  49244=>"111111111",
  49245=>"100000000",
  49246=>"001100111",
  49247=>"111011011",
  49248=>"111111111",
  49249=>"000000010",
  49250=>"111111111",
  49251=>"101001001",
  49252=>"000011010",
  49253=>"100101111",
  49254=>"111111111",
  49255=>"111000000",
  49256=>"111111011",
  49257=>"000000000",
  49258=>"000000111",
  49259=>"000000101",
  49260=>"100000000",
  49261=>"111110111",
  49262=>"001001111",
  49263=>"111011011",
  49264=>"000000000",
  49265=>"000100000",
  49266=>"000000000",
  49267=>"001111101",
  49268=>"101000000",
  49269=>"000000000",
  49270=>"000000000",
  49271=>"000000000",
  49272=>"111111000",
  49273=>"001101111",
  49274=>"000000000",
  49275=>"011000000",
  49276=>"000000000",
  49277=>"111111111",
  49278=>"111111001",
  49279=>"111111111",
  49280=>"000000000",
  49281=>"011010101",
  49282=>"000000000",
  49283=>"001011001",
  49284=>"000101001",
  49285=>"111101000",
  49286=>"101000000",
  49287=>"111111111",
  49288=>"111111111",
  49289=>"111111111",
  49290=>"101000000",
  49291=>"111111000",
  49292=>"111111111",
  49293=>"000000000",
  49294=>"000000000",
  49295=>"110111001",
  49296=>"100100111",
  49297=>"000110111",
  49298=>"011000000",
  49299=>"000000010",
  49300=>"011111110",
  49301=>"000000000",
  49302=>"111111111",
  49303=>"100100110",
  49304=>"001000000",
  49305=>"111111101",
  49306=>"111111111",
  49307=>"000111111",
  49308=>"000000000",
  49309=>"111110000",
  49310=>"011001111",
  49311=>"000000111",
  49312=>"000000000",
  49313=>"000000000",
  49314=>"111010111",
  49315=>"000000000",
  49316=>"100000001",
  49317=>"011011001",
  49318=>"111000000",
  49319=>"000011011",
  49320=>"111111100",
  49321=>"000000000",
  49322=>"001000000",
  49323=>"010011000",
  49324=>"111111111",
  49325=>"110101110",
  49326=>"111111111",
  49327=>"001001000",
  49328=>"000111111",
  49329=>"000001000",
  49330=>"111111111",
  49331=>"000000101",
  49332=>"000011111",
  49333=>"011100111",
  49334=>"000111100",
  49335=>"000000000",
  49336=>"111111111",
  49337=>"111111111",
  49338=>"011000100",
  49339=>"111000000",
  49340=>"001000000",
  49341=>"000000111",
  49342=>"111111111",
  49343=>"111110111",
  49344=>"001000001",
  49345=>"111111111",
  49346=>"000100100",
  49347=>"000000000",
  49348=>"110110000",
  49349=>"111111111",
  49350=>"000110010",
  49351=>"111000000",
  49352=>"111111100",
  49353=>"111000000",
  49354=>"000111011",
  49355=>"111111111",
  49356=>"111111111",
  49357=>"100110000",
  49358=>"000000000",
  49359=>"010000000",
  49360=>"111111111",
  49361=>"001001000",
  49362=>"000111110",
  49363=>"000010111",
  49364=>"110110111",
  49365=>"111111111",
  49366=>"101001000",
  49367=>"111111000",
  49368=>"000100000",
  49369=>"000011001",
  49370=>"111111111",
  49371=>"011111111",
  49372=>"111011111",
  49373=>"011000111",
  49374=>"110000010",
  49375=>"111000100",
  49376=>"000000111",
  49377=>"111111111",
  49378=>"000000000",
  49379=>"101000000",
  49380=>"001111111",
  49381=>"001000001",
  49382=>"001000000",
  49383=>"111111111",
  49384=>"100000000",
  49385=>"001011011",
  49386=>"100100111",
  49387=>"111111101",
  49388=>"000001000",
  49389=>"111111111",
  49390=>"011011111",
  49391=>"111101101",
  49392=>"100100100",
  49393=>"000000011",
  49394=>"111001111",
  49395=>"111111111",
  49396=>"000100111",
  49397=>"111000000",
  49398=>"000000001",
  49399=>"010011010",
  49400=>"000000000",
  49401=>"000101111",
  49402=>"111111110",
  49403=>"111110010",
  49404=>"110111111",
  49405=>"000000000",
  49406=>"000001111",
  49407=>"011000000",
  49408=>"011001111",
  49409=>"010011011",
  49410=>"011001000",
  49411=>"000000000",
  49412=>"111111111",
  49413=>"100110100",
  49414=>"100100000",
  49415=>"001111111",
  49416=>"000000101",
  49417=>"000000000",
  49418=>"111001000",
  49419=>"000000011",
  49420=>"000000000",
  49421=>"111111110",
  49422=>"000000000",
  49423=>"000000000",
  49424=>"101101111",
  49425=>"011100100",
  49426=>"111000100",
  49427=>"111111111",
  49428=>"000000000",
  49429=>"000000000",
  49430=>"100110111",
  49431=>"111111011",
  49432=>"010011111",
  49433=>"000000000",
  49434=>"000111111",
  49435=>"100110111",
  49436=>"000000010",
  49437=>"100000000",
  49438=>"000000000",
  49439=>"111001111",
  49440=>"110100111",
  49441=>"011111111",
  49442=>"111110110",
  49443=>"000010010",
  49444=>"001000100",
  49445=>"000001101",
  49446=>"111111111",
  49447=>"000100000",
  49448=>"000000000",
  49449=>"110111111",
  49450=>"010011111",
  49451=>"000101111",
  49452=>"001000010",
  49453=>"000010111",
  49454=>"101111111",
  49455=>"111111001",
  49456=>"000100100",
  49457=>"111110111",
  49458=>"111111000",
  49459=>"000000000",
  49460=>"000000000",
  49461=>"000100111",
  49462=>"111000101",
  49463=>"010001001",
  49464=>"100100010",
  49465=>"001111111",
  49466=>"001000000",
  49467=>"000000000",
  49468=>"000000000",
  49469=>"111110110",
  49470=>"000000000",
  49471=>"011111111",
  49472=>"000000001",
  49473=>"101101000",
  49474=>"001000000",
  49475=>"111111111",
  49476=>"111001001",
  49477=>"111111111",
  49478=>"000000000",
  49479=>"111101000",
  49480=>"000000000",
  49481=>"000000111",
  49482=>"011001111",
  49483=>"001100100",
  49484=>"000000111",
  49485=>"000110111",
  49486=>"000000101",
  49487=>"000000000",
  49488=>"111111111",
  49489=>"000001111",
  49490=>"011111000",
  49491=>"011111111",
  49492=>"111111111",
  49493=>"001001011",
  49494=>"000000000",
  49495=>"000000000",
  49496=>"111101111",
  49497=>"000000000",
  49498=>"000000000",
  49499=>"110110100",
  49500=>"111010000",
  49501=>"010111111",
  49502=>"111000110",
  49503=>"111111100",
  49504=>"111101100",
  49505=>"000000000",
  49506=>"111111111",
  49507=>"000000000",
  49508=>"000000000",
  49509=>"010000000",
  49510=>"111111111",
  49511=>"111000111",
  49512=>"100000000",
  49513=>"111111000",
  49514=>"000000000",
  49515=>"000100000",
  49516=>"100000100",
  49517=>"111111101",
  49518=>"000001000",
  49519=>"000001001",
  49520=>"100110111",
  49521=>"111101000",
  49522=>"000110100",
  49523=>"110100111",
  49524=>"000000000",
  49525=>"111111000",
  49526=>"111000000",
  49527=>"000000000",
  49528=>"000000000",
  49529=>"111111111",
  49530=>"000000010",
  49531=>"010000000",
  49532=>"100100110",
  49533=>"000100101",
  49534=>"111111111",
  49535=>"000000001",
  49536=>"000000100",
  49537=>"000000000",
  49538=>"111000000",
  49539=>"111111111",
  49540=>"000000111",
  49541=>"000100000",
  49542=>"000111111",
  49543=>"001000000",
  49544=>"111111100",
  49545=>"001000000",
  49546=>"011000000",
  49547=>"000000111",
  49548=>"000001111",
  49549=>"000000000",
  49550=>"000000001",
  49551=>"101111011",
  49552=>"011001000",
  49553=>"111111111",
  49554=>"110111111",
  49555=>"001001011",
  49556=>"111111111",
  49557=>"000000000",
  49558=>"111111111",
  49559=>"110100001",
  49560=>"111111100",
  49561=>"010010111",
  49562=>"100111111",
  49563=>"000000000",
  49564=>"000000000",
  49565=>"100100111",
  49566=>"000110100",
  49567=>"001111111",
  49568=>"000000001",
  49569=>"111111101",
  49570=>"111101111",
  49571=>"100000000",
  49572=>"111111111",
  49573=>"000100000",
  49574=>"000000000",
  49575=>"011000000",
  49576=>"111111100",
  49577=>"000110111",
  49578=>"111111111",
  49579=>"010010111",
  49580=>"011011111",
  49581=>"000100000",
  49582=>"111111111",
  49583=>"011011111",
  49584=>"111111111",
  49585=>"000111111",
  49586=>"000000100",
  49587=>"011000000",
  49588=>"001110110",
  49589=>"111111111",
  49590=>"100100101",
  49591=>"000111010",
  49592=>"100111111",
  49593=>"000000000",
  49594=>"110110000",
  49595=>"111111101",
  49596=>"000000000",
  49597=>"111111111",
  49598=>"100000100",
  49599=>"111010000",
  49600=>"001001011",
  49601=>"000111111",
  49602=>"000000000",
  49603=>"000000111",
  49604=>"000111111",
  49605=>"001000000",
  49606=>"000000000",
  49607=>"111111000",
  49608=>"111001000",
  49609=>"011000000",
  49610=>"001000000",
  49611=>"111111111",
  49612=>"111111000",
  49613=>"010000000",
  49614=>"111111111",
  49615=>"000100111",
  49616=>"100000111",
  49617=>"011000011",
  49618=>"111011011",
  49619=>"001001001",
  49620=>"001001000",
  49621=>"011001011",
  49622=>"001010010",
  49623=>"001001000",
  49624=>"111111100",
  49625=>"000000010",
  49626=>"000001011",
  49627=>"100000000",
  49628=>"000011011",
  49629=>"110000000",
  49630=>"000000000",
  49631=>"010111011",
  49632=>"111111000",
  49633=>"111111101",
  49634=>"000001000",
  49635=>"111000000",
  49636=>"111111111",
  49637=>"000001000",
  49638=>"111111111",
  49639=>"000000001",
  49640=>"110110000",
  49641=>"011011001",
  49642=>"110100000",
  49643=>"011111100",
  49644=>"111111111",
  49645=>"001001011",
  49646=>"000000000",
  49647=>"111111111",
  49648=>"001011000",
  49649=>"000000000",
  49650=>"111111111",
  49651=>"110111111",
  49652=>"001000000",
  49653=>"111000111",
  49654=>"111111000",
  49655=>"001111100",
  49656=>"101101100",
  49657=>"000000000",
  49658=>"111111111",
  49659=>"000001111",
  49660=>"111111111",
  49661=>"000000000",
  49662=>"111111110",
  49663=>"000000000",
  49664=>"000000000",
  49665=>"111111111",
  49666=>"111000000",
  49667=>"010000110",
  49668=>"111000000",
  49669=>"100100000",
  49670=>"000000000",
  49671=>"111111111",
  49672=>"111000000",
  49673=>"001111110",
  49674=>"111111111",
  49675=>"111111111",
  49676=>"100110111",
  49677=>"001001000",
  49678=>"000000000",
  49679=>"000000000",
  49680=>"000000011",
  49681=>"111000111",
  49682=>"000000000",
  49683=>"111111111",
  49684=>"111000000",
  49685=>"111101111",
  49686=>"000000000",
  49687=>"110100100",
  49688=>"000000000",
  49689=>"000001000",
  49690=>"000000000",
  49691=>"101111111",
  49692=>"000000111",
  49693=>"010000111",
  49694=>"001001101",
  49695=>"000110010",
  49696=>"010111111",
  49697=>"011000000",
  49698=>"111111011",
  49699=>"111111000",
  49700=>"111111111",
  49701=>"111111111",
  49702=>"110100100",
  49703=>"100111000",
  49704=>"000000000",
  49705=>"011011010",
  49706=>"111111100",
  49707=>"111111111",
  49708=>"000000000",
  49709=>"111111111",
  49710=>"100110000",
  49711=>"110111111",
  49712=>"100111111",
  49713=>"000000000",
  49714=>"000000000",
  49715=>"000000001",
  49716=>"001001000",
  49717=>"111111011",
  49718=>"110111111",
  49719=>"011000100",
  49720=>"101000000",
  49721=>"000111111",
  49722=>"111111111",
  49723=>"101111111",
  49724=>"111111111",
  49725=>"011101111",
  49726=>"000011001",
  49727=>"000000000",
  49728=>"000010011",
  49729=>"111111101",
  49730=>"000000100",
  49731=>"110111000",
  49732=>"000011011",
  49733=>"111111110",
  49734=>"000000100",
  49735=>"000000001",
  49736=>"111011011",
  49737=>"111111001",
  49738=>"111111110",
  49739=>"000000110",
  49740=>"110100100",
  49741=>"110000000",
  49742=>"101000000",
  49743=>"111101000",
  49744=>"001000000",
  49745=>"111111111",
  49746=>"100101111",
  49747=>"100000000",
  49748=>"000000000",
  49749=>"000000111",
  49750=>"001100001",
  49751=>"111111111",
  49752=>"101111111",
  49753=>"010111010",
  49754=>"000000111",
  49755=>"110100000",
  49756=>"000000000",
  49757=>"111111101",
  49758=>"000001101",
  49759=>"111111111",
  49760=>"010111010",
  49761=>"000001001",
  49762=>"111111111",
  49763=>"111111000",
  49764=>"011010000",
  49765=>"000000001",
  49766=>"000000001",
  49767=>"000000000",
  49768=>"110111100",
  49769=>"110110000",
  49770=>"110111000",
  49771=>"101001101",
  49772=>"010110100",
  49773=>"111111111",
  49774=>"100101111",
  49775=>"111000101",
  49776=>"111111010",
  49777=>"000111111",
  49778=>"111111111",
  49779=>"000000100",
  49780=>"110000000",
  49781=>"100000100",
  49782=>"111111111",
  49783=>"000000000",
  49784=>"010001011",
  49785=>"000000000",
  49786=>"000000000",
  49787=>"111100000",
  49788=>"000000000",
  49789=>"111111111",
  49790=>"000000000",
  49791=>"000000000",
  49792=>"000100100",
  49793=>"111111111",
  49794=>"111011000",
  49795=>"111111011",
  49796=>"110111111",
  49797=>"000000000",
  49798=>"010010111",
  49799=>"000000011",
  49800=>"000010100",
  49801=>"001000000",
  49802=>"000000000",
  49803=>"111111111",
  49804=>"000000101",
  49805=>"101101000",
  49806=>"000000100",
  49807=>"000000000",
  49808=>"001000111",
  49809=>"101001000",
  49810=>"111001011",
  49811=>"000110111",
  49812=>"000010000",
  49813=>"111110110",
  49814=>"111000001",
  49815=>"000101111",
  49816=>"000001111",
  49817=>"111111111",
  49818=>"111101110",
  49819=>"000000000",
  49820=>"111111100",
  49821=>"110000000",
  49822=>"111111110",
  49823=>"111111000",
  49824=>"111111111",
  49825=>"000111111",
  49826=>"000000000",
  49827=>"000000000",
  49828=>"000001001",
  49829=>"000000000",
  49830=>"010111110",
  49831=>"111110110",
  49832=>"000100111",
  49833=>"000000000",
  49834=>"010011000",
  49835=>"111101101",
  49836=>"011001111",
  49837=>"110111110",
  49838=>"111101111",
  49839=>"000111011",
  49840=>"000010000",
  49841=>"111111111",
  49842=>"000001011",
  49843=>"111111111",
  49844=>"111011010",
  49845=>"100111110",
  49846=>"000000111",
  49847=>"000000110",
  49848=>"111111011",
  49849=>"100000001",
  49850=>"111111111",
  49851=>"000001001",
  49852=>"000000000",
  49853=>"000000000",
  49854=>"100000111",
  49855=>"111111111",
  49856=>"000000001",
  49857=>"000110010",
  49858=>"000001001",
  49859=>"111111011",
  49860=>"111111111",
  49861=>"000000000",
  49862=>"000000000",
  49863=>"011011111",
  49864=>"000000000",
  49865=>"111111101",
  49866=>"110111111",
  49867=>"000000000",
  49868=>"000010000",
  49869=>"100100100",
  49870=>"000000000",
  49871=>"000100111",
  49872=>"011011111",
  49873=>"111111111",
  49874=>"000111010",
  49875=>"000000000",
  49876=>"000000000",
  49877=>"001011001",
  49878=>"000110111",
  49879=>"111111011",
  49880=>"000000000",
  49881=>"011001000",
  49882=>"000001000",
  49883=>"010101010",
  49884=>"000000000",
  49885=>"000001000",
  49886=>"000100111",
  49887=>"111111000",
  49888=>"000000000",
  49889=>"111100111",
  49890=>"000111111",
  49891=>"000000000",
  49892=>"100110011",
  49893=>"110100000",
  49894=>"110111011",
  49895=>"111001111",
  49896=>"000111111",
  49897=>"100111111",
  49898=>"101000000",
  49899=>"111111111",
  49900=>"000000000",
  49901=>"101111111",
  49902=>"000110000",
  49903=>"000000000",
  49904=>"111000000",
  49905=>"111111111",
  49906=>"111111111",
  49907=>"101101101",
  49908=>"000000000",
  49909=>"111111111",
  49910=>"110111111",
  49911=>"011011111",
  49912=>"111111111",
  49913=>"000000000",
  49914=>"000000000",
  49915=>"100110000",
  49916=>"111111111",
  49917=>"000100000",
  49918=>"000000111",
  49919=>"000000000",
  49920=>"110111111",
  49921=>"111110110",
  49922=>"111110000",
  49923=>"111111111",
  49924=>"000000001",
  49925=>"111000111",
  49926=>"001011000",
  49927=>"100111011",
  49928=>"111111111",
  49929=>"110110010",
  49930=>"000000100",
  49931=>"110100000",
  49932=>"110110100",
  49933=>"100111111",
  49934=>"111111000",
  49935=>"111111111",
  49936=>"000000100",
  49937=>"010011011",
  49938=>"010011011",
  49939=>"000000000",
  49940=>"000111111",
  49941=>"000000110",
  49942=>"111111001",
  49943=>"000000111",
  49944=>"111001000",
  49945=>"000010010",
  49946=>"000000000",
  49947=>"000010000",
  49948=>"000010111",
  49949=>"000000000",
  49950=>"111111111",
  49951=>"111001111",
  49952=>"000111000",
  49953=>"001111010",
  49954=>"101100000",
  49955=>"011111111",
  49956=>"000111111",
  49957=>"000000000",
  49958=>"000001000",
  49959=>"000000101",
  49960=>"100000000",
  49961=>"000111111",
  49962=>"101101111",
  49963=>"111111111",
  49964=>"111111000",
  49965=>"011011111",
  49966=>"111111010",
  49967=>"110111111",
  49968=>"011001000",
  49969=>"000000000",
  49970=>"110111111",
  49971=>"000001111",
  49972=>"000000000",
  49973=>"000000000",
  49974=>"000000101",
  49975=>"000000101",
  49976=>"000000111",
  49977=>"100111111",
  49978=>"000000100",
  49979=>"110100110",
  49980=>"010110001",
  49981=>"010111000",
  49982=>"000000111",
  49983=>"111010000",
  49984=>"000000000",
  49985=>"111111111",
  49986=>"111111111",
  49987=>"000000000",
  49988=>"111111111",
  49989=>"111111100",
  49990=>"111111111",
  49991=>"111111111",
  49992=>"110100111",
  49993=>"010010110",
  49994=>"110100100",
  49995=>"011011011",
  49996=>"111000000",
  49997=>"111001111",
  49998=>"000111100",
  49999=>"111111111",
  50000=>"011010000",
  50001=>"000000001",
  50002=>"111111111",
  50003=>"001001001",
  50004=>"111101111",
  50005=>"001011001",
  50006=>"010100111",
  50007=>"000000001",
  50008=>"001001011",
  50009=>"111111000",
  50010=>"000000000",
  50011=>"000000010",
  50012=>"111111100",
  50013=>"110000000",
  50014=>"011111011",
  50015=>"110011111",
  50016=>"000010000",
  50017=>"000000000",
  50018=>"000111111",
  50019=>"000011011",
  50020=>"110000000",
  50021=>"000001111",
  50022=>"110111111",
  50023=>"000000111",
  50024=>"100110110",
  50025=>"111111111",
  50026=>"000000000",
  50027=>"000000000",
  50028=>"011011011",
  50029=>"110110101",
  50030=>"111111011",
  50031=>"000000010",
  50032=>"111111111",
  50033=>"000000000",
  50034=>"111110000",
  50035=>"000000000",
  50036=>"100100000",
  50037=>"110110011",
  50038=>"000000000",
  50039=>"111100101",
  50040=>"101000000",
  50041=>"111111111",
  50042=>"010111111",
  50043=>"000000110",
  50044=>"000110100",
  50045=>"000000000",
  50046=>"111101001",
  50047=>"000000000",
  50048=>"111110000",
  50049=>"100000001",
  50050=>"111111111",
  50051=>"100101111",
  50052=>"111111010",
  50053=>"110111000",
  50054=>"111000000",
  50055=>"001001101",
  50056=>"000000000",
  50057=>"000011111",
  50058=>"000001000",
  50059=>"010010000",
  50060=>"000000001",
  50061=>"111110000",
  50062=>"000001000",
  50063=>"000000010",
  50064=>"111111111",
  50065=>"111111000",
  50066=>"100100111",
  50067=>"110000000",
  50068=>"111111111",
  50069=>"011000000",
  50070=>"100000000",
  50071=>"000000000",
  50072=>"111011000",
  50073=>"000110000",
  50074=>"000000001",
  50075=>"000000100",
  50076=>"101100111",
  50077=>"011000000",
  50078=>"000000000",
  50079=>"111101101",
  50080=>"111100111",
  50081=>"110110111",
  50082=>"000000000",
  50083=>"110100100",
  50084=>"111111111",
  50085=>"011111000",
  50086=>"111111010",
  50087=>"011011111",
  50088=>"000000000",
  50089=>"111111111",
  50090=>"100001001",
  50091=>"110110010",
  50092=>"010111111",
  50093=>"000000110",
  50094=>"111000000",
  50095=>"110110000",
  50096=>"000000000",
  50097=>"000000100",
  50098=>"111111111",
  50099=>"010111010",
  50100=>"000011000",
  50101=>"101000101",
  50102=>"111111111",
  50103=>"111101101",
  50104=>"000000000",
  50105=>"101001101",
  50106=>"000010011",
  50107=>"111000000",
  50108=>"000000000",
  50109=>"111110101",
  50110=>"101000000",
  50111=>"000010010",
  50112=>"001101000",
  50113=>"000011000",
  50114=>"111111111",
  50115=>"001001001",
  50116=>"111001111",
  50117=>"010110110",
  50118=>"000000000",
  50119=>"000000000",
  50120=>"000101111",
  50121=>"000110110",
  50122=>"000000000",
  50123=>"110110111",
  50124=>"000000000",
  50125=>"000000000",
  50126=>"010110111",
  50127=>"000000000",
  50128=>"010011000",
  50129=>"111111111",
  50130=>"111111111",
  50131=>"111000101",
  50132=>"110110000",
  50133=>"000000000",
  50134=>"000100100",
  50135=>"000101111",
  50136=>"000000000",
  50137=>"000000000",
  50138=>"111110111",
  50139=>"110110110",
  50140=>"110000000",
  50141=>"000000000",
  50142=>"111111111",
  50143=>"111011001",
  50144=>"111111110",
  50145=>"111110000",
  50146=>"111101000",
  50147=>"000111111",
  50148=>"000000001",
  50149=>"000001001",
  50150=>"000000000",
  50151=>"100100101",
  50152=>"111111111",
  50153=>"111111011",
  50154=>"000000000",
  50155=>"111101000",
  50156=>"110001011",
  50157=>"001001100",
  50158=>"111111111",
  50159=>"000000000",
  50160=>"000000000",
  50161=>"111111101",
  50162=>"011001111",
  50163=>"111110010",
  50164=>"000000001",
  50165=>"110110000",
  50166=>"001111000",
  50167=>"000111001",
  50168=>"111111111",
  50169=>"000010010",
  50170=>"000000000",
  50171=>"000000111",
  50172=>"000011000",
  50173=>"111101111",
  50174=>"000010011",
  50175=>"111101111",
  50176=>"001011001",
  50177=>"000001111",
  50178=>"001111111",
  50179=>"111111000",
  50180=>"000000000",
  50181=>"100110101",
  50182=>"111111111",
  50183=>"111001111",
  50184=>"000111000",
  50185=>"111111000",
  50186=>"000000000",
  50187=>"110000000",
  50188=>"111111000",
  50189=>"100000000",
  50190=>"111111111",
  50191=>"000000000",
  50192=>"110100110",
  50193=>"010111111",
  50194=>"000010111",
  50195=>"000000000",
  50196=>"101001100",
  50197=>"111111000",
  50198=>"000010000",
  50199=>"000011010",
  50200=>"001000111",
  50201=>"000000101",
  50202=>"111001000",
  50203=>"111111110",
  50204=>"111111001",
  50205=>"101111111",
  50206=>"000000000",
  50207=>"111011000",
  50208=>"010000000",
  50209=>"000100100",
  50210=>"000000111",
  50211=>"100110000",
  50212=>"000000000",
  50213=>"000000111",
  50214=>"100111111",
  50215=>"111111000",
  50216=>"000000110",
  50217=>"111000000",
  50218=>"000011111",
  50219=>"111111111",
  50220=>"000000000",
  50221=>"000111000",
  50222=>"000000000",
  50223=>"000000111",
  50224=>"101000000",
  50225=>"010011111",
  50226=>"000000111",
  50227=>"111000101",
  50228=>"000100111",
  50229=>"000110111",
  50230=>"000000110",
  50231=>"111100000",
  50232=>"111111000",
  50233=>"000001000",
  50234=>"000000001",
  50235=>"000000000",
  50236=>"111111000",
  50237=>"000000110",
  50238=>"011001000",
  50239=>"001101111",
  50240=>"111100000",
  50241=>"111101101",
  50242=>"101111111",
  50243=>"111011111",
  50244=>"111111000",
  50245=>"000000011",
  50246=>"001000000",
  50247=>"000110111",
  50248=>"110000000",
  50249=>"111101111",
  50250=>"111101000",
  50251=>"111111111",
  50252=>"001000000",
  50253=>"110011011",
  50254=>"001001001",
  50255=>"101000000",
  50256=>"000011010",
  50257=>"111111101",
  50258=>"000011111",
  50259=>"111110100",
  50260=>"000100110",
  50261=>"111111111",
  50262=>"101000111",
  50263=>"000000000",
  50264=>"000000001",
  50265=>"000000100",
  50266=>"111111111",
  50267=>"111100100",
  50268=>"111111110",
  50269=>"000000010",
  50270=>"111100100",
  50271=>"000001011",
  50272=>"001111111",
  50273=>"000000100",
  50274=>"110111111",
  50275=>"000000000",
  50276=>"000000001",
  50277=>"111111110",
  50278=>"111111111",
  50279=>"010110111",
  50280=>"000001111",
  50281=>"000000100",
  50282=>"111001001",
  50283=>"000011111",
  50284=>"111100101",
  50285=>"000111111",
  50286=>"100100111",
  50287=>"000000000",
  50288=>"110101100",
  50289=>"000000001",
  50290=>"111111111",
  50291=>"100000001",
  50292=>"111111111",
  50293=>"110110110",
  50294=>"111111100",
  50295=>"111011000",
  50296=>"000000111",
  50297=>"000000000",
  50298=>"111110000",
  50299=>"110000000",
  50300=>"100110111",
  50301=>"100100110",
  50302=>"010111000",
  50303=>"000000000",
  50304=>"101101111",
  50305=>"000000000",
  50306=>"000101111",
  50307=>"111000000",
  50308=>"101000001",
  50309=>"111111111",
  50310=>"100000000",
  50311=>"001001000",
  50312=>"000001111",
  50313=>"111101111",
  50314=>"100000011",
  50315=>"001000111",
  50316=>"000000000",
  50317=>"000000111",
  50318=>"000001011",
  50319=>"000011111",
  50320=>"000000001",
  50321=>"000000000",
  50322=>"000000001",
  50323=>"000011111",
  50324=>"000000011",
  50325=>"110111111",
  50326=>"100000001",
  50327=>"111111100",
  50328=>"111111111",
  50329=>"000000010",
  50330=>"111111011",
  50331=>"111000000",
  50332=>"000000000",
  50333=>"000000000",
  50334=>"000000110",
  50335=>"111111000",
  50336=>"111000000",
  50337=>"111110000",
  50338=>"111011010",
  50339=>"111110011",
  50340=>"111000000",
  50341=>"001000000",
  50342=>"110111111",
  50343=>"001011111",
  50344=>"111000111",
  50345=>"000000101",
  50346=>"110100100",
  50347=>"001000000",
  50348=>"111001111",
  50349=>"110111110",
  50350=>"000000000",
  50351=>"111110000",
  50352=>"111111011",
  50353=>"000110100",
  50354=>"111011010",
  50355=>"000111110",
  50356=>"001000100",
  50357=>"000000100",
  50358=>"000001111",
  50359=>"110100000",
  50360=>"000000011",
  50361=>"111101000",
  50362=>"000110010",
  50363=>"111100110",
  50364=>"111111111",
  50365=>"000010010",
  50366=>"111111101",
  50367=>"110111110",
  50368=>"111111111",
  50369=>"011000000",
  50370=>"000000000",
  50371=>"000000000",
  50372=>"000000100",
  50373=>"000001001",
  50374=>"000110110",
  50375=>"100100111",
  50376=>"000000011",
  50377=>"111000011",
  50378=>"000100111",
  50379=>"010011111",
  50380=>"111011000",
  50381=>"001001000",
  50382=>"111110101",
  50383=>"000110111",
  50384=>"001111110",
  50385=>"001111111",
  50386=>"000000000",
  50387=>"111101100",
  50388=>"001011111",
  50389=>"000000110",
  50390=>"001101111",
  50391=>"010110111",
  50392=>"101110000",
  50393=>"001000011",
  50394=>"000000000",
  50395=>"000001000",
  50396=>"111111111",
  50397=>"000000100",
  50398=>"111111111",
  50399=>"000000111",
  50400=>"001001011",
  50401=>"001000000",
  50402=>"000011111",
  50403=>"111000001",
  50404=>"110111111",
  50405=>"110000001",
  50406=>"111111110",
  50407=>"011011011",
  50408=>"111010000",
  50409=>"000010010",
  50410=>"111111001",
  50411=>"101000000",
  50412=>"011111001",
  50413=>"100100101",
  50414=>"111101000",
  50415=>"000000000",
  50416=>"111111111",
  50417=>"111011111",
  50418=>"000000000",
  50419=>"111000110",
  50420=>"111111111",
  50421=>"000000000",
  50422=>"001001001",
  50423=>"100110111",
  50424=>"111111011",
  50425=>"000000000",
  50426=>"000000011",
  50427=>"111111111",
  50428=>"100000000",
  50429=>"001011111",
  50430=>"100000000",
  50431=>"000000111",
  50432=>"100000000",
  50433=>"111111111",
  50434=>"001000000",
  50435=>"110000000",
  50436=>"111111111",
  50437=>"111001111",
  50438=>"001000000",
  50439=>"111011111",
  50440=>"111111111",
  50441=>"100011000",
  50442=>"000000000",
  50443=>"011000001",
  50444=>"000000111",
  50445=>"111111111",
  50446=>"000000000",
  50447=>"000111111",
  50448=>"110010110",
  50449=>"111111000",
  50450=>"110000000",
  50451=>"011011110",
  50452=>"000110010",
  50453=>"011101001",
  50454=>"111111100",
  50455=>"111111111",
  50456=>"111111111",
  50457=>"011101111",
  50458=>"000000000",
  50459=>"000001000",
  50460=>"010011111",
  50461=>"011001001",
  50462=>"000011000",
  50463=>"000000101",
  50464=>"000111111",
  50465=>"110000100",
  50466=>"101111111",
  50467=>"111011000",
  50468=>"101100111",
  50469=>"000000000",
  50470=>"111111000",
  50471=>"000000000",
  50472=>"001001111",
  50473=>"011111011",
  50474=>"000111111",
  50475=>"000000101",
  50476=>"111011001",
  50477=>"010011110",
  50478=>"000000000",
  50479=>"000111011",
  50480=>"000010000",
  50481=>"000000111",
  50482=>"000110110",
  50483=>"000111111",
  50484=>"000000000",
  50485=>"111001001",
  50486=>"111111111",
  50487=>"000000000",
  50488=>"000111111",
  50489=>"111110100",
  50490=>"010111111",
  50491=>"111000000",
  50492=>"111000000",
  50493=>"110000000",
  50494=>"000110011",
  50495=>"000000000",
  50496=>"001000000",
  50497=>"000000100",
  50498=>"111100000",
  50499=>"000000000",
  50500=>"111111111",
  50501=>"111011011",
  50502=>"111111100",
  50503=>"111111111",
  50504=>"000000000",
  50505=>"000000000",
  50506=>"000000111",
  50507=>"000010001",
  50508=>"001000000",
  50509=>"111111110",
  50510=>"101000000",
  50511=>"110100111",
  50512=>"111011011",
  50513=>"101000111",
  50514=>"101111111",
  50515=>"000000000",
  50516=>"000000000",
  50517=>"011011111",
  50518=>"000001001",
  50519=>"111000100",
  50520=>"100000000",
  50521=>"001000110",
  50522=>"000000001",
  50523=>"111110110",
  50524=>"111111110",
  50525=>"111111011",
  50526=>"001001100",
  50527=>"000010111",
  50528=>"000110110",
  50529=>"000111111",
  50530=>"000011011",
  50531=>"111000000",
  50532=>"000010111",
  50533=>"000000000",
  50534=>"000001001",
  50535=>"001000110",
  50536=>"001000110",
  50537=>"001111111",
  50538=>"111001001",
  50539=>"111000100",
  50540=>"011111110",
  50541=>"111110000",
  50542=>"000000111",
  50543=>"000000011",
  50544=>"000000000",
  50545=>"000111111",
  50546=>"110110011",
  50547=>"011111111",
  50548=>"101111111",
  50549=>"000011111",
  50550=>"001011000",
  50551=>"111000100",
  50552=>"111001000",
  50553=>"000000000",
  50554=>"111000110",
  50555=>"101101111",
  50556=>"110100101",
  50557=>"000110111",
  50558=>"000011011",
  50559=>"000100000",
  50560=>"000000110",
  50561=>"101111111",
  50562=>"000001001",
  50563=>"111100111",
  50564=>"000011011",
  50565=>"000000000",
  50566=>"001001000",
  50567=>"011011001",
  50568=>"101001000",
  50569=>"110000000",
  50570=>"110100000",
  50571=>"100100100",
  50572=>"011001111",
  50573=>"000100000",
  50574=>"000000000",
  50575=>"000000111",
  50576=>"000111000",
  50577=>"110100000",
  50578=>"000100111",
  50579=>"101001001",
  50580=>"000111111",
  50581=>"000011011",
  50582=>"100100110",
  50583=>"111111110",
  50584=>"111111111",
  50585=>"101000100",
  50586=>"111111111",
  50587=>"111100111",
  50588=>"111111111",
  50589=>"000010000",
  50590=>"000111111",
  50591=>"111000000",
  50592=>"100111111",
  50593=>"000111111",
  50594=>"000000110",
  50595=>"111101111",
  50596=>"111111111",
  50597=>"110101000",
  50598=>"000001000",
  50599=>"111111000",
  50600=>"111111011",
  50601=>"111111110",
  50602=>"101000000",
  50603=>"000101111",
  50604=>"000001111",
  50605=>"000000000",
  50606=>"000000100",
  50607=>"110001011",
  50608=>"111111001",
  50609=>"111101001",
  50610=>"111111000",
  50611=>"001000000",
  50612=>"101101000",
  50613=>"111000000",
  50614=>"000011010",
  50615=>"110100000",
  50616=>"111100110",
  50617=>"111111111",
  50618=>"000000000",
  50619=>"111000000",
  50620=>"000000000",
  50621=>"111111111",
  50622=>"100111111",
  50623=>"111110110",
  50624=>"111110000",
  50625=>"111111001",
  50626=>"111000000",
  50627=>"000000000",
  50628=>"101001111",
  50629=>"111000000",
  50630=>"000000110",
  50631=>"001101111",
  50632=>"110100110",
  50633=>"101001000",
  50634=>"100000100",
  50635=>"111111110",
  50636=>"111111001",
  50637=>"111110000",
  50638=>"001111110",
  50639=>"001000000",
  50640=>"001001101",
  50641=>"110110111",
  50642=>"111100110",
  50643=>"110111111",
  50644=>"001011111",
  50645=>"100100110",
  50646=>"000000000",
  50647=>"111111000",
  50648=>"111000001",
  50649=>"000111111",
  50650=>"000000010",
  50651=>"111111111",
  50652=>"000110110",
  50653=>"110111111",
  50654=>"000000000",
  50655=>"001011000",
  50656=>"011000000",
  50657=>"111110111",
  50658=>"000000000",
  50659=>"001000000",
  50660=>"000000101",
  50661=>"000100111",
  50662=>"111101001",
  50663=>"000000000",
  50664=>"111111111",
  50665=>"111111111",
  50666=>"110000100",
  50667=>"111000000",
  50668=>"000011011",
  50669=>"011111111",
  50670=>"001000000",
  50671=>"001001000",
  50672=>"111111111",
  50673=>"000010111",
  50674=>"111111100",
  50675=>"111000000",
  50676=>"111111111",
  50677=>"001001000",
  50678=>"000000000",
  50679=>"011010000",
  50680=>"000010000",
  50681=>"111001001",
  50682=>"001000000",
  50683=>"000000000",
  50684=>"100100100",
  50685=>"101100000",
  50686=>"101100110",
  50687=>"000000111",
  50688=>"001000000",
  50689=>"010000000",
  50690=>"000000111",
  50691=>"001111011",
  50692=>"000000101",
  50693=>"001000010",
  50694=>"011111111",
  50695=>"111111000",
  50696=>"000000000",
  50697=>"000000000",
  50698=>"001111111",
  50699=>"011110100",
  50700=>"001101111",
  50701=>"000000110",
  50702=>"000001111",
  50703=>"111111100",
  50704=>"010010000",
  50705=>"111011111",
  50706=>"000000000",
  50707=>"000111111",
  50708=>"110110010",
  50709=>"110100111",
  50710=>"111111000",
  50711=>"111111101",
  50712=>"011001101",
  50713=>"000000111",
  50714=>"111111110",
  50715=>"000000000",
  50716=>"111111111",
  50717=>"000000000",
  50718=>"111011000",
  50719=>"000000100",
  50720=>"000110010",
  50721=>"111111111",
  50722=>"100000000",
  50723=>"000100100",
  50724=>"000000000",
  50725=>"100000000",
  50726=>"110000000",
  50727=>"000000110",
  50728=>"000111111",
  50729=>"000000001",
  50730=>"111101000",
  50731=>"000111111",
  50732=>"111111000",
  50733=>"100111111",
  50734=>"111001000",
  50735=>"000111111",
  50736=>"000000000",
  50737=>"111111000",
  50738=>"111111111",
  50739=>"000000000",
  50740=>"100100000",
  50741=>"011011000",
  50742=>"111111100",
  50743=>"000000000",
  50744=>"000000011",
  50745=>"111111000",
  50746=>"000000000",
  50747=>"000000000",
  50748=>"000000011",
  50749=>"111111001",
  50750=>"000000100",
  50751=>"111011000",
  50752=>"000001001",
  50753=>"000000000",
  50754=>"000000000",
  50755=>"000011111",
  50756=>"110000010",
  50757=>"000100111",
  50758=>"111000100",
  50759=>"111000000",
  50760=>"000100111",
  50761=>"000000111",
  50762=>"111111111",
  50763=>"000000111",
  50764=>"100110111",
  50765=>"011001111",
  50766=>"010010110",
  50767=>"000011111",
  50768=>"000000111",
  50769=>"000001111",
  50770=>"000000000",
  50771=>"111111000",
  50772=>"001000000",
  50773=>"000110100",
  50774=>"111100000",
  50775=>"111111111",
  50776=>"111111000",
  50777=>"101000111",
  50778=>"111001001",
  50779=>"110000000",
  50780=>"000000000",
  50781=>"000010110",
  50782=>"100000000",
  50783=>"111011001",
  50784=>"000000000",
  50785=>"000000000",
  50786=>"110010000",
  50787=>"111111111",
  50788=>"000111000",
  50789=>"000000001",
  50790=>"110110111",
  50791=>"001001000",
  50792=>"110011010",
  50793=>"111000000",
  50794=>"000000001",
  50795=>"000000000",
  50796=>"111111111",
  50797=>"010000000",
  50798=>"111110111",
  50799=>"011011000",
  50800=>"000000011",
  50801=>"000000000",
  50802=>"011011000",
  50803=>"111111001",
  50804=>"110111111",
  50805=>"011001000",
  50806=>"100011111",
  50807=>"000111111",
  50808=>"000000000",
  50809=>"000111111",
  50810=>"001000000",
  50811=>"000000111",
  50812=>"111111111",
  50813=>"000011000",
  50814=>"001000000",
  50815=>"000000011",
  50816=>"000000000",
  50817=>"000000000",
  50818=>"111111111",
  50819=>"111111000",
  50820=>"000011111",
  50821=>"000000101",
  50822=>"110110110",
  50823=>"011000000",
  50824=>"111111011",
  50825=>"000111111",
  50826=>"111111111",
  50827=>"010110000",
  50828=>"000000100",
  50829=>"110111010",
  50830=>"110100111",
  50831=>"000000111",
  50832=>"111001000",
  50833=>"011111111",
  50834=>"000111001",
  50835=>"111111111",
  50836=>"000111111",
  50837=>"110110110",
  50838=>"111100000",
  50839=>"000001110",
  50840=>"000000000",
  50841=>"000111000",
  50842=>"111111110",
  50843=>"000100000",
  50844=>"111110000",
  50845=>"001000111",
  50846=>"001001000",
  50847=>"000101111",
  50848=>"010010011",
  50849=>"011011111",
  50850=>"001001000",
  50851=>"111000111",
  50852=>"011001001",
  50853=>"111110111",
  50854=>"111111011",
  50855=>"000100100",
  50856=>"000000000",
  50857=>"000000001",
  50858=>"000000000",
  50859=>"000111111",
  50860=>"000000000",
  50861=>"100100111",
  50862=>"000000000",
  50863=>"000000000",
  50864=>"000111111",
  50865=>"000000111",
  50866=>"010111010",
  50867=>"111111000",
  50868=>"000000000",
  50869=>"011010000",
  50870=>"011111001",
  50871=>"111111111",
  50872=>"111001000",
  50873=>"000000111",
  50874=>"011000000",
  50875=>"111110110",
  50876=>"000101001",
  50877=>"111111111",
  50878=>"000100100",
  50879=>"000000000",
  50880=>"110111001",
  50881=>"111010000",
  50882=>"111111010",
  50883=>"000001000",
  50884=>"110000000",
  50885=>"111111000",
  50886=>"000001000",
  50887=>"000000011",
  50888=>"000000000",
  50889=>"111111000",
  50890=>"010110000",
  50891=>"001111111",
  50892=>"000000101",
  50893=>"000000100",
  50894=>"110111000",
  50895=>"000000000",
  50896=>"010100100",
  50897=>"000000000",
  50898=>"111011111",
  50899=>"111000000",
  50900=>"001101111",
  50901=>"111111111",
  50902=>"111001111",
  50903=>"000000000",
  50904=>"111000000",
  50905=>"110100100",
  50906=>"000011111",
  50907=>"111111101",
  50908=>"000111111",
  50909=>"111111111",
  50910=>"000011000",
  50911=>"111110000",
  50912=>"000001111",
  50913=>"000000000",
  50914=>"000000111",
  50915=>"111111111",
  50916=>"000000110",
  50917=>"000000000",
  50918=>"111111000",
  50919=>"111111111",
  50920=>"000010111",
  50921=>"001000000",
  50922=>"011111000",
  50923=>"110011011",
  50924=>"100000111",
  50925=>"000110110",
  50926=>"111111111",
  50927=>"111111111",
  50928=>"111011111",
  50929=>"011011111",
  50930=>"001111111",
  50931=>"001100001",
  50932=>"000111111",
  50933=>"111111111",
  50934=>"001101001",
  50935=>"111000000",
  50936=>"100000000",
  50937=>"000000000",
  50938=>"111111010",
  50939=>"000000000",
  50940=>"010111011",
  50941=>"001001111",
  50942=>"111110111",
  50943=>"111111111",
  50944=>"000111111",
  50945=>"100111111",
  50946=>"111111111",
  50947=>"000000000",
  50948=>"110111111",
  50949=>"000111111",
  50950=>"110100100",
  50951=>"000001111",
  50952=>"000000000",
  50953=>"111111111",
  50954=>"000000000",
  50955=>"000101111",
  50956=>"101000000",
  50957=>"000000000",
  50958=>"100000000",
  50959=>"111000000",
  50960=>"111111010",
  50961=>"000000101",
  50962=>"000000010",
  50963=>"000000000",
  50964=>"000000111",
  50965=>"110111111",
  50966=>"000000000",
  50967=>"111111111",
  50968=>"000010000",
  50969=>"000000100",
  50970=>"110110100",
  50971=>"000010010",
  50972=>"011011001",
  50973=>"111111000",
  50974=>"000000111",
  50975=>"001111111",
  50976=>"100000000",
  50977=>"101101000",
  50978=>"010111000",
  50979=>"111111011",
  50980=>"111101001",
  50981=>"000000100",
  50982=>"000111011",
  50983=>"111111011",
  50984=>"111100111",
  50985=>"000010110",
  50986=>"010000000",
  50987=>"111111001",
  50988=>"111000000",
  50989=>"000001001",
  50990=>"111000111",
  50991=>"000000000",
  50992=>"110011111",
  50993=>"111010000",
  50994=>"000000111",
  50995=>"000000000",
  50996=>"000000000",
  50997=>"111111100",
  50998=>"010010000",
  50999=>"000001000",
  51000=>"000111000",
  51001=>"111000000",
  51002=>"111110111",
  51003=>"010000111",
  51004=>"011100111",
  51005=>"111111111",
  51006=>"001111111",
  51007=>"111111111",
  51008=>"000000001",
  51009=>"101001001",
  51010=>"000100111",
  51011=>"110110100",
  51012=>"100100000",
  51013=>"111111000",
  51014=>"111111000",
  51015=>"000000000",
  51016=>"110010000",
  51017=>"011000000",
  51018=>"111111110",
  51019=>"000111100",
  51020=>"000000000",
  51021=>"111000000",
  51022=>"111111111",
  51023=>"000001111",
  51024=>"011000000",
  51025=>"000000111",
  51026=>"000000000",
  51027=>"000000000",
  51028=>"100000000",
  51029=>"011011001",
  51030=>"110111000",
  51031=>"111000000",
  51032=>"010111111",
  51033=>"101101101",
  51034=>"110111111",
  51035=>"000010000",
  51036=>"000000000",
  51037=>"001001011",
  51038=>"000000111",
  51039=>"000110110",
  51040=>"111001111",
  51041=>"001000011",
  51042=>"110111111",
  51043=>"000100000",
  51044=>"100111111",
  51045=>"000000000",
  51046=>"111111111",
  51047=>"100111111",
  51048=>"100001001",
  51049=>"011111111",
  51050=>"111111111",
  51051=>"001001001",
  51052=>"000000000",
  51053=>"111111000",
  51054=>"000000000",
  51055=>"111101111",
  51056=>"000000000",
  51057=>"000000000",
  51058=>"000000000",
  51059=>"111111011",
  51060=>"111010010",
  51061=>"111111110",
  51062=>"101000101",
  51063=>"100111111",
  51064=>"110111111",
  51065=>"000000100",
  51066=>"110111000",
  51067=>"111111010",
  51068=>"111001000",
  51069=>"111111111",
  51070=>"000010010",
  51071=>"000000000",
  51072=>"010001000",
  51073=>"010011000",
  51074=>"110110111",
  51075=>"111111111",
  51076=>"000000111",
  51077=>"000000110",
  51078=>"000100111",
  51079=>"111111001",
  51080=>"010000000",
  51081=>"111011111",
  51082=>"000000010",
  51083=>"000000000",
  51084=>"111111111",
  51085=>"100100000",
  51086=>"110110110",
  51087=>"000000111",
  51088=>"000000000",
  51089=>"000000000",
  51090=>"000000001",
  51091=>"111111111",
  51092=>"000000000",
  51093=>"000111000",
  51094=>"000000000",
  51095=>"111111000",
  51096=>"000001111",
  51097=>"000000000",
  51098=>"000000001",
  51099=>"111111110",
  51100=>"110100000",
  51101=>"000000000",
  51102=>"011000000",
  51103=>"000000110",
  51104=>"000000010",
  51105=>"000000100",
  51106=>"000100111",
  51107=>"111111000",
  51108=>"000100111",
  51109=>"000000000",
  51110=>"010000111",
  51111=>"111111110",
  51112=>"000101101",
  51113=>"000110000",
  51114=>"000100111",
  51115=>"000001001",
  51116=>"111111000",
  51117=>"000110110",
  51118=>"000000000",
  51119=>"011011000",
  51120=>"000111111",
  51121=>"111111111",
  51122=>"000111111",
  51123=>"111100000",
  51124=>"000000000",
  51125=>"000000000",
  51126=>"000000110",
  51127=>"011001010",
  51128=>"000000111",
  51129=>"011000000",
  51130=>"110100111",
  51131=>"000110110",
  51132=>"111111111",
  51133=>"110111000",
  51134=>"111100000",
  51135=>"000000000",
  51136=>"110000001",
  51137=>"000000000",
  51138=>"110111111",
  51139=>"100000000",
  51140=>"100111111",
  51141=>"000010111",
  51142=>"111111111",
  51143=>"101101001",
  51144=>"001110000",
  51145=>"011011000",
  51146=>"000000110",
  51147=>"000000011",
  51148=>"000000010",
  51149=>"000000111",
  51150=>"000111111",
  51151=>"111111111",
  51152=>"111111111",
  51153=>"010010000",
  51154=>"000100000",
  51155=>"000000111",
  51156=>"011100101",
  51157=>"110111100",
  51158=>"000010111",
  51159=>"000111000",
  51160=>"000000000",
  51161=>"000000000",
  51162=>"000000010",
  51163=>"001111111",
  51164=>"111000000",
  51165=>"011111111",
  51166=>"111011000",
  51167=>"110100111",
  51168=>"100001001",
  51169=>"000110111",
  51170=>"000110111",
  51171=>"011111111",
  51172=>"001100000",
  51173=>"000001101",
  51174=>"101111111",
  51175=>"000011011",
  51176=>"001111111",
  51177=>"111111111",
  51178=>"000000000",
  51179=>"101001000",
  51180=>"011111110",
  51181=>"000000000",
  51182=>"011010110",
  51183=>"111111111",
  51184=>"001011010",
  51185=>"010000000",
  51186=>"011001010",
  51187=>"011000000",
  51188=>"111111011",
  51189=>"000000000",
  51190=>"111111111",
  51191=>"000110110",
  51192=>"111100000",
  51193=>"001000000",
  51194=>"111111011",
  51195=>"111111000",
  51196=>"000000010",
  51197=>"110110100",
  51198=>"111111010",
  51199=>"000000101",
  51200=>"001001111",
  51201=>"111111111",
  51202=>"111111111",
  51203=>"000000000",
  51204=>"001001001",
  51205=>"111111011",
  51206=>"000000000",
  51207=>"101000111",
  51208=>"111111111",
  51209=>"111111111",
  51210=>"000001111",
  51211=>"000000000",
  51212=>"100101000",
  51213=>"001011111",
  51214=>"100100000",
  51215=>"000000000",
  51216=>"111011111",
  51217=>"000000111",
  51218=>"011011111",
  51219=>"001101111",
  51220=>"000101111",
  51221=>"000000000",
  51222=>"111111111",
  51223=>"111111111",
  51224=>"000000000",
  51225=>"000000000",
  51226=>"111011111",
  51227=>"110110101",
  51228=>"111111001",
  51229=>"000111111",
  51230=>"111111110",
  51231=>"000000000",
  51232=>"000000001",
  51233=>"000000000",
  51234=>"111001100",
  51235=>"100111111",
  51236=>"111001011",
  51237=>"111111011",
  51238=>"111111111",
  51239=>"111000000",
  51240=>"111111001",
  51241=>"111100111",
  51242=>"111111111",
  51243=>"100110110",
  51244=>"100110001",
  51245=>"111000000",
  51246=>"110111011",
  51247=>"000000000",
  51248=>"111111111",
  51249=>"111111111",
  51250=>"111111101",
  51251=>"000000000",
  51252=>"001001111",
  51253=>"100100000",
  51254=>"101100000",
  51255=>"000010111",
  51256=>"011111000",
  51257=>"110111111",
  51258=>"000000100",
  51259=>"000110000",
  51260=>"111111111",
  51261=>"100110111",
  51262=>"000111101",
  51263=>"000101001",
  51264=>"111111110",
  51265=>"000000000",
  51266=>"111111111",
  51267=>"000000000",
  51268=>"000000000",
  51269=>"010000000",
  51270=>"111111111",
  51271=>"111111111",
  51272=>"000100111",
  51273=>"001001111",
  51274=>"111111111",
  51275=>"000000000",
  51276=>"101000000",
  51277=>"000000110",
  51278=>"010100110",
  51279=>"000000111",
  51280=>"111111111",
  51281=>"000000111",
  51282=>"000011010",
  51283=>"000000000",
  51284=>"000000000",
  51285=>"011011001",
  51286=>"000010110",
  51287=>"000000010",
  51288=>"001000000",
  51289=>"111100000",
  51290=>"110111111",
  51291=>"000000000",
  51292=>"000000011",
  51293=>"000000000",
  51294=>"010000000",
  51295=>"000000000",
  51296=>"000000000",
  51297=>"000010010",
  51298=>"100111001",
  51299=>"000000000",
  51300=>"000001001",
  51301=>"000000000",
  51302=>"111111111",
  51303=>"111000001",
  51304=>"111111110",
  51305=>"111111110",
  51306=>"111111111",
  51307=>"000010011",
  51308=>"011001000",
  51309=>"001000100",
  51310=>"011001111",
  51311=>"111111011",
  51312=>"000000000",
  51313=>"100010000",
  51314=>"111111111",
  51315=>"000000000",
  51316=>"110111111",
  51317=>"111111111",
  51318=>"000000000",
  51319=>"000000000",
  51320=>"000001000",
  51321=>"011111000",
  51322=>"000010000",
  51323=>"000000000",
  51324=>"110100000",
  51325=>"111111111",
  51326=>"000000111",
  51327=>"000000000",
  51328=>"111111110",
  51329=>"000000000",
  51330=>"001001011",
  51331=>"000000000",
  51332=>"110111111",
  51333=>"000000000",
  51334=>"000000000",
  51335=>"000010011",
  51336=>"000100111",
  51337=>"111111110",
  51338=>"000000000",
  51339=>"111101111",
  51340=>"011001001",
  51341=>"000000000",
  51342=>"011000000",
  51343=>"011000000",
  51344=>"010111111",
  51345=>"111111011",
  51346=>"000010010",
  51347=>"001001000",
  51348=>"100101111",
  51349=>"110111111",
  51350=>"111111111",
  51351=>"000000000",
  51352=>"111111100",
  51353=>"111111111",
  51354=>"000110111",
  51355=>"100110100",
  51356=>"011000111",
  51357=>"000000000",
  51358=>"110110111",
  51359=>"000000000",
  51360=>"110100100",
  51361=>"111001000",
  51362=>"000000000",
  51363=>"111111111",
  51364=>"001111111",
  51365=>"110110111",
  51366=>"111111111",
  51367=>"001001000",
  51368=>"100000000",
  51369=>"000010000",
  51370=>"000000000",
  51371=>"111111111",
  51372=>"110000000",
  51373=>"110000000",
  51374=>"000111111",
  51375=>"000000001",
  51376=>"000000000",
  51377=>"000000000",
  51378=>"100000000",
  51379=>"000000011",
  51380=>"000001000",
  51381=>"011011111",
  51382=>"011101111",
  51383=>"111110000",
  51384=>"001001000",
  51385=>"010000000",
  51386=>"000000000",
  51387=>"010000000",
  51388=>"011000000",
  51389=>"111111110",
  51390=>"111111000",
  51391=>"001011000",
  51392=>"000000000",
  51393=>"111111111",
  51394=>"011111011",
  51395=>"111000000",
  51396=>"000000000",
  51397=>"111111111",
  51398=>"000000000",
  51399=>"111111111",
  51400=>"000000000",
  51401=>"000000000",
  51402=>"000000000",
  51403=>"111110000",
  51404=>"000000000",
  51405=>"110000000",
  51406=>"000000000",
  51407=>"000000000",
  51408=>"111111001",
  51409=>"110111111",
  51410=>"000000000",
  51411=>"100110111",
  51412=>"000101111",
  51413=>"000000000",
  51414=>"111111111",
  51415=>"111001111",
  51416=>"111111111",
  51417=>"000111111",
  51418=>"000111111",
  51419=>"001100100",
  51420=>"111011111",
  51421=>"000000000",
  51422=>"000000001",
  51423=>"111111111",
  51424=>"111111111",
  51425=>"111111000",
  51426=>"111110100",
  51427=>"000000111",
  51428=>"110110111",
  51429=>"000000000",
  51430=>"111111000",
  51431=>"111111111",
  51432=>"101101001",
  51433=>"000010100",
  51434=>"111011111",
  51435=>"111000111",
  51436=>"010111010",
  51437=>"111111111",
  51438=>"111111111",
  51439=>"000111111",
  51440=>"111111111",
  51441=>"000110111",
  51442=>"010001000",
  51443=>"000000000",
  51444=>"111111111",
  51445=>"000000000",
  51446=>"001101001",
  51447=>"111111111",
  51448=>"010110110",
  51449=>"000000000",
  51450=>"000111110",
  51451=>"000000000",
  51452=>"111011111",
  51453=>"110111111",
  51454=>"111111111",
  51455=>"010110110",
  51456=>"000000000",
  51457=>"100110110",
  51458=>"000011000",
  51459=>"111111000",
  51460=>"000000000",
  51461=>"000000000",
  51462=>"111111111",
  51463=>"000000011",
  51464=>"100111111",
  51465=>"000000000",
  51466=>"111111011",
  51467=>"100000000",
  51468=>"110110000",
  51469=>"000000000",
  51470=>"111111111",
  51471=>"000000000",
  51472=>"000000000",
  51473=>"011111000",
  51474=>"000000000",
  51475=>"111111001",
  51476=>"000000000",
  51477=>"000000111",
  51478=>"111111001",
  51479=>"011111111",
  51480=>"000000000",
  51481=>"111111000",
  51482=>"111111111",
  51483=>"111000110",
  51484=>"111111111",
  51485=>"001011111",
  51486=>"000000100",
  51487=>"000000000",
  51488=>"000000111",
  51489=>"000000111",
  51490=>"100101001",
  51491=>"000000000",
  51492=>"111110110",
  51493=>"001011011",
  51494=>"111000011",
  51495=>"111010011",
  51496=>"010110001",
  51497=>"000000000",
  51498=>"111011011",
  51499=>"100001001",
  51500=>"010010000",
  51501=>"000110011",
  51502=>"101000010",
  51503=>"000000000",
  51504=>"100000000",
  51505=>"000100000",
  51506=>"111111111",
  51507=>"000000001",
  51508=>"010110110",
  51509=>"111011000",
  51510=>"111111111",
  51511=>"101001111",
  51512=>"101010010",
  51513=>"111111111",
  51514=>"011111011",
  51515=>"111110000",
  51516=>"111111011",
  51517=>"010000000",
  51518=>"000101001",
  51519=>"000000000",
  51520=>"000000000",
  51521=>"111100000",
  51522=>"000000111",
  51523=>"111011000",
  51524=>"011000000",
  51525=>"111111110",
  51526=>"000001011",
  51527=>"111111111",
  51528=>"001000000",
  51529=>"000000000",
  51530=>"100000010",
  51531=>"000000000",
  51532=>"000000000",
  51533=>"000000000",
  51534=>"111111111",
  51535=>"111111111",
  51536=>"110100100",
  51537=>"000000000",
  51538=>"000000000",
  51539=>"110100101",
  51540=>"000011000",
  51541=>"011011011",
  51542=>"111111111",
  51543=>"111111001",
  51544=>"111111111",
  51545=>"100000000",
  51546=>"001000000",
  51547=>"000000000",
  51548=>"111001001",
  51549=>"001000000",
  51550=>"111111111",
  51551=>"111111011",
  51552=>"000111111",
  51553=>"000000000",
  51554=>"111111011",
  51555=>"111000111",
  51556=>"111100100",
  51557=>"111110111",
  51558=>"111111111",
  51559=>"101000001",
  51560=>"000000000",
  51561=>"111111111",
  51562=>"000000000",
  51563=>"000000000",
  51564=>"111111111",
  51565=>"000110000",
  51566=>"111110000",
  51567=>"110000000",
  51568=>"111111111",
  51569=>"101001100",
  51570=>"111111111",
  51571=>"000000000",
  51572=>"000000000",
  51573=>"100000000",
  51574=>"000000000",
  51575=>"000100100",
  51576=>"111100100",
  51577=>"111111101",
  51578=>"000010111",
  51579=>"110110100",
  51580=>"111011010",
  51581=>"101001011",
  51582=>"000000001",
  51583=>"111111111",
  51584=>"111010000",
  51585=>"111000000",
  51586=>"011011011",
  51587=>"111101101",
  51588=>"111111100",
  51589=>"000000000",
  51590=>"000000000",
  51591=>"000010001",
  51592=>"111111111",
  51593=>"000000000",
  51594=>"111111111",
  51595=>"000100100",
  51596=>"100100111",
  51597=>"000000000",
  51598=>"111111111",
  51599=>"000000000",
  51600=>"000000000",
  51601=>"100100100",
  51602=>"000010001",
  51603=>"011111111",
  51604=>"111111111",
  51605=>"000000000",
  51606=>"111111111",
  51607=>"100100100",
  51608=>"000011100",
  51609=>"000000000",
  51610=>"111111111",
  51611=>"001001001",
  51612=>"000000000",
  51613=>"000000011",
  51614=>"000000000",
  51615=>"000110111",
  51616=>"101111111",
  51617=>"111111111",
  51618=>"011000000",
  51619=>"100000000",
  51620=>"000100000",
  51621=>"111110000",
  51622=>"000111111",
  51623=>"110100000",
  51624=>"000000000",
  51625=>"111111111",
  51626=>"000000100",
  51627=>"010100000",
  51628=>"000000000",
  51629=>"110100100",
  51630=>"111111001",
  51631=>"001000000",
  51632=>"000000000",
  51633=>"011000000",
  51634=>"110111100",
  51635=>"000000011",
  51636=>"011000011",
  51637=>"111111111",
  51638=>"000010100",
  51639=>"111111111",
  51640=>"011011011",
  51641=>"001111111",
  51642=>"000000000",
  51643=>"111111001",
  51644=>"001001111",
  51645=>"000000000",
  51646=>"000001111",
  51647=>"000000000",
  51648=>"000010000",
  51649=>"000000000",
  51650=>"000000000",
  51651=>"111100100",
  51652=>"111100100",
  51653=>"111111111",
  51654=>"000010111",
  51655=>"000011111",
  51656=>"010000000",
  51657=>"000011110",
  51658=>"100000000",
  51659=>"000000000",
  51660=>"001000000",
  51661=>"000111111",
  51662=>"111111111",
  51663=>"111010111",
  51664=>"000000000",
  51665=>"011001011",
  51666=>"001000000",
  51667=>"111001011",
  51668=>"000000000",
  51669=>"111111110",
  51670=>"010000000",
  51671=>"000101011",
  51672=>"010000000",
  51673=>"010010000",
  51674=>"000000111",
  51675=>"111000000",
  51676=>"000000111",
  51677=>"111011111",
  51678=>"011011000",
  51679=>"011011111",
  51680=>"011111111",
  51681=>"111011011",
  51682=>"000000000",
  51683=>"000000100",
  51684=>"000001000",
  51685=>"010000011",
  51686=>"001001000",
  51687=>"100000000",
  51688=>"111111111",
  51689=>"011001001",
  51690=>"111011111",
  51691=>"101011011",
  51692=>"111111111",
  51693=>"111001001",
  51694=>"111111111",
  51695=>"000001001",
  51696=>"000000000",
  51697=>"000011111",
  51698=>"000000000",
  51699=>"000100100",
  51700=>"000000000",
  51701=>"010000000",
  51702=>"011000000",
  51703=>"101001101",
  51704=>"000100111",
  51705=>"110010000",
  51706=>"000000000",
  51707=>"111111111",
  51708=>"100001111",
  51709=>"111111101",
  51710=>"111111111",
  51711=>"000000000",
  51712=>"000000000",
  51713=>"111111101",
  51714=>"001100000",
  51715=>"111101000",
  51716=>"000000011",
  51717=>"110110000",
  51718=>"111000000",
  51719=>"000000000",
  51720=>"100111111",
  51721=>"000010000",
  51722=>"110111111",
  51723=>"001001101",
  51724=>"110000000",
  51725=>"001001111",
  51726=>"000000000",
  51727=>"111111000",
  51728=>"100110000",
  51729=>"000001111",
  51730=>"000000000",
  51731=>"000001011",
  51732=>"111111111",
  51733=>"111001000",
  51734=>"111111111",
  51735=>"000000110",
  51736=>"000000000",
  51737=>"011111111",
  51738=>"011111001",
  51739=>"100100100",
  51740=>"111111110",
  51741=>"111100000",
  51742=>"000000000",
  51743=>"100110111",
  51744=>"001000111",
  51745=>"000111111",
  51746=>"111000001",
  51747=>"000000111",
  51748=>"111110110",
  51749=>"101111111",
  51750=>"111111100",
  51751=>"000110111",
  51752=>"111001000",
  51753=>"111110000",
  51754=>"111111000",
  51755=>"111000000",
  51756=>"000001000",
  51757=>"111111110",
  51758=>"111111001",
  51759=>"000000111",
  51760=>"000000000",
  51761=>"111111111",
  51762=>"111001001",
  51763=>"000000000",
  51764=>"000111111",
  51765=>"000000100",
  51766=>"111111001",
  51767=>"111111001",
  51768=>"000100111",
  51769=>"101111111",
  51770=>"111111111",
  51771=>"001100100",
  51772=>"000000111",
  51773=>"011000011",
  51774=>"000000000",
  51775=>"111111111",
  51776=>"111111100",
  51777=>"111111111",
  51778=>"111111011",
  51779=>"100111001",
  51780=>"000100000",
  51781=>"001000011",
  51782=>"101111110",
  51783=>"000000000",
  51784=>"000011011",
  51785=>"111111111",
  51786=>"000000000",
  51787=>"111111111",
  51788=>"000000011",
  51789=>"101111111",
  51790=>"110110011",
  51791=>"110111100",
  51792=>"111111111",
  51793=>"000101111",
  51794=>"011111110",
  51795=>"100000111",
  51796=>"101000000",
  51797=>"011000000",
  51798=>"111100111",
  51799=>"000000101",
  51800=>"111000100",
  51801=>"001000001",
  51802=>"001001111",
  51803=>"110111011",
  51804=>"111011001",
  51805=>"110111111",
  51806=>"111111111",
  51807=>"111011000",
  51808=>"000000000",
  51809=>"011111011",
  51810=>"110000000",
  51811=>"110010000",
  51812=>"000000000",
  51813=>"111101101",
  51814=>"111001001",
  51815=>"000000000",
  51816=>"000000000",
  51817=>"000111111",
  51818=>"111001111",
  51819=>"111111001",
  51820=>"000000000",
  51821=>"111111010",
  51822=>"111111111",
  51823=>"000000000",
  51824=>"000111111",
  51825=>"000111111",
  51826=>"000000111",
  51827=>"011111100",
  51828=>"111111011",
  51829=>"000000000",
  51830=>"000010111",
  51831=>"111111111",
  51832=>"000000000",
  51833=>"111111011",
  51834=>"000000000",
  51835=>"000000000",
  51836=>"010010000",
  51837=>"111111111",
  51838=>"100110100",
  51839=>"111001000",
  51840=>"111111111",
  51841=>"111011111",
  51842=>"001011100",
  51843=>"111000111",
  51844=>"111111111",
  51845=>"000001011",
  51846=>"001001111",
  51847=>"000000000",
  51848=>"111000000",
  51849=>"000000000",
  51850=>"111111111",
  51851=>"000010111",
  51852=>"111111111",
  51853=>"110000000",
  51854=>"010010000",
  51855=>"000001000",
  51856=>"111011011",
  51857=>"000000000",
  51858=>"111000000",
  51859=>"110100000",
  51860=>"000000000",
  51861=>"010111111",
  51862=>"000000000",
  51863=>"000011000",
  51864=>"111001011",
  51865=>"001000000",
  51866=>"100111111",
  51867=>"111111111",
  51868=>"000000000",
  51869=>"111000000",
  51870=>"001001111",
  51871=>"000001001",
  51872=>"000000000",
  51873=>"111100000",
  51874=>"111111101",
  51875=>"100110000",
  51876=>"100000000",
  51877=>"111111111",
  51878=>"000111011",
  51879=>"001001000",
  51880=>"100111111",
  51881=>"111001000",
  51882=>"000000000",
  51883=>"111111111",
  51884=>"100101111",
  51885=>"110110011",
  51886=>"000000000",
  51887=>"111111000",
  51888=>"111110000",
  51889=>"011111111",
  51890=>"000100000",
  51891=>"111111111",
  51892=>"111011011",
  51893=>"110001001",
  51894=>"111111001",
  51895=>"101000000",
  51896=>"000000000",
  51897=>"000000001",
  51898=>"000000000",
  51899=>"111111111",
  51900=>"000000000",
  51901=>"000000111",
  51902=>"000110000",
  51903=>"000111101",
  51904=>"011000000",
  51905=>"000000000",
  51906=>"000100111",
  51907=>"111111000",
  51908=>"000000000",
  51909=>"000111111",
  51910=>"011001111",
  51911=>"000111111",
  51912=>"000000100",
  51913=>"100000011",
  51914=>"111111110",
  51915=>"111111111",
  51916=>"111111000",
  51917=>"111111011",
  51918=>"110111110",
  51919=>"111111110",
  51920=>"111111010",
  51921=>"000000000",
  51922=>"111111100",
  51923=>"001111111",
  51924=>"111101001",
  51925=>"000011111",
  51926=>"001001111",
  51927=>"000000000",
  51928=>"000000000",
  51929=>"111110110",
  51930=>"000000000",
  51931=>"111111111",
  51932=>"111111000",
  51933=>"001111000",
  51934=>"111111011",
  51935=>"000000111",
  51936=>"111111111",
  51937=>"000000000",
  51938=>"111110000",
  51939=>"100100011",
  51940=>"001000001",
  51941=>"011000110",
  51942=>"000000111",
  51943=>"111111111",
  51944=>"000000000",
  51945=>"010011011",
  51946=>"011011111",
  51947=>"000100001",
  51948=>"010011000",
  51949=>"010000000",
  51950=>"100010111",
  51951=>"111111110",
  51952=>"111111111",
  51953=>"111110110",
  51954=>"000000001",
  51955=>"000000011",
  51956=>"111111111",
  51957=>"111111000",
  51958=>"000000100",
  51959=>"001000000",
  51960=>"100000000",
  51961=>"010111111",
  51962=>"100111001",
  51963=>"111111011",
  51964=>"000011000",
  51965=>"101000000",
  51966=>"101000000",
  51967=>"111110111",
  51968=>"111111111",
  51969=>"100110101",
  51970=>"100010000",
  51971=>"111100000",
  51972=>"010000000",
  51973=>"111100000",
  51974=>"000000000",
  51975=>"111110111",
  51976=>"111101001",
  51977=>"000000000",
  51978=>"100000000",
  51979=>"000001111",
  51980=>"000000110",
  51981=>"000000101",
  51982=>"000000000",
  51983=>"111111111",
  51984=>"100000001",
  51985=>"000000000",
  51986=>"000000011",
  51987=>"111000110",
  51988=>"000000101",
  51989=>"000000000",
  51990=>"000000000",
  51991=>"000000001",
  51992=>"111111111",
  51993=>"111111111",
  51994=>"111111111",
  51995=>"000000000",
  51996=>"111111111",
  51997=>"000000000",
  51998=>"000000000",
  51999=>"000100111",
  52000=>"111011111",
  52001=>"000000000",
  52002=>"000000000",
  52003=>"000000000",
  52004=>"000101111",
  52005=>"111111111",
  52006=>"011110110",
  52007=>"000000000",
  52008=>"000100100",
  52009=>"000000000",
  52010=>"111111001",
  52011=>"000011000",
  52012=>"100110111",
  52013=>"101001001",
  52014=>"101000001",
  52015=>"111111111",
  52016=>"000000000",
  52017=>"110111111",
  52018=>"110111111",
  52019=>"000000000",
  52020=>"111111100",
  52021=>"111111010",
  52022=>"000111011",
  52023=>"111000001",
  52024=>"011111111",
  52025=>"111001000",
  52026=>"110110110",
  52027=>"101111011",
  52028=>"001000000",
  52029=>"000000000",
  52030=>"111111000",
  52031=>"111111101",
  52032=>"111111000",
  52033=>"111000000",
  52034=>"111111000",
  52035=>"111001001",
  52036=>"000000100",
  52037=>"111101111",
  52038=>"000000011",
  52039=>"000000000",
  52040=>"000000000",
  52041=>"000000000",
  52042=>"000100000",
  52043=>"100100000",
  52044=>"000000000",
  52045=>"000000000",
  52046=>"111000000",
  52047=>"010011101",
  52048=>"011011011",
  52049=>"110110111",
  52050=>"101000000",
  52051=>"000000111",
  52052=>"000000000",
  52053=>"001000001",
  52054=>"000100100",
  52055=>"111100000",
  52056=>"000000000",
  52057=>"111111111",
  52058=>"110110010",
  52059=>"001000001",
  52060=>"000000000",
  52061=>"000000000",
  52062=>"000000000",
  52063=>"001011111",
  52064=>"111000000",
  52065=>"000101000",
  52066=>"000001000",
  52067=>"111001001",
  52068=>"000000000",
  52069=>"000000000",
  52070=>"000000000",
  52071=>"111001000",
  52072=>"011011001",
  52073=>"111110110",
  52074=>"000000000",
  52075=>"111111101",
  52076=>"100100000",
  52077=>"101011000",
  52078=>"111101111",
  52079=>"000000000",
  52080=>"000000000",
  52081=>"010110110",
  52082=>"000111111",
  52083=>"111111111",
  52084=>"000000000",
  52085=>"111111111",
  52086=>"111000000",
  52087=>"111000111",
  52088=>"111111111",
  52089=>"111111000",
  52090=>"000000000",
  52091=>"000000110",
  52092=>"111111111",
  52093=>"111111111",
  52094=>"000000001",
  52095=>"111111111",
  52096=>"011011011",
  52097=>"000100000",
  52098=>"000000000",
  52099=>"111111111",
  52100=>"001111111",
  52101=>"111111111",
  52102=>"011001000",
  52103=>"000111111",
  52104=>"001001011",
  52105=>"110100000",
  52106=>"000111000",
  52107=>"000000000",
  52108=>"001001111",
  52109=>"100100010",
  52110=>"000000000",
  52111=>"000100000",
  52112=>"000000000",
  52113=>"000101111",
  52114=>"111111111",
  52115=>"000000000",
  52116=>"111111111",
  52117=>"111111111",
  52118=>"111101001",
  52119=>"010000000",
  52120=>"000000000",
  52121=>"110111000",
  52122=>"011011111",
  52123=>"000000001",
  52124=>"000000000",
  52125=>"101000000",
  52126=>"000000100",
  52127=>"000000000",
  52128=>"110100110",
  52129=>"001011111",
  52130=>"111001111",
  52131=>"001011111",
  52132=>"110000111",
  52133=>"111111000",
  52134=>"000000000",
  52135=>"000000000",
  52136=>"111101000",
  52137=>"000010111",
  52138=>"100000000",
  52139=>"000000111",
  52140=>"000000000",
  52141=>"000000000",
  52142=>"111111111",
  52143=>"000011011",
  52144=>"111111111",
  52145=>"001011000",
  52146=>"100000000",
  52147=>"010000000",
  52148=>"011011011",
  52149=>"000001011",
  52150=>"000000011",
  52151=>"111111111",
  52152=>"111110000",
  52153=>"011111000",
  52154=>"111000000",
  52155=>"111100000",
  52156=>"111111111",
  52157=>"111111111",
  52158=>"111111010",
  52159=>"000001011",
  52160=>"000000111",
  52161=>"000000000",
  52162=>"111011111",
  52163=>"000111111",
  52164=>"100100111",
  52165=>"111111111",
  52166=>"001001111",
  52167=>"000110100",
  52168=>"111000000",
  52169=>"001011000",
  52170=>"111111001",
  52171=>"000000000",
  52172=>"000011000",
  52173=>"111111110",
  52174=>"000100000",
  52175=>"000000000",
  52176=>"111111111",
  52177=>"111111001",
  52178=>"000000001",
  52179=>"000000111",
  52180=>"000011001",
  52181=>"000000100",
  52182=>"000100100",
  52183=>"110000000",
  52184=>"011000000",
  52185=>"000000001",
  52186=>"000000000",
  52187=>"111101101",
  52188=>"000100000",
  52189=>"001100100",
  52190=>"000000000",
  52191=>"100100111",
  52192=>"000000000",
  52193=>"001001000",
  52194=>"111111111",
  52195=>"011011010",
  52196=>"111110110",
  52197=>"011111111",
  52198=>"010111111",
  52199=>"000000000",
  52200=>"000000100",
  52201=>"000000010",
  52202=>"111111111",
  52203=>"000000000",
  52204=>"011101001",
  52205=>"001011011",
  52206=>"110111111",
  52207=>"000000111",
  52208=>"111000001",
  52209=>"111111011",
  52210=>"000111111",
  52211=>"111111110",
  52212=>"100000000",
  52213=>"000000000",
  52214=>"111111111",
  52215=>"110110111",
  52216=>"000001111",
  52217=>"011001000",
  52218=>"111110000",
  52219=>"010000000",
  52220=>"111000100",
  52221=>"000000000",
  52222=>"111111100",
  52223=>"000000011",
  52224=>"001001101",
  52225=>"000000011",
  52226=>"000100111",
  52227=>"000000000",
  52228=>"111111010",
  52229=>"011101101",
  52230=>"100000000",
  52231=>"000000001",
  52232=>"000000001",
  52233=>"000010100",
  52234=>"111111111",
  52235=>"011111101",
  52236=>"110110100",
  52237=>"100000111",
  52238=>"110111011",
  52239=>"010010000",
  52240=>"100000100",
  52241=>"010111011",
  52242=>"000000000",
  52243=>"000000000",
  52244=>"101000000",
  52245=>"000001111",
  52246=>"110110010",
  52247=>"000111100",
  52248=>"000000001",
  52249=>"100111111",
  52250=>"111101000",
  52251=>"001110100",
  52252=>"001001101",
  52253=>"011111001",
  52254=>"110001000",
  52255=>"000000100",
  52256=>"001001000",
  52257=>"101001111",
  52258=>"110110000",
  52259=>"001000001",
  52260=>"111111011",
  52261=>"100000000",
  52262=>"111111111",
  52263=>"111101000",
  52264=>"111111111",
  52265=>"000110011",
  52266=>"101001001",
  52267=>"111110000",
  52268=>"000100000",
  52269=>"010000000",
  52270=>"000000001",
  52271=>"111111000",
  52272=>"110010111",
  52273=>"010010010",
  52274=>"000000000",
  52275=>"010011011",
  52276=>"001111111",
  52277=>"010010111",
  52278=>"011000000",
  52279=>"111111011",
  52280=>"000000100",
  52281=>"011011000",
  52282=>"111111111",
  52283=>"001000111",
  52284=>"000000001",
  52285=>"000000000",
  52286=>"100000000",
  52287=>"001001101",
  52288=>"000011001",
  52289=>"111111000",
  52290=>"001001000",
  52291=>"011011000",
  52292=>"000000010",
  52293=>"001100100",
  52294=>"111010000",
  52295=>"000000110",
  52296=>"100100100",
  52297=>"011001111",
  52298=>"111111111",
  52299=>"001001000",
  52300=>"000000001",
  52301=>"000001000",
  52302=>"101101111",
  52303=>"000000000",
  52304=>"111111010",
  52305=>"111111111",
  52306=>"111111111",
  52307=>"110110111",
  52308=>"011000000",
  52309=>"000000000",
  52310=>"000101101",
  52311=>"001001001",
  52312=>"110000000",
  52313=>"111101111",
  52314=>"000000000",
  52315=>"001000000",
  52316=>"000000000",
  52317=>"111111111",
  52318=>"110110000",
  52319=>"110000111",
  52320=>"000111111",
  52321=>"111110111",
  52322=>"000000000",
  52323=>"000000000",
  52324=>"110100000",
  52325=>"011000000",
  52326=>"100111100",
  52327=>"111101100",
  52328=>"111111111",
  52329=>"000000110",
  52330=>"110010000",
  52331=>"110100000",
  52332=>"001001000",
  52333=>"010010000",
  52334=>"011001011",
  52335=>"111111111",
  52336=>"111100101",
  52337=>"101111000",
  52338=>"111100100",
  52339=>"000000111",
  52340=>"111000000",
  52341=>"101001000",
  52342=>"000000000",
  52343=>"000000001",
  52344=>"001001100",
  52345=>"000101101",
  52346=>"000000000",
  52347=>"000000000",
  52348=>"000100101",
  52349=>"001011101",
  52350=>"000000100",
  52351=>"000000000",
  52352=>"111001101",
  52353=>"101111001",
  52354=>"010111111",
  52355=>"111111000",
  52356=>"111111111",
  52357=>"101001101",
  52358=>"001001111",
  52359=>"000100111",
  52360=>"110110110",
  52361=>"000000000",
  52362=>"111101111",
  52363=>"111110111",
  52364=>"000000011",
  52365=>"111111111",
  52366=>"101000000",
  52367=>"110110010",
  52368=>"000000101",
  52369=>"111110010",
  52370=>"000111000",
  52371=>"111111111",
  52372=>"010110000",
  52373=>"000100000",
  52374=>"111001111",
  52375=>"000000111",
  52376=>"001001001",
  52377=>"001001011",
  52378=>"110111111",
  52379=>"000000000",
  52380=>"000000011",
  52381=>"001000001",
  52382=>"101001101",
  52383=>"010110111",
  52384=>"000000000",
  52385=>"001101111",
  52386=>"000000000",
  52387=>"111111111",
  52388=>"001011011",
  52389=>"110110111",
  52390=>"111111111",
  52391=>"010111111",
  52392=>"011011111",
  52393=>"111111111",
  52394=>"111111111",
  52395=>"000000101",
  52396=>"010001000",
  52397=>"111101001",
  52398=>"111111010",
  52399=>"000110111",
  52400=>"001101001",
  52401=>"001000011",
  52402=>"110111110",
  52403=>"000100111",
  52404=>"001001001",
  52405=>"001001010",
  52406=>"010110111",
  52407=>"110100111",
  52408=>"000000001",
  52409=>"111111111",
  52410=>"001001001",
  52411=>"111110010",
  52412=>"101001001",
  52413=>"001001111",
  52414=>"111101100",
  52415=>"000110110",
  52416=>"101000101",
  52417=>"000000000",
  52418=>"001101111",
  52419=>"101000100",
  52420=>"111111111",
  52421=>"000000001",
  52422=>"111000101",
  52423=>"001011000",
  52424=>"111111011",
  52425=>"000000000",
  52426=>"001000000",
  52427=>"000000000",
  52428=>"011111111",
  52429=>"001111100",
  52430=>"000000000",
  52431=>"000101000",
  52432=>"100000011",
  52433=>"000010111",
  52434=>"000000010",
  52435=>"000000000",
  52436=>"000000111",
  52437=>"000000000",
  52438=>"111001001",
  52439=>"111111011",
  52440=>"111111000",
  52441=>"111111110",
  52442=>"111111111",
  52443=>"000000000",
  52444=>"111000000",
  52445=>"001001111",
  52446=>"110110000",
  52447=>"001101101",
  52448=>"000000000",
  52449=>"010000000",
  52450=>"000000000",
  52451=>"000000000",
  52452=>"111111111",
  52453=>"010110100",
  52454=>"111111100",
  52455=>"011111111",
  52456=>"001001101",
  52457=>"111110011",
  52458=>"110110010",
  52459=>"000110011",
  52460=>"111111000",
  52461=>"000001111",
  52462=>"111111111",
  52463=>"000001001",
  52464=>"111011111",
  52465=>"010000000",
  52466=>"110010000",
  52467=>"000000000",
  52468=>"110000100",
  52469=>"011111111",
  52470=>"011111011",
  52471=>"101101101",
  52472=>"111011111",
  52473=>"001001011",
  52474=>"010111011",
  52475=>"011111111",
  52476=>"001001001",
  52477=>"011011001",
  52478=>"010000000",
  52479=>"000000001",
  52480=>"001000101",
  52481=>"001001001",
  52482=>"000000001",
  52483=>"000100111",
  52484=>"110111000",
  52485=>"000000100",
  52486=>"111111111",
  52487=>"100001001",
  52488=>"000000000",
  52489=>"001000000",
  52490=>"001111111",
  52491=>"111111010",
  52492=>"100110111",
  52493=>"111111101",
  52494=>"111111111",
  52495=>"111000000",
  52496=>"100000010",
  52497=>"000111111",
  52498=>"101101111",
  52499=>"001101100",
  52500=>"000001101",
  52501=>"000010111",
  52502=>"010110110",
  52503=>"001001100",
  52504=>"111110010",
  52505=>"111001101",
  52506=>"011011111",
  52507=>"000000000",
  52508=>"001001001",
  52509=>"111111111",
  52510=>"101100101",
  52511=>"001111111",
  52512=>"110111000",
  52513=>"000001000",
  52514=>"111111000",
  52515=>"000000101",
  52516=>"000110111",
  52517=>"111111110",
  52518=>"011001000",
  52519=>"000000100",
  52520=>"000111111",
  52521=>"000000000",
  52522=>"000110110",
  52523=>"111100100",
  52524=>"000100000",
  52525=>"000000000",
  52526=>"101001001",
  52527=>"000000000",
  52528=>"110110111",
  52529=>"111011000",
  52530=>"011111111",
  52531=>"000000000",
  52532=>"010000000",
  52533=>"011011110",
  52534=>"010110000",
  52535=>"001011000",
  52536=>"000110110",
  52537=>"010000111",
  52538=>"001001001",
  52539=>"111001000",
  52540=>"111100100",
  52541=>"110111111",
  52542=>"001001101",
  52543=>"111111010",
  52544=>"000000000",
  52545=>"000001001",
  52546=>"000000110",
  52547=>"001001111",
  52548=>"111110010",
  52549=>"010001001",
  52550=>"000000000",
  52551=>"111110010",
  52552=>"010111011",
  52553=>"000000000",
  52554=>"000000001",
  52555=>"111111111",
  52556=>"110111101",
  52557=>"010011011",
  52558=>"000000001",
  52559=>"000010111",
  52560=>"000000110",
  52561=>"000001000",
  52562=>"111111111",
  52563=>"000000000",
  52564=>"111111001",
  52565=>"001011001",
  52566=>"000000111",
  52567=>"010010111",
  52568=>"111111111",
  52569=>"000000000",
  52570=>"000000000",
  52571=>"111111011",
  52572=>"000000000",
  52573=>"000001110",
  52574=>"111111111",
  52575=>"000100110",
  52576=>"000110111",
  52577=>"000000000",
  52578=>"111111011",
  52579=>"101001011",
  52580=>"101111111",
  52581=>"010110000",
  52582=>"000000000",
  52583=>"001001000",
  52584=>"111111110",
  52585=>"000000000",
  52586=>"000000000",
  52587=>"000001000",
  52588=>"110110110",
  52589=>"001001011",
  52590=>"111001000",
  52591=>"111100110",
  52592=>"001001000",
  52593=>"000000000",
  52594=>"111111111",
  52595=>"111111011",
  52596=>"000000000",
  52597=>"001001111",
  52598=>"001001001",
  52599=>"110110000",
  52600=>"111101111",
  52601=>"011000010",
  52602=>"000000000",
  52603=>"000001100",
  52604=>"010100100",
  52605=>"001001001",
  52606=>"111111000",
  52607=>"111111111",
  52608=>"100110110",
  52609=>"000000000",
  52610=>"000001001",
  52611=>"111111111",
  52612=>"000100111",
  52613=>"000011001",
  52614=>"000000000",
  52615=>"000101111",
  52616=>"001001111",
  52617=>"000000000",
  52618=>"000001101",
  52619=>"000000000",
  52620=>"000000011",
  52621=>"110111111",
  52622=>"001000100",
  52623=>"110111110",
  52624=>"111111001",
  52625=>"000000000",
  52626=>"101111001",
  52627=>"111011011",
  52628=>"111111011",
  52629=>"000000000",
  52630=>"000000000",
  52631=>"011111001",
  52632=>"000000001",
  52633=>"000000000",
  52634=>"011000000",
  52635=>"110111010",
  52636=>"000000000",
  52637=>"010010110",
  52638=>"000001001",
  52639=>"000000000",
  52640=>"000000101",
  52641=>"010110110",
  52642=>"100111111",
  52643=>"111001101",
  52644=>"111001000",
  52645=>"110111111",
  52646=>"000000000",
  52647=>"111011101",
  52648=>"111111111",
  52649=>"111111111",
  52650=>"110010001",
  52651=>"001110100",
  52652=>"000001001",
  52653=>"000000001",
  52654=>"111010000",
  52655=>"000000000",
  52656=>"000000000",
  52657=>"001000000",
  52658=>"010000110",
  52659=>"000000000",
  52660=>"000000001",
  52661=>"010000000",
  52662=>"111111100",
  52663=>"000000000",
  52664=>"001110110",
  52665=>"010111110",
  52666=>"101101111",
  52667=>"100110000",
  52668=>"000000001",
  52669=>"111011111",
  52670=>"000000000",
  52671=>"111001101",
  52672=>"010000101",
  52673=>"000000000",
  52674=>"000000101",
  52675=>"000111000",
  52676=>"000000000",
  52677=>"010011000",
  52678=>"010010000",
  52679=>"111111011",
  52680=>"111011000",
  52681=>"000010010",
  52682=>"101001111",
  52683=>"111111111",
  52684=>"110000000",
  52685=>"111111001",
  52686=>"000010011",
  52687=>"000000110",
  52688=>"000000000",
  52689=>"110111111",
  52690=>"111111111",
  52691=>"111110000",
  52692=>"111111000",
  52693=>"110100000",
  52694=>"000000000",
  52695=>"011111111",
  52696=>"010110010",
  52697=>"001001000",
  52698=>"001101110",
  52699=>"000000000",
  52700=>"000000001",
  52701=>"100111111",
  52702=>"001000000",
  52703=>"001001001",
  52704=>"000000000",
  52705=>"001001001",
  52706=>"000000000",
  52707=>"111111100",
  52708=>"001000000",
  52709=>"000001000",
  52710=>"000000111",
  52711=>"000000011",
  52712=>"111111010",
  52713=>"111111110",
  52714=>"111101100",
  52715=>"000111111",
  52716=>"111111111",
  52717=>"111010000",
  52718=>"000000010",
  52719=>"101000000",
  52720=>"000101101",
  52721=>"001111111",
  52722=>"101101100",
  52723=>"111110000",
  52724=>"000000001",
  52725=>"000010010",
  52726=>"011001111",
  52727=>"000110110",
  52728=>"000000000",
  52729=>"110010110",
  52730=>"111111011",
  52731=>"000000001",
  52732=>"001000000",
  52733=>"000000010",
  52734=>"111011000",
  52735=>"001001010",
  52736=>"000000000",
  52737=>"000000000",
  52738=>"000000000",
  52739=>"000000000",
  52740=>"000011111",
  52741=>"111111100",
  52742=>"000000000",
  52743=>"000000000",
  52744=>"000010101",
  52745=>"010110111",
  52746=>"000000000",
  52747=>"100100000",
  52748=>"000000001",
  52749=>"111111111",
  52750=>"111000111",
  52751=>"111111111",
  52752=>"110110100",
  52753=>"000111010",
  52754=>"000000101",
  52755=>"111111111",
  52756=>"000000000",
  52757=>"111001001",
  52758=>"000100100",
  52759=>"100111111",
  52760=>"100111111",
  52761=>"000000100",
  52762=>"111101101",
  52763=>"000000000",
  52764=>"101001001",
  52765=>"101100000",
  52766=>"001111111",
  52767=>"000001000",
  52768=>"101110111",
  52769=>"111111111",
  52770=>"000000000",
  52771=>"000000001",
  52772=>"000000000",
  52773=>"000000000",
  52774=>"000000000",
  52775=>"111111000",
  52776=>"001101100",
  52777=>"000000000",
  52778=>"000000000",
  52779=>"000000000",
  52780=>"000000000",
  52781=>"000000011",
  52782=>"110111111",
  52783=>"110010000",
  52784=>"000000000",
  52785=>"100100100",
  52786=>"001101110",
  52787=>"011011011",
  52788=>"000000001",
  52789=>"001111101",
  52790=>"000000000",
  52791=>"001111100",
  52792=>"111111111",
  52793=>"100110000",
  52794=>"000000000",
  52795=>"011000010",
  52796=>"000111111",
  52797=>"000100000",
  52798=>"111000000",
  52799=>"111000000",
  52800=>"100100111",
  52801=>"000111111",
  52802=>"000000000",
  52803=>"000000000",
  52804=>"100110110",
  52805=>"111111110",
  52806=>"000000011",
  52807=>"111111111",
  52808=>"011110111",
  52809=>"000000101",
  52810=>"111110111",
  52811=>"111111111",
  52812=>"011111100",
  52813=>"110110010",
  52814=>"000000001",
  52815=>"111111111",
  52816=>"000000000",
  52817=>"111111111",
  52818=>"000000110",
  52819=>"000000100",
  52820=>"000000000",
  52821=>"111111111",
  52822=>"100100000",
  52823=>"100100000",
  52824=>"000000111",
  52825=>"000000000",
  52826=>"111111110",
  52827=>"001000001",
  52828=>"010000111",
  52829=>"111111001",
  52830=>"000000000",
  52831=>"110110110",
  52832=>"111101111",
  52833=>"100100000",
  52834=>"000000000",
  52835=>"111111111",
  52836=>"111001111",
  52837=>"111000000",
  52838=>"000011111",
  52839=>"000000000",
  52840=>"111000000",
  52841=>"001111111",
  52842=>"001000000",
  52843=>"110011000",
  52844=>"110000000",
  52845=>"000000000",
  52846=>"111111001",
  52847=>"000010010",
  52848=>"111111011",
  52849=>"000000100",
  52850=>"000111111",
  52851=>"000001111",
  52852=>"000000000",
  52853=>"000000000",
  52854=>"000011111",
  52855=>"110110111",
  52856=>"000000000",
  52857=>"100001111",
  52858=>"100000000",
  52859=>"000100000",
  52860=>"111110110",
  52861=>"000000000",
  52862=>"110111111",
  52863=>"111111111",
  52864=>"011011111",
  52865=>"110000000",
  52866=>"000000011",
  52867=>"111111111",
  52868=>"111111010",
  52869=>"000000000",
  52870=>"000001000",
  52871=>"000000111",
  52872=>"000000111",
  52873=>"011000000",
  52874=>"111111111",
  52875=>"100000000",
  52876=>"000000000",
  52877=>"000000000",
  52878=>"001011000",
  52879=>"000000000",
  52880=>"000000011",
  52881=>"001000000",
  52882=>"000010000",
  52883=>"111110000",
  52884=>"100000000",
  52885=>"000000000",
  52886=>"010000000",
  52887=>"111111111",
  52888=>"000000000",
  52889=>"111111111",
  52890=>"111111111",
  52891=>"000111111",
  52892=>"000101001",
  52893=>"000000111",
  52894=>"000000000",
  52895=>"111111111",
  52896=>"000000000",
  52897=>"000111111",
  52898=>"000010111",
  52899=>"111111111",
  52900=>"000000100",
  52901=>"000111011",
  52902=>"000000001",
  52903=>"110110111",
  52904=>"100111111",
  52905=>"110000000",
  52906=>"000000000",
  52907=>"111111111",
  52908=>"000110111",
  52909=>"001111111",
  52910=>"011000000",
  52911=>"110011000",
  52912=>"000100000",
  52913=>"000001010",
  52914=>"111111111",
  52915=>"010001111",
  52916=>"110111111",
  52917=>"111111111",
  52918=>"111111111",
  52919=>"011001001",
  52920=>"000000000",
  52921=>"000000000",
  52922=>"000100100",
  52923=>"011011000",
  52924=>"100100000",
  52925=>"111111111",
  52926=>"111111111",
  52927=>"000000000",
  52928=>"101100001",
  52929=>"000001111",
  52930=>"011001001",
  52931=>"111001000",
  52932=>"111111111",
  52933=>"111011001",
  52934=>"001001000",
  52935=>"100111111",
  52936=>"000111110",
  52937=>"101000000",
  52938=>"100110000",
  52939=>"111111111",
  52940=>"111111000",
  52941=>"000000000",
  52942=>"000001111",
  52943=>"000000000",
  52944=>"111111111",
  52945=>"000000000",
  52946=>"100001111",
  52947=>"100100000",
  52948=>"000000000",
  52949=>"110110111",
  52950=>"001000000",
  52951=>"000000000",
  52952=>"000000110",
  52953=>"000000001",
  52954=>"000000110",
  52955=>"111011000",
  52956=>"111101111",
  52957=>"111111001",
  52958=>"111111111",
  52959=>"100110000",
  52960=>"000000000",
  52961=>"000000010",
  52962=>"000111111",
  52963=>"111111111",
  52964=>"110111111",
  52965=>"110110100",
  52966=>"000101111",
  52967=>"111111111",
  52968=>"111111111",
  52969=>"111000001",
  52970=>"111111111",
  52971=>"100000000",
  52972=>"110111111",
  52973=>"000000101",
  52974=>"000000000",
  52975=>"000000100",
  52976=>"110010010",
  52977=>"110111111",
  52978=>"111111001",
  52979=>"001001000",
  52980=>"000100111",
  52981=>"011111011",
  52982=>"000001111",
  52983=>"110001001",
  52984=>"000000000",
  52985=>"000000011",
  52986=>"001101000",
  52987=>"011001000",
  52988=>"011011111",
  52989=>"011001111",
  52990=>"000000001",
  52991=>"000000000",
  52992=>"000000000",
  52993=>"100100101",
  52994=>"000000000",
  52995=>"111111111",
  52996=>"000000011",
  52997=>"001011011",
  52998=>"000000000",
  52999=>"000100000",
  53000=>"000000111",
  53001=>"000000000",
  53002=>"111111111",
  53003=>"000000111",
  53004=>"111111111",
  53005=>"000011111",
  53006=>"001111111",
  53007=>"110000000",
  53008=>"110111111",
  53009=>"000000000",
  53010=>"000000000",
  53011=>"000111110",
  53012=>"111000000",
  53013=>"001000100",
  53014=>"100111001",
  53015=>"001111100",
  53016=>"111111111",
  53017=>"000000100",
  53018=>"111110010",
  53019=>"000000000",
  53020=>"001111011",
  53021=>"001001111",
  53022=>"000000000",
  53023=>"111011111",
  53024=>"000100011",
  53025=>"011001111",
  53026=>"011000000",
  53027=>"011000000",
  53028=>"111111111",
  53029=>"000100111",
  53030=>"111001000",
  53031=>"101101110",
  53032=>"000000000",
  53033=>"000000010",
  53034=>"001000000",
  53035=>"000000000",
  53036=>"111111000",
  53037=>"001001111",
  53038=>"101101000",
  53039=>"100000100",
  53040=>"111111110",
  53041=>"011111000",
  53042=>"000111010",
  53043=>"000000000",
  53044=>"000100000",
  53045=>"000000000",
  53046=>"000011011",
  53047=>"010011011",
  53048=>"111011000",
  53049=>"111000000",
  53050=>"000000010",
  53051=>"110000111",
  53052=>"100000000",
  53053=>"000111111",
  53054=>"000000000",
  53055=>"001111011",
  53056=>"111000000",
  53057=>"111111111",
  53058=>"000000101",
  53059=>"000001111",
  53060=>"101010111",
  53061=>"000000000",
  53062=>"000000000",
  53063=>"101100111",
  53064=>"000000000",
  53065=>"000000011",
  53066=>"100000111",
  53067=>"111011001",
  53068=>"000000000",
  53069=>"011011000",
  53070=>"111111111",
  53071=>"000000000",
  53072=>"110110000",
  53073=>"101111111",
  53074=>"110111111",
  53075=>"100111100",
  53076=>"000000111",
  53077=>"011011001",
  53078=>"111010000",
  53079=>"001001001",
  53080=>"001011001",
  53081=>"111111111",
  53082=>"111110111",
  53083=>"111111111",
  53084=>"000011001",
  53085=>"010111111",
  53086=>"111111011",
  53087=>"000000110",
  53088=>"111111111",
  53089=>"111011011",
  53090=>"001000101",
  53091=>"101000000",
  53092=>"111111111",
  53093=>"000000000",
  53094=>"010111111",
  53095=>"111111111",
  53096=>"101111001",
  53097=>"111011010",
  53098=>"000100111",
  53099=>"111001001",
  53100=>"000000110",
  53101=>"000000101",
  53102=>"110100000",
  53103=>"000000000",
  53104=>"110110110",
  53105=>"110010000",
  53106=>"111000000",
  53107=>"110111101",
  53108=>"000110110",
  53109=>"110110111",
  53110=>"100000111",
  53111=>"110110110",
  53112=>"111100000",
  53113=>"110111111",
  53114=>"000000011",
  53115=>"100111000",
  53116=>"011111111",
  53117=>"110111111",
  53118=>"000001011",
  53119=>"111001101",
  53120=>"111111111",
  53121=>"111111000",
  53122=>"111111111",
  53123=>"111111111",
  53124=>"000010111",
  53125=>"000001001",
  53126=>"011000000",
  53127=>"011000111",
  53128=>"000000000",
  53129=>"011011001",
  53130=>"000000000",
  53131=>"111111000",
  53132=>"111111110",
  53133=>"000000011",
  53134=>"111111111",
  53135=>"010000111",
  53136=>"000000000",
  53137=>"000000000",
  53138=>"000000001",
  53139=>"000001001",
  53140=>"111000000",
  53141=>"000010000",
  53142=>"110000000",
  53143=>"111111111",
  53144=>"000000000",
  53145=>"110111000",
  53146=>"111111111",
  53147=>"000000000",
  53148=>"110010110",
  53149=>"111111111",
  53150=>"111000000",
  53151=>"100000000",
  53152=>"000100110",
  53153=>"111110111",
  53154=>"001111111",
  53155=>"100111111",
  53156=>"001001111",
  53157=>"000000000",
  53158=>"001111011",
  53159=>"000111111",
  53160=>"010001001",
  53161=>"000000000",
  53162=>"000000000",
  53163=>"100100000",
  53164=>"000000000",
  53165=>"101101000",
  53166=>"110110000",
  53167=>"100101000",
  53168=>"111001000",
  53169=>"001001101",
  53170=>"100100000",
  53171=>"001011010",
  53172=>"111111111",
  53173=>"000000000",
  53174=>"000111111",
  53175=>"111001111",
  53176=>"110111011",
  53177=>"000001000",
  53178=>"000000111",
  53179=>"000011111",
  53180=>"011001001",
  53181=>"111111111",
  53182=>"111000000",
  53183=>"111111111",
  53184=>"111010000",
  53185=>"001000111",
  53186=>"111111111",
  53187=>"111000000",
  53188=>"000111000",
  53189=>"000110111",
  53190=>"111111111",
  53191=>"001001000",
  53192=>"000111111",
  53193=>"111111111",
  53194=>"000000000",
  53195=>"001111111",
  53196=>"000000000",
  53197=>"100000010",
  53198=>"111111111",
  53199=>"000111111",
  53200=>"111111000",
  53201=>"001000000",
  53202=>"000000011",
  53203=>"110110111",
  53204=>"011111001",
  53205=>"110111111",
  53206=>"000000000",
  53207=>"000000000",
  53208=>"000011111",
  53209=>"000000000",
  53210=>"111111110",
  53211=>"101111111",
  53212=>"011111111",
  53213=>"111111111",
  53214=>"100000001",
  53215=>"001111001",
  53216=>"101100111",
  53217=>"000111111",
  53218=>"111111101",
  53219=>"111111111",
  53220=>"111011000",
  53221=>"000000000",
  53222=>"001111111",
  53223=>"000000000",
  53224=>"111110110",
  53225=>"010000000",
  53226=>"111000000",
  53227=>"111111111",
  53228=>"111111111",
  53229=>"110111111",
  53230=>"000000001",
  53231=>"000000000",
  53232=>"110100000",
  53233=>"000111111",
  53234=>"101110110",
  53235=>"111111111",
  53236=>"000000000",
  53237=>"001000000",
  53238=>"111000000",
  53239=>"110010000",
  53240=>"100110000",
  53241=>"111111111",
  53242=>"111111111",
  53243=>"010000000",
  53244=>"001101111",
  53245=>"111111110",
  53246=>"000100001",
  53247=>"000111111",
  53248=>"100100111",
  53249=>"110110111",
  53250=>"101111111",
  53251=>"111111111",
  53252=>"111011000",
  53253=>"010111001",
  53254=>"111011110",
  53255=>"100111111",
  53256=>"101100100",
  53257=>"000000001",
  53258=>"000000101",
  53259=>"111001111",
  53260=>"111111111",
  53261=>"001000111",
  53262=>"000000111",
  53263=>"001111110",
  53264=>"001111100",
  53265=>"000000111",
  53266=>"001001001",
  53267=>"000000111",
  53268=>"110000111",
  53269=>"111110000",
  53270=>"100000000",
  53271=>"100111111",
  53272=>"000000100",
  53273=>"011111001",
  53274=>"110111000",
  53275=>"011011111",
  53276=>"000001111",
  53277=>"111011111",
  53278=>"000000001",
  53279=>"111111111",
  53280=>"111110110",
  53281=>"111110111",
  53282=>"011011000",
  53283=>"001000111",
  53284=>"000000111",
  53285=>"111110011",
  53286=>"100111111",
  53287=>"111000111",
  53288=>"111000000",
  53289=>"111011011",
  53290=>"111111111",
  53291=>"010010111",
  53292=>"111111010",
  53293=>"111111010",
  53294=>"000111111",
  53295=>"000000000",
  53296=>"100111111",
  53297=>"100000000",
  53298=>"100000000",
  53299=>"000000111",
  53300=>"011011000",
  53301=>"111111000",
  53302=>"111111011",
  53303=>"110010000",
  53304=>"000000011",
  53305=>"001001111",
  53306=>"111111111",
  53307=>"000000010",
  53308=>"000001111",
  53309=>"111111000",
  53310=>"000000111",
  53311=>"010111000",
  53312=>"000000000",
  53313=>"000001111",
  53314=>"111101000",
  53315=>"000011111",
  53316=>"001001000",
  53317=>"011011111",
  53318=>"000000001",
  53319=>"000000000",
  53320=>"110110000",
  53321=>"011101111",
  53322=>"000000011",
  53323=>"000000000",
  53324=>"011011100",
  53325=>"100100111",
  53326=>"011011011",
  53327=>"000000100",
  53328=>"111111000",
  53329=>"000000000",
  53330=>"000011011",
  53331=>"000000000",
  53332=>"010000000",
  53333=>"000000111",
  53334=>"111111010",
  53335=>"111100000",
  53336=>"111001001",
  53337=>"000100111",
  53338=>"110111000",
  53339=>"000000000",
  53340=>"000000011",
  53341=>"000110111",
  53342=>"000000101",
  53343=>"000000001",
  53344=>"011011111",
  53345=>"000000000",
  53346=>"100101111",
  53347=>"111111111",
  53348=>"011000000",
  53349=>"100000000",
  53350=>"001001111",
  53351=>"111001001",
  53352=>"111111111",
  53353=>"110100110",
  53354=>"111100011",
  53355=>"111110000",
  53356=>"000000111",
  53357=>"000011111",
  53358=>"000000101",
  53359=>"011111111",
  53360=>"001111000",
  53361=>"110000101",
  53362=>"101001000",
  53363=>"010010111",
  53364=>"000000000",
  53365=>"000000000",
  53366=>"100100000",
  53367=>"000000000",
  53368=>"000000000",
  53369=>"001101110",
  53370=>"000000101",
  53371=>"000000111",
  53372=>"100000000",
  53373=>"000000000",
  53374=>"100000000",
  53375=>"000000110",
  53376=>"111111000",
  53377=>"111000000",
  53378=>"100111111",
  53379=>"000000011",
  53380=>"000000111",
  53381=>"111111000",
  53382=>"000010100",
  53383=>"000111111",
  53384=>"111111100",
  53385=>"000000001",
  53386=>"111111111",
  53387=>"011111111",
  53388=>"101000000",
  53389=>"111111110",
  53390=>"111000000",
  53391=>"111111111",
  53392=>"000000100",
  53393=>"111000000",
  53394=>"111011000",
  53395=>"001000001",
  53396=>"000111111",
  53397=>"100110111",
  53398=>"000111111",
  53399=>"000000000",
  53400=>"101000000",
  53401=>"101001111",
  53402=>"000000111",
  53403=>"001100100",
  53404=>"111010000",
  53405=>"110010000",
  53406=>"111011000",
  53407=>"111001000",
  53408=>"000000000",
  53409=>"111111001",
  53410=>"110111111",
  53411=>"001001011",
  53412=>"000000000",
  53413=>"000111111",
  53414=>"000000111",
  53415=>"111111000",
  53416=>"000000111",
  53417=>"000000100",
  53418=>"111000000",
  53419=>"000000111",
  53420=>"111011011",
  53421=>"100100111",
  53422=>"010111110",
  53423=>"000111111",
  53424=>"111111111",
  53425=>"111101001",
  53426=>"010111111",
  53427=>"111111101",
  53428=>"100000000",
  53429=>"000000001",
  53430=>"000000001",
  53431=>"111111011",
  53432=>"110110111",
  53433=>"011011111",
  53434=>"000000000",
  53435=>"001000000",
  53436=>"000000000",
  53437=>"111011111",
  53438=>"000111111",
  53439=>"111000000",
  53440=>"101111111",
  53441=>"111111111",
  53442=>"011011000",
  53443=>"101111000",
  53444=>"111111110",
  53445=>"101000000",
  53446=>"110110000",
  53447=>"110010000",
  53448=>"000000010",
  53449=>"000000000",
  53450=>"100000001",
  53451=>"111000000",
  53452=>"000000000",
  53453=>"000000000",
  53454=>"000000000",
  53455=>"000111111",
  53456=>"111000000",
  53457=>"001110111",
  53458=>"000000110",
  53459=>"001000000",
  53460=>"000001011",
  53461=>"000000110",
  53462=>"001111111",
  53463=>"001001101",
  53464=>"111111011",
  53465=>"110111110",
  53466=>"111011111",
  53467=>"000010010",
  53468=>"111111111",
  53469=>"000000000",
  53470=>"000101111",
  53471=>"011000000",
  53472=>"111000001",
  53473=>"000000010",
  53474=>"111000000",
  53475=>"011011010",
  53476=>"111011000",
  53477=>"000000000",
  53478=>"000111111",
  53479=>"000000000",
  53480=>"111111011",
  53481=>"111011111",
  53482=>"001000000",
  53483=>"001000111",
  53484=>"000001001",
  53485=>"111111111",
  53486=>"111111111",
  53487=>"000111111",
  53488=>"000000000",
  53489=>"111111001",
  53490=>"000000000",
  53491=>"000010001",
  53492=>"111111111",
  53493=>"010000000",
  53494=>"001111000",
  53495=>"111001000",
  53496=>"001001111",
  53497=>"110111111",
  53498=>"001000000",
  53499=>"111111110",
  53500=>"001000000",
  53501=>"000010000",
  53502=>"000000001",
  53503=>"010111111",
  53504=>"111000000",
  53505=>"110110000",
  53506=>"111111111",
  53507=>"000000111",
  53508=>"001000000",
  53509=>"111111111",
  53510=>"100111000",
  53511=>"000011101",
  53512=>"100000000",
  53513=>"111010010",
  53514=>"000010100",
  53515=>"111111110",
  53516=>"110110110",
  53517=>"100000000",
  53518=>"100000000",
  53519=>"011111010",
  53520=>"000111111",
  53521=>"111000000",
  53522=>"000000000",
  53523=>"110110000",
  53524=>"111111000",
  53525=>"100100111",
  53526=>"111111111",
  53527=>"001100000",
  53528=>"000001000",
  53529=>"000000000",
  53530=>"111111010",
  53531=>"111000000",
  53532=>"111111111",
  53533=>"011011001",
  53534=>"000001000",
  53535=>"010111111",
  53536=>"000000101",
  53537=>"100000000",
  53538=>"000000000",
  53539=>"000000100",
  53540=>"000000111",
  53541=>"111100100",
  53542=>"111011011",
  53543=>"001011011",
  53544=>"000111111",
  53545=>"000000000",
  53546=>"111111000",
  53547=>"000000100",
  53548=>"000110111",
  53549=>"000110001",
  53550=>"111111000",
  53551=>"000000000",
  53552=>"110111111",
  53553=>"100000000",
  53554=>"111001111",
  53555=>"000001111",
  53556=>"000100000",
  53557=>"111000000",
  53558=>"011000000",
  53559=>"111011111",
  53560=>"010000000",
  53561=>"100100000",
  53562=>"000000001",
  53563=>"111100110",
  53564=>"000010011",
  53565=>"110111011",
  53566=>"011111111",
  53567=>"111111101",
  53568=>"111111000",
  53569=>"001111110",
  53570=>"011000111",
  53571=>"111011000",
  53572=>"001001111",
  53573=>"000000100",
  53574=>"100100011",
  53575=>"111111000",
  53576=>"000000001",
  53577=>"000000101",
  53578=>"100110110",
  53579=>"010000000",
  53580=>"110010001",
  53581=>"111111111",
  53582=>"000000111",
  53583=>"001011001",
  53584=>"000100111",
  53585=>"000000111",
  53586=>"000000000",
  53587=>"111011111",
  53588=>"000000000",
  53589=>"011011011",
  53590=>"000000111",
  53591=>"101110000",
  53592=>"000110110",
  53593=>"001111110",
  53594=>"000100101",
  53595=>"100100110",
  53596=>"100000000",
  53597=>"000101111",
  53598=>"111111111",
  53599=>"110001000",
  53600=>"000000000",
  53601=>"000000000",
  53602=>"000000100",
  53603=>"111000001",
  53604=>"111001001",
  53605=>"000000000",
  53606=>"111011111",
  53607=>"000000000",
  53608=>"000000001",
  53609=>"111011001",
  53610=>"010111111",
  53611=>"000000001",
  53612=>"111111111",
  53613=>"000000001",
  53614=>"111001111",
  53615=>"000000111",
  53616=>"000001111",
  53617=>"001111111",
  53618=>"110000000",
  53619=>"001000000",
  53620=>"000000000",
  53621=>"000000000",
  53622=>"000000000",
  53623=>"000000000",
  53624=>"011000000",
  53625=>"100111111",
  53626=>"111110000",
  53627=>"000000000",
  53628=>"111000111",
  53629=>"000111111",
  53630=>"000000110",
  53631=>"001111111",
  53632=>"100000111",
  53633=>"111111111",
  53634=>"100000000",
  53635=>"000000001",
  53636=>"000001111",
  53637=>"000111010",
  53638=>"010000100",
  53639=>"111011011",
  53640=>"010000000",
  53641=>"011011111",
  53642=>"000000000",
  53643=>"111111111",
  53644=>"111111111",
  53645=>"111100001",
  53646=>"111111111",
  53647=>"000111010",
  53648=>"000000111",
  53649=>"100100011",
  53650=>"111111111",
  53651=>"011111011",
  53652=>"111000000",
  53653=>"011011000",
  53654=>"111111010",
  53655=>"111011000",
  53656=>"111111000",
  53657=>"111011000",
  53658=>"011000000",
  53659=>"111000000",
  53660=>"110000000",
  53661=>"000000111",
  53662=>"110100000",
  53663=>"010111000",
  53664=>"000000111",
  53665=>"111110100",
  53666=>"111000000",
  53667=>"000000000",
  53668=>"000000100",
  53669=>"111111000",
  53670=>"000000000",
  53671=>"000000111",
  53672=>"111001101",
  53673=>"000000000",
  53674=>"111111111",
  53675=>"100100000",
  53676=>"111010000",
  53677=>"110000000",
  53678=>"111000101",
  53679=>"000011001",
  53680=>"000111111",
  53681=>"000000000",
  53682=>"111000110",
  53683=>"000000000",
  53684=>"000000011",
  53685=>"101000000",
  53686=>"101000000",
  53687=>"010010000",
  53688=>"000000000",
  53689=>"110111111",
  53690=>"011001000",
  53691=>"000011111",
  53692=>"001010010",
  53693=>"110111000",
  53694=>"100000000",
  53695=>"001111111",
  53696=>"000000000",
  53697=>"000000000",
  53698=>"111111111",
  53699=>"000000000",
  53700=>"111111000",
  53701=>"000000000",
  53702=>"000000000",
  53703=>"001001011",
  53704=>"110010000",
  53705=>"000111111",
  53706=>"111000000",
  53707=>"110110000",
  53708=>"111111100",
  53709=>"110000000",
  53710=>"000100111",
  53711=>"111010000",
  53712=>"000000111",
  53713=>"111001001",
  53714=>"110111111",
  53715=>"000000000",
  53716=>"001111111",
  53717=>"111111010",
  53718=>"001000000",
  53719=>"111101000",
  53720=>"111011000",
  53721=>"010000000",
  53722=>"000001111",
  53723=>"111111000",
  53724=>"101101001",
  53725=>"100000000",
  53726=>"111111011",
  53727=>"110001000",
  53728=>"001000000",
  53729=>"000000000",
  53730=>"000000001",
  53731=>"000000000",
  53732=>"000000011",
  53733=>"000010000",
  53734=>"110110111",
  53735=>"000000011",
  53736=>"000100000",
  53737=>"110001000",
  53738=>"011111111",
  53739=>"111111000",
  53740=>"001000001",
  53741=>"011011111",
  53742=>"000111100",
  53743=>"110111111",
  53744=>"100000110",
  53745=>"111011001",
  53746=>"000000000",
  53747=>"010010000",
  53748=>"111110111",
  53749=>"001000000",
  53750=>"001000010",
  53751=>"001000111",
  53752=>"000000000",
  53753=>"111011110",
  53754=>"010111010",
  53755=>"010000011",
  53756=>"001011011",
  53757=>"100100100",
  53758=>"100111111",
  53759=>"111111110",
  53760=>"000000000",
  53761=>"000000111",
  53762=>"001000000",
  53763=>"000011111",
  53764=>"000000000",
  53765=>"111010000",
  53766=>"001011111",
  53767=>"111111100",
  53768=>"111111111",
  53769=>"111111111",
  53770=>"111001101",
  53771=>"111110111",
  53772=>"000000000",
  53773=>"111010011",
  53774=>"111111111",
  53775=>"111111111",
  53776=>"010010010",
  53777=>"111111111",
  53778=>"000000100",
  53779=>"111111111",
  53780=>"111100111",
  53781=>"111111000",
  53782=>"000010111",
  53783=>"100000000",
  53784=>"001001101",
  53785=>"000000001",
  53786=>"000001001",
  53787=>"000100100",
  53788=>"000110110",
  53789=>"001000000",
  53790=>"001000001",
  53791=>"111111111",
  53792=>"111111111",
  53793=>"111111111",
  53794=>"101111111",
  53795=>"000000001",
  53796=>"000001000",
  53797=>"111110110",
  53798=>"111110111",
  53799=>"111101000",
  53800=>"110000011",
  53801=>"000000000",
  53802=>"000000000",
  53803=>"000000111",
  53804=>"000100100",
  53805=>"100000000",
  53806=>"000010000",
  53807=>"010011111",
  53808=>"111000100",
  53809=>"000000000",
  53810=>"100110110",
  53811=>"001111111",
  53812=>"000000000",
  53813=>"000000000",
  53814=>"011010111",
  53815=>"111111111",
  53816=>"000000001",
  53817=>"100100100",
  53818=>"000000001",
  53819=>"110110111",
  53820=>"111111111",
  53821=>"000000000",
  53822=>"000000000",
  53823=>"000000101",
  53824=>"100100100",
  53825=>"011000111",
  53826=>"001001011",
  53827=>"111000101",
  53828=>"111111011",
  53829=>"111111111",
  53830=>"101000110",
  53831=>"111111111",
  53832=>"001000000",
  53833=>"000000000",
  53834=>"111111111",
  53835=>"110101111",
  53836=>"000111111",
  53837=>"111011000",
  53838=>"011001011",
  53839=>"111111111",
  53840=>"000000100",
  53841=>"111111110",
  53842=>"011001001",
  53843=>"111111111",
  53844=>"000000000",
  53845=>"111101100",
  53846=>"000100111",
  53847=>"000000000",
  53848=>"000000000",
  53849=>"000000001",
  53850=>"100000000",
  53851=>"111111111",
  53852=>"000000000",
  53853=>"100000000",
  53854=>"000000000",
  53855=>"111111111",
  53856=>"000000000",
  53857=>"111111111",
  53858=>"000110111",
  53859=>"100111111",
  53860=>"100000000",
  53861=>"111111111",
  53862=>"111111000",
  53863=>"000000001",
  53864=>"000000000",
  53865=>"101100110",
  53866=>"000000000",
  53867=>"000000000",
  53868=>"000100100",
  53869=>"000001101",
  53870=>"111101001",
  53871=>"000000000",
  53872=>"000000010",
  53873=>"000010111",
  53874=>"110110100",
  53875=>"111111111",
  53876=>"111111111",
  53877=>"111000000",
  53878=>"000000000",
  53879=>"000010111",
  53880=>"111010000",
  53881=>"011000000",
  53882=>"000000000",
  53883=>"111001001",
  53884=>"111111100",
  53885=>"001000000",
  53886=>"000000000",
  53887=>"000000110",
  53888=>"111111111",
  53889=>"000100111",
  53890=>"110010000",
  53891=>"000000000",
  53892=>"000000000",
  53893=>"000000000",
  53894=>"111111000",
  53895=>"101000000",
  53896=>"111111001",
  53897=>"111000001",
  53898=>"100111111",
  53899=>"000011011",
  53900=>"110000110",
  53901=>"000010000",
  53902=>"000000010",
  53903=>"111111111",
  53904=>"111000000",
  53905=>"111111111",
  53906=>"000100101",
  53907=>"000001001",
  53908=>"000000010",
  53909=>"000010000",
  53910=>"111000000",
  53911=>"111111111",
  53912=>"000110110",
  53913=>"001111011",
  53914=>"111111111",
  53915=>"011111111",
  53916=>"001011111",
  53917=>"001000111",
  53918=>"101000000",
  53919=>"111111111",
  53920=>"000000000",
  53921=>"000000000",
  53922=>"111111110",
  53923=>"001001001",
  53924=>"000000100",
  53925=>"111111111",
  53926=>"111111111",
  53927=>"111001000",
  53928=>"001100000",
  53929=>"111111111",
  53930=>"111010000",
  53931=>"000010000",
  53932=>"111111111",
  53933=>"001101111",
  53934=>"000000111",
  53935=>"000000110",
  53936=>"111000011",
  53937=>"100000000",
  53938=>"111111110",
  53939=>"000000000",
  53940=>"111111111",
  53941=>"000110111",
  53942=>"111111111",
  53943=>"111111111",
  53944=>"001001000",
  53945=>"000000000",
  53946=>"000000000",
  53947=>"001101101",
  53948=>"111111111",
  53949=>"111011001",
  53950=>"000000000",
  53951=>"111111111",
  53952=>"000111111",
  53953=>"111011011",
  53954=>"110010111",
  53955=>"101111110",
  53956=>"111100000",
  53957=>"110000000",
  53958=>"111111111",
  53959=>"000001011",
  53960=>"000000000",
  53961=>"111111111",
  53962=>"000000000",
  53963=>"000100100",
  53964=>"110100110",
  53965=>"111111111",
  53966=>"111111111",
  53967=>"000000000",
  53968=>"111111111",
  53969=>"000000111",
  53970=>"000000000",
  53971=>"100000111",
  53972=>"110110000",
  53973=>"001001001",
  53974=>"000000000",
  53975=>"000110110",
  53976=>"100110111",
  53977=>"111101011",
  53978=>"101001111",
  53979=>"100100100",
  53980=>"111111111",
  53981=>"000000000",
  53982=>"100000100",
  53983=>"101101111",
  53984=>"000000000",
  53985=>"000000000",
  53986=>"000100000",
  53987=>"111111111",
  53988=>"000000001",
  53989=>"110110100",
  53990=>"111111111",
  53991=>"000000000",
  53992=>"111011111",
  53993=>"111111111",
  53994=>"000100100",
  53995=>"101100110",
  53996=>"101100000",
  53997=>"000000000",
  53998=>"000000000",
  53999=>"110000000",
  54000=>"011001001",
  54001=>"010010001",
  54002=>"000000000",
  54003=>"000100100",
  54004=>"000000000",
  54005=>"111111111",
  54006=>"100101111",
  54007=>"111111111",
  54008=>"110000000",
  54009=>"000000100",
  54010=>"111111101",
  54011=>"000000000",
  54012=>"011001000",
  54013=>"000000101",
  54014=>"101000000",
  54015=>"110000011",
  54016=>"110111111",
  54017=>"111110100",
  54018=>"000000000",
  54019=>"111011111",
  54020=>"111001001",
  54021=>"000000111",
  54022=>"111111111",
  54023=>"000000111",
  54024=>"111111111",
  54025=>"111111000",
  54026=>"111111111",
  54027=>"111111111",
  54028=>"111000000",
  54029=>"000000000",
  54030=>"111111011",
  54031=>"000000000",
  54032=>"000000111",
  54033=>"111000000",
  54034=>"001011011",
  54035=>"000111111",
  54036=>"111011011",
  54037=>"001001000",
  54038=>"111111111",
  54039=>"111111111",
  54040=>"110000000",
  54041=>"111111111",
  54042=>"000000000",
  54043=>"110100100",
  54044=>"111111111",
  54045=>"111111111",
  54046=>"000000000",
  54047=>"111111111",
  54048=>"111111111",
  54049=>"000000000",
  54050=>"011111110",
  54051=>"111111111",
  54052=>"000000111",
  54053=>"100100111",
  54054=>"110100000",
  54055=>"111000100",
  54056=>"000000000",
  54057=>"000011011",
  54058=>"111111111",
  54059=>"000000000",
  54060=>"000011111",
  54061=>"111101100",
  54062=>"111011111",
  54063=>"000000000",
  54064=>"000001111",
  54065=>"000000001",
  54066=>"111001100",
  54067=>"111111111",
  54068=>"000000000",
  54069=>"000000000",
  54070=>"111111111",
  54071=>"110010010",
  54072=>"011000000",
  54073=>"111111110",
  54074=>"101001001",
  54075=>"101111111",
  54076=>"110111001",
  54077=>"111111111",
  54078=>"000000000",
  54079=>"000000000",
  54080=>"100000000",
  54081=>"000111011",
  54082=>"000000000",
  54083=>"000111111",
  54084=>"111111111",
  54085=>"000000100",
  54086=>"100101001",
  54087=>"111111111",
  54088=>"000000000",
  54089=>"110110101",
  54090=>"000000000",
  54091=>"110110000",
  54092=>"000000000",
  54093=>"100111111",
  54094=>"000100111",
  54095=>"110110010",
  54096=>"000000000",
  54097=>"111011001",
  54098=>"111111111",
  54099=>"000000110",
  54100=>"111111111",
  54101=>"011011001",
  54102=>"000000000",
  54103=>"111010000",
  54104=>"000111111",
  54105=>"111111111",
  54106=>"010010111",
  54107=>"000000000",
  54108=>"111110111",
  54109=>"000000000",
  54110=>"111110111",
  54111=>"000000000",
  54112=>"100111010",
  54113=>"000000000",
  54114=>"000000100",
  54115=>"100000000",
  54116=>"111111111",
  54117=>"111000000",
  54118=>"000000000",
  54119=>"111011011",
  54120=>"111100100",
  54121=>"000000000",
  54122=>"000000000",
  54123=>"000000000",
  54124=>"111111111",
  54125=>"010000000",
  54126=>"000000001",
  54127=>"111101001",
  54128=>"111100100",
  54129=>"001001000",
  54130=>"000000111",
  54131=>"011011010",
  54132=>"001000000",
  54133=>"001101111",
  54134=>"111101100",
  54135=>"111101111",
  54136=>"101001001",
  54137=>"000000000",
  54138=>"000000000",
  54139=>"000000000",
  54140=>"000000000",
  54141=>"000011111",
  54142=>"111111111",
  54143=>"111111111",
  54144=>"010110000",
  54145=>"000000111",
  54146=>"111111011",
  54147=>"111000000",
  54148=>"000100111",
  54149=>"000011011",
  54150=>"001001101",
  54151=>"000001111",
  54152=>"011001000",
  54153=>"111110110",
  54154=>"111111110",
  54155=>"111111111",
  54156=>"111111100",
  54157=>"000000000",
  54158=>"111111111",
  54159=>"000001001",
  54160=>"110010000",
  54161=>"000000000",
  54162=>"011111000",
  54163=>"011101000",
  54164=>"000000000",
  54165=>"000000000",
  54166=>"000110100",
  54167=>"000000000",
  54168=>"000000000",
  54169=>"101000101",
  54170=>"111111111",
  54171=>"110111111",
  54172=>"111111111",
  54173=>"110110111",
  54174=>"000000000",
  54175=>"110111111",
  54176=>"111111111",
  54177=>"111011011",
  54178=>"110110111",
  54179=>"111001001",
  54180=>"000000101",
  54181=>"111111110",
  54182=>"000000000",
  54183=>"001111111",
  54184=>"000000111",
  54185=>"001100111",
  54186=>"111000000",
  54187=>"000000000",
  54188=>"000000000",
  54189=>"000000000",
  54190=>"111100000",
  54191=>"101000000",
  54192=>"110110000",
  54193=>"111111111",
  54194=>"110111111",
  54195=>"111000111",
  54196=>"111111111",
  54197=>"001000101",
  54198=>"110110111",
  54199=>"000000001",
  54200=>"111111111",
  54201=>"111111010",
  54202=>"110111111",
  54203=>"001011001",
  54204=>"111111111",
  54205=>"111111111",
  54206=>"000001000",
  54207=>"010110110",
  54208=>"110100110",
  54209=>"111111111",
  54210=>"000000000",
  54211=>"000000000",
  54212=>"110111111",
  54213=>"001000010",
  54214=>"110000000",
  54215=>"000000111",
  54216=>"000000000",
  54217=>"000000000",
  54218=>"101100000",
  54219=>"000000100",
  54220=>"111111111",
  54221=>"001000000",
  54222=>"000110110",
  54223=>"000000000",
  54224=>"000000000",
  54225=>"011000111",
  54226=>"111111111",
  54227=>"000000111",
  54228=>"011111011",
  54229=>"000000101",
  54230=>"000000100",
  54231=>"001011100",
  54232=>"111000000",
  54233=>"011000000",
  54234=>"111011001",
  54235=>"100101111",
  54236=>"011111111",
  54237=>"000000000",
  54238=>"111111111",
  54239=>"110000000",
  54240=>"111000000",
  54241=>"111111111",
  54242=>"000000000",
  54243=>"101101001",
  54244=>"000000000",
  54245=>"000110110",
  54246=>"111000100",
  54247=>"011001000",
  54248=>"000000111",
  54249=>"000000000",
  54250=>"100100100",
  54251=>"000000000",
  54252=>"010110111",
  54253=>"110110000",
  54254=>"111111111",
  54255=>"110000110",
  54256=>"000000000",
  54257=>"111010000",
  54258=>"110110111",
  54259=>"111110110",
  54260=>"000110111",
  54261=>"000000000",
  54262=>"100101111",
  54263=>"111111001",
  54264=>"000111111",
  54265=>"100000000",
  54266=>"001000001",
  54267=>"000000000",
  54268=>"000000000",
  54269=>"000000000",
  54270=>"000000000",
  54271=>"001000000",
  54272=>"101100000",
  54273=>"000111111",
  54274=>"000111111",
  54275=>"000000110",
  54276=>"001001000",
  54277=>"110000000",
  54278=>"111111110",
  54279=>"111111111",
  54280=>"110100100",
  54281=>"111101111",
  54282=>"101111111",
  54283=>"111101101",
  54284=>"111000000",
  54285=>"011000000",
  54286=>"111111111",
  54287=>"011111110",
  54288=>"111111110",
  54289=>"111111101",
  54290=>"010010110",
  54291=>"100110110",
  54292=>"000000010",
  54293=>"011111111",
  54294=>"111111111",
  54295=>"110111000",
  54296=>"000000000",
  54297=>"100100000",
  54298=>"001000111",
  54299=>"100000000",
  54300=>"111000001",
  54301=>"111111000",
  54302=>"111001000",
  54303=>"101001000",
  54304=>"001001000",
  54305=>"100000000",
  54306=>"111111111",
  54307=>"100001001",
  54308=>"000000000",
  54309=>"111100000",
  54310=>"000000000",
  54311=>"001001100",
  54312=>"000000000",
  54313=>"000000000",
  54314=>"000000000",
  54315=>"100111111",
  54316=>"111111111",
  54317=>"000000000",
  54318=>"111000000",
  54319=>"000000000",
  54320=>"111111001",
  54321=>"111011000",
  54322=>"100100000",
  54323=>"100100000",
  54324=>"111001101",
  54325=>"011011001",
  54326=>"111111111",
  54327=>"000000011",
  54328=>"001111111",
  54329=>"000000000",
  54330=>"000000000",
  54331=>"100000101",
  54332=>"000000000",
  54333=>"011001011",
  54334=>"110100111",
  54335=>"111111001",
  54336=>"100101111",
  54337=>"001001000",
  54338=>"101111000",
  54339=>"001001101",
  54340=>"011001000",
  54341=>"000000000",
  54342=>"111111100",
  54343=>"111111000",
  54344=>"000001000",
  54345=>"000000111",
  54346=>"000000111",
  54347=>"111001011",
  54348=>"111111111",
  54349=>"111001000",
  54350=>"100100000",
  54351=>"110100111",
  54352=>"100100000",
  54353=>"110111101",
  54354=>"001100100",
  54355=>"011001101",
  54356=>"011000000",
  54357=>"111001000",
  54358=>"110111111",
  54359=>"000000010",
  54360=>"000000000",
  54361=>"100000000",
  54362=>"000000101",
  54363=>"000001101",
  54364=>"001001001",
  54365=>"001111111",
  54366=>"110111000",
  54367=>"111111111",
  54368=>"000001001",
  54369=>"110111111",
  54370=>"000000010",
  54371=>"001000101",
  54372=>"001001000",
  54373=>"001000000",
  54374=>"010001000",
  54375=>"001111111",
  54376=>"111111111",
  54377=>"001001101",
  54378=>"010111111",
  54379=>"000000000",
  54380=>"010110111",
  54381=>"010110000",
  54382=>"000011111",
  54383=>"000001101",
  54384=>"000000001",
  54385=>"000000000",
  54386=>"111001000",
  54387=>"000000000",
  54388=>"111111111",
  54389=>"010000000",
  54390=>"000000000",
  54391=>"111111111",
  54392=>"000000000",
  54393=>"111111111",
  54394=>"010000000",
  54395=>"000000000",
  54396=>"001001000",
  54397=>"111111011",
  54398=>"000000000",
  54399=>"000111111",
  54400=>"011111111",
  54401=>"000000000",
  54402=>"000111111",
  54403=>"100110111",
  54404=>"000000111",
  54405=>"111111111",
  54406=>"111111000",
  54407=>"111000000",
  54408=>"111111111",
  54409=>"000110000",
  54410=>"111111101",
  54411=>"100111111",
  54412=>"111001000",
  54413=>"000110111",
  54414=>"110111101",
  54415=>"111111000",
  54416=>"111111111",
  54417=>"111111110",
  54418=>"000000000",
  54419=>"111111110",
  54420=>"111111111",
  54421=>"000011111",
  54422=>"000001111",
  54423=>"000000111",
  54424=>"011011001",
  54425=>"101111101",
  54426=>"000000110",
  54427=>"100100100",
  54428=>"110000000",
  54429=>"000111110",
  54430=>"111111111",
  54431=>"111100100",
  54432=>"011111111",
  54433=>"111001000",
  54434=>"000000000",
  54435=>"111111111",
  54436=>"011011011",
  54437=>"000010000",
  54438=>"011011010",
  54439=>"000000000",
  54440=>"000000111",
  54441=>"001001000",
  54442=>"101101100",
  54443=>"111111111",
  54444=>"110110110",
  54445=>"001000000",
  54446=>"001001111",
  54447=>"110110110",
  54448=>"000000110",
  54449=>"000000000",
  54450=>"111111110",
  54451=>"000000111",
  54452=>"010000000",
  54453=>"010000000",
  54454=>"011000000",
  54455=>"111000000",
  54456=>"111100101",
  54457=>"111111111",
  54458=>"000000000",
  54459=>"001000000",
  54460=>"010011011",
  54461=>"100111111",
  54462=>"000000000",
  54463=>"111111111",
  54464=>"000000000",
  54465=>"000000000",
  54466=>"110000000",
  54467=>"111001000",
  54468=>"000000000",
  54469=>"000000000",
  54470=>"000010010",
  54471=>"000001000",
  54472=>"000000111",
  54473=>"000000000",
  54474=>"000111111",
  54475=>"111111111",
  54476=>"100101101",
  54477=>"000000101",
  54478=>"111111000",
  54479=>"000000000",
  54480=>"000000000",
  54481=>"000011011",
  54482=>"111001000",
  54483=>"110110000",
  54484=>"000101000",
  54485=>"010111110",
  54486=>"000000000",
  54487=>"000000111",
  54488=>"111110000",
  54489=>"100101101",
  54490=>"000000000",
  54491=>"000101111",
  54492=>"111111111",
  54493=>"111111000",
  54494=>"000000000",
  54495=>"011011111",
  54496=>"111111111",
  54497=>"110000000",
  54498=>"111111111",
  54499=>"000000000",
  54500=>"111110100",
  54501=>"111110000",
  54502=>"100110110",
  54503=>"000000000",
  54504=>"111111110",
  54505=>"111111111",
  54506=>"000100101",
  54507=>"100111111",
  54508=>"000000000",
  54509=>"000000001",
  54510=>"000001111",
  54511=>"111111100",
  54512=>"010111111",
  54513=>"000111100",
  54514=>"001111111",
  54515=>"001101111",
  54516=>"111101101",
  54517=>"111111111",
  54518=>"000000011",
  54519=>"000000000",
  54520=>"000011111",
  54521=>"000000001",
  54522=>"000000000",
  54523=>"000001111",
  54524=>"000000111",
  54525=>"011111110",
  54526=>"000000111",
  54527=>"000000000",
  54528=>"111111111",
  54529=>"000010010",
  54530=>"100110111",
  54531=>"111000111",
  54532=>"101101001",
  54533=>"011111111",
  54534=>"111111111",
  54535=>"000010100",
  54536=>"010000000",
  54537=>"100100101",
  54538=>"111000000",
  54539=>"000000000",
  54540=>"111111111",
  54541=>"111111111",
  54542=>"000000000",
  54543=>"111111111",
  54544=>"100111111",
  54545=>"011000000",
  54546=>"000000000",
  54547=>"101111111",
  54548=>"100100111",
  54549=>"000000000",
  54550=>"011011111",
  54551=>"011100000",
  54552=>"111011011",
  54553=>"000000000",
  54554=>"000011010",
  54555=>"010010111",
  54556=>"111000000",
  54557=>"001000000",
  54558=>"111001001",
  54559=>"011111111",
  54560=>"000111000",
  54561=>"000100111",
  54562=>"000000111",
  54563=>"000000000",
  54564=>"000110000",
  54565=>"110111111",
  54566=>"111100000",
  54567=>"000000111",
  54568=>"000110100",
  54569=>"000000011",
  54570=>"000000000",
  54571=>"000010110",
  54572=>"000000100",
  54573=>"111111110",
  54574=>"000000000",
  54575=>"000001110",
  54576=>"110111111",
  54577=>"000000000",
  54578=>"101111111",
  54579=>"110000000",
  54580=>"000000000",
  54581=>"111111100",
  54582=>"000111111",
  54583=>"011001001",
  54584=>"000000111",
  54585=>"111100000",
  54586=>"010100111",
  54587=>"000000111",
  54588=>"001000000",
  54589=>"111111000",
  54590=>"111101000",
  54591=>"111111000",
  54592=>"101111111",
  54593=>"100000000",
  54594=>"010000000",
  54595=>"000000000",
  54596=>"011111101",
  54597=>"000001101",
  54598=>"011111010",
  54599=>"000000001",
  54600=>"000001011",
  54601=>"010000000",
  54602=>"111111111",
  54603=>"100100000",
  54604=>"000000101",
  54605=>"001001111",
  54606=>"110111111",
  54607=>"110110110",
  54608=>"000000100",
  54609=>"111111000",
  54610=>"001000101",
  54611=>"000000000",
  54612=>"000100111",
  54613=>"011011001",
  54614=>"111111111",
  54615=>"000000010",
  54616=>"111111101",
  54617=>"000000000",
  54618=>"000001000",
  54619=>"100000000",
  54620=>"000000000",
  54621=>"000000000",
  54622=>"111011010",
  54623=>"000110111",
  54624=>"001100100",
  54625=>"111111111",
  54626=>"100100100",
  54627=>"100000000",
  54628=>"110001111",
  54629=>"000000000",
  54630=>"000000000",
  54631=>"111111111",
  54632=>"000010100",
  54633=>"111101111",
  54634=>"111111000",
  54635=>"000001101",
  54636=>"011011011",
  54637=>"111111010",
  54638=>"101111111",
  54639=>"111111000",
  54640=>"000000000",
  54641=>"111111111",
  54642=>"011000000",
  54643=>"111100100",
  54644=>"111111100",
  54645=>"110111100",
  54646=>"001101101",
  54647=>"101101101",
  54648=>"111111111",
  54649=>"000101101",
  54650=>"111110110",
  54651=>"111011001",
  54652=>"000000000",
  54653=>"100111111",
  54654=>"011011001",
  54655=>"111000000",
  54656=>"010011010",
  54657=>"000000000",
  54658=>"000000000",
  54659=>"000000000",
  54660=>"000000100",
  54661=>"000000000",
  54662=>"000000001",
  54663=>"000111111",
  54664=>"000000000",
  54665=>"101100000",
  54666=>"100110000",
  54667=>"001101111",
  54668=>"000000000",
  54669=>"110010000",
  54670=>"000000001",
  54671=>"111111111",
  54672=>"000000000",
  54673=>"000101101",
  54674=>"000011110",
  54675=>"101001001",
  54676=>"000000000",
  54677=>"011000000",
  54678=>"100100000",
  54679=>"111111001",
  54680=>"000000000",
  54681=>"111011111",
  54682=>"111111111",
  54683=>"001011000",
  54684=>"011111111",
  54685=>"000000011",
  54686=>"111111111",
  54687=>"111011111",
  54688=>"000000000",
  54689=>"110001010",
  54690=>"000001101",
  54691=>"000000111",
  54692=>"011110000",
  54693=>"110100100",
  54694=>"100000000",
  54695=>"111101000",
  54696=>"111111101",
  54697=>"000000000",
  54698=>"001111111",
  54699=>"000000001",
  54700=>"110111010",
  54701=>"111110000",
  54702=>"011111111",
  54703=>"000000000",
  54704=>"000000000",
  54705=>"000000000",
  54706=>"111001001",
  54707=>"000000111",
  54708=>"111111111",
  54709=>"000111111",
  54710=>"100111111",
  54711=>"000000000",
  54712=>"000000000",
  54713=>"111111111",
  54714=>"100100111",
  54715=>"011011001",
  54716=>"101111111",
  54717=>"110110110",
  54718=>"111111110",
  54719=>"010011011",
  54720=>"111111111",
  54721=>"000000000",
  54722=>"000000000",
  54723=>"111010111",
  54724=>"110111000",
  54725=>"111100111",
  54726=>"000000001",
  54727=>"111111111",
  54728=>"011111011",
  54729=>"000000000",
  54730=>"000000000",
  54731=>"100000000",
  54732=>"000000000",
  54733=>"000000000",
  54734=>"000001111",
  54735=>"100111111",
  54736=>"111101101",
  54737=>"000100000",
  54738=>"000000000",
  54739=>"111111111",
  54740=>"100111011",
  54741=>"110111111",
  54742=>"000000001",
  54743=>"100000000",
  54744=>"100111111",
  54745=>"111111000",
  54746=>"110110000",
  54747=>"000001001",
  54748=>"111111111",
  54749=>"001111111",
  54750=>"111001000",
  54751=>"011110111",
  54752=>"101101111",
  54753=>"000000000",
  54754=>"000000000",
  54755=>"001000001",
  54756=>"111111111",
  54757=>"100111111",
  54758=>"100000111",
  54759=>"000000000",
  54760=>"001111110",
  54761=>"111101101",
  54762=>"000001001",
  54763=>"000111111",
  54764=>"111111111",
  54765=>"110111000",
  54766=>"000100111",
  54767=>"111111000",
  54768=>"111111111",
  54769=>"000000001",
  54770=>"000000000",
  54771=>"111111001",
  54772=>"111111000",
  54773=>"000000011",
  54774=>"101111111",
  54775=>"001001000",
  54776=>"111101000",
  54777=>"111001001",
  54778=>"101100110",
  54779=>"000000000",
  54780=>"000111100",
  54781=>"000000000",
  54782=>"111100100",
  54783=>"000000000",
  54784=>"111111100",
  54785=>"000001011",
  54786=>"101001000",
  54787=>"010000111",
  54788=>"001011000",
  54789=>"100101111",
  54790=>"111111111",
  54791=>"111111001",
  54792=>"000000001",
  54793=>"111111000",
  54794=>"111111000",
  54795=>"111111000",
  54796=>"001000000",
  54797=>"111011111",
  54798=>"111111111",
  54799=>"111111000",
  54800=>"001001001",
  54801=>"111111000",
  54802=>"000111111",
  54803=>"111111111",
  54804=>"000000000",
  54805=>"001000000",
  54806=>"011010000",
  54807=>"101001001",
  54808=>"111111001",
  54809=>"111100100",
  54810=>"001001111",
  54811=>"000110010",
  54812=>"001111111",
  54813=>"111111000",
  54814=>"111101111",
  54815=>"000000110",
  54816=>"101111111",
  54817=>"110110110",
  54818=>"110000000",
  54819=>"111111000",
  54820=>"000000111",
  54821=>"000001000",
  54822=>"101101101",
  54823=>"111000000",
  54824=>"101001001",
  54825=>"000000111",
  54826=>"000000000",
  54827=>"110111111",
  54828=>"111111000",
  54829=>"111111110",
  54830=>"000100000",
  54831=>"111010011",
  54832=>"110110111",
  54833=>"111111000",
  54834=>"001000001",
  54835=>"000101111",
  54836=>"000000111",
  54837=>"110110100",
  54838=>"001001011",
  54839=>"010011111",
  54840=>"000000000",
  54841=>"000000111",
  54842=>"000000001",
  54843=>"000000000",
  54844=>"111011000",
  54845=>"111111000",
  54846=>"111111111",
  54847=>"000000101",
  54848=>"000100111",
  54849=>"000000111",
  54850=>"000100000",
  54851=>"111001101",
  54852=>"110110000",
  54853=>"110011001",
  54854=>"000000111",
  54855=>"111111111",
  54856=>"111100000",
  54857=>"001000111",
  54858=>"111110000",
  54859=>"111000000",
  54860=>"001100100",
  54861=>"001011111",
  54862=>"010000000",
  54863=>"111110000",
  54864=>"000001011",
  54865=>"110000000",
  54866=>"111111110",
  54867=>"111111010",
  54868=>"000000100",
  54869=>"000000100",
  54870=>"000000000",
  54871=>"010000000",
  54872=>"000000000",
  54873=>"000011111",
  54874=>"110111111",
  54875=>"000000011",
  54876=>"110010000",
  54877=>"101111111",
  54878=>"100000000",
  54879=>"000001111",
  54880=>"111111111",
  54881=>"100001111",
  54882=>"111110100",
  54883=>"110110000",
  54884=>"000000000",
  54885=>"000001001",
  54886=>"111110000",
  54887=>"000011111",
  54888=>"000000111",
  54889=>"000000111",
  54890=>"000000111",
  54891=>"111111111",
  54892=>"110100000",
  54893=>"000000000",
  54894=>"001001111",
  54895=>"000001001",
  54896=>"000000100",
  54897=>"111010000",
  54898=>"011111000",
  54899=>"111111110",
  54900=>"100000000",
  54901=>"001000000",
  54902=>"000000000",
  54903=>"111111111",
  54904=>"110111100",
  54905=>"111111111",
  54906=>"001001001",
  54907=>"111101111",
  54908=>"000110000",
  54909=>"111111001",
  54910=>"001111101",
  54911=>"000000111",
  54912=>"111111000",
  54913=>"000000111",
  54914=>"001000111",
  54915=>"100100111",
  54916=>"111111111",
  54917=>"111111111",
  54918=>"110111010",
  54919=>"000000001",
  54920=>"001001001",
  54921=>"111111010",
  54922=>"110100000",
  54923=>"111011101",
  54924=>"011000000",
  54925=>"101000111",
  54926=>"111110000",
  54927=>"110000000",
  54928=>"000000111",
  54929=>"100100100",
  54930=>"000000000",
  54931=>"111111101",
  54932=>"100000111",
  54933=>"111111001",
  54934=>"000000001",
  54935=>"101001001",
  54936=>"000000000",
  54937=>"000000000",
  54938=>"111111111",
  54939=>"100000101",
  54940=>"000100000",
  54941=>"110111100",
  54942=>"001001111",
  54943=>"000110111",
  54944=>"000000100",
  54945=>"001000001",
  54946=>"111111011",
  54947=>"110110000",
  54948=>"001001101",
  54949=>"111111000",
  54950=>"111111000",
  54951=>"111111000",
  54952=>"000000000",
  54953=>"010010000",
  54954=>"011111000",
  54955=>"000000000",
  54956=>"110110000",
  54957=>"100100111",
  54958=>"111111111",
  54959=>"000001111",
  54960=>"110111111",
  54961=>"000001000",
  54962=>"110110010",
  54963=>"010000001",
  54964=>"000101111",
  54965=>"000000011",
  54966=>"010011000",
  54967=>"000000000",
  54968=>"110111111",
  54969=>"101001001",
  54970=>"000001101",
  54971=>"111010000",
  54972=>"000000111",
  54973=>"000001011",
  54974=>"000111000",
  54975=>"100000000",
  54976=>"001000000",
  54977=>"111011001",
  54978=>"101111111",
  54979=>"111111100",
  54980=>"000000011",
  54981=>"000000000",
  54982=>"111000000",
  54983=>"000110100",
  54984=>"111101101",
  54985=>"111111111",
  54986=>"000000000",
  54987=>"111011011",
  54988=>"100000100",
  54989=>"111111111",
  54990=>"001000000",
  54991=>"000001111",
  54992=>"101101110",
  54993=>"000000101",
  54994=>"000011000",
  54995=>"000000101",
  54996=>"111111110",
  54997=>"111001101",
  54998=>"111011001",
  54999=>"000000111",
  55000=>"111111000",
  55001=>"111111011",
  55002=>"000000000",
  55003=>"010111111",
  55004=>"111111111",
  55005=>"000000001",
  55006=>"111011001",
  55007=>"001011011",
  55008=>"111111000",
  55009=>"000000000",
  55010=>"000001110",
  55011=>"111000000",
  55012=>"111000000",
  55013=>"001001100",
  55014=>"001000000",
  55015=>"111111010",
  55016=>"111111000",
  55017=>"001001101",
  55018=>"111100100",
  55019=>"101000101",
  55020=>"010010000",
  55021=>"111010010",
  55022=>"000001001",
  55023=>"001111000",
  55024=>"111000000",
  55025=>"010111001",
  55026=>"001000000",
  55027=>"000100101",
  55028=>"010110000",
  55029=>"000000111",
  55030=>"110000101",
  55031=>"000000000",
  55032=>"111110000",
  55033=>"001000000",
  55034=>"010111000",
  55035=>"110111111",
  55036=>"001000111",
  55037=>"001000001",
  55038=>"111111111",
  55039=>"011111111",
  55040=>"000000000",
  55041=>"001000001",
  55042=>"110110111",
  55043=>"011011011",
  55044=>"101000000",
  55045=>"010110000",
  55046=>"000001000",
  55047=>"001001000",
  55048=>"111100000",
  55049=>"000101111",
  55050=>"011010000",
  55051=>"000000000",
  55052=>"000000110",
  55053=>"010111111",
  55054=>"001000000",
  55055=>"110010000",
  55056=>"111001111",
  55057=>"000000100",
  55058=>"000000000",
  55059=>"000000000",
  55060=>"111111000",
  55061=>"101111010",
  55062=>"101001011",
  55063=>"110110111",
  55064=>"111000000",
  55065=>"111111101",
  55066=>"000000111",
  55067=>"000001001",
  55068=>"000000000",
  55069=>"111110000",
  55070=>"011001000",
  55071=>"000000001",
  55072=>"110111000",
  55073=>"100111111",
  55074=>"111000111",
  55075=>"111111111",
  55076=>"000000000",
  55077=>"111000000",
  55078=>"100000000",
  55079=>"001000000",
  55080=>"000000111",
  55081=>"000000000",
  55082=>"110011001",
  55083=>"011111000",
  55084=>"001001001",
  55085=>"011001000",
  55086=>"111111000",
  55087=>"010010111",
  55088=>"001000111",
  55089=>"111111010",
  55090=>"010110110",
  55091=>"000110111",
  55092=>"011111111",
  55093=>"010011110",
  55094=>"000000001",
  55095=>"101000000",
  55096=>"111111111",
  55097=>"111111011",
  55098=>"111001001",
  55099=>"111111011",
  55100=>"000000000",
  55101=>"000000100",
  55102=>"000110100",
  55103=>"111111000",
  55104=>"000000111",
  55105=>"000100100",
  55106=>"000100000",
  55107=>"000000000",
  55108=>"110000111",
  55109=>"001001001",
  55110=>"011111010",
  55111=>"111110100",
  55112=>"000000000",
  55113=>"101001000",
  55114=>"111111101",
  55115=>"000000111",
  55116=>"000000000",
  55117=>"111111111",
  55118=>"000000001",
  55119=>"110111000",
  55120=>"001111101",
  55121=>"111111111",
  55122=>"001001110",
  55123=>"000000111",
  55124=>"000100111",
  55125=>"001001111",
  55126=>"111100111",
  55127=>"101001001",
  55128=>"101000000",
  55129=>"000110000",
  55130=>"110111111",
  55131=>"000000100",
  55132=>"000000100",
  55133=>"000010000",
  55134=>"100110000",
  55135=>"000000010",
  55136=>"111111000",
  55137=>"101111011",
  55138=>"001001111",
  55139=>"000000001",
  55140=>"111110011",
  55141=>"000000000",
  55142=>"010000010",
  55143=>"000000000",
  55144=>"001001111",
  55145=>"000000000",
  55146=>"000100100",
  55147=>"010011011",
  55148=>"000100111",
  55149=>"001110111",
  55150=>"111111000",
  55151=>"000000000",
  55152=>"000000000",
  55153=>"000111111",
  55154=>"000000000",
  55155=>"111111111",
  55156=>"101100000",
  55157=>"001000000",
  55158=>"101100111",
  55159=>"000000000",
  55160=>"011111000",
  55161=>"000000000",
  55162=>"111000000",
  55163=>"000100000",
  55164=>"111011000",
  55165=>"110110111",
  55166=>"001001001",
  55167=>"000001011",
  55168=>"011000000",
  55169=>"111101111",
  55170=>"010110000",
  55171=>"000000000",
  55172=>"000111010",
  55173=>"001001000",
  55174=>"000000000",
  55175=>"011010111",
  55176=>"111110000",
  55177=>"000110100",
  55178=>"001101101",
  55179=>"001011111",
  55180=>"100110000",
  55181=>"100110100",
  55182=>"111111111",
  55183=>"111111000",
  55184=>"000000110",
  55185=>"111111111",
  55186=>"001001111",
  55187=>"000000000",
  55188=>"000000000",
  55189=>"000011111",
  55190=>"101111011",
  55191=>"111001001",
  55192=>"000110111",
  55193=>"111101110",
  55194=>"000000000",
  55195=>"111111111",
  55196=>"010111111",
  55197=>"111001111",
  55198=>"000001101",
  55199=>"111111010",
  55200=>"000001101",
  55201=>"010011010",
  55202=>"111001111",
  55203=>"110111111",
  55204=>"000100000",
  55205=>"000110111",
  55206=>"111001000",
  55207=>"000001011",
  55208=>"101111111",
  55209=>"000010000",
  55210=>"111011000",
  55211=>"111110000",
  55212=>"000000000",
  55213=>"000000000",
  55214=>"000111111",
  55215=>"011001000",
  55216=>"001111111",
  55217=>"010010000",
  55218=>"110111000",
  55219=>"000000001",
  55220=>"011111000",
  55221=>"001001111",
  55222=>"111111000",
  55223=>"000000000",
  55224=>"000000111",
  55225=>"111011111",
  55226=>"111111000",
  55227=>"111111111",
  55228=>"000000100",
  55229=>"000000000",
  55230=>"001001111",
  55231=>"001100111",
  55232=>"111111101",
  55233=>"000000100",
  55234=>"100110000",
  55235=>"001000000",
  55236=>"000000000",
  55237=>"110110100",
  55238=>"001000100",
  55239=>"111011010",
  55240=>"000000111",
  55241=>"011100111",
  55242=>"000000000",
  55243=>"000000000",
  55244=>"000000000",
  55245=>"111111110",
  55246=>"000001111",
  55247=>"111111111",
  55248=>"000000111",
  55249=>"000111110",
  55250=>"001001111",
  55251=>"111001000",
  55252=>"111011000",
  55253=>"011000000",
  55254=>"000000011",
  55255=>"100100111",
  55256=>"000000110",
  55257=>"111111011",
  55258=>"011010000",
  55259=>"011000000",
  55260=>"000000000",
  55261=>"110110000",
  55262=>"100000001",
  55263=>"011111111",
  55264=>"001101111",
  55265=>"111000000",
  55266=>"000000000",
  55267=>"111110000",
  55268=>"111000000",
  55269=>"111111100",
  55270=>"000000000",
  55271=>"111111000",
  55272=>"111110110",
  55273=>"001001101",
  55274=>"000000000",
  55275=>"111110101",
  55276=>"011001000",
  55277=>"011000100",
  55278=>"111111010",
  55279=>"111011001",
  55280=>"000111101",
  55281=>"011111011",
  55282=>"110110000",
  55283=>"000000010",
  55284=>"001010111",
  55285=>"000000000",
  55286=>"000000110",
  55287=>"000111111",
  55288=>"101111110",
  55289=>"000000111",
  55290=>"111111001",
  55291=>"001001111",
  55292=>"110000111",
  55293=>"100000000",
  55294=>"000000110",
  55295=>"000100111",
  55296=>"110010010",
  55297=>"100110111",
  55298=>"001000000",
  55299=>"100100000",
  55300=>"101100110",
  55301=>"100010000",
  55302=>"110111110",
  55303=>"000000000",
  55304=>"111111010",
  55305=>"101111111",
  55306=>"111100000",
  55307=>"111111110",
  55308=>"100100100",
  55309=>"111110110",
  55310=>"001100000",
  55311=>"000000111",
  55312=>"001100111",
  55313=>"011110111",
  55314=>"001000100",
  55315=>"001001000",
  55316=>"110011111",
  55317=>"000000000",
  55318=>"111111111",
  55319=>"010111111",
  55320=>"101111111",
  55321=>"100001000",
  55322=>"100100101",
  55323=>"110010110",
  55324=>"000000000",
  55325=>"111111111",
  55326=>"100100100",
  55327=>"000000000",
  55328=>"001100110",
  55329=>"100010011",
  55330=>"000001000",
  55331=>"110000101",
  55332=>"001000101",
  55333=>"100111110",
  55334=>"010000000",
  55335=>"110110010",
  55336=>"000000000",
  55337=>"100110110",
  55338=>"111111111",
  55339=>"111001001",
  55340=>"000000000",
  55341=>"111001011",
  55342=>"000000000",
  55343=>"110110000",
  55344=>"001001111",
  55345=>"001000100",
  55346=>"111111011",
  55347=>"011101100",
  55348=>"011111111",
  55349=>"110010000",
  55350=>"001000000",
  55351=>"100000001",
  55352=>"111111000",
  55353=>"000000111",
  55354=>"010110010",
  55355=>"000101111",
  55356=>"001001111",
  55357=>"000000101",
  55358=>"111111111",
  55359=>"000000010",
  55360=>"000111111",
  55361=>"100101101",
  55362=>"110110111",
  55363=>"000001111",
  55364=>"000000000",
  55365=>"111111111",
  55366=>"110010010",
  55367=>"000000000",
  55368=>"000011010",
  55369=>"000111111",
  55370=>"110110000",
  55371=>"100111011",
  55372=>"000100111",
  55373=>"111100000",
  55374=>"000000101",
  55375=>"101111111",
  55376=>"011001001",
  55377=>"001001001",
  55378=>"111111111",
  55379=>"011000000",
  55380=>"000000100",
  55381=>"001000100",
  55382=>"110110110",
  55383=>"111111001",
  55384=>"011000000",
  55385=>"000000111",
  55386=>"111001001",
  55387=>"111011001",
  55388=>"111100000",
  55389=>"000000101",
  55390=>"000000110",
  55391=>"111011000",
  55392=>"000111111",
  55393=>"101111101",
  55394=>"000000000",
  55395=>"000000111",
  55396=>"110110000",
  55397=>"000000110",
  55398=>"100110110",
  55399=>"111000000",
  55400=>"000100111",
  55401=>"111111001",
  55402=>"000000010",
  55403=>"000110010",
  55404=>"110111010",
  55405=>"101101101",
  55406=>"101001001",
  55407=>"000111111",
  55408=>"100111111",
  55409=>"111000000",
  55410=>"101111000",
  55411=>"111111100",
  55412=>"110111010",
  55413=>"100110110",
  55414=>"111111000",
  55415=>"110110100",
  55416=>"001000111",
  55417=>"000000100",
  55418=>"111100101",
  55419=>"001000000",
  55420=>"000000000",
  55421=>"110100100",
  55422=>"110111110",
  55423=>"100010111",
  55424=>"010110010",
  55425=>"000000000",
  55426=>"110000000",
  55427=>"011000110",
  55428=>"000111111",
  55429=>"000000000",
  55430=>"100100010",
  55431=>"110010010",
  55432=>"010010000",
  55433=>"000000000",
  55434=>"111111111",
  55435=>"110110000",
  55436=>"110010001",
  55437=>"111111111",
  55438=>"000100111",
  55439=>"000000000",
  55440=>"001001101",
  55441=>"101101111",
  55442=>"000010110",
  55443=>"110000110",
  55444=>"010000000",
  55445=>"111110110",
  55446=>"000110111",
  55447=>"001001001",
  55448=>"001000001",
  55449=>"001001011",
  55450=>"101101110",
  55451=>"000000100",
  55452=>"010111110",
  55453=>"000000001",
  55454=>"010111000",
  55455=>"011111111",
  55456=>"010000000",
  55457=>"111111111",
  55458=>"111110000",
  55459=>"001001100",
  55460=>"010010110",
  55461=>"111010000",
  55462=>"001001111",
  55463=>"111111100",
  55464=>"110110010",
  55465=>"111001001",
  55466=>"000000000",
  55467=>"100111111",
  55468=>"111111111",
  55469=>"000000101",
  55470=>"101000000",
  55471=>"010011000",
  55472=>"000000000",
  55473=>"001100001",
  55474=>"111111111",
  55475=>"111111111",
  55476=>"111111111",
  55477=>"000000000",
  55478=>"111111000",
  55479=>"000000010",
  55480=>"111111011",
  55481=>"111111111",
  55482=>"011000100",
  55483=>"110110110",
  55484=>"000000000",
  55485=>"110110000",
  55486=>"111111010",
  55487=>"000000000",
  55488=>"111111010",
  55489=>"110000000",
  55490=>"011000111",
  55491=>"000000000",
  55492=>"111001111",
  55493=>"000000000",
  55494=>"001101001",
  55495=>"110000000",
  55496=>"111111111",
  55497=>"101001111",
  55498=>"000000101",
  55499=>"111111010",
  55500=>"001000000",
  55501=>"110111010",
  55502=>"000110011",
  55503=>"011011111",
  55504=>"111000000",
  55505=>"000000000",
  55506=>"000000000",
  55507=>"110000000",
  55508=>"000000110",
  55509=>"000001011",
  55510=>"001000001",
  55511=>"010000000",
  55512=>"111000000",
  55513=>"110110110",
  55514=>"111111110",
  55515=>"011110110",
  55516=>"111001001",
  55517=>"000000000",
  55518=>"000000000",
  55519=>"010000000",
  55520=>"000000000",
  55521=>"001111010",
  55522=>"100111111",
  55523=>"000000010",
  55524=>"000000000",
  55525=>"111110010",
  55526=>"111110111",
  55527=>"000000000",
  55528=>"000000100",
  55529=>"011011001",
  55530=>"101000001",
  55531=>"100001111",
  55532=>"111001111",
  55533=>"111001000",
  55534=>"100110111",
  55535=>"010011111",
  55536=>"000001000",
  55537=>"011111111",
  55538=>"000001010",
  55539=>"000000000",
  55540=>"111111010",
  55541=>"110100000",
  55542=>"111111110",
  55543=>"001001001",
  55544=>"110000111",
  55545=>"001001111",
  55546=>"110110111",
  55547=>"101111111",
  55548=>"111111100",
  55549=>"000100110",
  55550=>"111111010",
  55551=>"111111011",
  55552=>"110110100",
  55553=>"110100111",
  55554=>"101101111",
  55555=>"111111111",
  55556=>"000000001",
  55557=>"000000000",
  55558=>"011111000",
  55559=>"110010000",
  55560=>"001000000",
  55561=>"111111111",
  55562=>"110000000",
  55563=>"000001101",
  55564=>"111111111",
  55565=>"011010111",
  55566=>"110110010",
  55567=>"001001011",
  55568=>"000000000",
  55569=>"111111111",
  55570=>"111101111",
  55571=>"101111111",
  55572=>"000010110",
  55573=>"001111111",
  55574=>"111111001",
  55575=>"111010011",
  55576=>"001011011",
  55577=>"111111100",
  55578=>"111011111",
  55579=>"111001000",
  55580=>"110110110",
  55581=>"110110000",
  55582=>"000000000",
  55583=>"010110110",
  55584=>"111100100",
  55585=>"111111111",
  55586=>"000000010",
  55587=>"011011111",
  55588=>"110110110",
  55589=>"000000110",
  55590=>"101011001",
  55591=>"001001011",
  55592=>"111111111",
  55593=>"001001101",
  55594=>"111111110",
  55595=>"000000000",
  55596=>"111111111",
  55597=>"011010000",
  55598=>"001111111",
  55599=>"111111111",
  55600=>"001001111",
  55601=>"111001000",
  55602=>"111001111",
  55603=>"111111111",
  55604=>"111111001",
  55605=>"000000000",
  55606=>"011011011",
  55607=>"110110110",
  55608=>"000000000",
  55609=>"001000101",
  55610=>"111111111",
  55611=>"000000000",
  55612=>"100101100",
  55613=>"110100000",
  55614=>"110110110",
  55615=>"000001011",
  55616=>"000000000",
  55617=>"111001111",
  55618=>"000000111",
  55619=>"100100000",
  55620=>"001001111",
  55621=>"111001000",
  55622=>"000000000",
  55623=>"110000000",
  55624=>"111111111",
  55625=>"111010000",
  55626=>"111111101",
  55627=>"010011011",
  55628=>"010000000",
  55629=>"000011000",
  55630=>"000000000",
  55631=>"110010010",
  55632=>"011011011",
  55633=>"000000000",
  55634=>"010010110",
  55635=>"111111111",
  55636=>"101111111",
  55637=>"011000000",
  55638=>"101101111",
  55639=>"111111000",
  55640=>"000001111",
  55641=>"111101111",
  55642=>"000000110",
  55643=>"001011111",
  55644=>"000000000",
  55645=>"111000001",
  55646=>"011000001",
  55647=>"111110100",
  55648=>"011001000",
  55649=>"101000000",
  55650=>"000000000",
  55651=>"001001111",
  55652=>"110110100",
  55653=>"000000111",
  55654=>"000010110",
  55655=>"110110010",
  55656=>"101101100",
  55657=>"000000000",
  55658=>"110000000",
  55659=>"000110000",
  55660=>"111111000",
  55661=>"011011000",
  55662=>"110110111",
  55663=>"000000111",
  55664=>"101001001",
  55665=>"000000011",
  55666=>"000000000",
  55667=>"111111000",
  55668=>"000000000",
  55669=>"111111111",
  55670=>"000101111",
  55671=>"100111111",
  55672=>"111101111",
  55673=>"000000000",
  55674=>"111111111",
  55675=>"010110000",
  55676=>"100000000",
  55677=>"000001001",
  55678=>"011011000",
  55679=>"110111010",
  55680=>"110110100",
  55681=>"111011000",
  55682=>"010110110",
  55683=>"000000000",
  55684=>"001000001",
  55685=>"000000000",
  55686=>"111111111",
  55687=>"110111101",
  55688=>"101001111",
  55689=>"000010000",
  55690=>"000100101",
  55691=>"111111000",
  55692=>"111010000",
  55693=>"001000000",
  55694=>"110110010",
  55695=>"000000000",
  55696=>"001001111",
  55697=>"010000100",
  55698=>"111111000",
  55699=>"110011011",
  55700=>"011010111",
  55701=>"000110000",
  55702=>"000001101",
  55703=>"000000110",
  55704=>"010001000",
  55705=>"110100000",
  55706=>"101101001",
  55707=>"000000000",
  55708=>"001001111",
  55709=>"000000111",
  55710=>"001001111",
  55711=>"110110110",
  55712=>"000000110",
  55713=>"010000100",
  55714=>"111110110",
  55715=>"000000011",
  55716=>"000000001",
  55717=>"111111000",
  55718=>"000000101",
  55719=>"111000000",
  55720=>"100110000",
  55721=>"000000011",
  55722=>"110110010",
  55723=>"011001000",
  55724=>"000000111",
  55725=>"111111111",
  55726=>"011111111",
  55727=>"001000000",
  55728=>"000000001",
  55729=>"110111000",
  55730=>"111101001",
  55731=>"110110010",
  55732=>"000000001",
  55733=>"110010000",
  55734=>"100111111",
  55735=>"001001010",
  55736=>"000000111",
  55737=>"100111111",
  55738=>"110000000",
  55739=>"010110110",
  55740=>"001001111",
  55741=>"110010000",
  55742=>"111111000",
  55743=>"000000100",
  55744=>"000000101",
  55745=>"101000001",
  55746=>"001111111",
  55747=>"010111111",
  55748=>"001001001",
  55749=>"000001011",
  55750=>"000000001",
  55751=>"111101000",
  55752=>"000000000",
  55753=>"010100111",
  55754=>"111001111",
  55755=>"011011111",
  55756=>"001101110",
  55757=>"000000000",
  55758=>"110000000",
  55759=>"111111111",
  55760=>"011001000",
  55761=>"011111111",
  55762=>"000000110",
  55763=>"000000000",
  55764=>"000000000",
  55765=>"110010010",
  55766=>"111100111",
  55767=>"011111010",
  55768=>"000000100",
  55769=>"000000000",
  55770=>"000000110",
  55771=>"110010000",
  55772=>"011000101",
  55773=>"010011001",
  55774=>"111000111",
  55775=>"111011111",
  55776=>"111111001",
  55777=>"110010000",
  55778=>"010000011",
  55779=>"010110000",
  55780=>"000000000",
  55781=>"001100111",
  55782=>"111110100",
  55783=>"001000111",
  55784=>"110110110",
  55785=>"000000000",
  55786=>"100111001",
  55787=>"011011111",
  55788=>"000010110",
  55789=>"001001110",
  55790=>"001001001",
  55791=>"111000000",
  55792=>"001001111",
  55793=>"011111111",
  55794=>"101111100",
  55795=>"011011101",
  55796=>"110110000",
  55797=>"011111111",
  55798=>"110000001",
  55799=>"000001000",
  55800=>"000000001",
  55801=>"000100000",
  55802=>"001001001",
  55803=>"000000000",
  55804=>"000000000",
  55805=>"100000010",
  55806=>"000000000",
  55807=>"000000000",
  55808=>"111010110",
  55809=>"000000000",
  55810=>"000000011",
  55811=>"101101101",
  55812=>"101101101",
  55813=>"010000000",
  55814=>"000001001",
  55815=>"000000000",
  55816=>"111100101",
  55817=>"111011110",
  55818=>"100000000",
  55819=>"011001111",
  55820=>"000001001",
  55821=>"001101101",
  55822=>"111100110",
  55823=>"001101101",
  55824=>"101001001",
  55825=>"010000101",
  55826=>"011011001",
  55827=>"000000000",
  55828=>"000000000",
  55829=>"001000000",
  55830=>"000010111",
  55831=>"100000000",
  55832=>"000001111",
  55833=>"100100100",
  55834=>"101101111",
  55835=>"011011010",
  55836=>"001101101",
  55837=>"101000100",
  55838=>"100100100",
  55839=>"111000111",
  55840=>"000000011",
  55841=>"000000011",
  55842=>"110010110",
  55843=>"111111111",
  55844=>"101101111",
  55845=>"111110100",
  55846=>"000000000",
  55847=>"000000011",
  55848=>"000110000",
  55849=>"000000000",
  55850=>"111000111",
  55851=>"101100000",
  55852=>"100100101",
  55853=>"111101001",
  55854=>"101100001",
  55855=>"000111111",
  55856=>"111111111",
  55857=>"000001001",
  55858=>"100000000",
  55859=>"000100000",
  55860=>"101101101",
  55861=>"110110100",
  55862=>"111001011",
  55863=>"100100000",
  55864=>"111111111",
  55865=>"111111111",
  55866=>"001001101",
  55867=>"000000110",
  55868=>"001101000",
  55869=>"111111111",
  55870=>"110000000",
  55871=>"111101000",
  55872=>"001001110",
  55873=>"100100100",
  55874=>"000000000",
  55875=>"101111111",
  55876=>"000010011",
  55877=>"001001011",
  55878=>"101001000",
  55879=>"011000011",
  55880=>"101101100",
  55881=>"011000000",
  55882=>"100111111",
  55883=>"010010110",
  55884=>"111110110",
  55885=>"111110100",
  55886=>"000000101",
  55887=>"101101111",
  55888=>"000000011",
  55889=>"001101101",
  55890=>"111000000",
  55891=>"000000000",
  55892=>"100101001",
  55893=>"011010111",
  55894=>"110111111",
  55895=>"100100100",
  55896=>"100110111",
  55897=>"111101111",
  55898=>"100101001",
  55899=>"000000000",
  55900=>"100001101",
  55901=>"010000000",
  55902=>"111110110",
  55903=>"001001001",
  55904=>"111111111",
  55905=>"100111111",
  55906=>"111111111",
  55907=>"000100111",
  55908=>"111000000",
  55909=>"000000100",
  55910=>"101111000",
  55911=>"010010000",
  55912=>"111101101",
  55913=>"000000000",
  55914=>"000000010",
  55915=>"010011011",
  55916=>"001000000",
  55917=>"000000000",
  55918=>"100101101",
  55919=>"001001001",
  55920=>"000000001",
  55921=>"000101111",
  55922=>"000000001",
  55923=>"111110010",
  55924=>"011110100",
  55925=>"010010110",
  55926=>"100000000",
  55927=>"110010000",
  55928=>"000101101",
  55929=>"111111111",
  55930=>"110110111",
  55931=>"000000000",
  55932=>"100100100",
  55933=>"101111111",
  55934=>"111111100",
  55935=>"111111001",
  55936=>"000000000",
  55937=>"111111111",
  55938=>"011010110",
  55939=>"000011001",
  55940=>"100101100",
  55941=>"111001000",
  55942=>"000000000",
  55943=>"111110000",
  55944=>"000000000",
  55945=>"111101111",
  55946=>"001101111",
  55947=>"111111111",
  55948=>"110110111",
  55949=>"101111111",
  55950=>"001010000",
  55951=>"001111001",
  55952=>"101101101",
  55953=>"101100000",
  55954=>"010011011",
  55955=>"111001000",
  55956=>"111110100",
  55957=>"100000000",
  55958=>"101101100",
  55959=>"111111101",
  55960=>"101100000",
  55961=>"000001000",
  55962=>"101101100",
  55963=>"000000000",
  55964=>"101111111",
  55965=>"111111110",
  55966=>"101101001",
  55967=>"110110110",
  55968=>"111101000",
  55969=>"001000100",
  55970=>"001001001",
  55971=>"101000000",
  55972=>"010010000",
  55973=>"011000111",
  55974=>"000011011",
  55975=>"000001001",
  55976=>"111111111",
  55977=>"000001111",
  55978=>"111111011",
  55979=>"100101101",
  55980=>"010000000",
  55981=>"100100100",
  55982=>"111111111",
  55983=>"000000000",
  55984=>"010010000",
  55985=>"101101101",
  55986=>"000000000",
  55987=>"111111100",
  55988=>"111111111",
  55989=>"111111111",
  55990=>"000001000",
  55991=>"111111011",
  55992=>"101111111",
  55993=>"100101111",
  55994=>"100100001",
  55995=>"000010010",
  55996=>"011111111",
  55997=>"001001000",
  55998=>"010010000",
  55999=>"101100101",
  56000=>"000000100",
  56001=>"110110010",
  56002=>"000110110",
  56003=>"000000111",
  56004=>"111111111",
  56005=>"000000010",
  56006=>"010010010",
  56007=>"110010011",
  56008=>"010000001",
  56009=>"101100100",
  56010=>"010010010",
  56011=>"111111001",
  56012=>"111111111",
  56013=>"101101000",
  56014=>"101111111",
  56015=>"111001011",
  56016=>"000100111",
  56017=>"101001000",
  56018=>"011111111",
  56019=>"101100000",
  56020=>"101101100",
  56021=>"101100000",
  56022=>"000000000",
  56023=>"101100101",
  56024=>"001000000",
  56025=>"101100100",
  56026=>"010010110",
  56027=>"001001101",
  56028=>"000000110",
  56029=>"101101101",
  56030=>"000110000",
  56031=>"110110110",
  56032=>"000100101",
  56033=>"000000000",
  56034=>"000011101",
  56035=>"011011000",
  56036=>"010011111",
  56037=>"000000001",
  56038=>"010010010",
  56039=>"111111111",
  56040=>"101101111",
  56041=>"011011011",
  56042=>"111111111",
  56043=>"010010011",
  56044=>"011001111",
  56045=>"000000000",
  56046=>"000000111",
  56047=>"111111111",
  56048=>"111011111",
  56049=>"000000000",
  56050=>"111111111",
  56051=>"000010111",
  56052=>"111001011",
  56053=>"110110100",
  56054=>"101101111",
  56055=>"101101111",
  56056=>"111111111",
  56057=>"000000000",
  56058=>"100111111",
  56059=>"111111101",
  56060=>"000000100",
  56061=>"000000001",
  56062=>"110110011",
  56063=>"010010010",
  56064=>"000000101",
  56065=>"101001001",
  56066=>"000000001",
  56067=>"100001000",
  56068=>"000000000",
  56069=>"001000000",
  56070=>"011111010",
  56071=>"101001101",
  56072=>"100111010",
  56073=>"000000101",
  56074=>"100101101",
  56075=>"100111111",
  56076=>"001000001",
  56077=>"101101100",
  56078=>"111111000",
  56079=>"000011111",
  56080=>"111111110",
  56081=>"111111011",
  56082=>"101101101",
  56083=>"111001001",
  56084=>"111101000",
  56085=>"111111010",
  56086=>"100100100",
  56087=>"100000111",
  56088=>"000000110",
  56089=>"000000000",
  56090=>"111111111",
  56091=>"111111111",
  56092=>"001001001",
  56093=>"111111111",
  56094=>"101101101",
  56095=>"000000000",
  56096=>"000000111",
  56097=>"100000100",
  56098=>"000000010",
  56099=>"010110110",
  56100=>"010110110",
  56101=>"100110111",
  56102=>"011001000",
  56103=>"011110010",
  56104=>"000100000",
  56105=>"001000000",
  56106=>"100110110",
  56107=>"101100100",
  56108=>"100100100",
  56109=>"011111111",
  56110=>"101000111",
  56111=>"101101001",
  56112=>"111111110",
  56113=>"100000000",
  56114=>"110110000",
  56115=>"010010000",
  56116=>"111100010",
  56117=>"101101100",
  56118=>"111111101",
  56119=>"100100101",
  56120=>"110110110",
  56121=>"100100101",
  56122=>"001001001",
  56123=>"101101111",
  56124=>"111001001",
  56125=>"101101111",
  56126=>"110000111",
  56127=>"011011111",
  56128=>"101111111",
  56129=>"101101111",
  56130=>"000110111",
  56131=>"101101111",
  56132=>"101111111",
  56133=>"001111100",
  56134=>"000001111",
  56135=>"110100111",
  56136=>"111111111",
  56137=>"011000000",
  56138=>"000000100",
  56139=>"000000000",
  56140=>"000000000",
  56141=>"111111111",
  56142=>"111110010",
  56143=>"000000100",
  56144=>"001001001",
  56145=>"110010010",
  56146=>"100100110",
  56147=>"100100100",
  56148=>"100100100",
  56149=>"001001011",
  56150=>"000000000",
  56151=>"011011011",
  56152=>"001001111",
  56153=>"011000000",
  56154=>"011011011",
  56155=>"110111111",
  56156=>"000000000",
  56157=>"111111111",
  56158=>"010011111",
  56159=>"100010110",
  56160=>"111001001",
  56161=>"011111111",
  56162=>"001001001",
  56163=>"111111111",
  56164=>"100100100",
  56165=>"110000000",
  56166=>"000010111",
  56167=>"101101000",
  56168=>"000000000",
  56169=>"111011011",
  56170=>"100000101",
  56171=>"101101101",
  56172=>"111111111",
  56173=>"110110010",
  56174=>"111111111",
  56175=>"001110101",
  56176=>"111011010",
  56177=>"111111111",
  56178=>"010010011",
  56179=>"111011001",
  56180=>"011011010",
  56181=>"111101001",
  56182=>"000000000",
  56183=>"100000100",
  56184=>"000000000",
  56185=>"110111100",
  56186=>"010010000",
  56187=>"100100000",
  56188=>"010010010",
  56189=>"000000000",
  56190=>"000000000",
  56191=>"100000100",
  56192=>"000100110",
  56193=>"110100000",
  56194=>"110100000",
  56195=>"011001000",
  56196=>"001101100",
  56197=>"111111111",
  56198=>"011011111",
  56199=>"111100100",
  56200=>"000101111",
  56201=>"101000000",
  56202=>"011011000",
  56203=>"110010000",
  56204=>"100000000",
  56205=>"100100100",
  56206=>"000111111",
  56207=>"011000100",
  56208=>"101101000",
  56209=>"111001001",
  56210=>"001001100",
  56211=>"100100100",
  56212=>"000111111",
  56213=>"110010010",
  56214=>"111110111",
  56215=>"010011111",
  56216=>"111101000",
  56217=>"000010000",
  56218=>"101111111",
  56219=>"101100100",
  56220=>"111111111",
  56221=>"111111101",
  56222=>"110111110",
  56223=>"001001001",
  56224=>"000000000",
  56225=>"101111011",
  56226=>"001101111",
  56227=>"111111101",
  56228=>"100110111",
  56229=>"111111100",
  56230=>"101000000",
  56231=>"010000101",
  56232=>"111111111",
  56233=>"111111100",
  56234=>"000000000",
  56235=>"111111000",
  56236=>"000111000",
  56237=>"111010000",
  56238=>"000010010",
  56239=>"000010011",
  56240=>"010010110",
  56241=>"101111011",
  56242=>"000111101",
  56243=>"100100000",
  56244=>"000000100",
  56245=>"101101101",
  56246=>"000001101",
  56247=>"101100000",
  56248=>"001111001",
  56249=>"000110000",
  56250=>"001001000",
  56251=>"111111111",
  56252=>"111111101",
  56253=>"100100100",
  56254=>"100100100",
  56255=>"110100000",
  56256=>"111111111",
  56257=>"100100001",
  56258=>"101101101",
  56259=>"001000000",
  56260=>"110110100",
  56261=>"101100100",
  56262=>"100000000",
  56263=>"101101101",
  56264=>"110110011",
  56265=>"001000000",
  56266=>"000000100",
  56267=>"011011111",
  56268=>"001101000",
  56269=>"011011111",
  56270=>"100101100",
  56271=>"011011001",
  56272=>"000000000",
  56273=>"000000000",
  56274=>"000001111",
  56275=>"111111111",
  56276=>"000000000",
  56277=>"111000000",
  56278=>"000001001",
  56279=>"000000100",
  56280=>"111111111",
  56281=>"000000111",
  56282=>"111011010",
  56283=>"111101101",
  56284=>"110110101",
  56285=>"000000101",
  56286=>"111011011",
  56287=>"110100000",
  56288=>"100100100",
  56289=>"000000000",
  56290=>"111001011",
  56291=>"101111111",
  56292=>"110010000",
  56293=>"010000000",
  56294=>"101001000",
  56295=>"000000000",
  56296=>"100000000",
  56297=>"000000000",
  56298=>"011111010",
  56299=>"110111111",
  56300=>"101101101",
  56301=>"100110011",
  56302=>"111111010",
  56303=>"110100000",
  56304=>"011011011",
  56305=>"001011111",
  56306=>"111011001",
  56307=>"101101001",
  56308=>"001011111",
  56309=>"000010011",
  56310=>"011001100",
  56311=>"111111000",
  56312=>"001101011",
  56313=>"001001001",
  56314=>"000000100",
  56315=>"101101000",
  56316=>"101111101",
  56317=>"010110010",
  56318=>"011011011",
  56319=>"111000010",
  56320=>"000000000",
  56321=>"110110111",
  56322=>"000000101",
  56323=>"010000000",
  56324=>"011111111",
  56325=>"100110110",
  56326=>"110111011",
  56327=>"000000000",
  56328=>"000010000",
  56329=>"111111111",
  56330=>"011110111",
  56331=>"111111111",
  56332=>"011011111",
  56333=>"000000001",
  56334=>"100100111",
  56335=>"010000000",
  56336=>"000000000",
  56337=>"001001111",
  56338=>"111111010",
  56339=>"110110110",
  56340=>"000011000",
  56341=>"111111111",
  56342=>"111110110",
  56343=>"101101111",
  56344=>"101100100",
  56345=>"000001000",
  56346=>"100100111",
  56347=>"110111111",
  56348=>"000000001",
  56349=>"010111111",
  56350=>"011001000",
  56351=>"000000000",
  56352=>"001001001",
  56353=>"000000000",
  56354=>"000000000",
  56355=>"111111100",
  56356=>"111111111",
  56357=>"111011111",
  56358=>"000000000",
  56359=>"110111111",
  56360=>"111111111",
  56361=>"000111000",
  56362=>"101100000",
  56363=>"000000101",
  56364=>"101111100",
  56365=>"111111001",
  56366=>"111111110",
  56367=>"111111111",
  56368=>"011000000",
  56369=>"000000000",
  56370=>"011011011",
  56371=>"000110110",
  56372=>"000001001",
  56373=>"001000000",
  56374=>"011011011",
  56375=>"111000001",
  56376=>"000001111",
  56377=>"000000000",
  56378=>"111111111",
  56379=>"001011111",
  56380=>"000000000",
  56381=>"001000000",
  56382=>"111111001",
  56383=>"111111110",
  56384=>"011111100",
  56385=>"011011011",
  56386=>"010110111",
  56387=>"000100111",
  56388=>"000000100",
  56389=>"111000000",
  56390=>"100000100",
  56391=>"111111111",
  56392=>"011111111",
  56393=>"100110111",
  56394=>"111000000",
  56395=>"000000000",
  56396=>"110010001",
  56397=>"110110000",
  56398=>"101101000",
  56399=>"000000100",
  56400=>"100110110",
  56401=>"000000000",
  56402=>"111111010",
  56403=>"111101000",
  56404=>"000001001",
  56405=>"110111110",
  56406=>"001001011",
  56407=>"111000000",
  56408=>"100001011",
  56409=>"000000000",
  56410=>"000000000",
  56411=>"110110100",
  56412=>"111111111",
  56413=>"010111110",
  56414=>"111111110",
  56415=>"000110111",
  56416=>"001000111",
  56417=>"000111000",
  56418=>"111111111",
  56419=>"111111001",
  56420=>"111111111",
  56421=>"001001111",
  56422=>"110000000",
  56423=>"111111111",
  56424=>"110000101",
  56425=>"111111011",
  56426=>"111111011",
  56427=>"111111111",
  56428=>"110111011",
  56429=>"000000110",
  56430=>"001000001",
  56431=>"110111000",
  56432=>"000111111",
  56433=>"110111100",
  56434=>"000000001",
  56435=>"110000001",
  56436=>"100000000",
  56437=>"110111110",
  56438=>"000111011",
  56439=>"100000000",
  56440=>"111111111",
  56441=>"111111110",
  56442=>"111000000",
  56443=>"111111111",
  56444=>"000100000",
  56445=>"111111010",
  56446=>"100000000",
  56447=>"000110110",
  56448=>"111111111",
  56449=>"001111111",
  56450=>"000000000",
  56451=>"111011001",
  56452=>"101000000",
  56453=>"010010000",
  56454=>"000000000",
  56455=>"011101100",
  56456=>"000111110",
  56457=>"111111011",
  56458=>"011111000",
  56459=>"000001111",
  56460=>"111111111",
  56461=>"111110000",
  56462=>"000001001",
  56463=>"111110110",
  56464=>"000001111",
  56465=>"111001111",
  56466=>"001110011",
  56467=>"111110000",
  56468=>"111111000",
  56469=>"111111111",
  56470=>"100110111",
  56471=>"011001000",
  56472=>"000000001",
  56473=>"011000000",
  56474=>"111111011",
  56475=>"001011001",
  56476=>"111100100",
  56477=>"110110111",
  56478=>"011010000",
  56479=>"000001001",
  56480=>"000111100",
  56481=>"000000000",
  56482=>"001001111",
  56483=>"111000000",
  56484=>"000000000",
  56485=>"000110110",
  56486=>"001001111",
  56487=>"000000000",
  56488=>"110110111",
  56489=>"000001001",
  56490=>"000000000",
  56491=>"000000111",
  56492=>"111110101",
  56493=>"000000000",
  56494=>"111111111",
  56495=>"100001111",
  56496=>"000111011",
  56497=>"000000000",
  56498=>"111111111",
  56499=>"001111111",
  56500=>"111110110",
  56501=>"110100000",
  56502=>"000000000",
  56503=>"011000111",
  56504=>"000000001",
  56505=>"000000000",
  56506=>"101000110",
  56507=>"000000000",
  56508=>"011000101",
  56509=>"111111111",
  56510=>"111110111",
  56511=>"000000001",
  56512=>"001000000",
  56513=>"000000000",
  56514=>"000000111",
  56515=>"000111111",
  56516=>"000110110",
  56517=>"000000000",
  56518=>"000000000",
  56519=>"000101111",
  56520=>"000000010",
  56521=>"000000110",
  56522=>"111110110",
  56523=>"000000000",
  56524=>"000001001",
  56525=>"111111111",
  56526=>"110110000",
  56527=>"111111111",
  56528=>"110100110",
  56529=>"111111111",
  56530=>"111111111",
  56531=>"000000000",
  56532=>"001001111",
  56533=>"111111110",
  56534=>"000000000",
  56535=>"111001001",
  56536=>"011111100",
  56537=>"111111111",
  56538=>"000000000",
  56539=>"000000000",
  56540=>"000000011",
  56541=>"000110100",
  56542=>"000000000",
  56543=>"001100100",
  56544=>"000111111",
  56545=>"111111111",
  56546=>"000011111",
  56547=>"111111110",
  56548=>"111000000",
  56549=>"111111111",
  56550=>"000010000",
  56551=>"111001111",
  56552=>"011111000",
  56553=>"000000000",
  56554=>"001000111",
  56555=>"111001000",
  56556=>"000110000",
  56557=>"000000000",
  56558=>"111111101",
  56559=>"000000111",
  56560=>"111111000",
  56561=>"000000100",
  56562=>"111000111",
  56563=>"000000000",
  56564=>"111111111",
  56565=>"111111111",
  56566=>"000100100",
  56567=>"001011000",
  56568=>"001000111",
  56569=>"000000001",
  56570=>"000111010",
  56571=>"001000101",
  56572=>"000000111",
  56573=>"100100110",
  56574=>"111111000",
  56575=>"000110000",
  56576=>"000000000",
  56577=>"000000000",
  56578=>"000000000",
  56579=>"110100110",
  56580=>"100110111",
  56581=>"000000000",
  56582=>"001000001",
  56583=>"110110111",
  56584=>"011111011",
  56585=>"111111111",
  56586=>"110111111",
  56587=>"001001111",
  56588=>"001111111",
  56589=>"111000100",
  56590=>"000000111",
  56591=>"000111011",
  56592=>"000011011",
  56593=>"000000100",
  56594=>"101110110",
  56595=>"001010110",
  56596=>"111110000",
  56597=>"111111111",
  56598=>"001000000",
  56599=>"001011011",
  56600=>"001001100",
  56601=>"000100000",
  56602=>"110110000",
  56603=>"111110100",
  56604=>"000110110",
  56605=>"100000000",
  56606=>"011000011",
  56607=>"001001111",
  56608=>"100000000",
  56609=>"111110100",
  56610=>"111111111",
  56611=>"101111110",
  56612=>"000000000",
  56613=>"111111111",
  56614=>"001001111",
  56615=>"111111010",
  56616=>"000000000",
  56617=>"011111111",
  56618=>"101111110",
  56619=>"000000000",
  56620=>"000000000",
  56621=>"100110110",
  56622=>"111111000",
  56623=>"000000001",
  56624=>"000110100",
  56625=>"100000000",
  56626=>"000000000",
  56627=>"111011011",
  56628=>"011000000",
  56629=>"111110001",
  56630=>"101000000",
  56631=>"011011111",
  56632=>"111101000",
  56633=>"101000000",
  56634=>"000000010",
  56635=>"000011011",
  56636=>"000000000",
  56637=>"110010010",
  56638=>"111111111",
  56639=>"111101000",
  56640=>"111101100",
  56641=>"000000001",
  56642=>"111111111",
  56643=>"101101000",
  56644=>"000000110",
  56645=>"111000111",
  56646=>"100111111",
  56647=>"000011011",
  56648=>"011000111",
  56649=>"000010111",
  56650=>"001111111",
  56651=>"001111111",
  56652=>"110110110",
  56653=>"110000000",
  56654=>"011111111",
  56655=>"101111111",
  56656=>"111111111",
  56657=>"111111111",
  56658=>"111110110",
  56659=>"111110100",
  56660=>"000000000",
  56661=>"011011001",
  56662=>"000000000",
  56663=>"000000001",
  56664=>"000000000",
  56665=>"000000001",
  56666=>"010011000",
  56667=>"110111100",
  56668=>"111111000",
  56669=>"111111111",
  56670=>"011000001",
  56671=>"000100110",
  56672=>"101000000",
  56673=>"101001111",
  56674=>"000000000",
  56675=>"000000000",
  56676=>"010011111",
  56677=>"000000000",
  56678=>"000000110",
  56679=>"111110111",
  56680=>"000111011",
  56681=>"100111111",
  56682=>"111100100",
  56683=>"110110111",
  56684=>"000100110",
  56685=>"001010011",
  56686=>"100000000",
  56687=>"000000000",
  56688=>"000000000",
  56689=>"111111111",
  56690=>"110110010",
  56691=>"111011000",
  56692=>"110100000",
  56693=>"000000000",
  56694=>"111111111",
  56695=>"011000010",
  56696=>"111111111",
  56697=>"000001001",
  56698=>"110001001",
  56699=>"110111111",
  56700=>"000100111",
  56701=>"000100110",
  56702=>"011000110",
  56703=>"111101101",
  56704=>"001000000",
  56705=>"101100101",
  56706=>"000000000",
  56707=>"000000000",
  56708=>"100100100",
  56709=>"000000000",
  56710=>"111001001",
  56711=>"001001111",
  56712=>"101001101",
  56713=>"111111111",
  56714=>"111000100",
  56715=>"100000000",
  56716=>"111111111",
  56717=>"000110100",
  56718=>"111110100",
  56719=>"000000000",
  56720=>"000000000",
  56721=>"000010111",
  56722=>"000011000",
  56723=>"001000101",
  56724=>"000000000",
  56725=>"010110000",
  56726=>"011001000",
  56727=>"000100111",
  56728=>"000011111",
  56729=>"111111111",
  56730=>"110000000",
  56731=>"110000110",
  56732=>"000001011",
  56733=>"111111000",
  56734=>"000000000",
  56735=>"111111001",
  56736=>"100000000",
  56737=>"000000000",
  56738=>"000010001",
  56739=>"111111100",
  56740=>"000110111",
  56741=>"111111110",
  56742=>"000000101",
  56743=>"001001000",
  56744=>"011000011",
  56745=>"111111111",
  56746=>"011111111",
  56747=>"011111000",
  56748=>"010010010",
  56749=>"111111111",
  56750=>"001001001",
  56751=>"100001101",
  56752=>"111111111",
  56753=>"101011111",
  56754=>"000110111",
  56755=>"000011001",
  56756=>"001001101",
  56757=>"010110111",
  56758=>"000000101",
  56759=>"111110111",
  56760=>"100110111",
  56761=>"001010111",
  56762=>"110111111",
  56763=>"100000010",
  56764=>"000000000",
  56765=>"110000000",
  56766=>"101101001",
  56767=>"000000000",
  56768=>"111111011",
  56769=>"000000000",
  56770=>"000000111",
  56771=>"010111111",
  56772=>"000010111",
  56773=>"001001001",
  56774=>"001111000",
  56775=>"000100000",
  56776=>"011111001",
  56777=>"011001110",
  56778=>"100100111",
  56779=>"000110000",
  56780=>"111010000",
  56781=>"111111111",
  56782=>"111000000",
  56783=>"111111111",
  56784=>"001101001",
  56785=>"000000001",
  56786=>"001001001",
  56787=>"000000000",
  56788=>"000000000",
  56789=>"110100110",
  56790=>"000100110",
  56791=>"001001011",
  56792=>"000000110",
  56793=>"100110111",
  56794=>"111111110",
  56795=>"000000000",
  56796=>"110000111",
  56797=>"110000001",
  56798=>"111001011",
  56799=>"000011000",
  56800=>"111111111",
  56801=>"100000000",
  56802=>"111000000",
  56803=>"000000000",
  56804=>"000010111",
  56805=>"000000000",
  56806=>"000000000",
  56807=>"110110110",
  56808=>"111100111",
  56809=>"000000100",
  56810=>"100011001",
  56811=>"111111111",
  56812=>"011001111",
  56813=>"100110111",
  56814=>"111111111",
  56815=>"001111111",
  56816=>"000100110",
  56817=>"011001001",
  56818=>"101001000",
  56819=>"011001001",
  56820=>"000000100",
  56821=>"111111001",
  56822=>"111111111",
  56823=>"110110000",
  56824=>"010000000",
  56825=>"111001001",
  56826=>"000000000",
  56827=>"100000000",
  56828=>"111011000",
  56829=>"001001001",
  56830=>"000000111",
  56831=>"000000110",
  56832=>"000100110",
  56833=>"111111111",
  56834=>"000000101",
  56835=>"000000000",
  56836=>"011000000",
  56837=>"111100111",
  56838=>"000000110",
  56839=>"000000001",
  56840=>"000100111",
  56841=>"000110100",
  56842=>"111111011",
  56843=>"000000001",
  56844=>"000111111",
  56845=>"111111111",
  56846=>"000000000",
  56847=>"000000111",
  56848=>"000111111",
  56849=>"011000000",
  56850=>"110000000",
  56851=>"111111100",
  56852=>"000000000",
  56853=>"110000000",
  56854=>"000000000",
  56855=>"000100000",
  56856=>"111111000",
  56857=>"011001101",
  56858=>"000000000",
  56859=>"000000100",
  56860=>"000000011",
  56861=>"111111111",
  56862=>"110110110",
  56863=>"011111111",
  56864=>"111111111",
  56865=>"101111100",
  56866=>"000000000",
  56867=>"111111111",
  56868=>"000000000",
  56869=>"100111111",
  56870=>"000001000",
  56871=>"000100111",
  56872=>"111111111",
  56873=>"000111111",
  56874=>"000000111",
  56875=>"111111111",
  56876=>"000000000",
  56877=>"111111111",
  56878=>"010111111",
  56879=>"111011011",
  56880=>"000000000",
  56881=>"000000000",
  56882=>"111111001",
  56883=>"010000111",
  56884=>"110100100",
  56885=>"110110110",
  56886=>"000000000",
  56887=>"000010010",
  56888=>"101001000",
  56889=>"000001100",
  56890=>"111101001",
  56891=>"000010111",
  56892=>"100000000",
  56893=>"000000000",
  56894=>"000000000",
  56895=>"000001000",
  56896=>"001011111",
  56897=>"000000100",
  56898=>"000000001",
  56899=>"000111000",
  56900=>"111111111",
  56901=>"000000011",
  56902=>"000000000",
  56903=>"000000000",
  56904=>"100100000",
  56905=>"101101111",
  56906=>"000000000",
  56907=>"111111111",
  56908=>"101111111",
  56909=>"110000100",
  56910=>"000110111",
  56911=>"111111111",
  56912=>"000001011",
  56913=>"011111010",
  56914=>"111000000",
  56915=>"111011110",
  56916=>"111111001",
  56917=>"000111110",
  56918=>"000000000",
  56919=>"000000000",
  56920=>"100000000",
  56921=>"111001000",
  56922=>"000000110",
  56923=>"110111111",
  56924=>"111111111",
  56925=>"000111111",
  56926=>"101111111",
  56927=>"011011111",
  56928=>"000110101",
  56929=>"011111111",
  56930=>"011111111",
  56931=>"000111111",
  56932=>"001001001",
  56933=>"000000000",
  56934=>"101000001",
  56935=>"000100010",
  56936=>"111111111",
  56937=>"111111111",
  56938=>"000000000",
  56939=>"111010110",
  56940=>"110000001",
  56941=>"000000000",
  56942=>"000111111",
  56943=>"000000100",
  56944=>"111111011",
  56945=>"000111111",
  56946=>"000000000",
  56947=>"100110110",
  56948=>"001001000",
  56949=>"111111110",
  56950=>"000000000",
  56951=>"000000000",
  56952=>"111111001",
  56953=>"111111111",
  56954=>"000000000",
  56955=>"000001011",
  56956=>"110111111",
  56957=>"000000000",
  56958=>"000000110",
  56959=>"111111000",
  56960=>"000000000",
  56961=>"000000000",
  56962=>"000001101",
  56963=>"100000000",
  56964=>"000000111",
  56965=>"111111111",
  56966=>"100110000",
  56967=>"100000000",
  56968=>"100100111",
  56969=>"000000000",
  56970=>"101111111",
  56971=>"111101111",
  56972=>"000000000",
  56973=>"111111111",
  56974=>"000000000",
  56975=>"000011011",
  56976=>"000000000",
  56977=>"000100111",
  56978=>"001000000",
  56979=>"000000000",
  56980=>"111001101",
  56981=>"000000001",
  56982=>"111111111",
  56983=>"000000000",
  56984=>"111001111",
  56985=>"001000011",
  56986=>"111000000",
  56987=>"110100000",
  56988=>"000000100",
  56989=>"111111101",
  56990=>"111111111",
  56991=>"000111111",
  56992=>"000000000",
  56993=>"000101000",
  56994=>"100000000",
  56995=>"000111111",
  56996=>"011011001",
  56997=>"000110000",
  56998=>"011111111",
  56999=>"000100100",
  57000=>"000000100",
  57001=>"000000000",
  57002=>"000000000",
  57003=>"111111111",
  57004=>"011000000",
  57005=>"000110111",
  57006=>"001001101",
  57007=>"111011110",
  57008=>"000110110",
  57009=>"111111111",
  57010=>"000111111",
  57011=>"000000000",
  57012=>"111111111",
  57013=>"110110000",
  57014=>"010111011",
  57015=>"000000000",
  57016=>"111111111",
  57017=>"111111111",
  57018=>"101000001",
  57019=>"001000000",
  57020=>"000001111",
  57021=>"111111111",
  57022=>"110110110",
  57023=>"111111111",
  57024=>"000000000",
  57025=>"111111111",
  57026=>"111111111",
  57027=>"011001100",
  57028=>"000100000",
  57029=>"000000000",
  57030=>"001001111",
  57031=>"000000000",
  57032=>"111111111",
  57033=>"111111111",
  57034=>"111000101",
  57035=>"000000000",
  57036=>"111111111",
  57037=>"000000111",
  57038=>"110110111",
  57039=>"111111111",
  57040=>"000000000",
  57041=>"000010111",
  57042=>"010011111",
  57043=>"000010011",
  57044=>"011111111",
  57045=>"111111111",
  57046=>"111000000",
  57047=>"111111011",
  57048=>"001000000",
  57049=>"001111110",
  57050=>"111111110",
  57051=>"000100000",
  57052=>"010011011",
  57053=>"100110000",
  57054=>"100111111",
  57055=>"111111101",
  57056=>"111111111",
  57057=>"000000000",
  57058=>"010000000",
  57059=>"111111111",
  57060=>"001000000",
  57061=>"100110111",
  57062=>"111111000",
  57063=>"110000110",
  57064=>"011011101",
  57065=>"000000000",
  57066=>"111111111",
  57067=>"111111011",
  57068=>"000000000",
  57069=>"000000111",
  57070=>"000010100",
  57071=>"111001000",
  57072=>"000000000",
  57073=>"000000000",
  57074=>"111111111",
  57075=>"000001001",
  57076=>"000000000",
  57077=>"100110111",
  57078=>"111011001",
  57079=>"111000000",
  57080=>"111111011",
  57081=>"000011000",
  57082=>"000000111",
  57083=>"111111111",
  57084=>"111011001",
  57085=>"000000000",
  57086=>"000000011",
  57087=>"100110110",
  57088=>"111111010",
  57089=>"000000000",
  57090=>"000000000",
  57091=>"001000000",
  57092=>"000000000",
  57093=>"110111110",
  57094=>"111111111",
  57095=>"011011011",
  57096=>"110111111",
  57097=>"001000000",
  57098=>"111111111",
  57099=>"000000000",
  57100=>"101000000",
  57101=>"000001001",
  57102=>"111111111",
  57103=>"111111000",
  57104=>"000011111",
  57105=>"111111001",
  57106=>"111111001",
  57107=>"001100000",
  57108=>"111111111",
  57109=>"111111000",
  57110=>"111100000",
  57111=>"000110110",
  57112=>"011111011",
  57113=>"011110100",
  57114=>"111111111",
  57115=>"000000000",
  57116=>"110110111",
  57117=>"000000000",
  57118=>"000010000",
  57119=>"111111011",
  57120=>"100110000",
  57121=>"011111111",
  57122=>"111111100",
  57123=>"111001000",
  57124=>"111111000",
  57125=>"100000000",
  57126=>"101001000",
  57127=>"000000110",
  57128=>"111111111",
  57129=>"000000000",
  57130=>"011001111",
  57131=>"000000000",
  57132=>"111110110",
  57133=>"111111010",
  57134=>"000000000",
  57135=>"011000011",
  57136=>"000000000",
  57137=>"000000001",
  57138=>"000001111",
  57139=>"001111111",
  57140=>"000000000",
  57141=>"101100111",
  57142=>"000000000",
  57143=>"111111111",
  57144=>"111111111",
  57145=>"000000001",
  57146=>"000000011",
  57147=>"100000100",
  57148=>"000000000",
  57149=>"000000000",
  57150=>"011001000",
  57151=>"011001000",
  57152=>"111111100",
  57153=>"101111011",
  57154=>"110111001",
  57155=>"110111111",
  57156=>"110000111",
  57157=>"010010000",
  57158=>"011001000",
  57159=>"110100111",
  57160=>"000000000",
  57161=>"000000001",
  57162=>"110110000",
  57163=>"001000100",
  57164=>"100010000",
  57165=>"011000000",
  57166=>"111111111",
  57167=>"101111000",
  57168=>"000001011",
  57169=>"111110111",
  57170=>"000000111",
  57171=>"000000111",
  57172=>"100100111",
  57173=>"011011011",
  57174=>"111101000",
  57175=>"001111110",
  57176=>"000000111",
  57177=>"000100000",
  57178=>"111111111",
  57179=>"111100101",
  57180=>"111111111",
  57181=>"111111111",
  57182=>"111111111",
  57183=>"100110000",
  57184=>"010110010",
  57185=>"000000000",
  57186=>"011111001",
  57187=>"000000000",
  57188=>"101111111",
  57189=>"001000000",
  57190=>"000000000",
  57191=>"000000000",
  57192=>"000111111",
  57193=>"101000000",
  57194=>"000000000",
  57195=>"000000100",
  57196=>"000000000",
  57197=>"111111101",
  57198=>"100000001",
  57199=>"011111111",
  57200=>"000000000",
  57201=>"101100000",
  57202=>"000110101",
  57203=>"010110110",
  57204=>"000000000",
  57205=>"000000000",
  57206=>"000000000",
  57207=>"111110111",
  57208=>"000000000",
  57209=>"110111111",
  57210=>"111111111",
  57211=>"001101111",
  57212=>"111111111",
  57213=>"111111111",
  57214=>"011011111",
  57215=>"000000100",
  57216=>"111010000",
  57217=>"111111101",
  57218=>"000000000",
  57219=>"001101111",
  57220=>"110111100",
  57221=>"111111111",
  57222=>"011111000",
  57223=>"101111111",
  57224=>"000000010",
  57225=>"000000000",
  57226=>"000000111",
  57227=>"111100000",
  57228=>"111111111",
  57229=>"000110100",
  57230=>"000000000",
  57231=>"010110111",
  57232=>"111000000",
  57233=>"000101111",
  57234=>"111111111",
  57235=>"000000000",
  57236=>"000011011",
  57237=>"101000000",
  57238=>"011100100",
  57239=>"010000000",
  57240=>"100111111",
  57241=>"000100100",
  57242=>"001000000",
  57243=>"000000000",
  57244=>"110000011",
  57245=>"111111110",
  57246=>"000000000",
  57247=>"000000111",
  57248=>"000100110",
  57249=>"111110000",
  57250=>"000001111",
  57251=>"000000010",
  57252=>"000000000",
  57253=>"000000001",
  57254=>"000111111",
  57255=>"011111111",
  57256=>"000010111",
  57257=>"000111111",
  57258=>"100000111",
  57259=>"111011011",
  57260=>"000000000",
  57261=>"111111111",
  57262=>"000000110",
  57263=>"000000110",
  57264=>"111111111",
  57265=>"101111111",
  57266=>"110000000",
  57267=>"000000000",
  57268=>"001001001",
  57269=>"000000000",
  57270=>"111111111",
  57271=>"000000111",
  57272=>"000000000",
  57273=>"000111100",
  57274=>"000011111",
  57275=>"000000000",
  57276=>"000100000",
  57277=>"111111111",
  57278=>"111111111",
  57279=>"000000000",
  57280=>"111000011",
  57281=>"111101000",
  57282=>"111111111",
  57283=>"000100000",
  57284=>"111111111",
  57285=>"111110100",
  57286=>"000000000",
  57287=>"000111111",
  57288=>"111000001",
  57289=>"111111100",
  57290=>"011000000",
  57291=>"000000111",
  57292=>"100000000",
  57293=>"000000000",
  57294=>"000110100",
  57295=>"111110100",
  57296=>"000010111",
  57297=>"000000000",
  57298=>"100100111",
  57299=>"111111000",
  57300=>"111111111",
  57301=>"000000100",
  57302=>"011101111",
  57303=>"110000111",
  57304=>"000000111",
  57305=>"111111101",
  57306=>"000000000",
  57307=>"000000111",
  57308=>"000000100",
  57309=>"000000000",
  57310=>"000000000",
  57311=>"000001000",
  57312=>"111000000",
  57313=>"000000001",
  57314=>"111101101",
  57315=>"001111111",
  57316=>"001011000",
  57317=>"110110110",
  57318=>"000011011",
  57319=>"010010010",
  57320=>"000000011",
  57321=>"111111111",
  57322=>"001001111",
  57323=>"101111101",
  57324=>"111010000",
  57325=>"000000000",
  57326=>"111111111",
  57327=>"111111111",
  57328=>"000000000",
  57329=>"110111111",
  57330=>"111101000",
  57331=>"111111111",
  57332=>"101000111",
  57333=>"000000100",
  57334=>"011011001",
  57335=>"010111010",
  57336=>"111001000",
  57337=>"111111111",
  57338=>"001000000",
  57339=>"011111111",
  57340=>"000000000",
  57341=>"111001001",
  57342=>"111111111",
  57343=>"000000000",
  57344=>"000011001",
  57345=>"001000000",
  57346=>"001111111",
  57347=>"111111000",
  57348=>"111110000",
  57349=>"111100100",
  57350=>"000110000",
  57351=>"000100111",
  57352=>"000111111",
  57353=>"010000011",
  57354=>"000000000",
  57355=>"000000000",
  57356=>"111111111",
  57357=>"000000000",
  57358=>"001000000",
  57359=>"011111111",
  57360=>"000001001",
  57361=>"000001001",
  57362=>"111111001",
  57363=>"010000000",
  57364=>"100100000",
  57365=>"000000001",
  57366=>"000000000",
  57367=>"010100110",
  57368=>"000000110",
  57369=>"011000000",
  57370=>"000000011",
  57371=>"011011011",
  57372=>"000000100",
  57373=>"100000000",
  57374=>"011010000",
  57375=>"111111111",
  57376=>"000000000",
  57377=>"010000000",
  57378=>"000100111",
  57379=>"011000000",
  57380=>"000000000",
  57381=>"000000110",
  57382=>"111111111",
  57383=>"000000000",
  57384=>"011000000",
  57385=>"101000111",
  57386=>"000000000",
  57387=>"111111111",
  57388=>"111111111",
  57389=>"000000000",
  57390=>"111000000",
  57391=>"111101111",
  57392=>"110100100",
  57393=>"000000000",
  57394=>"000010111",
  57395=>"000000000",
  57396=>"111111111",
  57397=>"001111111",
  57398=>"111011000",
  57399=>"110111111",
  57400=>"000110010",
  57401=>"000000010",
  57402=>"000000001",
  57403=>"000000011",
  57404=>"000000000",
  57405=>"111000000",
  57406=>"101111111",
  57407=>"000000111",
  57408=>"000000000",
  57409=>"001100110",
  57410=>"000000111",
  57411=>"111111111",
  57412=>"000101111",
  57413=>"100000000",
  57414=>"000000000",
  57415=>"000000111",
  57416=>"111111100",
  57417=>"111110000",
  57418=>"111111111",
  57419=>"111111111",
  57420=>"111000000",
  57421=>"000100111",
  57422=>"110000000",
  57423=>"000000000",
  57424=>"111111111",
  57425=>"001000001",
  57426=>"000000010",
  57427=>"011011001",
  57428=>"000110110",
  57429=>"000000000",
  57430=>"001000001",
  57431=>"111001000",
  57432=>"111111000",
  57433=>"000100111",
  57434=>"111111111",
  57435=>"011001001",
  57436=>"000000000",
  57437=>"000001000",
  57438=>"001110100",
  57439=>"110110110",
  57440=>"000101111",
  57441=>"110111111",
  57442=>"000000000",
  57443=>"000000000",
  57444=>"000000111",
  57445=>"000110000",
  57446=>"001001000",
  57447=>"000000001",
  57448=>"111111111",
  57449=>"110110111",
  57450=>"001000111",
  57451=>"000111111",
  57452=>"001111111",
  57453=>"100111111",
  57454=>"000000000",
  57455=>"000111111",
  57456=>"000011001",
  57457=>"101111001",
  57458=>"111011011",
  57459=>"000000011",
  57460=>"000000000",
  57461=>"111001000",
  57462=>"001100000",
  57463=>"000000111",
  57464=>"000110100",
  57465=>"000111111",
  57466=>"000100111",
  57467=>"111111111",
  57468=>"001001001",
  57469=>"000000000",
  57470=>"000000111",
  57471=>"000000000",
  57472=>"111111011",
  57473=>"001000011",
  57474=>"111010011",
  57475=>"011000000",
  57476=>"001000000",
  57477=>"110000111",
  57478=>"111000000",
  57479=>"111111111",
  57480=>"111000000",
  57481=>"111011111",
  57482=>"000000000",
  57483=>"111000000",
  57484=>"100000000",
  57485=>"111111000",
  57486=>"111111111",
  57487=>"111110000",
  57488=>"000001111",
  57489=>"110111111",
  57490=>"111111111",
  57491=>"000110111",
  57492=>"000100110",
  57493=>"010110000",
  57494=>"111111100",
  57495=>"111111000",
  57496=>"000000110",
  57497=>"100100101",
  57498=>"001000000",
  57499=>"100000000",
  57500=>"100000000",
  57501=>"000100110",
  57502=>"000101101",
  57503=>"111111111",
  57504=>"100000000",
  57505=>"000000101",
  57506=>"111111111",
  57507=>"011011011",
  57508=>"000001001",
  57509=>"000100000",
  57510=>"000110110",
  57511=>"000100110",
  57512=>"001001000",
  57513=>"000000001",
  57514=>"111000000",
  57515=>"000000011",
  57516=>"111111111",
  57517=>"001001000",
  57518=>"001000000",
  57519=>"000000000",
  57520=>"000000011",
  57521=>"110110000",
  57522=>"110110110",
  57523=>"111110000",
  57524=>"101101100",
  57525=>"111111101",
  57526=>"000011101",
  57527=>"111111100",
  57528=>"111001000",
  57529=>"100000000",
  57530=>"001111111",
  57531=>"100111111",
  57532=>"001011111",
  57533=>"101000000",
  57534=>"100110000",
  57535=>"000000111",
  57536=>"010000000",
  57537=>"111111111",
  57538=>"101101000",
  57539=>"111111111",
  57540=>"011011011",
  57541=>"000000110",
  57542=>"110111111",
  57543=>"100000100",
  57544=>"111101110",
  57545=>"010000101",
  57546=>"011000000",
  57547=>"110110000",
  57548=>"000000000",
  57549=>"111111111",
  57550=>"100000101",
  57551=>"000000001",
  57552=>"111111100",
  57553=>"111110100",
  57554=>"110000100",
  57555=>"000000000",
  57556=>"001001000",
  57557=>"100100110",
  57558=>"111111111",
  57559=>"111111111",
  57560=>"111111110",
  57561=>"001000111",
  57562=>"111111000",
  57563=>"111111100",
  57564=>"111111111",
  57565=>"111111000",
  57566=>"000000111",
  57567=>"101111001",
  57568=>"111111111",
  57569=>"001000000",
  57570=>"111000000",
  57571=>"111111000",
  57572=>"000000000",
  57573=>"110110100",
  57574=>"001101111",
  57575=>"100000000",
  57576=>"111111000",
  57577=>"100010000",
  57578=>"111000000",
  57579=>"000000000",
  57580=>"001111011",
  57581=>"000100110",
  57582=>"000000000",
  57583=>"000111111",
  57584=>"000000000",
  57585=>"111110000",
  57586=>"111111011",
  57587=>"100111000",
  57588=>"111110111",
  57589=>"001001010",
  57590=>"010011000",
  57591=>"100111111",
  57592=>"111001000",
  57593=>"100111110",
  57594=>"001001111",
  57595=>"000111111",
  57596=>"110111111",
  57597=>"111110010",
  57598=>"000011111",
  57599=>"111000100",
  57600=>"111001000",
  57601=>"011010001",
  57602=>"000111111",
  57603=>"000001000",
  57604=>"001111111",
  57605=>"100100000",
  57606=>"111111100",
  57607=>"000100111",
  57608=>"111101101",
  57609=>"101111111",
  57610=>"111111000",
  57611=>"001001000",
  57612=>"000000111",
  57613=>"111011000",
  57614=>"111000111",
  57615=>"111111000",
  57616=>"100100000",
  57617=>"000001111",
  57618=>"111110100",
  57619=>"111000000",
  57620=>"111111111",
  57621=>"001001011",
  57622=>"111111001",
  57623=>"001000000",
  57624=>"111001001",
  57625=>"000000000",
  57626=>"000000000",
  57627=>"110111100",
  57628=>"111110000",
  57629=>"000000000",
  57630=>"000010000",
  57631=>"000000000",
  57632=>"000100110",
  57633=>"110100000",
  57634=>"111000000",
  57635=>"001111111",
  57636=>"000000110",
  57637=>"000011111",
  57638=>"011111111",
  57639=>"101111111",
  57640=>"000000000",
  57641=>"111111000",
  57642=>"111111100",
  57643=>"111111000",
  57644=>"000000100",
  57645=>"000001001",
  57646=>"000000000",
  57647=>"001000000",
  57648=>"100010111",
  57649=>"010000101",
  57650=>"000000000",
  57651=>"111111111",
  57652=>"000000000",
  57653=>"100111111",
  57654=>"111110110",
  57655=>"111111000",
  57656=>"010111000",
  57657=>"000000000",
  57658=>"110000000",
  57659=>"111000000",
  57660=>"000000000",
  57661=>"000000111",
  57662=>"000110000",
  57663=>"100101110",
  57664=>"000000000",
  57665=>"111110111",
  57666=>"110110000",
  57667=>"111100100",
  57668=>"001111110",
  57669=>"000001000",
  57670=>"000111111",
  57671=>"000000000",
  57672=>"000000011",
  57673=>"111111000",
  57674=>"001111101",
  57675=>"110110110",
  57676=>"000000011",
  57677=>"111111000",
  57678=>"001111111",
  57679=>"110110110",
  57680=>"110110010",
  57681=>"001011111",
  57682=>"111111111",
  57683=>"000110111",
  57684=>"000000000",
  57685=>"100110111",
  57686=>"110011110",
  57687=>"011001000",
  57688=>"111000000",
  57689=>"100000100",
  57690=>"000000111",
  57691=>"111100111",
  57692=>"000011011",
  57693=>"010011001",
  57694=>"100100101",
  57695=>"111111001",
  57696=>"000001111",
  57697=>"100000101",
  57698=>"111110000",
  57699=>"000000100",
  57700=>"110111000",
  57701=>"001101001",
  57702=>"111111000",
  57703=>"000000100",
  57704=>"111011001",
  57705=>"111011011",
  57706=>"111111111",
  57707=>"011011011",
  57708=>"111010000",
  57709=>"011001001",
  57710=>"001101110",
  57711=>"011111111",
  57712=>"000010110",
  57713=>"000100111",
  57714=>"111011111",
  57715=>"111110110",
  57716=>"000000110",
  57717=>"111111100",
  57718=>"000100111",
  57719=>"000100000",
  57720=>"100000000",
  57721=>"100000000",
  57722=>"110000000",
  57723=>"000001000",
  57724=>"110111111",
  57725=>"000000000",
  57726=>"111111111",
  57727=>"000000001",
  57728=>"000001000",
  57729=>"000001000",
  57730=>"000000000",
  57731=>"000000000",
  57732=>"000000111",
  57733=>"111000100",
  57734=>"111111111",
  57735=>"000101001",
  57736=>"010000001",
  57737=>"011111111",
  57738=>"100100111",
  57739=>"111111000",
  57740=>"000101111",
  57741=>"011011011",
  57742=>"001001101",
  57743=>"000010000",
  57744=>"111111111",
  57745=>"111001011",
  57746=>"111001000",
  57747=>"000000000",
  57748=>"111110110",
  57749=>"000000000",
  57750=>"111111001",
  57751=>"001001001",
  57752=>"111000000",
  57753=>"111010110",
  57754=>"111111100",
  57755=>"111111111",
  57756=>"100100000",
  57757=>"000101011",
  57758=>"110110111",
  57759=>"000000000",
  57760=>"111111111",
  57761=>"000000001",
  57762=>"000000110",
  57763=>"111111111",
  57764=>"001000111",
  57765=>"011111111",
  57766=>"000000111",
  57767=>"111111111",
  57768=>"011111110",
  57769=>"000000110",
  57770=>"111111110",
  57771=>"110111111",
  57772=>"000010000",
  57773=>"100111000",
  57774=>"111111111",
  57775=>"100000000",
  57776=>"000000111",
  57777=>"000000000",
  57778=>"000000110",
  57779=>"010111100",
  57780=>"110000101",
  57781=>"101100100",
  57782=>"000000000",
  57783=>"000000111",
  57784=>"100000011",
  57785=>"000000000",
  57786=>"000000001",
  57787=>"000001111",
  57788=>"000000000",
  57789=>"000000111",
  57790=>"010111111",
  57791=>"111111001",
  57792=>"001111010",
  57793=>"000000111",
  57794=>"111111111",
  57795=>"111100100",
  57796=>"011001101",
  57797=>"001001111",
  57798=>"111110000",
  57799=>"000111111",
  57800=>"000001111",
  57801=>"010000110",
  57802=>"101111110",
  57803=>"111111000",
  57804=>"001111000",
  57805=>"000010111",
  57806=>"000001100",
  57807=>"110000000",
  57808=>"111000001",
  57809=>"000000111",
  57810=>"111111110",
  57811=>"000000000",
  57812=>"111111000",
  57813=>"000101111",
  57814=>"000000111",
  57815=>"011111111",
  57816=>"010111110",
  57817=>"000000000",
  57818=>"111101001",
  57819=>"000001000",
  57820=>"000111010",
  57821=>"000000000",
  57822=>"111111111",
  57823=>"000000011",
  57824=>"000000111",
  57825=>"111111111",
  57826=>"111111111",
  57827=>"111111111",
  57828=>"100000000",
  57829=>"101111111",
  57830=>"000000111",
  57831=>"111111000",
  57832=>"101101100",
  57833=>"000110111",
  57834=>"000000100",
  57835=>"000000100",
  57836=>"100011110",
  57837=>"010010100",
  57838=>"000000000",
  57839=>"000010011",
  57840=>"000000111",
  57841=>"111111000",
  57842=>"111111111",
  57843=>"000111111",
  57844=>"001011011",
  57845=>"111111111",
  57846=>"111011000",
  57847=>"111000000",
  57848=>"000000000",
  57849=>"111110110",
  57850=>"110111000",
  57851=>"111111111",
  57852=>"111000111",
  57853=>"110111111",
  57854=>"111001011",
  57855=>"100000111",
  57856=>"000110100",
  57857=>"000010011",
  57858=>"000001101",
  57859=>"111111111",
  57860=>"010110110",
  57861=>"000000000",
  57862=>"000000001",
  57863=>"111111111",
  57864=>"000000000",
  57865=>"011111111",
  57866=>"000000101",
  57867=>"011000000",
  57868=>"000100000",
  57869=>"000000100",
  57870=>"111111111",
  57871=>"111111111",
  57872=>"101111011",
  57873=>"011111111",
  57874=>"000000000",
  57875=>"000000000",
  57876=>"111111111",
  57877=>"111111111",
  57878=>"111111111",
  57879=>"000000100",
  57880=>"000000000",
  57881=>"001001000",
  57882=>"111100101",
  57883=>"000000011",
  57884=>"111001000",
  57885=>"110111011",
  57886=>"110111110",
  57887=>"111111111",
  57888=>"111001011",
  57889=>"100101100",
  57890=>"000000000",
  57891=>"111111001",
  57892=>"000000000",
  57893=>"111111111",
  57894=>"000000000",
  57895=>"000000000",
  57896=>"000000100",
  57897=>"011011011",
  57898=>"111000000",
  57899=>"111111101",
  57900=>"000000000",
  57901=>"000000000",
  57902=>"111100000",
  57903=>"101111000",
  57904=>"111111100",
  57905=>"111111111",
  57906=>"110100100",
  57907=>"101111111",
  57908=>"111111000",
  57909=>"111111111",
  57910=>"111111001",
  57911=>"110111000",
  57912=>"111101000",
  57913=>"000000000",
  57914=>"111111111",
  57915=>"111111111",
  57916=>"111001001",
  57917=>"000100110",
  57918=>"001001011",
  57919=>"000000000",
  57920=>"000000001",
  57921=>"111111100",
  57922=>"000000000",
  57923=>"000000000",
  57924=>"100100100",
  57925=>"000000111",
  57926=>"001000000",
  57927=>"111111111",
  57928=>"101100100",
  57929=>"000000011",
  57930=>"110111100",
  57931=>"000010000",
  57932=>"111111111",
  57933=>"001111111",
  57934=>"111111111",
  57935=>"111111011",
  57936=>"000000111",
  57937=>"111111111",
  57938=>"111111000",
  57939=>"101100100",
  57940=>"111111111",
  57941=>"000111110",
  57942=>"100000001",
  57943=>"011001001",
  57944=>"110000000",
  57945=>"000000000",
  57946=>"111111111",
  57947=>"011011010",
  57948=>"111111111",
  57949=>"111111111",
  57950=>"000000110",
  57951=>"011111110",
  57952=>"000111111",
  57953=>"000000000",
  57954=>"011111111",
  57955=>"001000101",
  57956=>"111111011",
  57957=>"111001111",
  57958=>"111100110",
  57959=>"000000000",
  57960=>"011010000",
  57961=>"000000000",
  57962=>"000000000",
  57963=>"110110000",
  57964=>"110000000",
  57965=>"111111111",
  57966=>"100100111",
  57967=>"000001111",
  57968=>"000000000",
  57969=>"110111110",
  57970=>"111100100",
  57971=>"011111111",
  57972=>"000000000",
  57973=>"011111100",
  57974=>"000011010",
  57975=>"000111101",
  57976=>"000000000",
  57977=>"001001000",
  57978=>"100100000",
  57979=>"000000110",
  57980=>"101101101",
  57981=>"001000000",
  57982=>"000000000",
  57983=>"000000000",
  57984=>"000000000",
  57985=>"000011011",
  57986=>"111000111",
  57987=>"111111111",
  57988=>"000000000",
  57989=>"101000001",
  57990=>"111111001",
  57991=>"110110111",
  57992=>"000000001",
  57993=>"110111111",
  57994=>"110111111",
  57995=>"000000000",
  57996=>"011111111",
  57997=>"000100000",
  57998=>"111100110",
  57999=>"011111111",
  58000=>"101001000",
  58001=>"000010000",
  58002=>"001111111",
  58003=>"000000100",
  58004=>"001011111",
  58005=>"000000001",
  58006=>"000000000",
  58007=>"000000000",
  58008=>"000000000",
  58009=>"011001001",
  58010=>"011001001",
  58011=>"000000000",
  58012=>"000000000",
  58013=>"111011001",
  58014=>"111101000",
  58015=>"000000000",
  58016=>"111111111",
  58017=>"001000001",
  58018=>"111111111",
  58019=>"000000000",
  58020=>"110110111",
  58021=>"000111111",
  58022=>"000000000",
  58023=>"100110110",
  58024=>"000111111",
  58025=>"011000000",
  58026=>"000000000",
  58027=>"111101111",
  58028=>"100000001",
  58029=>"000000110",
  58030=>"111111111",
  58031=>"111110100",
  58032=>"110111110",
  58033=>"011000000",
  58034=>"010111010",
  58035=>"000000111",
  58036=>"111110011",
  58037=>"111111111",
  58038=>"001001001",
  58039=>"111111000",
  58040=>"111100100",
  58041=>"111101111",
  58042=>"011000001",
  58043=>"001011111",
  58044=>"101001111",
  58045=>"000010010",
  58046=>"111000001",
  58047=>"000000000",
  58048=>"111111111",
  58049=>"111111100",
  58050=>"000000001",
  58051=>"000000000",
  58052=>"000111111",
  58053=>"000000000",
  58054=>"000000000",
  58055=>"011000000",
  58056=>"111111111",
  58057=>"100100100",
  58058=>"001001000",
  58059=>"111001011",
  58060=>"100000000",
  58061=>"111111111",
  58062=>"111111111",
  58063=>"000000011",
  58064=>"000000000",
  58065=>"000110111",
  58066=>"111000111",
  58067=>"010111011",
  58068=>"001111110",
  58069=>"100100000",
  58070=>"000000000",
  58071=>"000000000",
  58072=>"000000000",
  58073=>"000100111",
  58074=>"000000110",
  58075=>"000011111",
  58076=>"110000001",
  58077=>"001000000",
  58078=>"010111100",
  58079=>"000000000",
  58080=>"000000000",
  58081=>"000111100",
  58082=>"000010010",
  58083=>"000000000",
  58084=>"001000000",
  58085=>"100100100",
  58086=>"000000000",
  58087=>"111111111",
  58088=>"111101111",
  58089=>"000000100",
  58090=>"000001001",
  58091=>"111011000",
  58092=>"111111011",
  58093=>"111001000",
  58094=>"010010011",
  58095=>"111011111",
  58096=>"000000000",
  58097=>"000000000",
  58098=>"000000111",
  58099=>"010010111",
  58100=>"111111011",
  58101=>"000000000",
  58102=>"000110000",
  58103=>"000100000",
  58104=>"111111111",
  58105=>"000000000",
  58106=>"111111111",
  58107=>"111011110",
  58108=>"000000000",
  58109=>"011011001",
  58110=>"000011011",
  58111=>"111101000",
  58112=>"110111011",
  58113=>"111101101",
  58114=>"011001000",
  58115=>"001000001",
  58116=>"000100100",
  58117=>"111011001",
  58118=>"101000101",
  58119=>"000000001",
  58120=>"100110111",
  58121=>"001111111",
  58122=>"111111111",
  58123=>"000000000",
  58124=>"000000000",
  58125=>"000000000",
  58126=>"000000000",
  58127=>"111111000",
  58128=>"000011111",
  58129=>"111111111",
  58130=>"000001011",
  58131=>"001001001",
  58132=>"000001000",
  58133=>"111111001",
  58134=>"100100111",
  58135=>"101101001",
  58136=>"111111111",
  58137=>"111111111",
  58138=>"000000000",
  58139=>"100100100",
  58140=>"000000000",
  58141=>"110000010",
  58142=>"010111110",
  58143=>"111111111",
  58144=>"001100111",
  58145=>"011111111",
  58146=>"000000000",
  58147=>"000000001",
  58148=>"011001011",
  58149=>"001101111",
  58150=>"000100000",
  58151=>"010111111",
  58152=>"001000000",
  58153=>"000001001",
  58154=>"111111111",
  58155=>"111111111",
  58156=>"001001110",
  58157=>"000000000",
  58158=>"100111111",
  58159=>"111111111",
  58160=>"000000000",
  58161=>"111011111",
  58162=>"111010000",
  58163=>"000000000",
  58164=>"000000000",
  58165=>"000011011",
  58166=>"000000010",
  58167=>"000000000",
  58168=>"000000000",
  58169=>"000000111",
  58170=>"000011011",
  58171=>"110111111",
  58172=>"000000000",
  58173=>"111111111",
  58174=>"110000000",
  58175=>"100000000",
  58176=>"100100000",
  58177=>"000000000",
  58178=>"111111111",
  58179=>"111111111",
  58180=>"000000000",
  58181=>"011000001",
  58182=>"000000000",
  58183=>"100100000",
  58184=>"111111111",
  58185=>"000000011",
  58186=>"111111101",
  58187=>"110000000",
  58188=>"111101101",
  58189=>"000001000",
  58190=>"001001111",
  58191=>"110110110",
  58192=>"111001101",
  58193=>"110111111",
  58194=>"001001011",
  58195=>"000000000",
  58196=>"000000001",
  58197=>"011000000",
  58198=>"111111111",
  58199=>"111111111",
  58200=>"000000000",
  58201=>"010010111",
  58202=>"000001111",
  58203=>"000000100",
  58204=>"001001000",
  58205=>"111111111",
  58206=>"010111111",
  58207=>"100101101",
  58208=>"010000000",
  58209=>"111111111",
  58210=>"000000000",
  58211=>"000000001",
  58212=>"000000000",
  58213=>"011000000",
  58214=>"000100110",
  58215=>"101101000",
  58216=>"111111111",
  58217=>"111100100",
  58218=>"000000001",
  58219=>"001001000",
  58220=>"000000000",
  58221=>"000000000",
  58222=>"001001010",
  58223=>"111111101",
  58224=>"011111001",
  58225=>"000000000",
  58226=>"000011111",
  58227=>"110111111",
  58228=>"000000000",
  58229=>"011000000",
  58230=>"111111111",
  58231=>"000001000",
  58232=>"000000111",
  58233=>"000011010",
  58234=>"111011011",
  58235=>"011011011",
  58236=>"011111111",
  58237=>"111111111",
  58238=>"001000011",
  58239=>"000000111",
  58240=>"000000001",
  58241=>"111111111",
  58242=>"101000000",
  58243=>"111111011",
  58244=>"000000000",
  58245=>"110100001",
  58246=>"001001011",
  58247=>"000000000",
  58248=>"000000001",
  58249=>"011011111",
  58250=>"001011111",
  58251=>"000000000",
  58252=>"111111111",
  58253=>"111111111",
  58254=>"110111111",
  58255=>"000000000",
  58256=>"000000000",
  58257=>"101001001",
  58258=>"000100001",
  58259=>"000000000",
  58260=>"000011111",
  58261=>"000010010",
  58262=>"011011110",
  58263=>"000000000",
  58264=>"110111111",
  58265=>"111111111",
  58266=>"010111001",
  58267=>"111111111",
  58268=>"000000010",
  58269=>"000010011",
  58270=>"011001011",
  58271=>"111100111",
  58272=>"111111010",
  58273=>"111001111",
  58274=>"111101101",
  58275=>"000000000",
  58276=>"111101111",
  58277=>"000000000",
  58278=>"111111111",
  58279=>"000110100",
  58280=>"000000000",
  58281=>"000000000",
  58282=>"111111111",
  58283=>"011001011",
  58284=>"000010000",
  58285=>"000111010",
  58286=>"000000100",
  58287=>"001000000",
  58288=>"000000111",
  58289=>"000101111",
  58290=>"000000111",
  58291=>"111111111",
  58292=>"100000100",
  58293=>"111000000",
  58294=>"111111111",
  58295=>"000000001",
  58296=>"111111001",
  58297=>"000100111",
  58298=>"000000000",
  58299=>"111111111",
  58300=>"000011001",
  58301=>"000000100",
  58302=>"111111000",
  58303=>"101101101",
  58304=>"111111011",
  58305=>"111111111",
  58306=>"111111111",
  58307=>"010000000",
  58308=>"111111111",
  58309=>"001001000",
  58310=>"000000000",
  58311=>"110110110",
  58312=>"000100111",
  58313=>"000000000",
  58314=>"000000000",
  58315=>"000000000",
  58316=>"011011000",
  58317=>"100000000",
  58318=>"100110000",
  58319=>"000111111",
  58320=>"111101000",
  58321=>"101001100",
  58322=>"000100111",
  58323=>"111111110",
  58324=>"111101100",
  58325=>"111111111",
  58326=>"000011111",
  58327=>"000000000",
  58328=>"000010000",
  58329=>"000001110",
  58330=>"000111111",
  58331=>"011001000",
  58332=>"011111111",
  58333=>"111111111",
  58334=>"000000000",
  58335=>"100000000",
  58336=>"001000000",
  58337=>"011011111",
  58338=>"001000000",
  58339=>"010001000",
  58340=>"111111111",
  58341=>"001001000",
  58342=>"111000001",
  58343=>"000000000",
  58344=>"111111111",
  58345=>"111111111",
  58346=>"111111011",
  58347=>"001001000",
  58348=>"111000001",
  58349=>"000000000",
  58350=>"111111111",
  58351=>"110111111",
  58352=>"000000000",
  58353=>"000000000",
  58354=>"111110101",
  58355=>"111011000",
  58356=>"001001001",
  58357=>"011111111",
  58358=>"100100100",
  58359=>"111111001",
  58360=>"100111000",
  58361=>"100101000",
  58362=>"000000000",
  58363=>"001001001",
  58364=>"000000001",
  58365=>"111111111",
  58366=>"111111010",
  58367=>"000000111",
  58368=>"001011111",
  58369=>"000011111",
  58370=>"111000001",
  58371=>"001111000",
  58372=>"000001001",
  58373=>"000000110",
  58374=>"101100000",
  58375=>"100111111",
  58376=>"111010000",
  58377=>"000000000",
  58378=>"000000100",
  58379=>"000000000",
  58380=>"000001001",
  58381=>"101000000",
  58382=>"111111101",
  58383=>"000111111",
  58384=>"000001011",
  58385=>"000110111",
  58386=>"111111001",
  58387=>"000000000",
  58388=>"000000000",
  58389=>"101011111",
  58390=>"000000000",
  58391=>"000001000",
  58392=>"100110000",
  58393=>"111111111",
  58394=>"000011011",
  58395=>"000000000",
  58396=>"001000111",
  58397=>"000000000",
  58398=>"000101111",
  58399=>"111111111",
  58400=>"011011001",
  58401=>"000111001",
  58402=>"000000000",
  58403=>"000000000",
  58404=>"000000000",
  58405=>"001011111",
  58406=>"000000001",
  58407=>"100100000",
  58408=>"100110101",
  58409=>"000000000",
  58410=>"000000000",
  58411=>"111111001",
  58412=>"000000111",
  58413=>"000111000",
  58414=>"000000111",
  58415=>"111110100",
  58416=>"000110000",
  58417=>"000000111",
  58418=>"000000000",
  58419=>"000111000",
  58420=>"000011011",
  58421=>"101111100",
  58422=>"101000101",
  58423=>"000000000",
  58424=>"011011000",
  58425=>"001001011",
  58426=>"000111000",
  58427=>"111111111",
  58428=>"111111111",
  58429=>"100100000",
  58430=>"111000000",
  58431=>"000000000",
  58432=>"100000110",
  58433=>"000000001",
  58434=>"000000000",
  58435=>"000100111",
  58436=>"100111011",
  58437=>"000000000",
  58438=>"111101111",
  58439=>"111111111",
  58440=>"110110000",
  58441=>"111100111",
  58442=>"111111010",
  58443=>"111111111",
  58444=>"011110000",
  58445=>"111011111",
  58446=>"111111110",
  58447=>"000111111",
  58448=>"000000000",
  58449=>"101000100",
  58450=>"000001111",
  58451=>"000100000",
  58452=>"000000000",
  58453=>"001111111",
  58454=>"000000000",
  58455=>"000000000",
  58456=>"111001111",
  58457=>"000000111",
  58458=>"101100000",
  58459=>"111111000",
  58460=>"111101011",
  58461=>"000000000",
  58462=>"000000100",
  58463=>"111100000",
  58464=>"000111111",
  58465=>"000000000",
  58466=>"000000001",
  58467=>"111111111",
  58468=>"111100000",
  58469=>"000001000",
  58470=>"000000000",
  58471=>"111111000",
  58472=>"001000101",
  58473=>"000111111",
  58474=>"111110111",
  58475=>"110111011",
  58476=>"111000000",
  58477=>"000000000",
  58478=>"111111011",
  58479=>"000000100",
  58480=>"111110000",
  58481=>"111000000",
  58482=>"000110111",
  58483=>"000000101",
  58484=>"000000011",
  58485=>"111111111",
  58486=>"000111111",
  58487=>"111101001",
  58488=>"100000111",
  58489=>"111111111",
  58490=>"000000000",
  58491=>"111110111",
  58492=>"100001111",
  58493=>"000110000",
  58494=>"111111111",
  58495=>"111001111",
  58496=>"111111111",
  58497=>"000110111",
  58498=>"111111111",
  58499=>"101110100",
  58500=>"000000000",
  58501=>"011111000",
  58502=>"110000000",
  58503=>"000000001",
  58504=>"100011111",
  58505=>"000000111",
  58506=>"100111100",
  58507=>"000000000",
  58508=>"100110111",
  58509=>"001111111",
  58510=>"111000000",
  58511=>"111111010",
  58512=>"000111111",
  58513=>"000000000",
  58514=>"000000000",
  58515=>"000011111",
  58516=>"000011111",
  58517=>"011011111",
  58518=>"100111001",
  58519=>"000001001",
  58520=>"000000111",
  58521=>"111111100",
  58522=>"000000000",
  58523=>"001001111",
  58524=>"110000001",
  58525=>"001001011",
  58526=>"111111000",
  58527=>"111110000",
  58528=>"000000000",
  58529=>"000111111",
  58530=>"111111111",
  58531=>"111111000",
  58532=>"011001011",
  58533=>"100000100",
  58534=>"000000111",
  58535=>"110100000",
  58536=>"000000111",
  58537=>"111000111",
  58538=>"111111111",
  58539=>"000001001",
  58540=>"000000111",
  58541=>"110111100",
  58542=>"000000011",
  58543=>"000111111",
  58544=>"100100111",
  58545=>"101100101",
  58546=>"010001000",
  58547=>"111111000",
  58548=>"000011110",
  58549=>"011011000",
  58550=>"000001111",
  58551=>"000000111",
  58552=>"000000111",
  58553=>"000100111",
  58554=>"001000100",
  58555=>"111111011",
  58556=>"111000000",
  58557=>"111100000",
  58558=>"000111111",
  58559=>"111111111",
  58560=>"111100100",
  58561=>"001011011",
  58562=>"001111111",
  58563=>"000000000",
  58564=>"000000000",
  58565=>"001011011",
  58566=>"000100000",
  58567=>"011011000",
  58568=>"000000000",
  58569=>"000000000",
  58570=>"000100111",
  58571=>"111010000",
  58572=>"000000000",
  58573=>"001001111",
  58574=>"000110110",
  58575=>"000000000",
  58576=>"111111000",
  58577=>"111000000",
  58578=>"101100111",
  58579=>"000000000",
  58580=>"111000100",
  58581=>"100000000",
  58582=>"101001111",
  58583=>"000000111",
  58584=>"000000111",
  58585=>"000000111",
  58586=>"110000000",
  58587=>"111001000",
  58588=>"111101011",
  58589=>"011000001",
  58590=>"000000000",
  58591=>"010100000",
  58592=>"000000111",
  58593=>"001000000",
  58594=>"100110111",
  58595=>"001011111",
  58596=>"111001000",
  58597=>"000100000",
  58598=>"001010011",
  58599=>"110111111",
  58600=>"111111011",
  58601=>"011000000",
  58602=>"000000000",
  58603=>"110110000",
  58604=>"111011001",
  58605=>"000000110",
  58606=>"000101111",
  58607=>"000001001",
  58608=>"011011010",
  58609=>"111111110",
  58610=>"000000011",
  58611=>"000000000",
  58612=>"111111111",
  58613=>"111111001",
  58614=>"111111000",
  58615=>"000110111",
  58616=>"000000111",
  58617=>"000000001",
  58618=>"000000000",
  58619=>"111001001",
  58620=>"100100000",
  58621=>"001011011",
  58622=>"000000000",
  58623=>"100000011",
  58624=>"101001001",
  58625=>"011001001",
  58626=>"111000111",
  58627=>"000000001",
  58628=>"110111111",
  58629=>"111111110",
  58630=>"000000000",
  58631=>"111001000",
  58632=>"110110111",
  58633=>"000000111",
  58634=>"100111100",
  58635=>"000000000",
  58636=>"100000100",
  58637=>"000000011",
  58638=>"111111000",
  58639=>"111111000",
  58640=>"011010000",
  58641=>"000000000",
  58642=>"100001111",
  58643=>"000000000",
  58644=>"000000100",
  58645=>"000000100",
  58646=>"110110000",
  58647=>"111111011",
  58648=>"011011000",
  58649=>"111011011",
  58650=>"000000000",
  58651=>"111111111",
  58652=>"011000000",
  58653=>"000000010",
  58654=>"100000111",
  58655=>"000000111",
  58656=>"011000100",
  58657=>"000000111",
  58658=>"111111111",
  58659=>"000101101",
  58660=>"011001001",
  58661=>"111111111",
  58662=>"000000101",
  58663=>"001000000",
  58664=>"000010111",
  58665=>"111111011",
  58666=>"000000000",
  58667=>"001001000",
  58668=>"111111000",
  58669=>"000000000",
  58670=>"111001011",
  58671=>"000000111",
  58672=>"000000000",
  58673=>"111111010",
  58674=>"110110110",
  58675=>"111111000",
  58676=>"000000111",
  58677=>"111111000",
  58678=>"000000111",
  58679=>"111101111",
  58680=>"000000000",
  58681=>"000000001",
  58682=>"000000000",
  58683=>"110110111",
  58684=>"000000000",
  58685=>"111111000",
  58686=>"000011111",
  58687=>"100000000",
  58688=>"000000000",
  58689=>"000001000",
  58690=>"000010111",
  58691=>"000000000",
  58692=>"000000000",
  58693=>"010110000",
  58694=>"111111111",
  58695=>"101001000",
  58696=>"000000000",
  58697=>"011101101",
  58698=>"000111111",
  58699=>"110000000",
  58700=>"111101000",
  58701=>"110000001",
  58702=>"000000111",
  58703=>"000110111",
  58704=>"111100000",
  58705=>"100111111",
  58706=>"110011111",
  58707=>"100111110",
  58708=>"110111111",
  58709=>"011011001",
  58710=>"110010000",
  58711=>"111111010",
  58712=>"111111111",
  58713=>"000000000",
  58714=>"010000000",
  58715=>"000111111",
  58716=>"000000000",
  58717=>"111111111",
  58718=>"111111000",
  58719=>"000000000",
  58720=>"011000001",
  58721=>"000000000",
  58722=>"000000000",
  58723=>"001000001",
  58724=>"011000000",
  58725=>"000000011",
  58726=>"000000000",
  58727=>"111111111",
  58728=>"111111011",
  58729=>"111110000",
  58730=>"001011000",
  58731=>"111000100",
  58732=>"000100001",
  58733=>"000000100",
  58734=>"000000111",
  58735=>"000001000",
  58736=>"110000011",
  58737=>"110111111",
  58738=>"111111111",
  58739=>"000111011",
  58740=>"111111101",
  58741=>"111111111",
  58742=>"000001111",
  58743=>"000000000",
  58744=>"111111000",
  58745=>"111111111",
  58746=>"110000110",
  58747=>"111111011",
  58748=>"111011000",
  58749=>"111111111",
  58750=>"111011000",
  58751=>"000000111",
  58752=>"000000111",
  58753=>"001000000",
  58754=>"000001001",
  58755=>"010101000",
  58756=>"111100110",
  58757=>"000111111",
  58758=>"111111111",
  58759=>"000000000",
  58760=>"000000000",
  58761=>"111100111",
  58762=>"000000000",
  58763=>"000000111",
  58764=>"001011111",
  58765=>"100100100",
  58766=>"101100000",
  58767=>"000001111",
  58768=>"011000001",
  58769=>"111110110",
  58770=>"110100000",
  58771=>"000000111",
  58772=>"000000111",
  58773=>"000111111",
  58774=>"000101111",
  58775=>"111111000",
  58776=>"111000000",
  58777=>"000000001",
  58778=>"111000001",
  58779=>"111100111",
  58780=>"110111000",
  58781=>"011111111",
  58782=>"111000111",
  58783=>"011111111",
  58784=>"111111110",
  58785=>"001001100",
  58786=>"011011000",
  58787=>"000000000",
  58788=>"000001111",
  58789=>"000000000",
  58790=>"000101101",
  58791=>"111111111",
  58792=>"000000011",
  58793=>"000000000",
  58794=>"011011111",
  58795=>"111011111",
  58796=>"000000000",
  58797=>"000000111",
  58798=>"000000011",
  58799=>"111111000",
  58800=>"000011111",
  58801=>"010111101",
  58802=>"011011111",
  58803=>"111111111",
  58804=>"001000000",
  58805=>"110111111",
  58806=>"100111000",
  58807=>"000001001",
  58808=>"011001011",
  58809=>"000000000",
  58810=>"000000001",
  58811=>"000000000",
  58812=>"000000001",
  58813=>"111011100",
  58814=>"000000000",
  58815=>"111001000",
  58816=>"111111011",
  58817=>"000100111",
  58818=>"111111111",
  58819=>"110000000",
  58820=>"000000000",
  58821=>"000000000",
  58822=>"111001001",
  58823=>"000000000",
  58824=>"100001101",
  58825=>"000000000",
  58826=>"000000000",
  58827=>"011011000",
  58828=>"010000000",
  58829=>"000100111",
  58830=>"111111111",
  58831=>"010111111",
  58832=>"111110000",
  58833=>"000100101",
  58834=>"101110000",
  58835=>"000001111",
  58836=>"011001001",
  58837=>"111111111",
  58838=>"000000000",
  58839=>"110100100",
  58840=>"000000110",
  58841=>"111000000",
  58842=>"000000111",
  58843=>"000001001",
  58844=>"011111111",
  58845=>"110110000",
  58846=>"000100000",
  58847=>"101100101",
  58848=>"000000000",
  58849=>"111111111",
  58850=>"000000101",
  58851=>"000000000",
  58852=>"010000000",
  58853=>"101111111",
  58854=>"000000000",
  58855=>"000000011",
  58856=>"111011011",
  58857=>"100001011",
  58858=>"000000000",
  58859=>"010111111",
  58860=>"011111111",
  58861=>"011111000",
  58862=>"000000000",
  58863=>"111000000",
  58864=>"111111111",
  58865=>"110111111",
  58866=>"000111111",
  58867=>"000000000",
  58868=>"001001010",
  58869=>"000000000",
  58870=>"000000110",
  58871=>"000111011",
  58872=>"000011000",
  58873=>"000000000",
  58874=>"110101011",
  58875=>"000000000",
  58876=>"111111111",
  58877=>"111011011",
  58878=>"000111111",
  58879=>"010110111",
  58880=>"011000000",
  58881=>"000000010",
  58882=>"111000111",
  58883=>"110110111",
  58884=>"111111111",
  58885=>"000000101",
  58886=>"111111111",
  58887=>"101101101",
  58888=>"111111111",
  58889=>"010111111",
  58890=>"000000000",
  58891=>"110001001",
  58892=>"100111111",
  58893=>"110110111",
  58894=>"100000000",
  58895=>"001111011",
  58896=>"111111111",
  58897=>"011110001",
  58898=>"000011111",
  58899=>"100000100",
  58900=>"011111111",
  58901=>"000000000",
  58902=>"110100001",
  58903=>"000000100",
  58904=>"011001000",
  58905=>"100100111",
  58906=>"101000000",
  58907=>"001000011",
  58908=>"001001011",
  58909=>"111011000",
  58910=>"100111011",
  58911=>"000000001",
  58912=>"000000110",
  58913=>"111101100",
  58914=>"111001000",
  58915=>"000000000",
  58916=>"000000000",
  58917=>"100110010",
  58918=>"000000000",
  58919=>"000000000",
  58920=>"010011111",
  58921=>"000011111",
  58922=>"000000000",
  58923=>"111010010",
  58924=>"000000111",
  58925=>"000000000",
  58926=>"101100110",
  58927=>"100111111",
  58928=>"001111111",
  58929=>"101001001",
  58930=>"001001100",
  58931=>"000000100",
  58932=>"000101011",
  58933=>"110000110",
  58934=>"000000000",
  58935=>"000110000",
  58936=>"101111000",
  58937=>"111001000",
  58938=>"011111011",
  58939=>"000000011",
  58940=>"100000000",
  58941=>"110001111",
  58942=>"000000011",
  58943=>"000000000",
  58944=>"010010011",
  58945=>"000000011",
  58946=>"111111111",
  58947=>"111100000",
  58948=>"110000111",
  58949=>"001101111",
  58950=>"011000000",
  58951=>"111111100",
  58952=>"000000011",
  58953=>"000010010",
  58954=>"111111000",
  58955=>"111111011",
  58956=>"011010111",
  58957=>"001001000",
  58958=>"111111100",
  58959=>"100110111",
  58960=>"000000000",
  58961=>"000000000",
  58962=>"100100110",
  58963=>"111111011",
  58964=>"111111111",
  58965=>"100000000",
  58966=>"111111110",
  58967=>"100111111",
  58968=>"001000000",
  58969=>"110100110",
  58970=>"111111010",
  58971=>"111011001",
  58972=>"001011001",
  58973=>"110000000",
  58974=>"111000000",
  58975=>"111110000",
  58976=>"110001001",
  58977=>"001000001",
  58978=>"111111111",
  58979=>"100111111",
  58980=>"011000001",
  58981=>"011001111",
  58982=>"011000011",
  58983=>"000000100",
  58984=>"000000000",
  58985=>"111101111",
  58986=>"011111111",
  58987=>"000000000",
  58988=>"111111100",
  58989=>"000000000",
  58990=>"111111111",
  58991=>"111111111",
  58992=>"010000110",
  58993=>"110000111",
  58994=>"101001001",
  58995=>"111111111",
  58996=>"000000000",
  58997=>"011001001",
  58998=>"010011111",
  58999=>"111111111",
  59000=>"000000100",
  59001=>"001000000",
  59002=>"111100100",
  59003=>"100110001",
  59004=>"111101111",
  59005=>"000110111",
  59006=>"000111110",
  59007=>"001011000",
  59008=>"111111111",
  59009=>"111111111",
  59010=>"000000111",
  59011=>"001000001",
  59012=>"000000111",
  59013=>"000100000",
  59014=>"000100000",
  59015=>"000000000",
  59016=>"111111011",
  59017=>"000000000",
  59018=>"111111111",
  59019=>"111111111",
  59020=>"100000000",
  59021=>"000000000",
  59022=>"111111011",
  59023=>"000000000",
  59024=>"000000000",
  59025=>"000001011",
  59026=>"011000000",
  59027=>"111111111",
  59028=>"111110000",
  59029=>"011111111",
  59030=>"001000000",
  59031=>"111100000",
  59032=>"000000000",
  59033=>"110111110",
  59034=>"000110111",
  59035=>"001000011",
  59036=>"111001000",
  59037=>"100100110",
  59038=>"110000111",
  59039=>"100010000",
  59040=>"000011110",
  59041=>"010001001",
  59042=>"000001111",
  59043=>"100110111",
  59044=>"110000000",
  59045=>"000000000",
  59046=>"100101000",
  59047=>"000010011",
  59048=>"000000110",
  59049=>"011001001",
  59050=>"001101101",
  59051=>"011010110",
  59052=>"111111110",
  59053=>"101011011",
  59054=>"000000000",
  59055=>"101111111",
  59056=>"111111111",
  59057=>"111001000",
  59058=>"000110000",
  59059=>"111000000",
  59060=>"000000000",
  59061=>"101100110",
  59062=>"000011011",
  59063=>"000000111",
  59064=>"111110110",
  59065=>"000111011",
  59066=>"110000000",
  59067=>"110110110",
  59068=>"000000000",
  59069=>"111111110",
  59070=>"111111111",
  59071=>"111111111",
  59072=>"111101110",
  59073=>"011001000",
  59074=>"000000000",
  59075=>"000000000",
  59076=>"000000000",
  59077=>"000010000",
  59078=>"100110111",
  59079=>"100100110",
  59080=>"000000000",
  59081=>"000100000",
  59082=>"111111111",
  59083=>"000111111",
  59084=>"000111111",
  59085=>"011001011",
  59086=>"000000000",
  59087=>"111010001",
  59088=>"111011111",
  59089=>"001111100",
  59090=>"111001000",
  59091=>"110111111",
  59092=>"111001001",
  59093=>"000000101",
  59094=>"000000001",
  59095=>"111111111",
  59096=>"000000000",
  59097=>"111111000",
  59098=>"100111111",
  59099=>"111111010",
  59100=>"000000001",
  59101=>"111001000",
  59102=>"000001111",
  59103=>"110100000",
  59104=>"000001000",
  59105=>"000000000",
  59106=>"000000001",
  59107=>"101000010",
  59108=>"111110111",
  59109=>"110110110",
  59110=>"000000100",
  59111=>"000000000",
  59112=>"001101111",
  59113=>"111111011",
  59114=>"111111111",
  59115=>"011001101",
  59116=>"101001001",
  59117=>"000000000",
  59118=>"111001101",
  59119=>"111111000",
  59120=>"000110010",
  59121=>"110110111",
  59122=>"111111111",
  59123=>"000000000",
  59124=>"111100000",
  59125=>"100000001",
  59126=>"000000001",
  59127=>"000000000",
  59128=>"000000111",
  59129=>"010000000",
  59130=>"000000000",
  59131=>"000000001",
  59132=>"000010010",
  59133=>"111101101",
  59134=>"000000000",
  59135=>"000000000",
  59136=>"100000111",
  59137=>"000000001",
  59138=>"111111100",
  59139=>"000000100",
  59140=>"101001001",
  59141=>"011111111",
  59142=>"111101001",
  59143=>"111110001",
  59144=>"111110111",
  59145=>"001000000",
  59146=>"000000000",
  59147=>"111011000",
  59148=>"110000000",
  59149=>"111111011",
  59150=>"111110110",
  59151=>"000000000",
  59152=>"010111111",
  59153=>"100111111",
  59154=>"000000000",
  59155=>"111011010",
  59156=>"111111111",
  59157=>"011111111",
  59158=>"000000000",
  59159=>"110110000",
  59160=>"010111111",
  59161=>"111001101",
  59162=>"100110110",
  59163=>"011111011",
  59164=>"001000000",
  59165=>"111000011",
  59166=>"000000000",
  59167=>"001001011",
  59168=>"100000000",
  59169=>"001000000",
  59170=>"111110110",
  59171=>"111111111",
  59172=>"111000010",
  59173=>"111111111",
  59174=>"000000000",
  59175=>"111011011",
  59176=>"011101100",
  59177=>"000000000",
  59178=>"110000000",
  59179=>"000000000",
  59180=>"111111000",
  59181=>"000010000",
  59182=>"111111111",
  59183=>"010010000",
  59184=>"001001001",
  59185=>"000110000",
  59186=>"000001111",
  59187=>"111111111",
  59188=>"010010110",
  59189=>"111100000",
  59190=>"111011000",
  59191=>"000111110",
  59192=>"111010000",
  59193=>"110000000",
  59194=>"111111111",
  59195=>"111111111",
  59196=>"111000000",
  59197=>"100000000",
  59198=>"000011111",
  59199=>"111111010",
  59200=>"101000100",
  59201=>"100110111",
  59202=>"111000110",
  59203=>"011111110",
  59204=>"011111111",
  59205=>"010010000",
  59206=>"100100111",
  59207=>"111111000",
  59208=>"100000000",
  59209=>"111111011",
  59210=>"011011100",
  59211=>"000000001",
  59212=>"100000000",
  59213=>"110000000",
  59214=>"111011011",
  59215=>"000000000",
  59216=>"010011111",
  59217=>"000000101",
  59218=>"111111111",
  59219=>"011000000",
  59220=>"000001000",
  59221=>"001001001",
  59222=>"110000000",
  59223=>"000000000",
  59224=>"111111111",
  59225=>"000000000",
  59226=>"100000000",
  59227=>"000000000",
  59228=>"000011000",
  59229=>"000000101",
  59230=>"011001011",
  59231=>"110111010",
  59232=>"000001000",
  59233=>"111111000",
  59234=>"011010111",
  59235=>"000000000",
  59236=>"100010000",
  59237=>"111101111",
  59238=>"000000100",
  59239=>"100111000",
  59240=>"111011110",
  59241=>"110110111",
  59242=>"111000000",
  59243=>"001000000",
  59244=>"111111111",
  59245=>"011011010",
  59246=>"010000000",
  59247=>"000000001",
  59248=>"000000000",
  59249=>"111111111",
  59250=>"000100110",
  59251=>"111111111",
  59252=>"111000001",
  59253=>"000000000",
  59254=>"111000000",
  59255=>"000000000",
  59256=>"111111111",
  59257=>"001011111",
  59258=>"000011111",
  59259=>"010010011",
  59260=>"111111000",
  59261=>"111111111",
  59262=>"011111110",
  59263=>"111111000",
  59264=>"000010000",
  59265=>"000111111",
  59266=>"110111111",
  59267=>"001001000",
  59268=>"000000011",
  59269=>"000000000",
  59270=>"000010110",
  59271=>"001001001",
  59272=>"011011011",
  59273=>"010010111",
  59274=>"111111111",
  59275=>"110111110",
  59276=>"111111111",
  59277=>"000000001",
  59278=>"110111110",
  59279=>"100111111",
  59280=>"111100111",
  59281=>"110111110",
  59282=>"111000000",
  59283=>"000000110",
  59284=>"000000000",
  59285=>"000110000",
  59286=>"000001101",
  59287=>"111100101",
  59288=>"000111101",
  59289=>"111111011",
  59290=>"111110010",
  59291=>"101111111",
  59292=>"000000111",
  59293=>"111000011",
  59294=>"110100110",
  59295=>"000111111",
  59296=>"000100011",
  59297=>"000001001",
  59298=>"111100010",
  59299=>"110110010",
  59300=>"110000000",
  59301=>"000000000",
  59302=>"000000000",
  59303=>"011000000",
  59304=>"111111001",
  59305=>"111111000",
  59306=>"111111111",
  59307=>"111111110",
  59308=>"000000000",
  59309=>"000100001",
  59310=>"000000100",
  59311=>"111000111",
  59312=>"010000000",
  59313=>"111111111",
  59314=>"000000000",
  59315=>"000000000",
  59316=>"101000000",
  59317=>"000000000",
  59318=>"111111011",
  59319=>"000000111",
  59320=>"000000000",
  59321=>"100111111",
  59322=>"000000100",
  59323=>"000111111",
  59324=>"110111011",
  59325=>"011000000",
  59326=>"000000000",
  59327=>"110110010",
  59328=>"000000000",
  59329=>"111111000",
  59330=>"111111010",
  59331=>"111111011",
  59332=>"110100110",
  59333=>"110010110",
  59334=>"000000000",
  59335=>"000000011",
  59336=>"000000000",
  59337=>"000110111",
  59338=>"101000000",
  59339=>"000000000",
  59340=>"101000000",
  59341=>"000000001",
  59342=>"010000001",
  59343=>"000001101",
  59344=>"111111111",
  59345=>"100100010",
  59346=>"110111111",
  59347=>"000001111",
  59348=>"101100001",
  59349=>"001011011",
  59350=>"111111111",
  59351=>"001111111",
  59352=>"101101001",
  59353=>"111111111",
  59354=>"000000111",
  59355=>"111110100",
  59356=>"000000001",
  59357=>"100000000",
  59358=>"001000000",
  59359=>"111111111",
  59360=>"001001000",
  59361=>"000000110",
  59362=>"111111010",
  59363=>"111111110",
  59364=>"000011111",
  59365=>"000100101",
  59366=>"111111111",
  59367=>"011111000",
  59368=>"100000000",
  59369=>"000000110",
  59370=>"000011111",
  59371=>"110110100",
  59372=>"001000111",
  59373=>"000110011",
  59374=>"100001011",
  59375=>"010000001",
  59376=>"111111010",
  59377=>"001001001",
  59378=>"111001000",
  59379=>"111111111",
  59380=>"111111111",
  59381=>"000000011",
  59382=>"001001001",
  59383=>"001000000",
  59384=>"000000000",
  59385=>"000000000",
  59386=>"011001011",
  59387=>"000000000",
  59388=>"000000000",
  59389=>"000000101",
  59390=>"000000001",
  59391=>"000000000",
  59392=>"001000000",
  59393=>"000000001",
  59394=>"011001111",
  59395=>"000000111",
  59396=>"111111001",
  59397=>"100000001",
  59398=>"000000000",
  59399=>"101000101",
  59400=>"000011111",
  59401=>"111111111",
  59402=>"111111111",
  59403=>"111111111",
  59404=>"000011111",
  59405=>"100111000",
  59406=>"100111011",
  59407=>"111111111",
  59408=>"001110111",
  59409=>"110100000",
  59410=>"000000000",
  59411=>"100000000",
  59412=>"000100000",
  59413=>"011001001",
  59414=>"010000001",
  59415=>"111100000",
  59416=>"111110100",
  59417=>"111100100",
  59418=>"011001000",
  59419=>"000000001",
  59420=>"111010111",
  59421=>"010111111",
  59422=>"111100000",
  59423=>"110010100",
  59424=>"001001000",
  59425=>"001001000",
  59426=>"101111101",
  59427=>"111111011",
  59428=>"000000000",
  59429=>"110111111",
  59430=>"111111000",
  59431=>"111110100",
  59432=>"000100111",
  59433=>"000000000",
  59434=>"000000000",
  59435=>"111111010",
  59436=>"011111101",
  59437=>"111111110",
  59438=>"000001111",
  59439=>"011011011",
  59440=>"000000100",
  59441=>"101001111",
  59442=>"110110100",
  59443=>"111000000",
  59444=>"101111011",
  59445=>"011011101",
  59446=>"000011000",
  59447=>"111111001",
  59448=>"000000001",
  59449=>"111001000",
  59450=>"000000110",
  59451=>"101101101",
  59452=>"111111111",
  59453=>"110000000",
  59454=>"111110100",
  59455=>"000100111",
  59456=>"001111111",
  59457=>"001011010",
  59458=>"000111101",
  59459=>"001000000",
  59460=>"011111001",
  59461=>"000111111",
  59462=>"011011000",
  59463=>"101100111",
  59464=>"101111011",
  59465=>"000000000",
  59466=>"000000000",
  59467=>"000000000",
  59468=>"000001011",
  59469=>"100000100",
  59470=>"111101111",
  59471=>"001011001",
  59472=>"100100000",
  59473=>"000000111",
  59474=>"001000001",
  59475=>"000100111",
  59476=>"111111111",
  59477=>"110010111",
  59478=>"011010000",
  59479=>"000000000",
  59480=>"000000000",
  59481=>"101000000",
  59482=>"010111111",
  59483=>"000001001",
  59484=>"000110111",
  59485=>"010010110",
  59486=>"110110100",
  59487=>"001001011",
  59488=>"000111111",
  59489=>"010011111",
  59490=>"011111000",
  59491=>"110101101",
  59492=>"100000001",
  59493=>"001011011",
  59494=>"011111000",
  59495=>"000000010",
  59496=>"000000000",
  59497=>"000000000",
  59498=>"001111111",
  59499=>"011111100",
  59500=>"011011011",
  59501=>"110010000",
  59502=>"111111111",
  59503=>"000001011",
  59504=>"111111001",
  59505=>"101101111",
  59506=>"100000001",
  59507=>"000000000",
  59508=>"111111111",
  59509=>"001001001",
  59510=>"001000000",
  59511=>"101000000",
  59512=>"000110111",
  59513=>"110110111",
  59514=>"000000000",
  59515=>"000111111",
  59516=>"100110110",
  59517=>"000000000",
  59518=>"000000000",
  59519=>"111111011",
  59520=>"111101111",
  59521=>"001000000",
  59522=>"000000000",
  59523=>"110111111",
  59524=>"000000000",
  59525=>"000000000",
  59526=>"111111110",
  59527=>"000111111",
  59528=>"000000000",
  59529=>"000100111",
  59530=>"111011011",
  59531=>"111010011",
  59532=>"001111011",
  59533=>"001011001",
  59534=>"101000110",
  59535=>"110110000",
  59536=>"000000100",
  59537=>"001000100",
  59538=>"000000001",
  59539=>"001000010",
  59540=>"000110100",
  59541=>"111111111",
  59542=>"111111111",
  59543=>"001001000",
  59544=>"000000000",
  59545=>"000000000",
  59546=>"100101001",
  59547=>"000110100",
  59548=>"111111111",
  59549=>"000000001",
  59550=>"000000111",
  59551=>"000000000",
  59552=>"000000000",
  59553=>"100001001",
  59554=>"111111101",
  59555=>"000000000",
  59556=>"111001011",
  59557=>"110110111",
  59558=>"111000000",
  59559=>"110110111",
  59560=>"011011010",
  59561=>"111000000",
  59562=>"000000000",
  59563=>"111111111",
  59564=>"111111111",
  59565=>"111111111",
  59566=>"000001111",
  59567=>"000000000",
  59568=>"111111011",
  59569=>"100100100",
  59570=>"111011111",
  59571=>"111000000",
  59572=>"001000000",
  59573=>"000000000",
  59574=>"000000000",
  59575=>"000000000",
  59576=>"000100101",
  59577=>"101001000",
  59578=>"111000000",
  59579=>"111000000",
  59580=>"011111111",
  59581=>"000000100",
  59582=>"000011011",
  59583=>"010000000",
  59584=>"101000111",
  59585=>"000000000",
  59586=>"100000000",
  59587=>"111000000",
  59588=>"000000001",
  59589=>"000000111",
  59590=>"101000010",
  59591=>"000000101",
  59592=>"000000100",
  59593=>"111000000",
  59594=>"111111111",
  59595=>"000000000",
  59596=>"111101101",
  59597=>"110000111",
  59598=>"000000000",
  59599=>"111111010",
  59600=>"111111001",
  59601=>"111111000",
  59602=>"111011011",
  59603=>"000000000",
  59604=>"101110111",
  59605=>"111101101",
  59606=>"000000000",
  59607=>"011111111",
  59608=>"001000101",
  59609=>"100111111",
  59610=>"110111101",
  59611=>"111111111",
  59612=>"000000000",
  59613=>"000001001",
  59614=>"111100111",
  59615=>"111111111",
  59616=>"100000000",
  59617=>"010010000",
  59618=>"000000000",
  59619=>"001000000",
  59620=>"000000110",
  59621=>"000000000",
  59622=>"111111111",
  59623=>"111110100",
  59624=>"111111010",
  59625=>"110110111",
  59626=>"000001000",
  59627=>"000000000",
  59628=>"010000111",
  59629=>"000000000",
  59630=>"111110111",
  59631=>"001000000",
  59632=>"011111111",
  59633=>"111100101",
  59634=>"111000001",
  59635=>"001001101",
  59636=>"111111111",
  59637=>"111010000",
  59638=>"000000000",
  59639=>"111001000",
  59640=>"111111111",
  59641=>"011000000",
  59642=>"000000100",
  59643=>"100100001",
  59644=>"000000110",
  59645=>"000000100",
  59646=>"000000111",
  59647=>"000000010",
  59648=>"000111110",
  59649=>"101101100",
  59650=>"111111101",
  59651=>"001000000",
  59652=>"110111111",
  59653=>"111111011",
  59654=>"111111100",
  59655=>"011011011",
  59656=>"110111110",
  59657=>"111111111",
  59658=>"000111111",
  59659=>"111000100",
  59660=>"111111011",
  59661=>"011000111",
  59662=>"111111111",
  59663=>"000101101",
  59664=>"111111111",
  59665=>"000111001",
  59666=>"101111111",
  59667=>"111001011",
  59668=>"000000001",
  59669=>"000110111",
  59670=>"111001100",
  59671=>"111111101",
  59672=>"001000111",
  59673=>"000000111",
  59674=>"000000001",
  59675=>"000000000",
  59676=>"001111111",
  59677=>"000000000",
  59678=>"000000000",
  59679=>"001000000",
  59680=>"111111111",
  59681=>"001101111",
  59682=>"100110010",
  59683=>"111111000",
  59684=>"111011011",
  59685=>"000000001",
  59686=>"000001000",
  59687=>"100100111",
  59688=>"110110000",
  59689=>"111111111",
  59690=>"000101111",
  59691=>"000110000",
  59692=>"100100110",
  59693=>"111111111",
  59694=>"000000000",
  59695=>"111111111",
  59696=>"001001101",
  59697=>"000110111",
  59698=>"000000001",
  59699=>"111000000",
  59700=>"000111110",
  59701=>"000010000",
  59702=>"000000000",
  59703=>"100111001",
  59704=>"000000000",
  59705=>"000000000",
  59706=>"111000000",
  59707=>"000011010",
  59708=>"000000001",
  59709=>"111110100",
  59710=>"011111111",
  59711=>"111110000",
  59712=>"100101000",
  59713=>"001000000",
  59714=>"101111001",
  59715=>"111111111",
  59716=>"111111111",
  59717=>"100000000",
  59718=>"000000100",
  59719=>"111000000",
  59720=>"111111000",
  59721=>"000000000",
  59722=>"000000001",
  59723=>"111011001",
  59724=>"100000100",
  59725=>"000100000",
  59726=>"000111100",
  59727=>"001001001",
  59728=>"111000000",
  59729=>"100110110",
  59730=>"000000000",
  59731=>"000010111",
  59732=>"111111111",
  59733=>"011010010",
  59734=>"110110111",
  59735=>"111111000",
  59736=>"111111111",
  59737=>"111111010",
  59738=>"000100111",
  59739=>"111000000",
  59740=>"000000000",
  59741=>"000001111",
  59742=>"000001001",
  59743=>"110010010",
  59744=>"111111111",
  59745=>"001011111",
  59746=>"101001100",
  59747=>"111111111",
  59748=>"000000000",
  59749=>"000000001",
  59750=>"000000000",
  59751=>"000001101",
  59752=>"101101101",
  59753=>"000000001",
  59754=>"111111100",
  59755=>"110111001",
  59756=>"000000000",
  59757=>"100000101",
  59758=>"000111000",
  59759=>"111111111",
  59760=>"000000000",
  59761=>"111111111",
  59762=>"101000000",
  59763=>"101111111",
  59764=>"000000000",
  59765=>"000000000",
  59766=>"000000001",
  59767=>"000000000",
  59768=>"000111011",
  59769=>"110111111",
  59770=>"111111011",
  59771=>"001000100",
  59772=>"011001011",
  59773=>"111111111",
  59774=>"011011011",
  59775=>"111100000",
  59776=>"100111110",
  59777=>"000000000",
  59778=>"000011111",
  59779=>"111000000",
  59780=>"000000000",
  59781=>"111010000",
  59782=>"000111111",
  59783=>"001011011",
  59784=>"001001000",
  59785=>"111110000",
  59786=>"000000100",
  59787=>"101000100",
  59788=>"100000111",
  59789=>"111001101",
  59790=>"000000100",
  59791=>"001000000",
  59792=>"000000000",
  59793=>"001111001",
  59794=>"000000000",
  59795=>"111111111",
  59796=>"111111111",
  59797=>"000000010",
  59798=>"011011000",
  59799=>"100110110",
  59800=>"001000000",
  59801=>"010010000",
  59802=>"110111111",
  59803=>"101101111",
  59804=>"001111111",
  59805=>"000000101",
  59806=>"111111111",
  59807=>"011000000",
  59808=>"000000000",
  59809=>"110110110",
  59810=>"101111111",
  59811=>"000000111",
  59812=>"101010000",
  59813=>"000110111",
  59814=>"111100000",
  59815=>"010000000",
  59816=>"000001001",
  59817=>"000000000",
  59818=>"001011000",
  59819=>"111111111",
  59820=>"000000000",
  59821=>"000110100",
  59822=>"000000101",
  59823=>"001000011",
  59824=>"111011000",
  59825=>"101111111",
  59826=>"000000000",
  59827=>"000111011",
  59828=>"001000000",
  59829=>"111000000",
  59830=>"000100111",
  59831=>"001000000",
  59832=>"111111111",
  59833=>"111111111",
  59834=>"011111000",
  59835=>"000111111",
  59836=>"001100100",
  59837=>"000000010",
  59838=>"000000000",
  59839=>"100101101",
  59840=>"110100111",
  59841=>"011001011",
  59842=>"000000000",
  59843=>"111111001",
  59844=>"001001001",
  59845=>"111000000",
  59846=>"000000000",
  59847=>"000111101",
  59848=>"101000000",
  59849=>"000000110",
  59850=>"001100110",
  59851=>"000000011",
  59852=>"111111111",
  59853=>"011011000",
  59854=>"101100000",
  59855=>"010110000",
  59856=>"111100101",
  59857=>"111111111",
  59858=>"111010000",
  59859=>"011001101",
  59860=>"000000001",
  59861=>"000000000",
  59862=>"000100100",
  59863=>"000000000",
  59864=>"111101000",
  59865=>"000100110",
  59866=>"111011000",
  59867=>"111111111",
  59868=>"110100001",
  59869=>"001001111",
  59870=>"000000000",
  59871=>"110100000",
  59872=>"000111111",
  59873=>"111111011",
  59874=>"000000011",
  59875=>"000000000",
  59876=>"001111111",
  59877=>"101111111",
  59878=>"000000000",
  59879=>"111011000",
  59880=>"101001001",
  59881=>"000000000",
  59882=>"111100111",
  59883=>"101001000",
  59884=>"111001001",
  59885=>"111111011",
  59886=>"000000110",
  59887=>"111001000",
  59888=>"001001111",
  59889=>"111101101",
  59890=>"111000000",
  59891=>"011111001",
  59892=>"000001001",
  59893=>"011011111",
  59894=>"110000000",
  59895=>"011111011",
  59896=>"000000000",
  59897=>"011001011",
  59898=>"000000000",
  59899=>"111111001",
  59900=>"001011111",
  59901=>"000001111",
  59902=>"100000000",
  59903=>"111000000",
  59904=>"110111011",
  59905=>"111110100",
  59906=>"111011011",
  59907=>"110000000",
  59908=>"011000100",
  59909=>"111000000",
  59910=>"111111000",
  59911=>"111111111",
  59912=>"111000111",
  59913=>"000101111",
  59914=>"111111111",
  59915=>"111101111",
  59916=>"001111111",
  59917=>"010111001",
  59918=>"110010010",
  59919=>"000110111",
  59920=>"110111111",
  59921=>"111000101",
  59922=>"000000110",
  59923=>"110111111",
  59924=>"000111111",
  59925=>"110111111",
  59926=>"111111110",
  59927=>"000111011",
  59928=>"100100100",
  59929=>"110000000",
  59930=>"100000000",
  59931=>"000000000",
  59932=>"111111111",
  59933=>"111000001",
  59934=>"001000111",
  59935=>"011001111",
  59936=>"100000111",
  59937=>"000000111",
  59938=>"001100100",
  59939=>"000000000",
  59940=>"000001000",
  59941=>"001111111",
  59942=>"110000000",
  59943=>"000110000",
  59944=>"110000000",
  59945=>"000000000",
  59946=>"111111000",
  59947=>"001000000",
  59948=>"111111110",
  59949=>"110010000",
  59950=>"011000000",
  59951=>"000000111",
  59952=>"111000010",
  59953=>"010000001",
  59954=>"111111011",
  59955=>"001001111",
  59956=>"000000111",
  59957=>"011001011",
  59958=>"000011011",
  59959=>"011011111",
  59960=>"110111111",
  59961=>"001010000",
  59962=>"000000001",
  59963=>"100110011",
  59964=>"001000000",
  59965=>"000000010",
  59966=>"111111000",
  59967=>"000000000",
  59968=>"100000010",
  59969=>"100000001",
  59970=>"011011011",
  59971=>"111111010",
  59972=>"000111000",
  59973=>"001101100",
  59974=>"000000110",
  59975=>"111000000",
  59976=>"000010000",
  59977=>"100000000",
  59978=>"110110000",
  59979=>"000000000",
  59980=>"001101111",
  59981=>"101000000",
  59982=>"000000111",
  59983=>"111111111",
  59984=>"000000111",
  59985=>"111111011",
  59986=>"000100111",
  59987=>"000000010",
  59988=>"111111111",
  59989=>"000000110",
  59990=>"001111111",
  59991=>"000000100",
  59992=>"000010111",
  59993=>"000000000",
  59994=>"111111000",
  59995=>"001111111",
  59996=>"110010000",
  59997=>"111111111",
  59998=>"001011001",
  59999=>"100101110",
  60000=>"110000100",
  60001=>"101111111",
  60002=>"111101000",
  60003=>"111011000",
  60004=>"000000110",
  60005=>"111001000",
  60006=>"100001001",
  60007=>"000111111",
  60008=>"111110111",
  60009=>"000011001",
  60010=>"000111111",
  60011=>"111001000",
  60012=>"100110011",
  60013=>"000000100",
  60014=>"111000000",
  60015=>"001000110",
  60016=>"111111001",
  60017=>"000000000",
  60018=>"001001011",
  60019=>"101011000",
  60020=>"001100000",
  60021=>"000000000",
  60022=>"000000000",
  60023=>"000000111",
  60024=>"111000100",
  60025=>"001101001",
  60026=>"000111111",
  60027=>"000000011",
  60028=>"000000111",
  60029=>"000010100",
  60030=>"000000000",
  60031=>"000000000",
  60032=>"000000001",
  60033=>"001011000",
  60034=>"000000000",
  60035=>"001011011",
  60036=>"000000011",
  60037=>"110000000",
  60038=>"111011111",
  60039=>"111011111",
  60040=>"000000000",
  60041=>"101011010",
  60042=>"000000000",
  60043=>"010011111",
  60044=>"111111011",
  60045=>"000000011",
  60046=>"011011001",
  60047=>"000011000",
  60048=>"000111111",
  60049=>"111010011",
  60050=>"111111110",
  60051=>"000000001",
  60052=>"101100110",
  60053=>"000000000",
  60054=>"000000101",
  60055=>"000000111",
  60056=>"111111111",
  60057=>"000000000",
  60058=>"111111111",
  60059=>"000000000",
  60060=>"111001000",
  60061=>"111111000",
  60062=>"111111111",
  60063=>"111111111",
  60064=>"000000110",
  60065=>"000000000",
  60066=>"011111000",
  60067=>"001111000",
  60068=>"001000111",
  60069=>"001001101",
  60070=>"111111111",
  60071=>"000100111",
  60072=>"000111111",
  60073=>"100110111",
  60074=>"111000100",
  60075=>"000000111",
  60076=>"111111111",
  60077=>"011011111",
  60078=>"111111100",
  60079=>"000010000",
  60080=>"011111010",
  60081=>"011000010",
  60082=>"110111010",
  60083=>"100111111",
  60084=>"100000000",
  60085=>"100110111",
  60086=>"000000111",
  60087=>"000000000",
  60088=>"000000000",
  60089=>"000000000",
  60090=>"111100111",
  60091=>"111111111",
  60092=>"000110111",
  60093=>"000000111",
  60094=>"000111111",
  60095=>"000000000",
  60096=>"000000000",
  60097=>"000111111",
  60098=>"111110110",
  60099=>"111110111",
  60100=>"100111111",
  60101=>"111000000",
  60102=>"000111111",
  60103=>"000111011",
  60104=>"111111111",
  60105=>"000000000",
  60106=>"000000111",
  60107=>"111001000",
  60108=>"001011110",
  60109=>"000110110",
  60110=>"010011111",
  60111=>"000000000",
  60112=>"011010000",
  60113=>"110110111",
  60114=>"111111000",
  60115=>"000000000",
  60116=>"111100000",
  60117=>"111111111",
  60118=>"110010000",
  60119=>"110111000",
  60120=>"000010111",
  60121=>"011011111",
  60122=>"000110101",
  60123=>"001110100",
  60124=>"000000111",
  60125=>"000110000",
  60126=>"111011000",
  60127=>"000000111",
  60128=>"110110111",
  60129=>"100111111",
  60130=>"000000000",
  60131=>"000001111",
  60132=>"000000111",
  60133=>"010111011",
  60134=>"001000000",
  60135=>"111000000",
  60136=>"000000000",
  60137=>"110110101",
  60138=>"000001000",
  60139=>"001000100",
  60140=>"111111001",
  60141=>"010111000",
  60142=>"111111111",
  60143=>"111000000",
  60144=>"000001111",
  60145=>"000111111",
  60146=>"111001111",
  60147=>"111010010",
  60148=>"000000000",
  60149=>"000111111",
  60150=>"110010000",
  60151=>"110010010",
  60152=>"111000110",
  60153=>"000000000",
  60154=>"100110111",
  60155=>"110000111",
  60156=>"001011011",
  60157=>"100100000",
  60158=>"111111100",
  60159=>"000111110",
  60160=>"100101100",
  60161=>"001000110",
  60162=>"111101111",
  60163=>"101000110",
  60164=>"000000011",
  60165=>"111001001",
  60166=>"000100101",
  60167=>"010110000",
  60168=>"000000000",
  60169=>"000111000",
  60170=>"111111111",
  60171=>"011010010",
  60172=>"001000111",
  60173=>"000001111",
  60174=>"000010111",
  60175=>"110000000",
  60176=>"111111001",
  60177=>"110010011",
  60178=>"010000111",
  60179=>"111000100",
  60180=>"001000000",
  60181=>"110000111",
  60182=>"100000000",
  60183=>"000011000",
  60184=>"000001111",
  60185=>"001000111",
  60186=>"000000010",
  60187=>"000000000",
  60188=>"111111110",
  60189=>"001000111",
  60190=>"111111111",
  60191=>"111110000",
  60192=>"011011001",
  60193=>"000111000",
  60194=>"000001001",
  60195=>"110011000",
  60196=>"000000111",
  60197=>"001000000",
  60198=>"110000000",
  60199=>"110111001",
  60200=>"001000111",
  60201=>"110111111",
  60202=>"011010110",
  60203=>"111010000",
  60204=>"000000000",
  60205=>"110100100",
  60206=>"000000011",
  60207=>"000000010",
  60208=>"111111111",
  60209=>"000010000",
  60210=>"000000110",
  60211=>"111000111",
  60212=>"000110100",
  60213=>"011011010",
  60214=>"000000001",
  60215=>"110110000",
  60216=>"000111000",
  60217=>"000000111",
  60218=>"111111110",
  60219=>"111100000",
  60220=>"100110110",
  60221=>"111111100",
  60222=>"101001111",
  60223=>"000000101",
  60224=>"111100000",
  60225=>"111000100",
  60226=>"111111111",
  60227=>"000000111",
  60228=>"000000000",
  60229=>"111111111",
  60230=>"000000100",
  60231=>"001001000",
  60232=>"000000111",
  60233=>"111000110",
  60234=>"110111010",
  60235=>"100011001",
  60236=>"000000000",
  60237=>"111000000",
  60238=>"000100000",
  60239=>"000000001",
  60240=>"000011011",
  60241=>"000000000",
  60242=>"110101111",
  60243=>"000000000",
  60244=>"000000011",
  60245=>"011000000",
  60246=>"111111111",
  60247=>"011011010",
  60248=>"000111111",
  60249=>"100000111",
  60250=>"000000000",
  60251=>"100000000",
  60252=>"000110110",
  60253=>"000001101",
  60254=>"010000111",
  60255=>"101001011",
  60256=>"111111100",
  60257=>"000100000",
  60258=>"001101111",
  60259=>"111111000",
  60260=>"101001000",
  60261=>"000000000",
  60262=>"110110111",
  60263=>"000000000",
  60264=>"000100000",
  60265=>"111111000",
  60266=>"001000000",
  60267=>"110110000",
  60268=>"001100000",
  60269=>"000000000",
  60270=>"101000001",
  60271=>"001111111",
  60272=>"000101001",
  60273=>"111111111",
  60274=>"000100111",
  60275=>"000100100",
  60276=>"111101100",
  60277=>"101111000",
  60278=>"111111001",
  60279=>"011111001",
  60280=>"111111111",
  60281=>"110110111",
  60282=>"000111111",
  60283=>"111001111",
  60284=>"000000111",
  60285=>"000110111",
  60286=>"000111111",
  60287=>"111000000",
  60288=>"111111110",
  60289=>"001001111",
  60290=>"111111011",
  60291=>"000110110",
  60292=>"000010110",
  60293=>"000000111",
  60294=>"110111111",
  60295=>"000000111",
  60296=>"000001111",
  60297=>"111111000",
  60298=>"001000000",
  60299=>"111111000",
  60300=>"001011111",
  60301=>"000000000",
  60302=>"000001011",
  60303=>"111111111",
  60304=>"000000111",
  60305=>"001000000",
  60306=>"010110001",
  60307=>"111001001",
  60308=>"000110111",
  60309=>"000000000",
  60310=>"110111001",
  60311=>"111111111",
  60312=>"111011001",
  60313=>"111001101",
  60314=>"111111111",
  60315=>"000000000",
  60316=>"001000000",
  60317=>"100100000",
  60318=>"111000000",
  60319=>"000000111",
  60320=>"000001000",
  60321=>"001001111",
  60322=>"000000000",
  60323=>"011000000",
  60324=>"111110000",
  60325=>"100000000",
  60326=>"000101001",
  60327=>"111000000",
  60328=>"111110110",
  60329=>"111111000",
  60330=>"111100101",
  60331=>"000000000",
  60332=>"000000001",
  60333=>"101101000",
  60334=>"111111110",
  60335=>"000000110",
  60336=>"111110110",
  60337=>"000010110",
  60338=>"011001111",
  60339=>"000010010",
  60340=>"111001111",
  60341=>"100111110",
  60342=>"110111011",
  60343=>"110111110",
  60344=>"000000000",
  60345=>"111011011",
  60346=>"000000110",
  60347=>"000000111",
  60348=>"111111111",
  60349=>"111111100",
  60350=>"000111111",
  60351=>"100100000",
  60352=>"000000111",
  60353=>"001001000",
  60354=>"000011000",
  60355=>"000000111",
  60356=>"111111111",
  60357=>"011111111",
  60358=>"111111010",
  60359=>"000000011",
  60360=>"101111001",
  60361=>"000000001",
  60362=>"000000100",
  60363=>"000000001",
  60364=>"000000000",
  60365=>"001001001",
  60366=>"001111010",
  60367=>"000111111",
  60368=>"000000111",
  60369=>"111111010",
  60370=>"000111111",
  60371=>"000001001",
  60372=>"001011000",
  60373=>"111111111",
  60374=>"111000000",
  60375=>"101000000",
  60376=>"001000000",
  60377=>"000000101",
  60378=>"111111000",
  60379=>"100000000",
  60380=>"111111111",
  60381=>"110110011",
  60382=>"000000001",
  60383=>"111110000",
  60384=>"110110110",
  60385=>"000001111",
  60386=>"111111111",
  60387=>"111111111",
  60388=>"111000000",
  60389=>"100100000",
  60390=>"111000000",
  60391=>"000011111",
  60392=>"010111111",
  60393=>"111111011",
  60394=>"100000000",
  60395=>"111111000",
  60396=>"111111111",
  60397=>"100110111",
  60398=>"100000001",
  60399=>"111100100",
  60400=>"000000110",
  60401=>"111111110",
  60402=>"111011111",
  60403=>"011001000",
  60404=>"000100111",
  60405=>"000000000",
  60406=>"111001000",
  60407=>"001000000",
  60408=>"111000000",
  60409=>"011010000",
  60410=>"000000000",
  60411=>"110110000",
  60412=>"000000001",
  60413=>"111001001",
  60414=>"000000000",
  60415=>"000000000",
  60416=>"000001000",
  60417=>"110000000",
  60418=>"000000111",
  60419=>"000110010",
  60420=>"111111001",
  60421=>"100000000",
  60422=>"100110111",
  60423=>"011111111",
  60424=>"101110100",
  60425=>"111100100",
  60426=>"000000001",
  60427=>"101011001",
  60428=>"110000100",
  60429=>"011111111",
  60430=>"011011111",
  60431=>"000010000",
  60432=>"110111111",
  60433=>"111111001",
  60434=>"111111111",
  60435=>"111111111",
  60436=>"000000000",
  60437=>"110011110",
  60438=>"000001111",
  60439=>"100100001",
  60440=>"101111111",
  60441=>"111111101",
  60442=>"011001001",
  60443=>"111010000",
  60444=>"000011001",
  60445=>"000000000",
  60446=>"111101111",
  60447=>"111111111",
  60448=>"000000000",
  60449=>"001001111",
  60450=>"011011001",
  60451=>"000000000",
  60452=>"111111001",
  60453=>"111111000",
  60454=>"000010111",
  60455=>"000000111",
  60456=>"110011111",
  60457=>"111010000",
  60458=>"111110100",
  60459=>"110100000",
  60460=>"000110100",
  60461=>"111110011",
  60462=>"000000000",
  60463=>"000000000",
  60464=>"001000101",
  60465=>"000000000",
  60466=>"000000000",
  60467=>"000000000",
  60468=>"000000000",
  60469=>"010000000",
  60470=>"111111111",
  60471=>"111111111",
  60472=>"111111110",
  60473=>"000110100",
  60474=>"000000111",
  60475=>"000000111",
  60476=>"000000000",
  60477=>"011011011",
  60478=>"100000000",
  60479=>"000000000",
  60480=>"001111110",
  60481=>"110011000",
  60482=>"110111111",
  60483=>"101101001",
  60484=>"001100000",
  60485=>"101001111",
  60486=>"011011000",
  60487=>"000000000",
  60488=>"000000010",
  60489=>"000000000",
  60490=>"010111101",
  60491=>"111111111",
  60492=>"101000111",
  60493=>"011111111",
  60494=>"110000111",
  60495=>"101000000",
  60496=>"111111111",
  60497=>"111111011",
  60498=>"111000010",
  60499=>"000000100",
  60500=>"001001000",
  60501=>"001110100",
  60502=>"000110100",
  60503=>"000000000",
  60504=>"000101100",
  60505=>"000100110",
  60506=>"001000010",
  60507=>"000110110",
  60508=>"000000000",
  60509=>"111111110",
  60510=>"000100100",
  60511=>"110110110",
  60512=>"110100000",
  60513=>"101101111",
  60514=>"000000000",
  60515=>"000000000",
  60516=>"111110111",
  60517=>"001101101",
  60518=>"010110100",
  60519=>"111101101",
  60520=>"000100000",
  60521=>"000110111",
  60522=>"110111111",
  60523=>"000000011",
  60524=>"000001000",
  60525=>"100111111",
  60526=>"111111011",
  60527=>"000000000",
  60528=>"100000000",
  60529=>"000011000",
  60530=>"000000000",
  60531=>"110101100",
  60532=>"000001001",
  60533=>"000000000",
  60534=>"001001001",
  60535=>"000000000",
  60536=>"000000000",
  60537=>"000000000",
  60538=>"000000000",
  60539=>"111111111",
  60540=>"011011111",
  60541=>"000010000",
  60542=>"000111100",
  60543=>"000001111",
  60544=>"000001111",
  60545=>"000000000",
  60546=>"001000001",
  60547=>"000000110",
  60548=>"111111111",
  60549=>"000000110",
  60550=>"000000000",
  60551=>"111111111",
  60552=>"000000000",
  60553=>"011000000",
  60554=>"000000111",
  60555=>"011111111",
  60556=>"111111101",
  60557=>"011000000",
  60558=>"111111010",
  60559=>"000000000",
  60560=>"000100000",
  60561=>"000000000",
  60562=>"011011111",
  60563=>"001100100",
  60564=>"000110110",
  60565=>"110111011",
  60566=>"000000000",
  60567=>"111000111",
  60568=>"000000100",
  60569=>"111111111",
  60570=>"111111111",
  60571=>"111111111",
  60572=>"100100100",
  60573=>"111011111",
  60574=>"000111111",
  60575=>"100111010",
  60576=>"000110100",
  60577=>"111111101",
  60578=>"111111111",
  60579=>"111111111",
  60580=>"011110100",
  60581=>"100000101",
  60582=>"010111110",
  60583=>"101100100",
  60584=>"110111100",
  60585=>"111111111",
  60586=>"111111100",
  60587=>"000110110",
  60588=>"111000000",
  60589=>"110110110",
  60590=>"001100110",
  60591=>"000000000",
  60592=>"000110111",
  60593=>"110010010",
  60594=>"000011011",
  60595=>"000111011",
  60596=>"010100000",
  60597=>"111100100",
  60598=>"000110100",
  60599=>"101111110",
  60600=>"001001111",
  60601=>"001000000",
  60602=>"100111110",
  60603=>"001101101",
  60604=>"111101111",
  60605=>"010111111",
  60606=>"000110000",
  60607=>"001111111",
  60608=>"000000001",
  60609=>"111111111",
  60610=>"110111111",
  60611=>"110111111",
  60612=>"011000001",
  60613=>"000000100",
  60614=>"010111110",
  60615=>"100101000",
  60616=>"111111111",
  60617=>"000000000",
  60618=>"000000000",
  60619=>"001000000",
  60620=>"000000000",
  60621=>"111111000",
  60622=>"111100111",
  60623=>"000110100",
  60624=>"110100001",
  60625=>"111111111",
  60626=>"111000001",
  60627=>"100110110",
  60628=>"111011001",
  60629=>"111001111",
  60630=>"111000000",
  60631=>"000000000",
  60632=>"000000101",
  60633=>"110110100",
  60634=>"000000000",
  60635=>"011011111",
  60636=>"111111111",
  60637=>"000100101",
  60638=>"111111111",
  60639=>"000100100",
  60640=>"111101101",
  60641=>"111111010",
  60642=>"110000000",
  60643=>"011111110",
  60644=>"100100100",
  60645=>"100110111",
  60646=>"000000000",
  60647=>"111111111",
  60648=>"111111110",
  60649=>"001011111",
  60650=>"100100111",
  60651=>"000000000",
  60652=>"000000000",
  60653=>"000000100",
  60654=>"111000000",
  60655=>"111000000",
  60656=>"000111111",
  60657=>"000000001",
  60658=>"011011111",
  60659=>"011010000",
  60660=>"001011000",
  60661=>"111111011",
  60662=>"111101000",
  60663=>"001000000",
  60664=>"111000000",
  60665=>"000000101",
  60666=>"010110110",
  60667=>"100000000",
  60668=>"000000000",
  60669=>"000000000",
  60670=>"001111111",
  60671=>"000000110",
  60672=>"111110110",
  60673=>"110110000",
  60674=>"001000100",
  60675=>"000000000",
  60676=>"000111111",
  60677=>"011111111",
  60678=>"111111111",
  60679=>"001000000",
  60680=>"000000110",
  60681=>"111111110",
  60682=>"101000011",
  60683=>"110000110",
  60684=>"000000000",
  60685=>"000000000",
  60686=>"111111111",
  60687=>"111111000",
  60688=>"010000001",
  60689=>"111111111",
  60690=>"000011111",
  60691=>"111011011",
  60692=>"000111100",
  60693=>"110100100",
  60694=>"000000100",
  60695=>"110100110",
  60696=>"111111111",
  60697=>"000000100",
  60698=>"000000001",
  60699=>"111111110",
  60700=>"001100000",
  60701=>"111111111",
  60702=>"110111111",
  60703=>"000000111",
  60704=>"111111111",
  60705=>"111011001",
  60706=>"011111100",
  60707=>"010110110",
  60708=>"111111011",
  60709=>"000000000",
  60710=>"001000011",
  60711=>"111111111",
  60712=>"111001001",
  60713=>"000000000",
  60714=>"000010110",
  60715=>"000000000",
  60716=>"110111111",
  60717=>"111111111",
  60718=>"110111111",
  60719=>"000100111",
  60720=>"000001001",
  60721=>"001000000",
  60722=>"111100100",
  60723=>"000000000",
  60724=>"110000000",
  60725=>"000001000",
  60726=>"011000000",
  60727=>"001111111",
  60728=>"111111111",
  60729=>"000000110",
  60730=>"000000000",
  60731=>"110110000",
  60732=>"111111111",
  60733=>"000100110",
  60734=>"000100100",
  60735=>"000100110",
  60736=>"111001000",
  60737=>"011111111",
  60738=>"001011011",
  60739=>"000000000",
  60740=>"110100110",
  60741=>"000000100",
  60742=>"111111101",
  60743=>"000001111",
  60744=>"000000000",
  60745=>"010010000",
  60746=>"100110110",
  60747=>"000000000",
  60748=>"000000111",
  60749=>"111110110",
  60750=>"010110111",
  60751=>"000000101",
  60752=>"001111111",
  60753=>"111111100",
  60754=>"111111111",
  60755=>"000000000",
  60756=>"000110110",
  60757=>"111111111",
  60758=>"001100100",
  60759=>"001000111",
  60760=>"111111111",
  60761=>"000000000",
  60762=>"111001001",
  60763=>"000011111",
  60764=>"011010000",
  60765=>"000000000",
  60766=>"000000000",
  60767=>"111111111",
  60768=>"000000000",
  60769=>"111111111",
  60770=>"001111111",
  60771=>"000000000",
  60772=>"010110100",
  60773=>"001001101",
  60774=>"000001111",
  60775=>"110010000",
  60776=>"101101101",
  60777=>"011110111",
  60778=>"100111000",
  60779=>"000100000",
  60780=>"111110111",
  60781=>"111111110",
  60782=>"111110110",
  60783=>"111111111",
  60784=>"001001111",
  60785=>"111111000",
  60786=>"000101101",
  60787=>"111011011",
  60788=>"111111011",
  60789=>"000000111",
  60790=>"011111100",
  60791=>"000000100",
  60792=>"111100100",
  60793=>"011001000",
  60794=>"000000001",
  60795=>"011000000",
  60796=>"000000111",
  60797=>"100100100",
  60798=>"011000000",
  60799=>"111111101",
  60800=>"000000000",
  60801=>"110110111",
  60802=>"000000000",
  60803=>"000000000",
  60804=>"100111100",
  60805=>"110100000",
  60806=>"111111111",
  60807=>"111111100",
  60808=>"111111101",
  60809=>"101001001",
  60810=>"101101111",
  60811=>"000000111",
  60812=>"111010010",
  60813=>"000000000",
  60814=>"000000111",
  60815=>"111010000",
  60816=>"111111011",
  60817=>"110100110",
  60818=>"111111111",
  60819=>"000110111",
  60820=>"111111111",
  60821=>"000000000",
  60822=>"011111011",
  60823=>"000000110",
  60824=>"111100100",
  60825=>"111001000",
  60826=>"000000000",
  60827=>"000000000",
  60828=>"000000011",
  60829=>"100100000",
  60830=>"000000000",
  60831=>"000000000",
  60832=>"101111100",
  60833=>"000100100",
  60834=>"000111111",
  60835=>"010000000",
  60836=>"000000010",
  60837=>"111110100",
  60838=>"110111111",
  60839=>"111111101",
  60840=>"000000000",
  60841=>"110010000",
  60842=>"111111100",
  60843=>"111110100",
  60844=>"000000000",
  60845=>"111000100",
  60846=>"111011010",
  60847=>"100000000",
  60848=>"011111111",
  60849=>"001001000",
  60850=>"001011111",
  60851=>"011111111",
  60852=>"000111111",
  60853=>"000000001",
  60854=>"000000000",
  60855=>"110000000",
  60856=>"111111000",
  60857=>"000000011",
  60858=>"111111111",
  60859=>"001000000",
  60860=>"110000111",
  60861=>"110110000",
  60862=>"000000000",
  60863=>"010100100",
  60864=>"000000111",
  60865=>"111100000",
  60866=>"110000111",
  60867=>"000111001",
  60868=>"110110110",
  60869=>"001000000",
  60870=>"001000000",
  60871=>"000100000",
  60872=>"101000110",
  60873=>"000110110",
  60874=>"000000000",
  60875=>"000000000",
  60876=>"000000111",
  60877=>"000000100",
  60878=>"000000000",
  60879=>"011011111",
  60880=>"011111111",
  60881=>"111111111",
  60882=>"111111111",
  60883=>"000011000",
  60884=>"000011011",
  60885=>"110010010",
  60886=>"100000000",
  60887=>"000011011",
  60888=>"000110001",
  60889=>"111111010",
  60890=>"010010000",
  60891=>"100110100",
  60892=>"011111011",
  60893=>"000000000",
  60894=>"111111111",
  60895=>"000000000",
  60896=>"000100000",
  60897=>"000000000",
  60898=>"111111111",
  60899=>"000000000",
  60900=>"011111011",
  60901=>"000000000",
  60902=>"000000111",
  60903=>"000000000",
  60904=>"110111010",
  60905=>"001111111",
  60906=>"011111110",
  60907=>"111000100",
  60908=>"000000000",
  60909=>"111111011",
  60910=>"111111111",
  60911=>"000100100",
  60912=>"000000000",
  60913=>"111111101",
  60914=>"101100101",
  60915=>"000000000",
  60916=>"110110111",
  60917=>"000000011",
  60918=>"001001011",
  60919=>"000001001",
  60920=>"110000000",
  60921=>"000000000",
  60922=>"000000000",
  60923=>"111111111",
  60924=>"000000100",
  60925=>"111001000",
  60926=>"000000001",
  60927=>"000000000",
  60928=>"100001111",
  60929=>"111001001",
  60930=>"111010111",
  60931=>"000000001",
  60932=>"111000000",
  60933=>"011000000",
  60934=>"000000000",
  60935=>"000000000",
  60936=>"100001000",
  60937=>"111111000",
  60938=>"111111111",
  60939=>"000111111",
  60940=>"110100000",
  60941=>"011001001",
  60942=>"000000111",
  60943=>"110110010",
  60944=>"000000110",
  60945=>"000011011",
  60946=>"011011111",
  60947=>"010000001",
  60948=>"000000111",
  60949=>"000000000",
  60950=>"000000000",
  60951=>"011011011",
  60952=>"000000000",
  60953=>"100100100",
  60954=>"111111111",
  60955=>"001000000",
  60956=>"000000000",
  60957=>"110100000",
  60958=>"000001001",
  60959=>"110010000",
  60960=>"000000110",
  60961=>"111101111",
  60962=>"000110111",
  60963=>"000111111",
  60964=>"000000000",
  60965=>"111010000",
  60966=>"111000111",
  60967=>"000000000",
  60968=>"000011100",
  60969=>"000111101",
  60970=>"000001000",
  60971=>"000000111",
  60972=>"000111111",
  60973=>"000001000",
  60974=>"110110000",
  60975=>"011011111",
  60976=>"001011001",
  60977=>"000111111",
  60978=>"111111000",
  60979=>"000100111",
  60980=>"111110000",
  60981=>"110110000",
  60982=>"111000000",
  60983=>"000111011",
  60984=>"000000111",
  60985=>"100100111",
  60986=>"000000000",
  60987=>"110110000",
  60988=>"111111000",
  60989=>"011111110",
  60990=>"000110000",
  60991=>"111101001",
  60992=>"000110111",
  60993=>"111111000",
  60994=>"000000001",
  60995=>"111111010",
  60996=>"100000100",
  60997=>"100000000",
  60998=>"000000000",
  60999=>"111111001",
  61000=>"011111011",
  61001=>"111111111",
  61002=>"111111000",
  61003=>"111000010",
  61004=>"000000000",
  61005=>"111011010",
  61006=>"111000100",
  61007=>"000101111",
  61008=>"111011111",
  61009=>"000011111",
  61010=>"110111111",
  61011=>"000001101",
  61012=>"111100000",
  61013=>"110111111",
  61014=>"111111111",
  61015=>"111111010",
  61016=>"111000000",
  61017=>"101000000",
  61018=>"001000011",
  61019=>"111111110",
  61020=>"000000111",
  61021=>"110111111",
  61022=>"110110100",
  61023=>"000100110",
  61024=>"000000011",
  61025=>"100100100",
  61026=>"000000111",
  61027=>"000010000",
  61028=>"000000011",
  61029=>"000000111",
  61030=>"111100000",
  61031=>"110000000",
  61032=>"111111000",
  61033=>"000000000",
  61034=>"000000111",
  61035=>"000000000",
  61036=>"010110000",
  61037=>"000000110",
  61038=>"111111111",
  61039=>"000001000",
  61040=>"101000001",
  61041=>"001000000",
  61042=>"010000000",
  61043=>"000000110",
  61044=>"111101000",
  61045=>"111111110",
  61046=>"110010111",
  61047=>"000111000",
  61048=>"110001111",
  61049=>"100000000",
  61050=>"001111111",
  61051=>"000100000",
  61052=>"111110110",
  61053=>"111111000",
  61054=>"111111110",
  61055=>"011110010",
  61056=>"001001000",
  61057=>"111111100",
  61058=>"111011111",
  61059=>"000000111",
  61060=>"000000000",
  61061=>"011001000",
  61062=>"100001111",
  61063=>"110100101",
  61064=>"000000000",
  61065=>"000010000",
  61066=>"000000000",
  61067=>"111111011",
  61068=>"011111011",
  61069=>"010000111",
  61070=>"000111110",
  61071=>"000000111",
  61072=>"000000101",
  61073=>"111101000",
  61074=>"110000100",
  61075=>"111111001",
  61076=>"000100101",
  61077=>"100110111",
  61078=>"000000000",
  61079=>"111111111",
  61080=>"111100111",
  61081=>"000100000",
  61082=>"111000000",
  61083=>"111111000",
  61084=>"111110111",
  61085=>"000001111",
  61086=>"111111000",
  61087=>"000000000",
  61088=>"000001000",
  61089=>"000100001",
  61090=>"110111111",
  61091=>"000000000",
  61092=>"100100000",
  61093=>"100100000",
  61094=>"001011111",
  61095=>"001011011",
  61096=>"111111000",
  61097=>"101000001",
  61098=>"000010011",
  61099=>"110110000",
  61100=>"010110000",
  61101=>"000000000",
  61102=>"100100000",
  61103=>"000000111",
  61104=>"000011111",
  61105=>"011010000",
  61106=>"011011111",
  61107=>"011010010",
  61108=>"100101110",
  61109=>"111111111",
  61110=>"000000000",
  61111=>"000000000",
  61112=>"000000000",
  61113=>"011011000",
  61114=>"000000010",
  61115=>"100001001",
  61116=>"111110000",
  61117=>"001000000",
  61118=>"011111010",
  61119=>"111000011",
  61120=>"010111111",
  61121=>"000000111",
  61122=>"110111000",
  61123=>"000000111",
  61124=>"000000111",
  61125=>"000111111",
  61126=>"000001111",
  61127=>"000000000",
  61128=>"001000111",
  61129=>"001000110",
  61130=>"100100000",
  61131=>"000000110",
  61132=>"000000111",
  61133=>"010111111",
  61134=>"110000000",
  61135=>"100000000",
  61136=>"011000000",
  61137=>"111110000",
  61138=>"011010000",
  61139=>"011000000",
  61140=>"100101011",
  61141=>"000000001",
  61142=>"111111011",
  61143=>"110111111",
  61144=>"000000100",
  61145=>"000111111",
  61146=>"101001000",
  61147=>"010000000",
  61148=>"111001100",
  61149=>"111000000",
  61150=>"001101111",
  61151=>"000000100",
  61152=>"001000000",
  61153=>"011001111",
  61154=>"001111001",
  61155=>"111110000",
  61156=>"110111101",
  61157=>"001111001",
  61158=>"111111100",
  61159=>"110110111",
  61160=>"000000000",
  61161=>"000011111",
  61162=>"110000111",
  61163=>"111111100",
  61164=>"111111111",
  61165=>"000111111",
  61166=>"000011001",
  61167=>"011001101",
  61168=>"111111101",
  61169=>"111000000",
  61170=>"001000000",
  61171=>"000000111",
  61172=>"111111111",
  61173=>"000110001",
  61174=>"111111111",
  61175=>"000110111",
  61176=>"001001000",
  61177=>"000000000",
  61178=>"000000000",
  61179=>"111111000",
  61180=>"011111100",
  61181=>"100001011",
  61182=>"110100000",
  61183=>"000010000",
  61184=>"111010001",
  61185=>"111100000",
  61186=>"000000000",
  61187=>"110100000",
  61188=>"000000001",
  61189=>"111010000",
  61190=>"001000110",
  61191=>"000000000",
  61192=>"010110111",
  61193=>"011011000",
  61194=>"111011001",
  61195=>"111000111",
  61196=>"111111111",
  61197=>"010000000",
  61198=>"000001000",
  61199=>"000000000",
  61200=>"111000000",
  61201=>"100100111",
  61202=>"000111111",
  61203=>"011011000",
  61204=>"010000000",
  61205=>"111101001",
  61206=>"011011001",
  61207=>"000001000",
  61208=>"100110111",
  61209=>"100001001",
  61210=>"111110100",
  61211=>"111111111",
  61212=>"100100000",
  61213=>"111111111",
  61214=>"011000010",
  61215=>"111101111",
  61216=>"000100111",
  61217=>"010000000",
  61218=>"000000101",
  61219=>"111111111",
  61220=>"111000110",
  61221=>"001000010",
  61222=>"111111111",
  61223=>"000001110",
  61224=>"001111111",
  61225=>"111111011",
  61226=>"111001000",
  61227=>"111000111",
  61228=>"001111100",
  61229=>"110000000",
  61230=>"111011010",
  61231=>"110111110",
  61232=>"110110110",
  61233=>"000000000",
  61234=>"111111111",
  61235=>"111111111",
  61236=>"111111111",
  61237=>"001000111",
  61238=>"000000000",
  61239=>"111001011",
  61240=>"100011111",
  61241=>"000001001",
  61242=>"111111111",
  61243=>"000011011",
  61244=>"111111111",
  61245=>"101000000",
  61246=>"110100101",
  61247=>"000000000",
  61248=>"111111111",
  61249=>"011111111",
  61250=>"110100110",
  61251=>"111000000",
  61252=>"000000000",
  61253=>"000001111",
  61254=>"001001111",
  61255=>"000000000",
  61256=>"000000000",
  61257=>"111000000",
  61258=>"001100000",
  61259=>"111111110",
  61260=>"111101111",
  61261=>"101111111",
  61262=>"111111111",
  61263=>"001001000",
  61264=>"110000100",
  61265=>"111000000",
  61266=>"000100101",
  61267=>"000100110",
  61268=>"000000100",
  61269=>"001001011",
  61270=>"111001001",
  61271=>"000000111",
  61272=>"000000110",
  61273=>"110111111",
  61274=>"101100100",
  61275=>"010111111",
  61276=>"001011011",
  61277=>"000000000",
  61278=>"000000000",
  61279=>"111111111",
  61280=>"100001001",
  61281=>"111111111",
  61282=>"111110100",
  61283=>"111111000",
  61284=>"110100100",
  61285=>"000000100",
  61286=>"000000111",
  61287=>"000000000",
  61288=>"111111000",
  61289=>"000000111",
  61290=>"110100001",
  61291=>"011100110",
  61292=>"000000111",
  61293=>"111011010",
  61294=>"000000000",
  61295=>"000000111",
  61296=>"000000110",
  61297=>"011111111",
  61298=>"001001000",
  61299=>"111011100",
  61300=>"000000101",
  61301=>"111111000",
  61302=>"110000111",
  61303=>"000000000",
  61304=>"111001000",
  61305=>"111101001",
  61306=>"111111000",
  61307=>"100100000",
  61308=>"011000001",
  61309=>"111000000",
  61310=>"111110000",
  61311=>"000000011",
  61312=>"110110000",
  61313=>"111101000",
  61314=>"111111000",
  61315=>"111000000",
  61316=>"100110000",
  61317=>"010010000",
  61318=>"000101101",
  61319=>"111111111",
  61320=>"111111000",
  61321=>"000000000",
  61322=>"111110110",
  61323=>"000001001",
  61324=>"111000111",
  61325=>"011000000",
  61326=>"000001001",
  61327=>"000011111",
  61328=>"011000000",
  61329=>"111110000",
  61330=>"000000000",
  61331=>"111111111",
  61332=>"110001011",
  61333=>"000010010",
  61334=>"100101001",
  61335=>"110000000",
  61336=>"101000111",
  61337=>"000000000",
  61338=>"111110110",
  61339=>"000000000",
  61340=>"111111000",
  61341=>"111000000",
  61342=>"000000000",
  61343=>"001000000",
  61344=>"000000000",
  61345=>"100100101",
  61346=>"111111000",
  61347=>"111000000",
  61348=>"000000000",
  61349=>"000010110",
  61350=>"001011111",
  61351=>"000000000",
  61352=>"100000000",
  61353=>"101101000",
  61354=>"100000110",
  61355=>"000000100",
  61356=>"000000111",
  61357=>"000100111",
  61358=>"000000000",
  61359=>"010000011",
  61360=>"111111111",
  61361=>"110110000",
  61362=>"110000000",
  61363=>"011111111",
  61364=>"000000000",
  61365=>"111111111",
  61366=>"100111111",
  61367=>"000001001",
  61368=>"111001111",
  61369=>"000010111",
  61370=>"101000000",
  61371=>"111111110",
  61372=>"101111011",
  61373=>"111111001",
  61374=>"111000001",
  61375=>"011000100",
  61376=>"111001000",
  61377=>"111111000",
  61378=>"111111111",
  61379=>"000011001",
  61380=>"110000000",
  61381=>"110110100",
  61382=>"100100111",
  61383=>"000001000",
  61384=>"111111101",
  61385=>"000000000",
  61386=>"111000000",
  61387=>"111110111",
  61388=>"101000111",
  61389=>"000100100",
  61390=>"111001000",
  61391=>"000001011",
  61392=>"100000000",
  61393=>"111111111",
  61394=>"110000111",
  61395=>"001001101",
  61396=>"011011011",
  61397=>"110100000",
  61398=>"111111110",
  61399=>"111010000",
  61400=>"001000000",
  61401=>"111111111",
  61402=>"111111111",
  61403=>"000000000",
  61404=>"011111111",
  61405=>"100001111",
  61406=>"000000000",
  61407=>"000000001",
  61408=>"111000000",
  61409=>"011111110",
  61410=>"000000000",
  61411=>"000000000",
  61412=>"001111111",
  61413=>"000110000",
  61414=>"110110111",
  61415=>"000000101",
  61416=>"100100100",
  61417=>"000001000",
  61418=>"000111111",
  61419=>"111111111",
  61420=>"010001111",
  61421=>"011011011",
  61422=>"111001000",
  61423=>"001111111",
  61424=>"000010001",
  61425=>"100100100",
  61426=>"000000111",
  61427=>"110110000",
  61428=>"000000001",
  61429=>"100111111",
  61430=>"111000000",
  61431=>"111111111",
  61432=>"011011111",
  61433=>"000000000",
  61434=>"010000111",
  61435=>"111111011",
  61436=>"111000000",
  61437=>"111111100",
  61438=>"010000110",
  61439=>"000000000",
  61440=>"001000111",
  61441=>"111000000",
  61442=>"111111111",
  61443=>"111100111",
  61444=>"000000100",
  61445=>"010000000",
  61446=>"011001000",
  61447=>"000000000",
  61448=>"111111111",
  61449=>"001010000",
  61450=>"011000000",
  61451=>"101111111",
  61452=>"111101111",
  61453=>"001000011",
  61454=>"000011010",
  61455=>"111100100",
  61456=>"110111001",
  61457=>"110011111",
  61458=>"111000000",
  61459=>"111111111",
  61460=>"110111111",
  61461=>"111110000",
  61462=>"110000001",
  61463=>"111110000",
  61464=>"110000000",
  61465=>"100110111",
  61466=>"101101000",
  61467=>"111000000",
  61468=>"001000111",
  61469=>"000000111",
  61470=>"111111001",
  61471=>"111110110",
  61472=>"100100000",
  61473=>"100111001",
  61474=>"110110011",
  61475=>"000001101",
  61476=>"111111001",
  61477=>"000101000",
  61478=>"001000000",
  61479=>"111100000",
  61480=>"000000000",
  61481=>"000001000",
  61482=>"010000000",
  61483=>"111011000",
  61484=>"111111111",
  61485=>"111001111",
  61486=>"000000111",
  61487=>"111111111",
  61488=>"111111111",
  61489=>"000000100",
  61490=>"011100100",
  61491=>"111111111",
  61492=>"111111011",
  61493=>"110110100",
  61494=>"111111111",
  61495=>"000110110",
  61496=>"000011111",
  61497=>"000000111",
  61498=>"000000001",
  61499=>"111000000",
  61500=>"111111100",
  61501=>"111011111",
  61502=>"000111111",
  61503=>"100000110",
  61504=>"111111000",
  61505=>"000000111",
  61506=>"100100111",
  61507=>"000111111",
  61508=>"100111011",
  61509=>"110100111",
  61510=>"111111000",
  61511=>"111111111",
  61512=>"001100110",
  61513=>"111111111",
  61514=>"111111000",
  61515=>"101100111",
  61516=>"000000010",
  61517=>"000000000",
  61518=>"101000000",
  61519=>"000000100",
  61520=>"000000101",
  61521=>"111111000",
  61522=>"111111110",
  61523=>"100100000",
  61524=>"111111111",
  61525=>"111111111",
  61526=>"111111100",
  61527=>"000100101",
  61528=>"111011111",
  61529=>"100000111",
  61530=>"000000111",
  61531=>"000000111",
  61532=>"111111000",
  61533=>"001000000",
  61534=>"110000000",
  61535=>"111000000",
  61536=>"100100000",
  61537=>"111110110",
  61538=>"111001001",
  61539=>"111100111",
  61540=>"111011010",
  61541=>"111000101",
  61542=>"000000000",
  61543=>"000001000",
  61544=>"111111111",
  61545=>"111111111",
  61546=>"000000111",
  61547=>"111111010",
  61548=>"000111111",
  61549=>"000001000",
  61550=>"000111100",
  61551=>"110111000",
  61552=>"011001000",
  61553=>"000010111",
  61554=>"100111000",
  61555=>"111100000",
  61556=>"011000000",
  61557=>"111100000",
  61558=>"111001000",
  61559=>"000000000",
  61560=>"000000000",
  61561=>"111111111",
  61562=>"000000011",
  61563=>"100000000",
  61564=>"100100000",
  61565=>"000010000",
  61566=>"011001111",
  61567=>"000000000",
  61568=>"000000000",
  61569=>"000000111",
  61570=>"111000000",
  61571=>"100000000",
  61572=>"111111111",
  61573=>"000000000",
  61574=>"000000111",
  61575=>"111111010",
  61576=>"000000000",
  61577=>"000000000",
  61578=>"000000000",
  61579=>"111111000",
  61580=>"000000000",
  61581=>"000000000",
  61582=>"111111111",
  61583=>"100111111",
  61584=>"000000101",
  61585=>"000000000",
  61586=>"000111111",
  61587=>"111101000",
  61588=>"110110111",
  61589=>"111111000",
  61590=>"101111111",
  61591=>"111111000",
  61592=>"111001011",
  61593=>"010100001",
  61594=>"000000111",
  61595=>"000111100",
  61596=>"111111111",
  61597=>"000111111",
  61598=>"111110111",
  61599=>"111000000",
  61600=>"111001000",
  61601=>"100111011",
  61602=>"111001000",
  61603=>"000000000",
  61604=>"000110111",
  61605=>"111110111",
  61606=>"111111111",
  61607=>"111111111",
  61608=>"011011110",
  61609=>"000000111",
  61610=>"111111000",
  61611=>"000100110",
  61612=>"111111111",
  61613=>"110001001",
  61614=>"111001000",
  61615=>"000000111",
  61616=>"000000111",
  61617=>"011000100",
  61618=>"101101111",
  61619=>"111100000",
  61620=>"000000000",
  61621=>"111111001",
  61622=>"000000000",
  61623=>"101111111",
  61624=>"111111000",
  61625=>"000000111",
  61626=>"011111011",
  61627=>"111001001",
  61628=>"111111111",
  61629=>"000000000",
  61630=>"011011111",
  61631=>"001001111",
  61632=>"111000000",
  61633=>"000000000",
  61634=>"100000000",
  61635=>"000000111",
  61636=>"111101111",
  61637=>"111111001",
  61638=>"111111111",
  61639=>"110111100",
  61640=>"000000000",
  61641=>"111110110",
  61642=>"000000001",
  61643=>"000010000",
  61644=>"000000000",
  61645=>"000000000",
  61646=>"111001111",
  61647=>"011000000",
  61648=>"001011000",
  61649=>"100100111",
  61650=>"001000001",
  61651=>"001000100",
  61652=>"100110000",
  61653=>"111111111",
  61654=>"000101000",
  61655=>"010111111",
  61656=>"111000000",
  61657=>"111111111",
  61658=>"111011000",
  61659=>"111111001",
  61660=>"111100000",
  61661=>"100100111",
  61662=>"000001001",
  61663=>"111011000",
  61664=>"000000111",
  61665=>"001011000",
  61666=>"111000000",
  61667=>"111001101",
  61668=>"111111111",
  61669=>"000000100",
  61670=>"111000101",
  61671=>"111111011",
  61672=>"101001010",
  61673=>"111111111",
  61674=>"101111111",
  61675=>"011111111",
  61676=>"001001111",
  61677=>"111111110",
  61678=>"000000111",
  61679=>"111111111",
  61680=>"111111111",
  61681=>"011111000",
  61682=>"000001001",
  61683=>"000000000",
  61684=>"000000000",
  61685=>"111011001",
  61686=>"101111000",
  61687=>"100000000",
  61688=>"011111111",
  61689=>"111111111",
  61690=>"000000111",
  61691=>"001000000",
  61692=>"111110110",
  61693=>"111111111",
  61694=>"111000111",
  61695=>"000000000",
  61696=>"111001101",
  61697=>"111111000",
  61698=>"111110110",
  61699=>"011111111",
  61700=>"110000111",
  61701=>"000110011",
  61702=>"111111111",
  61703=>"110111111",
  61704=>"000000000",
  61705=>"000000110",
  61706=>"111111101",
  61707=>"011111001",
  61708=>"000000001",
  61709=>"000000000",
  61710=>"000000001",
  61711=>"000000000",
  61712=>"000000001",
  61713=>"000100000",
  61714=>"111100000",
  61715=>"000000001",
  61716=>"111111001",
  61717=>"100100000",
  61718=>"100100000",
  61719=>"111000000",
  61720=>"000000100",
  61721=>"111100100",
  61722=>"111000000",
  61723=>"000111000",
  61724=>"001000001",
  61725=>"000100111",
  61726=>"000000001",
  61727=>"111111010",
  61728=>"000000000",
  61729=>"111000000",
  61730=>"000000000",
  61731=>"000011000",
  61732=>"000000100",
  61733=>"111100000",
  61734=>"000000000",
  61735=>"000001011",
  61736=>"111111100",
  61737=>"111100000",
  61738=>"011000011",
  61739=>"000111111",
  61740=>"111000000",
  61741=>"000001011",
  61742=>"001000000",
  61743=>"010111111",
  61744=>"000000110",
  61745=>"000000000",
  61746=>"000011001",
  61747=>"011111111",
  61748=>"000000000",
  61749=>"111000000",
  61750=>"000000000",
  61751=>"111101001",
  61752=>"000111000",
  61753=>"111111000",
  61754=>"000000111",
  61755=>"100111111",
  61756=>"000000100",
  61757=>"000000000",
  61758=>"000000000",
  61759=>"111000111",
  61760=>"000100111",
  61761=>"111101111",
  61762=>"101000000",
  61763=>"000000000",
  61764=>"000000100",
  61765=>"100111111",
  61766=>"111111000",
  61767=>"000001001",
  61768=>"000000100",
  61769=>"011111111",
  61770=>"110011111",
  61771=>"000110111",
  61772=>"111111000",
  61773=>"000100000",
  61774=>"111001001",
  61775=>"111111000",
  61776=>"111001000",
  61777=>"000100100",
  61778=>"111110110",
  61779=>"000111111",
  61780=>"011111111",
  61781=>"011011011",
  61782=>"111111111",
  61783=>"111111111",
  61784=>"111100110",
  61785=>"101101111",
  61786=>"100111111",
  61787=>"111111110",
  61788=>"000001000",
  61789=>"111111001",
  61790=>"100000000",
  61791=>"110111000",
  61792=>"000111111",
  61793=>"111000000",
  61794=>"001000100",
  61795=>"111000000",
  61796=>"000000111",
  61797=>"000000000",
  61798=>"111111111",
  61799=>"111000000",
  61800=>"011001111",
  61801=>"111111111",
  61802=>"000000100",
  61803=>"011111111",
  61804=>"111100000",
  61805=>"000001111",
  61806=>"000111111",
  61807=>"000111111",
  61808=>"001011111",
  61809=>"000110111",
  61810=>"101000100",
  61811=>"000001100",
  61812=>"111111111",
  61813=>"111111000",
  61814=>"100011101",
  61815=>"111111000",
  61816=>"111000000",
  61817=>"000101111",
  61818=>"111001000",
  61819=>"111111111",
  61820=>"111111010",
  61821=>"111011000",
  61822=>"111111111",
  61823=>"111111111",
  61824=>"000000000",
  61825=>"010010111",
  61826=>"111111111",
  61827=>"000000111",
  61828=>"000000111",
  61829=>"000000111",
  61830=>"111111111",
  61831=>"001000100",
  61832=>"111111111",
  61833=>"110000111",
  61834=>"111110111",
  61835=>"111111111",
  61836=>"111000000",
  61837=>"010001001",
  61838=>"000000101",
  61839=>"111111000",
  61840=>"111110111",
  61841=>"000000000",
  61842=>"000001011",
  61843=>"000000111",
  61844=>"111000000",
  61845=>"111011000",
  61846=>"111111011",
  61847=>"100100001",
  61848=>"000111111",
  61849=>"000000001",
  61850=>"000000111",
  61851=>"111000000",
  61852=>"111111000",
  61853=>"111001111",
  61854=>"000101001",
  61855=>"000000000",
  61856=>"001001000",
  61857=>"110110000",
  61858=>"100000000",
  61859=>"000111111",
  61860=>"000100110",
  61861=>"000000000",
  61862=>"000000001",
  61863=>"111011001",
  61864=>"001111111",
  61865=>"000000000",
  61866=>"101000101",
  61867=>"000000011",
  61868=>"111111010",
  61869=>"111110110",
  61870=>"111111111",
  61871=>"111000000",
  61872=>"010011111",
  61873=>"000000001",
  61874=>"000000000",
  61875=>"111111111",
  61876=>"000000110",
  61877=>"111000000",
  61878=>"011111111",
  61879=>"001001110",
  61880=>"011111111",
  61881=>"101001001",
  61882=>"101000000",
  61883=>"000000101",
  61884=>"111111111",
  61885=>"100000100",
  61886=>"111001001",
  61887=>"000000000",
  61888=>"111111111",
  61889=>"111000110",
  61890=>"000000111",
  61891=>"011000000",
  61892=>"111111111",
  61893=>"111111111",
  61894=>"000000000",
  61895=>"000000101",
  61896=>"111011001",
  61897=>"111111000",
  61898=>"011000000",
  61899=>"000000000",
  61900=>"000000000",
  61901=>"001010100",
  61902=>"000000000",
  61903=>"111111000",
  61904=>"111011011",
  61905=>"000000100",
  61906=>"111111111",
  61907=>"000000100",
  61908=>"011111000",
  61909=>"111001000",
  61910=>"111111111",
  61911=>"000000000",
  61912=>"111001111",
  61913=>"100100111",
  61914=>"111110000",
  61915=>"001001001",
  61916=>"100111111",
  61917=>"111111111",
  61918=>"100000000",
  61919=>"111000001",
  61920=>"000000100",
  61921=>"000111111",
  61922=>"000000000",
  61923=>"001111111",
  61924=>"001111111",
  61925=>"111111111",
  61926=>"111010110",
  61927=>"011000000",
  61928=>"110110000",
  61929=>"000000000",
  61930=>"000000100",
  61931=>"111111111",
  61932=>"111111001",
  61933=>"000001011",
  61934=>"111101000",
  61935=>"011111011",
  61936=>"000011001",
  61937=>"111000000",
  61938=>"011111111",
  61939=>"111111111",
  61940=>"000000111",
  61941=>"111111000",
  61942=>"011111000",
  61943=>"110010011",
  61944=>"000000111",
  61945=>"111101100",
  61946=>"111111001",
  61947=>"111011000",
  61948=>"110000111",
  61949=>"001000000",
  61950=>"000000000",
  61951=>"000000000",
  61952=>"000000100",
  61953=>"000000000",
  61954=>"111001000",
  61955=>"111111111",
  61956=>"111111011",
  61957=>"000001011",
  61958=>"001111111",
  61959=>"111111111",
  61960=>"111000001",
  61961=>"100100111",
  61962=>"111111010",
  61963=>"111001000",
  61964=>"011011011",
  61965=>"000000000",
  61966=>"111111000",
  61967=>"000000000",
  61968=>"110000000",
  61969=>"011000000",
  61970=>"001001111",
  61971=>"000111111",
  61972=>"000100000",
  61973=>"111111111",
  61974=>"111111001",
  61975=>"111111111",
  61976=>"000000000",
  61977=>"011111110",
  61978=>"111111111",
  61979=>"100101110",
  61980=>"000000000",
  61981=>"000111111",
  61982=>"000000001",
  61983=>"001000000",
  61984=>"001001000",
  61985=>"111111111",
  61986=>"111011111",
  61987=>"101001001",
  61988=>"111111111",
  61989=>"010011001",
  61990=>"111101000",
  61991=>"111111000",
  61992=>"111111010",
  61993=>"000000000",
  61994=>"000000000",
  61995=>"111111111",
  61996=>"000000000",
  61997=>"000000000",
  61998=>"000100000",
  61999=>"000100111",
  62000=>"101101000",
  62001=>"000000000",
  62002=>"101001001",
  62003=>"110111111",
  62004=>"000000000",
  62005=>"111011011",
  62006=>"110000000",
  62007=>"000000111",
  62008=>"001000111",
  62009=>"001111101",
  62010=>"111111111",
  62011=>"000000000",
  62012=>"000101101",
  62013=>"001001111",
  62014=>"000001001",
  62015=>"111111000",
  62016=>"111101000",
  62017=>"011011111",
  62018=>"111000000",
  62019=>"111111101",
  62020=>"100000001",
  62021=>"000000000",
  62022=>"000000000",
  62023=>"111111111",
  62024=>"100100100",
  62025=>"000000000",
  62026=>"111101000",
  62027=>"111111111",
  62028=>"000000000",
  62029=>"110111111",
  62030=>"000000000",
  62031=>"000000000",
  62032=>"100110000",
  62033=>"110110000",
  62034=>"000000000",
  62035=>"111000111",
  62036=>"000111111",
  62037=>"111111011",
  62038=>"111111111",
  62039=>"000000000",
  62040=>"000000100",
  62041=>"000000111",
  62042=>"111111111",
  62043=>"000000001",
  62044=>"100100111",
  62045=>"001000111",
  62046=>"001011111",
  62047=>"000010000",
  62048=>"000000110",
  62049=>"000000000",
  62050=>"000000000",
  62051=>"000000000",
  62052=>"111111111",
  62053=>"111101000",
  62054=>"000000000",
  62055=>"000110010",
  62056=>"000000000",
  62057=>"000000000",
  62058=>"111111111",
  62059=>"111000000",
  62060=>"000000111",
  62061=>"111110111",
  62062=>"101000000",
  62063=>"000000000",
  62064=>"111111111",
  62065=>"101111111",
  62066=>"011001011",
  62067=>"000001111",
  62068=>"111011111",
  62069=>"000000111",
  62070=>"000000000",
  62071=>"000000000",
  62072=>"010010110",
  62073=>"111111111",
  62074=>"111111111",
  62075=>"000101111",
  62076=>"000000001",
  62077=>"000000000",
  62078=>"001000000",
  62079=>"000000000",
  62080=>"000010000",
  62081=>"000011111",
  62082=>"100000100",
  62083=>"100110111",
  62084=>"111111000",
  62085=>"000001111",
  62086=>"000000000",
  62087=>"000000100",
  62088=>"111001000",
  62089=>"000110000",
  62090=>"000000000",
  62091=>"011000010",
  62092=>"000000110",
  62093=>"110111111",
  62094=>"111001000",
  62095=>"000000110",
  62096=>"000000000",
  62097=>"000000100",
  62098=>"000001000",
  62099=>"000110000",
  62100=>"110001111",
  62101=>"001000000",
  62102=>"111111111",
  62103=>"001001000",
  62104=>"010111000",
  62105=>"000000000",
  62106=>"000000000",
  62107=>"110110000",
  62108=>"011111011",
  62109=>"100100000",
  62110=>"100110000",
  62111=>"111111000",
  62112=>"000000100",
  62113=>"100000000",
  62114=>"111111111",
  62115=>"000000000",
  62116=>"111101001",
  62117=>"100000000",
  62118=>"000000000",
  62119=>"000011011",
  62120=>"110100000",
  62121=>"000000000",
  62122=>"111011000",
  62123=>"111111111",
  62124=>"001011011",
  62125=>"111111111",
  62126=>"111111111",
  62127=>"111111111",
  62128=>"000000000",
  62129=>"110100100",
  62130=>"111111110",
  62131=>"000000100",
  62132=>"000000000",
  62133=>"111111001",
  62134=>"011111100",
  62135=>"111000000",
  62136=>"011110100",
  62137=>"111111111",
  62138=>"111111111",
  62139=>"111111011",
  62140=>"111111101",
  62141=>"111111111",
  62142=>"111111111",
  62143=>"000000000",
  62144=>"101100000",
  62145=>"100111111",
  62146=>"000001000",
  62147=>"111111001",
  62148=>"111111111",
  62149=>"000000000",
  62150=>"010110011",
  62151=>"111101100",
  62152=>"111010000",
  62153=>"100101011",
  62154=>"111111011",
  62155=>"000000000",
  62156=>"111001001",
  62157=>"000110000",
  62158=>"000000000",
  62159=>"111111001",
  62160=>"000000010",
  62161=>"010111000",
  62162=>"000111111",
  62163=>"010111111",
  62164=>"111111111",
  62165=>"111111111",
  62166=>"000001000",
  62167=>"000110110",
  62168=>"111111000",
  62169=>"100100000",
  62170=>"111111111",
  62171=>"111111111",
  62172=>"000000110",
  62173=>"000000000",
  62174=>"000001111",
  62175=>"000000000",
  62176=>"000000000",
  62177=>"000000011",
  62178=>"000000000",
  62179=>"000101001",
  62180=>"000011011",
  62181=>"000000000",
  62182=>"111111001",
  62183=>"000000100",
  62184=>"010000010",
  62185=>"000101100",
  62186=>"011111000",
  62187=>"100100111",
  62188=>"000100100",
  62189=>"000000000",
  62190=>"100111111",
  62191=>"111100000",
  62192=>"100000000",
  62193=>"000000000",
  62194=>"000000000",
  62195=>"111101000",
  62196=>"111111010",
  62197=>"011011010",
  62198=>"001000000",
  62199=>"000011011",
  62200=>"111111111",
  62201=>"111111111",
  62202=>"000000000",
  62203=>"111111111",
  62204=>"000100101",
  62205=>"100101100",
  62206=>"000000100",
  62207=>"111111111",
  62208=>"000000000",
  62209=>"011111000",
  62210=>"111000000",
  62211=>"000000000",
  62212=>"111011001",
  62213=>"011010000",
  62214=>"111111111",
  62215=>"101000000",
  62216=>"100101001",
  62217=>"100100000",
  62218=>"011011111",
  62219=>"111111111",
  62220=>"111101000",
  62221=>"100111111",
  62222=>"010110111",
  62223=>"000000000",
  62224=>"000010000",
  62225=>"111011000",
  62226=>"111010000",
  62227=>"000000000",
  62228=>"010010000",
  62229=>"111111011",
  62230=>"001111111",
  62231=>"001000000",
  62232=>"101000111",
  62233=>"111100001",
  62234=>"000000100",
  62235=>"010000000",
  62236=>"111111101",
  62237=>"111111111",
  62238=>"000000000",
  62239=>"101111110",
  62240=>"111111011",
  62241=>"000000000",
  62242=>"101100000",
  62243=>"111111111",
  62244=>"000000000",
  62245=>"110110000",
  62246=>"111111110",
  62247=>"111111111",
  62248=>"111111111",
  62249=>"000000000",
  62250=>"111110110",
  62251=>"000000000",
  62252=>"000000100",
  62253=>"011100100",
  62254=>"000000000",
  62255=>"110010000",
  62256=>"001111110",
  62257=>"000111011",
  62258=>"000000000",
  62259=>"000111111",
  62260=>"000000000",
  62261=>"000000000",
  62262=>"111111111",
  62263=>"000000000",
  62264=>"111011000",
  62265=>"001000000",
  62266=>"000000000",
  62267=>"111000000",
  62268=>"001000000",
  62269=>"111111111",
  62270=>"000000000",
  62271=>"000011110",
  62272=>"010111111",
  62273=>"011101000",
  62274=>"001111111",
  62275=>"000100111",
  62276=>"100111000",
  62277=>"010100000",
  62278=>"110100100",
  62279=>"111000000",
  62280=>"000000000",
  62281=>"000000000",
  62282=>"111011001",
  62283=>"000111000",
  62284=>"000001111",
  62285=>"111011000",
  62286=>"101101100",
  62287=>"000111111",
  62288=>"000000111",
  62289=>"111111000",
  62290=>"111111010",
  62291=>"111111111",
  62292=>"111111111",
  62293=>"011001001",
  62294=>"000000000",
  62295=>"100111111",
  62296=>"100101101",
  62297=>"000000000",
  62298=>"000100000",
  62299=>"111111111",
  62300=>"111111010",
  62301=>"111111111",
  62302=>"101000000",
  62303=>"000100000",
  62304=>"000000010",
  62305=>"000000001",
  62306=>"011001101",
  62307=>"111111000",
  62308=>"001001001",
  62309=>"000000000",
  62310=>"000000100",
  62311=>"010000000",
  62312=>"000000000",
  62313=>"000000000",
  62314=>"000000000",
  62315=>"001111111",
  62316=>"111111100",
  62317=>"111000000",
  62318=>"000000000",
  62319=>"000000000",
  62320=>"000000000",
  62321=>"111111111",
  62322=>"100100110",
  62323=>"111111011",
  62324=>"011011001",
  62325=>"000000000",
  62326=>"000000000",
  62327=>"000100111",
  62328=>"000000000",
  62329=>"111010010",
  62330=>"111000100",
  62331=>"000010010",
  62332=>"000001011",
  62333=>"000000000",
  62334=>"100110111",
  62335=>"100111111",
  62336=>"000000000",
  62337=>"001000001",
  62338=>"100000000",
  62339=>"011001001",
  62340=>"110110000",
  62341=>"110111000",
  62342=>"000001011",
  62343=>"111001000",
  62344=>"111111110",
  62345=>"100101000",
  62346=>"000010010",
  62347=>"111111111",
  62348=>"111111111",
  62349=>"111110000",
  62350=>"000000011",
  62351=>"000000000",
  62352=>"111111111",
  62353=>"111111001",
  62354=>"111111111",
  62355=>"100100000",
  62356=>"111111111",
  62357=>"000011111",
  62358=>"111111111",
  62359=>"101101000",
  62360=>"111111111",
  62361=>"000011111",
  62362=>"111111111",
  62363=>"111111111",
  62364=>"000101000",
  62365=>"111001000",
  62366=>"000000101",
  62367=>"111111111",
  62368=>"000000000",
  62369=>"000011011",
  62370=>"111000000",
  62371=>"000000000",
  62372=>"100000001",
  62373=>"111111111",
  62374=>"000000000",
  62375=>"000000000",
  62376=>"111111111",
  62377=>"111111110",
  62378=>"111111011",
  62379=>"001000111",
  62380=>"110111111",
  62381=>"111111111",
  62382=>"111111100",
  62383=>"000000000",
  62384=>"100111111",
  62385=>"111011000",
  62386=>"000000000",
  62387=>"111000100",
  62388=>"000000000",
  62389=>"110000000",
  62390=>"000000000",
  62391=>"000000000",
  62392=>"101110110",
  62393=>"111111011",
  62394=>"000111011",
  62395=>"000010000",
  62396=>"000000000",
  62397=>"111110000",
  62398=>"101000000",
  62399=>"001011001",
  62400=>"000000000",
  62401=>"111111011",
  62402=>"111111010",
  62403=>"000100000",
  62404=>"001000111",
  62405=>"101111111",
  62406=>"001101110",
  62407=>"000000000",
  62408=>"000000000",
  62409=>"101101000",
  62410=>"000101111",
  62411=>"000000111",
  62412=>"111000001",
  62413=>"100000000",
  62414=>"111001111",
  62415=>"111111111",
  62416=>"000000010",
  62417=>"000111111",
  62418=>"111111001",
  62419=>"001000001",
  62420=>"001000000",
  62421=>"011011000",
  62422=>"111111000",
  62423=>"100100110",
  62424=>"000000000",
  62425=>"000110110",
  62426=>"000000000",
  62427=>"111111111",
  62428=>"111101101",
  62429=>"000000000",
  62430=>"000000000",
  62431=>"100011000",
  62432=>"000000100",
  62433=>"000000000",
  62434=>"000000000",
  62435=>"101000000",
  62436=>"100111111",
  62437=>"111111000",
  62438=>"000000000",
  62439=>"100100110",
  62440=>"111111000",
  62441=>"011011001",
  62442=>"100111111",
  62443=>"000000000",
  62444=>"011011000",
  62445=>"111111111",
  62446=>"111111111",
  62447=>"111111111",
  62448=>"111101111",
  62449=>"000000010",
  62450=>"111111011",
  62451=>"000000000",
  62452=>"111111111",
  62453=>"101111111",
  62454=>"100111110",
  62455=>"000001000",
  62456=>"011011111",
  62457=>"011111111",
  62458=>"011011000",
  62459=>"000000111",
  62460=>"011011111",
  62461=>"110110111",
  62462=>"001111111",
  62463=>"100100111",
  62464=>"000000000",
  62465=>"000000000",
  62466=>"111111111",
  62467=>"000100000",
  62468=>"110111111",
  62469=>"111110100",
  62470=>"111111111",
  62471=>"111111111",
  62472=>"110100100",
  62473=>"000000000",
  62474=>"000001001",
  62475=>"000011001",
  62476=>"011011011",
  62477=>"000000000",
  62478=>"111111111",
  62479=>"001000000",
  62480=>"000000000",
  62481=>"000000101",
  62482=>"111111111",
  62483=>"000000000",
  62484=>"000111111",
  62485=>"000000111",
  62486=>"111111000",
  62487=>"100100100",
  62488=>"001011011",
  62489=>"011011111",
  62490=>"000000011",
  62491=>"111111111",
  62492=>"111111111",
  62493=>"000000000",
  62494=>"001000000",
  62495=>"111010111",
  62496=>"000001000",
  62497=>"000000000",
  62498=>"111111111",
  62499=>"111011000",
  62500=>"000111010",
  62501=>"110000000",
  62502=>"111110111",
  62503=>"000000000",
  62504=>"000000111",
  62505=>"111111000",
  62506=>"111111111",
  62507=>"111011111",
  62508=>"001000111",
  62509=>"111111111",
  62510=>"111000000",
  62511=>"000000000",
  62512=>"011001001",
  62513=>"000000000",
  62514=>"111110100",
  62515=>"000000000",
  62516=>"110100000",
  62517=>"110000000",
  62518=>"000111111",
  62519=>"000010001",
  62520=>"100001001",
  62521=>"000000000",
  62522=>"101101111",
  62523=>"111111111",
  62524=>"111101001",
  62525=>"000000000",
  62526=>"000000000",
  62527=>"000001111",
  62528=>"100100000",
  62529=>"010000000",
  62530=>"110001000",
  62531=>"110111111",
  62532=>"000010110",
  62533=>"000000000",
  62534=>"111111111",
  62535=>"110110100",
  62536=>"111111000",
  62537=>"111111111",
  62538=>"110000100",
  62539=>"111111111",
  62540=>"000000000",
  62541=>"000010001",
  62542=>"000000001",
  62543=>"000000000",
  62544=>"111111111",
  62545=>"000000000",
  62546=>"111110111",
  62547=>"111000000",
  62548=>"000011000",
  62549=>"110111111",
  62550=>"111111111",
  62551=>"111001000",
  62552=>"111111111",
  62553=>"111111111",
  62554=>"100101100",
  62555=>"111111111",
  62556=>"000011011",
  62557=>"000000010",
  62558=>"000111111",
  62559=>"000000110",
  62560=>"001111111",
  62561=>"000000000",
  62562=>"010000011",
  62563=>"000000000",
  62564=>"001001111",
  62565=>"000000000",
  62566=>"000000000",
  62567=>"000111010",
  62568=>"111111111",
  62569=>"111111011",
  62570=>"000000000",
  62571=>"000000000",
  62572=>"000000000",
  62573=>"111111111",
  62574=>"111111000",
  62575=>"000000100",
  62576=>"111111111",
  62577=>"111010000",
  62578=>"000000000",
  62579=>"111100010",
  62580=>"100100111",
  62581=>"000000000",
  62582=>"111111111",
  62583=>"000000011",
  62584=>"000000000",
  62585=>"001100101",
  62586=>"001011011",
  62587=>"000010111",
  62588=>"000000000",
  62589=>"000000000",
  62590=>"111111111",
  62591=>"111111011",
  62592=>"100000000",
  62593=>"111010000",
  62594=>"000110111",
  62595=>"000110111",
  62596=>"010010111",
  62597=>"111111111",
  62598=>"111111010",
  62599=>"000101000",
  62600=>"000100000",
  62601=>"100000000",
  62602=>"000000000",
  62603=>"000000000",
  62604=>"111111111",
  62605=>"111111111",
  62606=>"111111111",
  62607=>"000000000",
  62608=>"111111111",
  62609=>"000000000",
  62610=>"110100000",
  62611=>"111000000",
  62612=>"000000000",
  62613=>"000000000",
  62614=>"000000000",
  62615=>"111111111",
  62616=>"101101111",
  62617=>"110111111",
  62618=>"111001001",
  62619=>"110110000",
  62620=>"111111111",
  62621=>"100000001",
  62622=>"000000000",
  62623=>"111111100",
  62624=>"000000100",
  62625=>"000000000",
  62626=>"111111111",
  62627=>"000000000",
  62628=>"001111111",
  62629=>"110110111",
  62630=>"111111111",
  62631=>"011011001",
  62632=>"000000111",
  62633=>"000001111",
  62634=>"111000000",
  62635=>"001000000",
  62636=>"111110100",
  62637=>"110000000",
  62638=>"000000100",
  62639=>"000000000",
  62640=>"111111111",
  62641=>"110110010",
  62642=>"111111100",
  62643=>"101101101",
  62644=>"011000000",
  62645=>"110000000",
  62646=>"000011111",
  62647=>"000000000",
  62648=>"010000111",
  62649=>"000000000",
  62650=>"000000000",
  62651=>"111111111",
  62652=>"010110000",
  62653=>"111010000",
  62654=>"111111111",
  62655=>"100100111",
  62656=>"111111111",
  62657=>"100111011",
  62658=>"000000000",
  62659=>"111111111",
  62660=>"111101001",
  62661=>"111111111",
  62662=>"111111111",
  62663=>"000000000",
  62664=>"000111011",
  62665=>"111101100",
  62666=>"010110000",
  62667=>"000000000",
  62668=>"000000000",
  62669=>"000101111",
  62670=>"111111111",
  62671=>"011111111",
  62672=>"000000000",
  62673=>"000000000",
  62674=>"010011010",
  62675=>"000000000",
  62676=>"111111000",
  62677=>"000000000",
  62678=>"000000000",
  62679=>"110000000",
  62680=>"000000000",
  62681=>"111111111",
  62682=>"110110010",
  62683=>"110111111",
  62684=>"111110111",
  62685=>"000111111",
  62686=>"000111011",
  62687=>"110110000",
  62688=>"111011111",
  62689=>"111111111",
  62690=>"000110111",
  62691=>"111111111",
  62692=>"111111000",
  62693=>"110110110",
  62694=>"111111111",
  62695=>"110011011",
  62696=>"010111111",
  62697=>"000000001",
  62698=>"000000001",
  62699=>"000000011",
  62700=>"101000001",
  62701=>"010010000",
  62702=>"000000001",
  62703=>"000001111",
  62704=>"000000000",
  62705=>"111111110",
  62706=>"111111111",
  62707=>"111000000",
  62708=>"010000000",
  62709=>"000000001",
  62710=>"100100100",
  62711=>"111111111",
  62712=>"001000000",
  62713=>"001000001",
  62714=>"000000000",
  62715=>"101000000",
  62716=>"011001000",
  62717=>"011011001",
  62718=>"111101111",
  62719=>"111111111",
  62720=>"000000000",
  62721=>"001011001",
  62722=>"011111011",
  62723=>"110110000",
  62724=>"111111111",
  62725=>"000011111",
  62726=>"100000111",
  62727=>"111000000",
  62728=>"111111111",
  62729=>"000000000",
  62730=>"111111101",
  62731=>"011000111",
  62732=>"001000100",
  62733=>"000110110",
  62734=>"110110111",
  62735=>"111111111",
  62736=>"010011000",
  62737=>"111111111",
  62738=>"111111111",
  62739=>"111100000",
  62740=>"011111111",
  62741=>"110111111",
  62742=>"111011010",
  62743=>"111001000",
  62744=>"000000000",
  62745=>"100010011",
  62746=>"111111111",
  62747=>"000000000",
  62748=>"111111111",
  62749=>"111111111",
  62750=>"111100000",
  62751=>"101111111",
  62752=>"011111000",
  62753=>"000000000",
  62754=>"100000000",
  62755=>"111111111",
  62756=>"000000011",
  62757=>"111000000",
  62758=>"111111111",
  62759=>"111111101",
  62760=>"111111111",
  62761=>"111111100",
  62762=>"100100100",
  62763=>"111011000",
  62764=>"011111001",
  62765=>"010010000",
  62766=>"111000111",
  62767=>"000000000",
  62768=>"110110110",
  62769=>"000000000",
  62770=>"110001111",
  62771=>"110110111",
  62772=>"000000000",
  62773=>"000000010",
  62774=>"111000110",
  62775=>"000111111",
  62776=>"000010000",
  62777=>"111000111",
  62778=>"000101111",
  62779=>"110111111",
  62780=>"000000000",
  62781=>"000000000",
  62782=>"000111011",
  62783=>"000000000",
  62784=>"000000000",
  62785=>"111111000",
  62786=>"110111111",
  62787=>"011001001",
  62788=>"111111111",
  62789=>"111111111",
  62790=>"000000110",
  62791=>"001000000",
  62792=>"000000000",
  62793=>"111111111",
  62794=>"111110111",
  62795=>"111111100",
  62796=>"000000000",
  62797=>"100000111",
  62798=>"111111111",
  62799=>"011000000",
  62800=>"000000000",
  62801=>"111111111",
  62802=>"111111111",
  62803=>"000000110",
  62804=>"011011000",
  62805=>"011011011",
  62806=>"000000000",
  62807=>"000100000",
  62808=>"110110100",
  62809=>"000000000",
  62810=>"110110000",
  62811=>"000000000",
  62812=>"010111111",
  62813=>"000000000",
  62814=>"000000000",
  62815=>"111111111",
  62816=>"000000000",
  62817=>"011111110",
  62818=>"001010000",
  62819=>"111111111",
  62820=>"001001001",
  62821=>"000000000",
  62822=>"111111111",
  62823=>"011011111",
  62824=>"011111001",
  62825=>"111111111",
  62826=>"000000000",
  62827=>"000000000",
  62828=>"101101111",
  62829=>"000000001",
  62830=>"111011000",
  62831=>"111111111",
  62832=>"100000000",
  62833=>"000000000",
  62834=>"001111111",
  62835=>"111011011",
  62836=>"100111110",
  62837=>"111111111",
  62838=>"000000000",
  62839=>"000000111",
  62840=>"000000000",
  62841=>"000000000",
  62842=>"000000000",
  62843=>"000010000",
  62844=>"111111111",
  62845=>"111110111",
  62846=>"000000000",
  62847=>"000000000",
  62848=>"001111011",
  62849=>"110100001",
  62850=>"000100000",
  62851=>"000000001",
  62852=>"000000111",
  62853=>"111111000",
  62854=>"111011011",
  62855=>"111111111",
  62856=>"000000000",
  62857=>"000000000",
  62858=>"110000111",
  62859=>"010011010",
  62860=>"001000000",
  62861=>"001001000",
  62862=>"110111010",
  62863=>"011011000",
  62864=>"000000011",
  62865=>"111111000",
  62866=>"010110111",
  62867=>"000100000",
  62868=>"000000111",
  62869=>"000000000",
  62870=>"110000001",
  62871=>"110100000",
  62872=>"111100111",
  62873=>"000100100",
  62874=>"011000000",
  62875=>"000000000",
  62876=>"000100100",
  62877=>"111111111",
  62878=>"000010000",
  62879=>"100000000",
  62880=>"111111111",
  62881=>"000000000",
  62882=>"011000000",
  62883=>"111111111",
  62884=>"111111111",
  62885=>"000000000",
  62886=>"101111111",
  62887=>"000000000",
  62888=>"110110100",
  62889=>"000000100",
  62890=>"000000000",
  62891=>"000000000",
  62892=>"000110000",
  62893=>"111100110",
  62894=>"010000000",
  62895=>"111111111",
  62896=>"000000000",
  62897=>"000001000",
  62898=>"111111111",
  62899=>"000111111",
  62900=>"011000000",
  62901=>"111111111",
  62902=>"011001101",
  62903=>"011111100",
  62904=>"110111111",
  62905=>"111111000",
  62906=>"101100110",
  62907=>"110011011",
  62908=>"000011111",
  62909=>"111011000",
  62910=>"000000000",
  62911=>"111011001",
  62912=>"111111111",
  62913=>"000000000",
  62914=>"111111111",
  62915=>"000000000",
  62916=>"000000110",
  62917=>"000000100",
  62918=>"000000000",
  62919=>"111111001",
  62920=>"011011000",
  62921=>"000000000",
  62922=>"111000001",
  62923=>"111111010",
  62924=>"111111000",
  62925=>"100100000",
  62926=>"000000000",
  62927=>"111100000",
  62928=>"000000000",
  62929=>"111111111",
  62930=>"111111000",
  62931=>"100100111",
  62932=>"000000000",
  62933=>"000000000",
  62934=>"000000110",
  62935=>"110000100",
  62936=>"000000111",
  62937=>"000111110",
  62938=>"000000000",
  62939=>"110111111",
  62940=>"000000000",
  62941=>"000000000",
  62942=>"101101101",
  62943=>"001001001",
  62944=>"000000000",
  62945=>"110000010",
  62946=>"110111111",
  62947=>"100000110",
  62948=>"000000000",
  62949=>"111111110",
  62950=>"000000000",
  62951=>"000000000",
  62952=>"111111111",
  62953=>"000000000",
  62954=>"110110010",
  62955=>"101101000",
  62956=>"111111111",
  62957=>"011000000",
  62958=>"111111101",
  62959=>"000000000",
  62960=>"000000000",
  62961=>"000000000",
  62962=>"000000000",
  62963=>"111000000",
  62964=>"011000000",
  62965=>"000000000",
  62966=>"111000000",
  62967=>"110100111",
  62968=>"111000000",
  62969=>"000000000",
  62970=>"001101111",
  62971=>"000000000",
  62972=>"111001111",
  62973=>"111000101",
  62974=>"000000000",
  62975=>"100111111",
  62976=>"000000000",
  62977=>"000000001",
  62978=>"111011111",
  62979=>"110110100",
  62980=>"110110000",
  62981=>"000000100",
  62982=>"100100111",
  62983=>"011111111",
  62984=>"111110111",
  62985=>"010110010",
  62986=>"000110001",
  62987=>"111000000",
  62988=>"001001011",
  62989=>"000000001",
  62990=>"110110111",
  62991=>"000000111",
  62992=>"000000000",
  62993=>"000100111",
  62994=>"001111111",
  62995=>"001100101",
  62996=>"000000001",
  62997=>"001000111",
  62998=>"010110111",
  62999=>"000001101",
  63000=>"011011011",
  63001=>"001001011",
  63002=>"101101101",
  63003=>"000001111",
  63004=>"000000000",
  63005=>"100110110",
  63006=>"100000000",
  63007=>"101101001",
  63008=>"000000000",
  63009=>"001000000",
  63010=>"000001111",
  63011=>"110010000",
  63012=>"111111111",
  63013=>"000000000",
  63014=>"111100000",
  63015=>"000000000",
  63016=>"000000001",
  63017=>"000000000",
  63018=>"000000000",
  63019=>"111000000",
  63020=>"000000100",
  63021=>"100101101",
  63022=>"111001000",
  63023=>"000100100",
  63024=>"111000000",
  63025=>"000000000",
  63026=>"011000001",
  63027=>"100101111",
  63028=>"001001000",
  63029=>"110110000",
  63030=>"101101101",
  63031=>"000000010",
  63032=>"100110111",
  63033=>"000000001",
  63034=>"000000100",
  63035=>"011001111",
  63036=>"111111000",
  63037=>"111111111",
  63038=>"110110110",
  63039=>"000000000",
  63040=>"000000111",
  63041=>"111111111",
  63042=>"101111111",
  63043=>"111111111",
  63044=>"010000000",
  63045=>"001001001",
  63046=>"001000111",
  63047=>"111111111",
  63048=>"000100000",
  63049=>"111101110",
  63050=>"111111111",
  63051=>"011000000",
  63052=>"001000000",
  63053=>"101001001",
  63054=>"011001100",
  63055=>"000000101",
  63056=>"000111111",
  63057=>"101101111",
  63058=>"000000001",
  63059=>"010001001",
  63060=>"101001001",
  63061=>"111111111",
  63062=>"000000001",
  63063=>"000000000",
  63064=>"001000001",
  63065=>"001101001",
  63066=>"110110111",
  63067=>"000000100",
  63068=>"010000000",
  63069=>"111101101",
  63070=>"111111110",
  63071=>"001001011",
  63072=>"111111011",
  63073=>"101001101",
  63074=>"010000010",
  63075=>"000000000",
  63076=>"000000110",
  63077=>"101001111",
  63078=>"000010100",
  63079=>"101111111",
  63080=>"000001001",
  63081=>"111101000",
  63082=>"101100111",
  63083=>"111111101",
  63084=>"010011111",
  63085=>"000001011",
  63086=>"110110110",
  63087=>"000000000",
  63088=>"001000010",
  63089=>"010110111",
  63090=>"111111011",
  63091=>"000010110",
  63092=>"000000000",
  63093=>"000000100",
  63094=>"000000000",
  63095=>"001000101",
  63096=>"111101000",
  63097=>"000111111",
  63098=>"101000000",
  63099=>"001000111",
  63100=>"110110100",
  63101=>"110110000",
  63102=>"101001001",
  63103=>"001001000",
  63104=>"110110010",
  63105=>"001101111",
  63106=>"111101000",
  63107=>"110000010",
  63108=>"100100101",
  63109=>"101101101",
  63110=>"010000110",
  63111=>"111111111",
  63112=>"011001101",
  63113=>"111111010",
  63114=>"111111001",
  63115=>"111011111",
  63116=>"000001111",
  63117=>"000001000",
  63118=>"000000000",
  63119=>"010000111",
  63120=>"000010111",
  63121=>"000000000",
  63122=>"111011111",
  63123=>"000000000",
  63124=>"111001001",
  63125=>"111110111",
  63126=>"111111101",
  63127=>"111111000",
  63128=>"101001101",
  63129=>"000000000",
  63130=>"110100110",
  63131=>"000000000",
  63132=>"001000110",
  63133=>"111111110",
  63134=>"111111111",
  63135=>"000100111",
  63136=>"111001000",
  63137=>"011001001",
  63138=>"000000000",
  63139=>"111111110",
  63140=>"001001011",
  63141=>"100001111",
  63142=>"111111000",
  63143=>"110110000",
  63144=>"110000000",
  63145=>"001001000",
  63146=>"110110110",
  63147=>"000000010",
  63148=>"111100000",
  63149=>"101100110",
  63150=>"000000001",
  63151=>"000100111",
  63152=>"000000111",
  63153=>"100110111",
  63154=>"100100101",
  63155=>"111111000",
  63156=>"001101101",
  63157=>"000000000",
  63158=>"110101000",
  63159=>"000000000",
  63160=>"000000011",
  63161=>"000101111",
  63162=>"000000100",
  63163=>"000001011",
  63164=>"111001001",
  63165=>"100101111",
  63166=>"001010000",
  63167=>"100100000",
  63168=>"110110100",
  63169=>"011111101",
  63170=>"011111110",
  63171=>"101111111",
  63172=>"011010110",
  63173=>"000000000",
  63174=>"010010010",
  63175=>"001001001",
  63176=>"001001001",
  63177=>"111110111",
  63178=>"010010111",
  63179=>"101111111",
  63180=>"110000000",
  63181=>"101100110",
  63182=>"111111111",
  63183=>"101101111",
  63184=>"111110100",
  63185=>"000000000",
  63186=>"111111111",
  63187=>"000000000",
  63188=>"010010000",
  63189=>"001101001",
  63190=>"010010000",
  63191=>"001001101",
  63192=>"001001000",
  63193=>"111110110",
  63194=>"000000000",
  63195=>"011111111",
  63196=>"111100000",
  63197=>"111111111",
  63198=>"111011111",
  63199=>"011011111",
  63200=>"100111011",
  63201=>"000000011",
  63202=>"010011111",
  63203=>"111111000",
  63204=>"000000000",
  63205=>"001001001",
  63206=>"111111111",
  63207=>"111111111",
  63208=>"110110111",
  63209=>"101101001",
  63210=>"000000000",
  63211=>"000000001",
  63212=>"011011000",
  63213=>"111000000",
  63214=>"110111101",
  63215=>"111111010",
  63216=>"101001001",
  63217=>"111111000",
  63218=>"101101111",
  63219=>"010111111",
  63220=>"110000111",
  63221=>"110110110",
  63222=>"100000000",
  63223=>"000100111",
  63224=>"111111111",
  63225=>"000000000",
  63226=>"100000000",
  63227=>"010011111",
  63228=>"110111110",
  63229=>"100000000",
  63230=>"000000001",
  63231=>"110100110",
  63232=>"000000000",
  63233=>"011011011",
  63234=>"000011111",
  63235=>"111111111",
  63236=>"111111010",
  63237=>"111110010",
  63238=>"110110101",
  63239=>"110010000",
  63240=>"001000000",
  63241=>"111111101",
  63242=>"111101001",
  63243=>"110111111",
  63244=>"010000000",
  63245=>"001000010",
  63246=>"111111000",
  63247=>"000000111",
  63248=>"000100100",
  63249=>"110110010",
  63250=>"111001000",
  63251=>"011001111",
  63252=>"001101000",
  63253=>"111111111",
  63254=>"001001101",
  63255=>"110111010",
  63256=>"000000000",
  63257=>"111001000",
  63258=>"111111111",
  63259=>"101111111",
  63260=>"000000110",
  63261=>"010000000",
  63262=>"000000000",
  63263=>"000000010",
  63264=>"000100111",
  63265=>"001111011",
  63266=>"111111111",
  63267=>"111101101",
  63268=>"000111111",
  63269=>"110110111",
  63270=>"111111110",
  63271=>"011001001",
  63272=>"110010111",
  63273=>"000010011",
  63274=>"111100000",
  63275=>"111111111",
  63276=>"000000000",
  63277=>"000001000",
  63278=>"110010000",
  63279=>"111110000",
  63280=>"001000000",
  63281=>"110110010",
  63282=>"000110110",
  63283=>"110010011",
  63284=>"010010000",
  63285=>"011011011",
  63286=>"101001000",
  63287=>"000101111",
  63288=>"100110110",
  63289=>"101101000",
  63290=>"000000000",
  63291=>"111101100",
  63292=>"110010000",
  63293=>"001111110",
  63294=>"000010111",
  63295=>"100010000",
  63296=>"001000001",
  63297=>"001000100",
  63298=>"110000000",
  63299=>"111000011",
  63300=>"000000001",
  63301=>"000111111",
  63302=>"110111111",
  63303=>"000000000",
  63304=>"000000000",
  63305=>"001101000",
  63306=>"110001000",
  63307=>"101001001",
  63308=>"111101111",
  63309=>"110111111",
  63310=>"001001111",
  63311=>"110110100",
  63312=>"000000000",
  63313=>"000001011",
  63314=>"000101111",
  63315=>"010000000",
  63316=>"110111010",
  63317=>"011011000",
  63318=>"000000111",
  63319=>"000000000",
  63320=>"010000000",
  63321=>"011111111",
  63322=>"100111111",
  63323=>"111000000",
  63324=>"111111010",
  63325=>"001001001",
  63326=>"110110010",
  63327=>"111111011",
  63328=>"110001000",
  63329=>"111111111",
  63330=>"001000001",
  63331=>"111111010",
  63332=>"010011111",
  63333=>"000000000",
  63334=>"000000100",
  63335=>"111101101",
  63336=>"001000101",
  63337=>"100010010",
  63338=>"111110111",
  63339=>"001001001",
  63340=>"000001001",
  63341=>"001001110",
  63342=>"110110110",
  63343=>"000000000",
  63344=>"000000000",
  63345=>"111111111",
  63346=>"000000000",
  63347=>"000111111",
  63348=>"111101101",
  63349=>"000000000",
  63350=>"111000000",
  63351=>"011000000",
  63352=>"000000000",
  63353=>"000000011",
  63354=>"001110110",
  63355=>"000101000",
  63356=>"101000000",
  63357=>"101101111",
  63358=>"110111111",
  63359=>"000000111",
  63360=>"011011111",
  63361=>"111101011",
  63362=>"110100100",
  63363=>"111111111",
  63364=>"110110111",
  63365=>"110111111",
  63366=>"000001000",
  63367=>"011011101",
  63368=>"110110010",
  63369=>"011001011",
  63370=>"001101101",
  63371=>"101000010",
  63372=>"111111011",
  63373=>"100100100",
  63374=>"110000010",
  63375=>"000000001",
  63376=>"000000000",
  63377=>"000000001",
  63378=>"000000000",
  63379=>"000110100",
  63380=>"000000000",
  63381=>"010010000",
  63382=>"011001000",
  63383=>"001001001",
  63384=>"001001000",
  63385=>"001001110",
  63386=>"101001111",
  63387=>"111000000",
  63388=>"101101001",
  63389=>"101100000",
  63390=>"000000001",
  63391=>"101101101",
  63392=>"000001111",
  63393=>"011111011",
  63394=>"111100000",
  63395=>"010000001",
  63396=>"000000000",
  63397=>"000010000",
  63398=>"111011000",
  63399=>"111001000",
  63400=>"000001001",
  63401=>"000000000",
  63402=>"010011000",
  63403=>"111111111",
  63404=>"010110111",
  63405=>"011111111",
  63406=>"010000000",
  63407=>"000000010",
  63408=>"001001101",
  63409=>"001001110",
  63410=>"011011001",
  63411=>"111101111",
  63412=>"000000111",
  63413=>"111111111",
  63414=>"000110110",
  63415=>"001000000",
  63416=>"111101111",
  63417=>"111111110",
  63418=>"010010011",
  63419=>"010110110",
  63420=>"101101001",
  63421=>"110110100",
  63422=>"111101101",
  63423=>"000000100",
  63424=>"001000111",
  63425=>"000000001",
  63426=>"101001001",
  63427=>"000101111",
  63428=>"000000000",
  63429=>"110110000",
  63430=>"001101111",
  63431=>"111111101",
  63432=>"100100000",
  63433=>"000000000",
  63434=>"000000000",
  63435=>"010111010",
  63436=>"111001111",
  63437=>"111111110",
  63438=>"001001000",
  63439=>"110111010",
  63440=>"011000000",
  63441=>"100111111",
  63442=>"011110111",
  63443=>"100000001",
  63444=>"111100000",
  63445=>"111111111",
  63446=>"000000000",
  63447=>"000100100",
  63448=>"101000000",
  63449=>"111111100",
  63450=>"010000000",
  63451=>"000010010",
  63452=>"110111111",
  63453=>"110110111",
  63454=>"111000000",
  63455=>"011011111",
  63456=>"111111001",
  63457=>"000000110",
  63458=>"111101111",
  63459=>"111111100",
  63460=>"111111000",
  63461=>"110110010",
  63462=>"100000000",
  63463=>"111111001",
  63464=>"011011011",
  63465=>"100010111",
  63466=>"010011010",
  63467=>"111111011",
  63468=>"100000000",
  63469=>"001001001",
  63470=>"110110010",
  63471=>"111001100",
  63472=>"111111101",
  63473=>"111111111",
  63474=>"111110110",
  63475=>"000010111",
  63476=>"000000111",
  63477=>"111100000",
  63478=>"111111110",
  63479=>"111110000",
  63480=>"001111011",
  63481=>"000000001",
  63482=>"000110111",
  63483=>"101101111",
  63484=>"111010000",
  63485=>"111111111",
  63486=>"011011111",
  63487=>"001001111",
  63488=>"111111011",
  63489=>"111111010",
  63490=>"000000000",
  63491=>"100111111",
  63492=>"010010011",
  63493=>"110100000",
  63494=>"111011111",
  63495=>"000000000",
  63496=>"111101000",
  63497=>"101000100",
  63498=>"111110000",
  63499=>"001111111",
  63500=>"000110110",
  63501=>"011111000",
  63502=>"010111111",
  63503=>"111111111",
  63504=>"110011011",
  63505=>"111111111",
  63506=>"101100000",
  63507=>"100111111",
  63508=>"010111011",
  63509=>"111100100",
  63510=>"010110111",
  63511=>"111110101",
  63512=>"010011011",
  63513=>"100000001",
  63514=>"000000000",
  63515=>"111111000",
  63516=>"000000000",
  63517=>"111110010",
  63518=>"011001000",
  63519=>"111001111",
  63520=>"000111011",
  63521=>"000110100",
  63522=>"110111000",
  63523=>"010110010",
  63524=>"111111111",
  63525=>"111111111",
  63526=>"011111111",
  63527=>"000110101",
  63528=>"000110000",
  63529=>"000000000",
  63530=>"011011000",
  63531=>"000000000",
  63532=>"000000001",
  63533=>"000000010",
  63534=>"000001001",
  63535=>"101111111",
  63536=>"000000000",
  63537=>"111111111",
  63538=>"111110111",
  63539=>"110110110",
  63540=>"111101000",
  63541=>"111100101",
  63542=>"000011000",
  63543=>"000010000",
  63544=>"110011111",
  63545=>"000010110",
  63546=>"011000000",
  63547=>"100000000",
  63548=>"000000000",
  63549=>"000011111",
  63550=>"000011011",
  63551=>"101101101",
  63552=>"110010010",
  63553=>"000110111",
  63554=>"010010001",
  63555=>"000000000",
  63556=>"111111110",
  63557=>"001111111",
  63558=>"000111011",
  63559=>"000000000",
  63560=>"000000001",
  63561=>"111111010",
  63562=>"000111011",
  63563=>"010111011",
  63564=>"110110100",
  63565=>"100000100",
  63566=>"111111000",
  63567=>"100101100",
  63568=>"001111111",
  63569=>"000110000",
  63570=>"011111111",
  63571=>"110110111",
  63572=>"001101101",
  63573=>"111111111",
  63574=>"000010010",
  63575=>"000100100",
  63576=>"000100100",
  63577=>"000000000",
  63578=>"000000000",
  63579=>"110011110",
  63580=>"111111001",
  63581=>"000001001",
  63582=>"000110000",
  63583=>"110111111",
  63584=>"000000110",
  63585=>"111111010",
  63586=>"000000000",
  63587=>"101100000",
  63588=>"100111000",
  63589=>"011111111",
  63590=>"011011111",
  63591=>"111111100",
  63592=>"110110111",
  63593=>"000000000",
  63594=>"000110111",
  63595=>"001011111",
  63596=>"100000000",
  63597=>"111111111",
  63598=>"111101101",
  63599=>"111111111",
  63600=>"010010111",
  63601=>"000011111",
  63602=>"011011001",
  63603=>"111111111",
  63604=>"011111111",
  63605=>"110010111",
  63606=>"111001001",
  63607=>"000010000",
  63608=>"111111111",
  63609=>"111111110",
  63610=>"111111011",
  63611=>"111111111",
  63612=>"001001001",
  63613=>"000000000",
  63614=>"011111000",
  63615=>"111111011",
  63616=>"100111111",
  63617=>"111111111",
  63618=>"000000000",
  63619=>"000010111",
  63620=>"101100000",
  63621=>"000000000",
  63622=>"000010000",
  63623=>"000000000",
  63624=>"000000000",
  63625=>"011111111",
  63626=>"001101101",
  63627=>"000000000",
  63628=>"011111111",
  63629=>"101111000",
  63630=>"000111000",
  63631=>"011111111",
  63632=>"111111000",
  63633=>"000000100",
  63634=>"100111111",
  63635=>"111111111",
  63636=>"001011001",
  63637=>"111111101",
  63638=>"000100000",
  63639=>"000000000",
  63640=>"010000101",
  63641=>"000110000",
  63642=>"010000010",
  63643=>"111011000",
  63644=>"000000000",
  63645=>"111111110",
  63646=>"000000000",
  63647=>"000000000",
  63648=>"111010011",
  63649=>"000010010",
  63650=>"111111110",
  63651=>"100000000",
  63652=>"110110110",
  63653=>"011010111",
  63654=>"000000000",
  63655=>"111001001",
  63656=>"000000000",
  63657=>"101001001",
  63658=>"111101111",
  63659=>"100100111",
  63660=>"010011011",
  63661=>"000001001",
  63662=>"000010000",
  63663=>"000000100",
  63664=>"000000000",
  63665=>"001101111",
  63666=>"000000000",
  63667=>"000000000",
  63668=>"111111111",
  63669=>"010010000",
  63670=>"111111111",
  63671=>"111110100",
  63672=>"000111111",
  63673=>"000000000",
  63674=>"000000111",
  63675=>"000111111",
  63676=>"000101001",
  63677=>"010110000",
  63678=>"000110000",
  63679=>"111111111",
  63680=>"000000000",
  63681=>"011111011",
  63682=>"001000000",
  63683=>"000000000",
  63684=>"101101000",
  63685=>"000000010",
  63686=>"010110010",
  63687=>"111111111",
  63688=>"000000000",
  63689=>"111111111",
  63690=>"000000000",
  63691=>"001111111",
  63692=>"010011010",
  63693=>"001000000",
  63694=>"011111111",
  63695=>"111111111",
  63696=>"111110100",
  63697=>"011011001",
  63698=>"111111000",
  63699=>"111111111",
  63700=>"100000101",
  63701=>"100111111",
  63702=>"000000000",
  63703=>"010011000",
  63704=>"000000000",
  63705=>"000000000",
  63706=>"000111111",
  63707=>"001000000",
  63708=>"000000001",
  63709=>"000010000",
  63710=>"101111111",
  63711=>"001111001",
  63712=>"101011001",
  63713=>"000000011",
  63714=>"000000010",
  63715=>"100110010",
  63716=>"111111101",
  63717=>"011110110",
  63718=>"010011011",
  63719=>"111111000",
  63720=>"000000011",
  63721=>"101010000",
  63722=>"111011001",
  63723=>"111111111",
  63724=>"010010011",
  63725=>"111110111",
  63726=>"101100000",
  63727=>"000000000",
  63728=>"111110000",
  63729=>"111110100",
  63730=>"000000111",
  63731=>"110110110",
  63732=>"000100111",
  63733=>"111011111",
  63734=>"000011111",
  63735=>"000000000",
  63736=>"110000000",
  63737=>"101100000",
  63738=>"000000111",
  63739=>"010111000",
  63740=>"111111111",
  63741=>"000000000",
  63742=>"111111111",
  63743=>"111111110",
  63744=>"000000111",
  63745=>"001001000",
  63746=>"000000000",
  63747=>"111111110",
  63748=>"010010010",
  63749=>"000010000",
  63750=>"000010000",
  63751=>"000111000",
  63752=>"110110011",
  63753=>"000000000",
  63754=>"100001000",
  63755=>"000000000",
  63756=>"000000000",
  63757=>"000100010",
  63758=>"000000000",
  63759=>"000011000",
  63760=>"101000000",
  63761=>"000010111",
  63762=>"000000000",
  63763=>"000011011",
  63764=>"111111111",
  63765=>"000000001",
  63766=>"111111111",
  63767=>"111111111",
  63768=>"111111000",
  63769=>"111001001",
  63770=>"001001001",
  63771=>"000000000",
  63772=>"001001011",
  63773=>"111000000",
  63774=>"011001000",
  63775=>"101111110",
  63776=>"010011100",
  63777=>"000000000",
  63778=>"110111101",
  63779=>"110111010",
  63780=>"000110000",
  63781=>"111111011",
  63782=>"010111010",
  63783=>"111111111",
  63784=>"001010000",
  63785=>"111111111",
  63786=>"000010000",
  63787=>"111011011",
  63788=>"111111111",
  63789=>"001000100",
  63790=>"000000000",
  63791=>"111111111",
  63792=>"000111001",
  63793=>"111111101",
  63794=>"000000000",
  63795=>"001111111",
  63796=>"000000000",
  63797=>"000100000",
  63798=>"100000000",
  63799=>"000001000",
  63800=>"000000010",
  63801=>"000010000",
  63802=>"111111111",
  63803=>"000000111",
  63804=>"001011001",
  63805=>"000000010",
  63806=>"111011101",
  63807=>"000011000",
  63808=>"000001001",
  63809=>"000010000",
  63810=>"000000111",
  63811=>"000011000",
  63812=>"011111001",
  63813=>"000000000",
  63814=>"011011011",
  63815=>"011001001",
  63816=>"000101101",
  63817=>"000010000",
  63818=>"010010010",
  63819=>"010110000",
  63820=>"000111110",
  63821=>"010111111",
  63822=>"111111111",
  63823=>"100110100",
  63824=>"111101001",
  63825=>"000101010",
  63826=>"111110110",
  63827=>"111111010",
  63828=>"110000010",
  63829=>"001000111",
  63830=>"111111010",
  63831=>"011011111",
  63832=>"000000000",
  63833=>"000000000",
  63834=>"000000101",
  63835=>"010010000",
  63836=>"100000010",
  63837=>"111111111",
  63838=>"100000000",
  63839=>"011011011",
  63840=>"111111000",
  63841=>"111011111",
  63842=>"010010010",
  63843=>"000000000",
  63844=>"011001001",
  63845=>"000001001",
  63846=>"100000000",
  63847=>"000000000",
  63848=>"011011000",
  63849=>"000110000",
  63850=>"111111000",
  63851=>"000101000",
  63852=>"111011011",
  63853=>"010010000",
  63854=>"111111110",
  63855=>"000000000",
  63856=>"010011111",
  63857=>"111000001",
  63858=>"000000100",
  63859=>"100110110",
  63860=>"000000111",
  63861=>"000000000",
  63862=>"111100100",
  63863=>"111111111",
  63864=>"001111111",
  63865=>"111111111",
  63866=>"001000000",
  63867=>"000000000",
  63868=>"110101101",
  63869=>"010011011",
  63870=>"000000000",
  63871=>"111111110",
  63872=>"001001001",
  63873=>"110110110",
  63874=>"111111111",
  63875=>"000111011",
  63876=>"110110110",
  63877=>"000000000",
  63878=>"111111000",
  63879=>"010011010",
  63880=>"000010000",
  63881=>"111100011",
  63882=>"001010000",
  63883=>"000000000",
  63884=>"111100001",
  63885=>"100011111",
  63886=>"111111100",
  63887=>"000000001",
  63888=>"000000100",
  63889=>"000000000",
  63890=>"001000000",
  63891=>"111001100",
  63892=>"011010000",
  63893=>"111111111",
  63894=>"000000010",
  63895=>"000000111",
  63896=>"010111111",
  63897=>"111011010",
  63898=>"000000000",
  63899=>"000111001",
  63900=>"101100111",
  63901=>"111111100",
  63902=>"100100100",
  63903=>"111111111",
  63904=>"111111111",
  63905=>"111001001",
  63906=>"000100000",
  63907=>"000111111",
  63908=>"000010000",
  63909=>"000000000",
  63910=>"000000000",
  63911=>"100111000",
  63912=>"111111001",
  63913=>"000000001",
  63914=>"000000000",
  63915=>"000000000",
  63916=>"010110111",
  63917=>"000110111",
  63918=>"000001011",
  63919=>"101000000",
  63920=>"000000010",
  63921=>"000000000",
  63922=>"010000000",
  63923=>"111001111",
  63924=>"000010000",
  63925=>"000010000",
  63926=>"000010000",
  63927=>"111101101",
  63928=>"000000000",
  63929=>"000000101",
  63930=>"101000111",
  63931=>"000110000",
  63932=>"111111110",
  63933=>"000000000",
  63934=>"110111000",
  63935=>"000001000",
  63936=>"000000000",
  63937=>"000000000",
  63938=>"000000000",
  63939=>"000000000",
  63940=>"000000000",
  63941=>"000110111",
  63942=>"000111111",
  63943=>"111111000",
  63944=>"010000000",
  63945=>"011000101",
  63946=>"111111111",
  63947=>"000000000",
  63948=>"000000000",
  63949=>"000000000",
  63950=>"010000000",
  63951=>"111000000",
  63952=>"111111010",
  63953=>"000110100",
  63954=>"011111111",
  63955=>"111101101",
  63956=>"110111111",
  63957=>"100100110",
  63958=>"000111101",
  63959=>"011011111",
  63960=>"000010000",
  63961=>"000000000",
  63962=>"110101101",
  63963=>"111111111",
  63964=>"101101100",
  63965=>"001111111",
  63966=>"000111000",
  63967=>"111111111",
  63968=>"000001001",
  63969=>"111111111",
  63970=>"000010010",
  63971=>"000000000",
  63972=>"000110111",
  63973=>"111111111",
  63974=>"000111010",
  63975=>"000100101",
  63976=>"010011011",
  63977=>"001111011",
  63978=>"110010000",
  63979=>"000000000",
  63980=>"011111000",
  63981=>"001000000",
  63982=>"101101001",
  63983=>"110110000",
  63984=>"111101101",
  63985=>"000000000",
  63986=>"011001000",
  63987=>"000000000",
  63988=>"111101001",
  63989=>"101111111",
  63990=>"010111000",
  63991=>"011011011",
  63992=>"000000000",
  63993=>"100100100",
  63994=>"111001001",
  63995=>"010000000",
  63996=>"000011000",
  63997=>"111011001",
  63998=>"000010001",
  63999=>"111111111",
  64000=>"111000000",
  64001=>"000000111",
  64002=>"000000000",
  64003=>"000000000",
  64004=>"011011011",
  64005=>"000000000",
  64006=>"011111001",
  64007=>"111111000",
  64008=>"111111101",
  64009=>"110011011",
  64010=>"001001111",
  64011=>"110000000",
  64012=>"111101001",
  64013=>"101111111",
  64014=>"000000111",
  64015=>"111111100",
  64016=>"100111000",
  64017=>"111111111",
  64018=>"111111000",
  64019=>"000000000",
  64020=>"000000111",
  64021=>"000000000",
  64022=>"111111111",
  64023=>"000100110",
  64024=>"001111111",
  64025=>"001000000",
  64026=>"110110111",
  64027=>"011011111",
  64028=>"111111111",
  64029=>"000001111",
  64030=>"010110110",
  64031=>"001111111",
  64032=>"110111111",
  64033=>"111110000",
  64034=>"111110111",
  64035=>"011011111",
  64036=>"111111101",
  64037=>"001000000",
  64038=>"111111110",
  64039=>"000000111",
  64040=>"000010010",
  64041=>"111111111",
  64042=>"001000111",
  64043=>"101111111",
  64044=>"000000100",
  64045=>"111111000",
  64046=>"010000000",
  64047=>"111111011",
  64048=>"111111111",
  64049=>"111111000",
  64050=>"100000100",
  64051=>"111000000",
  64052=>"110111111",
  64053=>"111110100",
  64054=>"001001000",
  64055=>"000000000",
  64056=>"000000111",
  64057=>"111000111",
  64058=>"001000000",
  64059=>"100000111",
  64060=>"000010111",
  64061=>"111111001",
  64062=>"000000001",
  64063=>"111111000",
  64064=>"000000000",
  64065=>"000000001",
  64066=>"001000000",
  64067=>"000000111",
  64068=>"001000110",
  64069=>"000000000",
  64070=>"000000111",
  64071=>"111111111",
  64072=>"111000000",
  64073=>"000000111",
  64074=>"111100010",
  64075=>"000000010",
  64076=>"100111111",
  64077=>"111111111",
  64078=>"100110111",
  64079=>"000000101",
  64080=>"000010111",
  64081=>"111111110",
  64082=>"111111110",
  64083=>"111111100",
  64084=>"001001000",
  64085=>"000010111",
  64086=>"101111110",
  64087=>"000111111",
  64088=>"111111111",
  64089=>"111111111",
  64090=>"110110111",
  64091=>"110100110",
  64092=>"000000000",
  64093=>"111111000",
  64094=>"001101110",
  64095=>"001001001",
  64096=>"000111111",
  64097=>"000000000",
  64098=>"111011111",
  64099=>"111000000",
  64100=>"000000000",
  64101=>"000000001",
  64102=>"100010110",
  64103=>"000101100",
  64104=>"000000000",
  64105=>"000000000",
  64106=>"000000000",
  64107=>"111000000",
  64108=>"110110100",
  64109=>"111111111",
  64110=>"111111111",
  64111=>"111111010",
  64112=>"000001000",
  64113=>"001001100",
  64114=>"101111101",
  64115=>"111110000",
  64116=>"000010111",
  64117=>"111111110",
  64118=>"000000000",
  64119=>"101001111",
  64120=>"001001000",
  64121=>"011111000",
  64122=>"000000000",
  64123=>"000000001",
  64124=>"110100100",
  64125=>"110010000",
  64126=>"000000000",
  64127=>"000000000",
  64128=>"000111111",
  64129=>"000000100",
  64130=>"101000000",
  64131=>"110010000",
  64132=>"000001111",
  64133=>"011001111",
  64134=>"000000000",
  64135=>"110110111",
  64136=>"111111111",
  64137=>"000000000",
  64138=>"000000000",
  64139=>"000000000",
  64140=>"100111111",
  64141=>"000000000",
  64142=>"111111000",
  64143=>"000000111",
  64144=>"000111111",
  64145=>"000000000",
  64146=>"100000000",
  64147=>"100110111",
  64148=>"000111111",
  64149=>"111111110",
  64150=>"111111100",
  64151=>"100000000",
  64152=>"000000000",
  64153=>"000000000",
  64154=>"111111110",
  64155=>"011111000",
  64156=>"111100110",
  64157=>"111110111",
  64158=>"111111111",
  64159=>"000000110",
  64160=>"000000000",
  64161=>"000000111",
  64162=>"001000000",
  64163=>"110110111",
  64164=>"111110010",
  64165=>"111111101",
  64166=>"111111110",
  64167=>"111110000",
  64168=>"000111111",
  64169=>"111111010",
  64170=>"000111111",
  64171=>"000110110",
  64172=>"001011001",
  64173=>"000110110",
  64174=>"011001000",
  64175=>"000111111",
  64176=>"000111111",
  64177=>"111111000",
  64178=>"011111010",
  64179=>"111111100",
  64180=>"000000000",
  64181=>"110111000",
  64182=>"101111011",
  64183=>"110110111",
  64184=>"111101110",
  64185=>"111111110",
  64186=>"001001001",
  64187=>"100100111",
  64188=>"001111111",
  64189=>"110110010",
  64190=>"100100100",
  64191=>"111000000",
  64192=>"000000000",
  64193=>"001101111",
  64194=>"101111000",
  64195=>"000000011",
  64196=>"110110110",
  64197=>"001000011",
  64198=>"111111010",
  64199=>"000000000",
  64200=>"000000111",
  64201=>"000001111",
  64202=>"111111111",
  64203=>"111100001",
  64204=>"000000000",
  64205=>"101111111",
  64206=>"001110111",
  64207=>"011101111",
  64208=>"000000011",
  64209=>"000010111",
  64210=>"111111111",
  64211=>"010000111",
  64212=>"100111110",
  64213=>"111110110",
  64214=>"000100101",
  64215=>"001111000",
  64216=>"000000000",
  64217=>"111100101",
  64218=>"111111111",
  64219=>"110111001",
  64220=>"110101100",
  64221=>"000000011",
  64222=>"111111111",
  64223=>"000000000",
  64224=>"000000001",
  64225=>"000001111",
  64226=>"001101111",
  64227=>"110100000",
  64228=>"100000000",
  64229=>"001000111",
  64230=>"111111111",
  64231=>"111111111",
  64232=>"101000100",
  64233=>"011000010",
  64234=>"110100101",
  64235=>"000100111",
  64236=>"110000010",
  64237=>"000000101",
  64238=>"110111111",
  64239=>"101111111",
  64240=>"101000000",
  64241=>"111010000",
  64242=>"111111111",
  64243=>"001001001",
  64244=>"001100111",
  64245=>"100000001",
  64246=>"000001111",
  64247=>"000000001",
  64248=>"011111111",
  64249=>"001111101",
  64250=>"111111110",
  64251=>"000101111",
  64252=>"110011000",
  64253=>"000001000",
  64254=>"000000000",
  64255=>"111111100",
  64256=>"111111111",
  64257=>"000000111",
  64258=>"000101001",
  64259=>"000000100",
  64260=>"111111111",
  64261=>"000110111",
  64262=>"111111111",
  64263=>"001000000",
  64264=>"000000000",
  64265=>"111111111",
  64266=>"000000111",
  64267=>"000000000",
  64268=>"000110110",
  64269=>"100111011",
  64270=>"001010110",
  64271=>"000100100",
  64272=>"001101001",
  64273=>"000100111",
  64274=>"100001000",
  64275=>"011000000",
  64276=>"000000010",
  64277=>"111100111",
  64278=>"000000000",
  64279=>"011111000",
  64280=>"111000000",
  64281=>"111111000",
  64282=>"100111110",
  64283=>"111011111",
  64284=>"111010000",
  64285=>"000000001",
  64286=>"000000000",
  64287=>"000100111",
  64288=>"110000001",
  64289=>"111000000",
  64290=>"000001000",
  64291=>"000111111",
  64292=>"010000010",
  64293=>"011111111",
  64294=>"100000111",
  64295=>"011001110",
  64296=>"000010111",
  64297=>"111111111",
  64298=>"000111111",
  64299=>"101001011",
  64300=>"111000000",
  64301=>"000000001",
  64302=>"111111111",
  64303=>"111000111",
  64304=>"111100100",
  64305=>"000000000",
  64306=>"111111111",
  64307=>"000000111",
  64308=>"000000111",
  64309=>"000000000",
  64310=>"000000000",
  64311=>"011001111",
  64312=>"111111111",
  64313=>"000000000",
  64314=>"000000001",
  64315=>"110111111",
  64316=>"000001111",
  64317=>"110010000",
  64318=>"000000000",
  64319=>"000000000",
  64320=>"100110000",
  64321=>"111111110",
  64322=>"100000000",
  64323=>"000001111",
  64324=>"000000000",
  64325=>"000000001",
  64326=>"111111111",
  64327=>"111111101",
  64328=>"000000000",
  64329=>"001000111",
  64330=>"000000000",
  64331=>"100100110",
  64332=>"010111111",
  64333=>"100111110",
  64334=>"111111111",
  64335=>"100101101",
  64336=>"001101100",
  64337=>"000000111",
  64338=>"111111111",
  64339=>"000000001",
  64340=>"111000000",
  64341=>"011001001",
  64342=>"111111111",
  64343=>"111111000",
  64344=>"111111111",
  64345=>"111111111",
  64346=>"111110010",
  64347=>"000000010",
  64348=>"010001001",
  64349=>"000011001",
  64350=>"111111111",
  64351=>"110100000",
  64352=>"110111111",
  64353=>"001000000",
  64354=>"100000001",
  64355=>"111111111",
  64356=>"111111111",
  64357=>"001000011",
  64358=>"100000000",
  64359=>"000000001",
  64360=>"111000000",
  64361=>"000000000",
  64362=>"111111111",
  64363=>"000000000",
  64364=>"111111001",
  64365=>"000000000",
  64366=>"001001101",
  64367=>"001001000",
  64368=>"000000100",
  64369=>"111000000",
  64370=>"010000111",
  64371=>"111111011",
  64372=>"111111111",
  64373=>"011001100",
  64374=>"111100111",
  64375=>"000000000",
  64376=>"111111111",
  64377=>"000100111",
  64378=>"000110111",
  64379=>"001011000",
  64380=>"111011000",
  64381=>"011111111",
  64382=>"000100111",
  64383=>"011100111",
  64384=>"101111110",
  64385=>"000010110",
  64386=>"000000110",
  64387=>"000000011",
  64388=>"000000000",
  64389=>"111111111",
  64390=>"000011011",
  64391=>"011010011",
  64392=>"000111111",
  64393=>"111111111",
  64394=>"111111000",
  64395=>"101101111",
  64396=>"111111111",
  64397=>"110111111",
  64398=>"111111010",
  64399=>"000000000",
  64400=>"000000000",
  64401=>"000000000",
  64402=>"100111111",
  64403=>"000000111",
  64404=>"000000000",
  64405=>"000000000",
  64406=>"011000000",
  64407=>"001001100",
  64408=>"000000110",
  64409=>"100111111",
  64410=>"100111000",
  64411=>"111110000",
  64412=>"101111000",
  64413=>"100100000",
  64414=>"000000000",
  64415=>"101100111",
  64416=>"011011000",
  64417=>"111111111",
  64418=>"001000000",
  64419=>"110111111",
  64420=>"000101000",
  64421=>"111111111",
  64422=>"111001000",
  64423=>"101111111",
  64424=>"000000000",
  64425=>"000000001",
  64426=>"100100000",
  64427=>"111111000",
  64428=>"000101111",
  64429=>"111111100",
  64430=>"111000000",
  64431=>"111111111",
  64432=>"101111111",
  64433=>"111000000",
  64434=>"111111101",
  64435=>"011001000",
  64436=>"001000000",
  64437=>"111000000",
  64438=>"111110000",
  64439=>"000100000",
  64440=>"001110111",
  64441=>"000000000",
  64442=>"111100111",
  64443=>"101111111",
  64444=>"000001000",
  64445=>"000000111",
  64446=>"111111111",
  64447=>"000000000",
  64448=>"111111000",
  64449=>"000111001",
  64450=>"000000000",
  64451=>"111111111",
  64452=>"111100101",
  64453=>"000001101",
  64454=>"111000000",
  64455=>"111111001",
  64456=>"111001000",
  64457=>"011000000",
  64458=>"000000111",
  64459=>"000010111",
  64460=>"011111000",
  64461=>"000000000",
  64462=>"000000110",
  64463=>"000000000",
  64464=>"100000000",
  64465=>"000010111",
  64466=>"100100000",
  64467=>"011010011",
  64468=>"001111010",
  64469=>"100100100",
  64470=>"000000011",
  64471=>"101001001",
  64472=>"000000100",
  64473=>"111111111",
  64474=>"101001000",
  64475=>"000000111",
  64476=>"011011000",
  64477=>"111111111",
  64478=>"111111111",
  64479=>"000100110",
  64480=>"000000000",
  64481=>"010011111",
  64482=>"000000000",
  64483=>"110000111",
  64484=>"010000111",
  64485=>"000101111",
  64486=>"100010010",
  64487=>"001000000",
  64488=>"111111111",
  64489=>"111111001",
  64490=>"000111001",
  64491=>"111101000",
  64492=>"111101111",
  64493=>"000000111",
  64494=>"011111111",
  64495=>"011010000",
  64496=>"111111000",
  64497=>"000000111",
  64498=>"000000000",
  64499=>"000111111",
  64500=>"111110110",
  64501=>"000000001",
  64502=>"111000000",
  64503=>"000011011",
  64504=>"000111000",
  64505=>"001000011",
  64506=>"000000101",
  64507=>"100110110",
  64508=>"001000000",
  64509=>"111101100",
  64510=>"111111110",
  64511=>"000000000",
  64512=>"101101100",
  64513=>"000000000",
  64514=>"100000111",
  64515=>"111111111",
  64516=>"111111010",
  64517=>"111000011",
  64518=>"111111111",
  64519=>"111111111",
  64520=>"111111111",
  64521=>"100000000",
  64522=>"001000000",
  64523=>"000111110",
  64524=>"001000000",
  64525=>"100000100",
  64526=>"111000001",
  64527=>"001000000",
  64528=>"000000000",
  64529=>"000000101",
  64530=>"111000001",
  64531=>"001001001",
  64532=>"110111010",
  64533=>"000000000",
  64534=>"001000000",
  64535=>"011110000",
  64536=>"001000111",
  64537=>"001111111",
  64538=>"110000000",
  64539=>"111111000",
  64540=>"100001001",
  64541=>"000001101",
  64542=>"010011011",
  64543=>"111111011",
  64544=>"011110110",
  64545=>"111111010",
  64546=>"011111111",
  64547=>"100110110",
  64548=>"100011011",
  64549=>"000000000",
  64550=>"011010000",
  64551=>"100110111",
  64552=>"000100100",
  64553=>"000111000",
  64554=>"001000110",
  64555=>"000000111",
  64556=>"000100111",
  64557=>"000000010",
  64558=>"000000111",
  64559=>"011111111",
  64560=>"010001000",
  64561=>"000000000",
  64562=>"100100000",
  64563=>"111111111",
  64564=>"000000001",
  64565=>"111110100",
  64566=>"111111101",
  64567=>"000110111",
  64568=>"100000001",
  64569=>"000000100",
  64570=>"001000011",
  64571=>"001101111",
  64572=>"111111100",
  64573=>"111100100",
  64574=>"000000000",
  64575=>"000000001",
  64576=>"000000111",
  64577=>"000000010",
  64578=>"000111111",
  64579=>"111111111",
  64580=>"000000000",
  64581=>"111111110",
  64582=>"100000000",
  64583=>"110111111",
  64584=>"011001000",
  64585=>"100000001",
  64586=>"100000111",
  64587=>"111111010",
  64588=>"011011001",
  64589=>"010010000",
  64590=>"000110111",
  64591=>"110100000",
  64592=>"000000000",
  64593=>"011001001",
  64594=>"000010111",
  64595=>"001000100",
  64596=>"001001111",
  64597=>"111110110",
  64598=>"001000000",
  64599=>"000110110",
  64600=>"011001000",
  64601=>"111000101",
  64602=>"111111100",
  64603=>"110100000",
  64604=>"111111111",
  64605=>"001001001",
  64606=>"110000000",
  64607=>"110000000",
  64608=>"000000000",
  64609=>"111111010",
  64610=>"000000011",
  64611=>"000000000",
  64612=>"000000011",
  64613=>"111111111",
  64614=>"111111000",
  64615=>"000100111",
  64616=>"000011111",
  64617=>"111010010",
  64618=>"111111111",
  64619=>"110111001",
  64620=>"001001010",
  64621=>"010000000",
  64622=>"111111000",
  64623=>"100001000",
  64624=>"010011011",
  64625=>"111011011",
  64626=>"001001111",
  64627=>"101000000",
  64628=>"001000000",
  64629=>"110110110",
  64630=>"100111111",
  64631=>"111111111",
  64632=>"111111111",
  64633=>"001011111",
  64634=>"000000000",
  64635=>"100000100",
  64636=>"000001011",
  64637=>"100100100",
  64638=>"111011000",
  64639=>"011111011",
  64640=>"001000000",
  64641=>"010000000",
  64642=>"000000000",
  64643=>"111111011",
  64644=>"000000001",
  64645=>"000000111",
  64646=>"000000000",
  64647=>"000000000",
  64648=>"001111111",
  64649=>"000000011",
  64650=>"001000000",
  64651=>"111010110",
  64652=>"111111000",
  64653=>"100101111",
  64654=>"000000011",
  64655=>"000000111",
  64656=>"111101111",
  64657=>"111111001",
  64658=>"110100000",
  64659=>"111000000",
  64660=>"111111110",
  64661=>"000111111",
  64662=>"000111111",
  64663=>"111011000",
  64664=>"000000000",
  64665=>"111111011",
  64666=>"000100100",
  64667=>"011111111",
  64668=>"011011011",
  64669=>"110100111",
  64670=>"110001000",
  64671=>"111111111",
  64672=>"111111111",
  64673=>"111111111",
  64674=>"111111111",
  64675=>"000000000",
  64676=>"010000000",
  64677=>"111111111",
  64678=>"000011000",
  64679=>"000111111",
  64680=>"110000000",
  64681=>"001000000",
  64682=>"111111000",
  64683=>"000000000",
  64684=>"111111100",
  64685=>"110010010",
  64686=>"111111000",
  64687=>"101111111",
  64688=>"111111111",
  64689=>"111111011",
  64690=>"001011011",
  64691=>"000000000",
  64692=>"000111111",
  64693=>"000001000",
  64694=>"101001111",
  64695=>"100000111",
  64696=>"111101101",
  64697=>"001001111",
  64698=>"001110110",
  64699=>"000000111",
  64700=>"000000000",
  64701=>"111110100",
  64702=>"000000100",
  64703=>"000000000",
  64704=>"000001111",
  64705=>"101000110",
  64706=>"000110110",
  64707=>"000011111",
  64708=>"111111111",
  64709=>"000000010",
  64710=>"101011111",
  64711=>"000001011",
  64712=>"110110000",
  64713=>"111111111",
  64714=>"110110000",
  64715=>"011001000",
  64716=>"001000000",
  64717=>"000111111",
  64718=>"000000000",
  64719=>"000000000",
  64720=>"110110100",
  64721=>"000001101",
  64722=>"101000000",
  64723=>"000000000",
  64724=>"101001000",
  64725=>"111111110",
  64726=>"000000111",
  64727=>"000000001",
  64728=>"000111111",
  64729=>"001001111",
  64730=>"000000000",
  64731=>"101101111",
  64732=>"000000100",
  64733=>"000000100",
  64734=>"000001010",
  64735=>"000010110",
  64736=>"001011011",
  64737=>"000010010",
  64738=>"111111110",
  64739=>"111000000",
  64740=>"000000011",
  64741=>"111111010",
  64742=>"011000000",
  64743=>"111111011",
  64744=>"011011011",
  64745=>"111111110",
  64746=>"001001011",
  64747=>"000010010",
  64748=>"101101111",
  64749=>"111011000",
  64750=>"001111111",
  64751=>"000000000",
  64752=>"100000111",
  64753=>"001000000",
  64754=>"111111001",
  64755=>"100100110",
  64756=>"000000000",
  64757=>"111100000",
  64758=>"001001111",
  64759=>"001111111",
  64760=>"000110111",
  64761=>"001011111",
  64762=>"111110110",
  64763=>"111111111",
  64764=>"111111111",
  64765=>"100100111",
  64766=>"100000111",
  64767=>"000000000",
  64768=>"100111111",
  64769=>"000000000",
  64770=>"000100100",
  64771=>"100100000",
  64772=>"000000011",
  64773=>"000001001",
  64774=>"000000001",
  64775=>"111001000",
  64776=>"000010111",
  64777=>"000000000",
  64778=>"001000111",
  64779=>"011001011",
  64780=>"111000111",
  64781=>"011001000",
  64782=>"111111010",
  64783=>"000110111",
  64784=>"000000111",
  64785=>"000000110",
  64786=>"110111110",
  64787=>"000000001",
  64788=>"000000110",
  64789=>"111111110",
  64790=>"000000000",
  64791=>"000000000",
  64792=>"001101111",
  64793=>"111111000",
  64794=>"111111111",
  64795=>"010000000",
  64796=>"000000000",
  64797=>"000000000",
  64798=>"111110000",
  64799=>"111101001",
  64800=>"000100110",
  64801=>"000000011",
  64802=>"111111111",
  64803=>"000000100",
  64804=>"111111111",
  64805=>"111000000",
  64806=>"000000000",
  64807=>"111111110",
  64808=>"111111011",
  64809=>"000000111",
  64810=>"010110110",
  64811=>"111000000",
  64812=>"100111111",
  64813=>"000000111",
  64814=>"111111111",
  64815=>"111111000",
  64816=>"111111011",
  64817=>"010011010",
  64818=>"001000111",
  64819=>"100111101",
  64820=>"011011010",
  64821=>"100010111",
  64822=>"000011111",
  64823=>"111011011",
  64824=>"000000000",
  64825=>"101110111",
  64826=>"000111111",
  64827=>"000111111",
  64828=>"000000000",
  64829=>"101001111",
  64830=>"000011111",
  64831=>"111011011",
  64832=>"000000011",
  64833=>"000100000",
  64834=>"000110110",
  64835=>"000000000",
  64836=>"001000000",
  64837=>"101111111",
  64838=>"000001111",
  64839=>"000001000",
  64840=>"000000000",
  64841=>"000000000",
  64842=>"000000000",
  64843=>"110100000",
  64844=>"000000000",
  64845=>"000110100",
  64846=>"001000000",
  64847=>"000111111",
  64848=>"011011000",
  64849=>"100000000",
  64850=>"111100000",
  64851=>"111111011",
  64852=>"001111011",
  64853=>"001001011",
  64854=>"011000000",
  64855=>"111000000",
  64856=>"101000000",
  64857=>"000000111",
  64858=>"001000000",
  64859=>"101000000",
  64860=>"111100000",
  64861=>"111111111",
  64862=>"000111111",
  64863=>"111111001",
  64864=>"000000000",
  64865=>"000110111",
  64866=>"111111111",
  64867=>"000011000",
  64868=>"111111111",
  64869=>"000101111",
  64870=>"000000000",
  64871=>"000000011",
  64872=>"000000000",
  64873=>"000000101",
  64874=>"000000110",
  64875=>"110000000",
  64876=>"010100110",
  64877=>"100100101",
  64878=>"111011000",
  64879=>"001000001",
  64880=>"100111111",
  64881=>"100110010",
  64882=>"000000000",
  64883=>"001001001",
  64884=>"111111000",
  64885=>"111110100",
  64886=>"100000000",
  64887=>"011000000",
  64888=>"000000011",
  64889=>"000000000",
  64890=>"111111111",
  64891=>"111111011",
  64892=>"000100110",
  64893=>"000011001",
  64894=>"000000000",
  64895=>"111111111",
  64896=>"001000100",
  64897=>"000000000",
  64898=>"110110110",
  64899=>"000000000",
  64900=>"100110111",
  64901=>"010111010",
  64902=>"111110111",
  64903=>"001000100",
  64904=>"001000001",
  64905=>"000000010",
  64906=>"101000000",
  64907=>"111011001",
  64908=>"111111111",
  64909=>"000001100",
  64910=>"011001001",
  64911=>"000111111",
  64912=>"000000101",
  64913=>"000000000",
  64914=>"000001001",
  64915=>"000000000",
  64916=>"000111011",
  64917=>"000000011",
  64918=>"100000000",
  64919=>"001000000",
  64920=>"000000001",
  64921=>"110110100",
  64922=>"001000000",
  64923=>"001000000",
  64924=>"001000000",
  64925=>"111111111",
  64926=>"001011111",
  64927=>"000000000",
  64928=>"010011001",
  64929=>"000100111",
  64930=>"111111111",
  64931=>"110111010",
  64932=>"001111101",
  64933=>"111001000",
  64934=>"111001000",
  64935=>"010111111",
  64936=>"000000000",
  64937=>"010010011",
  64938=>"111111100",
  64939=>"000000001",
  64940=>"000001011",
  64941=>"111111111",
  64942=>"100101101",
  64943=>"001000001",
  64944=>"100111111",
  64945=>"000000000",
  64946=>"111111110",
  64947=>"110111111",
  64948=>"001000000",
  64949=>"111111111",
  64950=>"011000111",
  64951=>"111110000",
  64952=>"100010000",
  64953=>"001000000",
  64954=>"111111100",
  64955=>"111011111",
  64956=>"000000111",
  64957=>"001111000",
  64958=>"000000000",
  64959=>"000000000",
  64960=>"111111010",
  64961=>"000001111",
  64962=>"000011111",
  64963=>"111101000",
  64964=>"011111011",
  64965=>"001000000",
  64966=>"011011000",
  64967=>"000000001",
  64968=>"111011011",
  64969=>"011111111",
  64970=>"100100111",
  64971=>"000000000",
  64972=>"111000000",
  64973=>"001011111",
  64974=>"000000110",
  64975=>"111111111",
  64976=>"011000000",
  64977=>"000000000",
  64978=>"000001111",
  64979=>"111111111",
  64980=>"011011001",
  64981=>"111101111",
  64982=>"111111111",
  64983=>"001000010",
  64984=>"001000000",
  64985=>"000000001",
  64986=>"111110000",
  64987=>"111111000",
  64988=>"111111111",
  64989=>"111111111",
  64990=>"101000000",
  64991=>"011011111",
  64992=>"111001111",
  64993=>"000000011",
  64994=>"001000000",
  64995=>"000000011",
  64996=>"000000100",
  64997=>"111111111",
  64998=>"000000111",
  64999=>"111111000",
  65000=>"111111111",
  65001=>"000100000",
  65002=>"100000000",
  65003=>"111111111",
  65004=>"111111111",
  65005=>"000000000",
  65006=>"000000111",
  65007=>"111100111",
  65008=>"100000000",
  65009=>"000000101",
  65010=>"111111110",
  65011=>"000010000",
  65012=>"000001000",
  65013=>"111111101",
  65014=>"111111100",
  65015=>"010001000",
  65016=>"000000000",
  65017=>"011011000",
  65018=>"111001001",
  65019=>"111111000",
  65020=>"011011011",
  65021=>"011011100",
  65022=>"000001000",
  65023=>"000110111",
  65024=>"111111111",
  65025=>"101111111",
  65026=>"000000101",
  65027=>"110110111",
  65028=>"110110110",
  65029=>"100000000",
  65030=>"000000000",
  65031=>"101000000",
  65032=>"111110100",
  65033=>"000000000",
  65034=>"111111000",
  65035=>"110110110",
  65036=>"111111110",
  65037=>"010011001",
  65038=>"000000000",
  65039=>"000000000",
  65040=>"110000000",
  65041=>"011111111",
  65042=>"111111111",
  65043=>"111111111",
  65044=>"011101101",
  65045=>"111111111",
  65046=>"110111000",
  65047=>"000011111",
  65048=>"111001101",
  65049=>"110111010",
  65050=>"000000111",
  65051=>"001011011",
  65052=>"000101111",
  65053=>"100000001",
  65054=>"011111011",
  65055=>"001111000",
  65056=>"011011111",
  65057=>"111110100",
  65058=>"111111110",
  65059=>"000000000",
  65060=>"000000000",
  65061=>"111111111",
  65062=>"111111110",
  65063=>"111111111",
  65064=>"111110000",
  65065=>"000000000",
  65066=>"001001011",
  65067=>"111111111",
  65068=>"111111111",
  65069=>"000111111",
  65070=>"000000111",
  65071=>"011011001",
  65072=>"000000000",
  65073=>"000100100",
  65074=>"111111110",
  65075=>"100000000",
  65076=>"000000111",
  65077=>"100000000",
  65078=>"000000111",
  65079=>"001001000",
  65080=>"001000000",
  65081=>"001001111",
  65082=>"010111110",
  65083=>"000000000",
  65084=>"001000000",
  65085=>"000000000",
  65086=>"000000000",
  65087=>"000000000",
  65088=>"111111111",
  65089=>"000001001",
  65090=>"111111111",
  65091=>"000000111",
  65092=>"100100000",
  65093=>"000000000",
  65094=>"001111111",
  65095=>"000000000",
  65096=>"100100110",
  65097=>"000000000",
  65098=>"000000000",
  65099=>"110111000",
  65100=>"000000000",
  65101=>"000010111",
  65102=>"110000000",
  65103=>"001001000",
  65104=>"111111100",
  65105=>"111011011",
  65106=>"001001001",
  65107=>"000000000",
  65108=>"110111111",
  65109=>"000000000",
  65110=>"110110110",
  65111=>"111111111",
  65112=>"111111111",
  65113=>"000000000",
  65114=>"000000111",
  65115=>"100111111",
  65116=>"000001011",
  65117=>"111111111",
  65118=>"001011000",
  65119=>"001111111",
  65120=>"000000000",
  65121=>"100001111",
  65122=>"000000000",
  65123=>"001001001",
  65124=>"111110110",
  65125=>"100000000",
  65126=>"110111000",
  65127=>"111111111",
  65128=>"111111111",
  65129=>"111101111",
  65130=>"000000000",
  65131=>"000000000",
  65132=>"000000000",
  65133=>"000000000",
  65134=>"000000000",
  65135=>"101000011",
  65136=>"000000000",
  65137=>"010111111",
  65138=>"110110011",
  65139=>"100000000",
  65140=>"101101110",
  65141=>"011000000",
  65142=>"001000000",
  65143=>"000000000",
  65144=>"100100100",
  65145=>"000000000",
  65146=>"000000000",
  65147=>"001001011",
  65148=>"100110110",
  65149=>"000100100",
  65150=>"000010000",
  65151=>"100000000",
  65152=>"111111000",
  65153=>"000011111",
  65154=>"000111111",
  65155=>"110000000",
  65156=>"000000000",
  65157=>"111111111",
  65158=>"011111010",
  65159=>"000001011",
  65160=>"100000000",
  65161=>"011111001",
  65162=>"000000000",
  65163=>"111100100",
  65164=>"000000000",
  65165=>"010000000",
  65166=>"100000110",
  65167=>"110100110",
  65168=>"001001011",
  65169=>"000000000",
  65170=>"011111110",
  65171=>"111111111",
  65172=>"011000001",
  65173=>"101100110",
  65174=>"101111111",
  65175=>"001001000",
  65176=>"000110101",
  65177=>"111111111",
  65178=>"100000000",
  65179=>"000010000",
  65180=>"111111111",
  65181=>"000000001",
  65182=>"110100101",
  65183=>"111111111",
  65184=>"110000001",
  65185=>"010111111",
  65186=>"000001000",
  65187=>"110111111",
  65188=>"000010000",
  65189=>"110011000",
  65190=>"000000101",
  65191=>"011011111",
  65192=>"100111111",
  65193=>"000000001",
  65194=>"000000000",
  65195=>"000000000",
  65196=>"101011011",
  65197=>"000000001",
  65198=>"100100000",
  65199=>"111111111",
  65200=>"010011000",
  65201=>"111100110",
  65202=>"111111111",
  65203=>"000000001",
  65204=>"110000000",
  65205=>"111000000",
  65206=>"000000000",
  65207=>"111111111",
  65208=>"101101000",
  65209=>"011000000",
  65210=>"000000100",
  65211=>"000000011",
  65212=>"000000111",
  65213=>"111111110",
  65214=>"000000000",
  65215=>"111111111",
  65216=>"000100110",
  65217=>"111111111",
  65218=>"000001000",
  65219=>"110110000",
  65220=>"111111111",
  65221=>"000000001",
  65222=>"111000000",
  65223=>"000000011",
  65224=>"010110111",
  65225=>"111001000",
  65226=>"000000000",
  65227=>"010100110",
  65228=>"011011001",
  65229=>"000000110",
  65230=>"110111111",
  65231=>"000111111",
  65232=>"000100110",
  65233=>"011111011",
  65234=>"110111111",
  65235=>"100000111",
  65236=>"101111100",
  65237=>"111111111",
  65238=>"000000000",
  65239=>"000000000",
  65240=>"011110000",
  65241=>"011001000",
  65242=>"111001011",
  65243=>"010111110",
  65244=>"100100100",
  65245=>"111111111",
  65246=>"111111111",
  65247=>"000000000",
  65248=>"000000000",
  65249=>"000011011",
  65250=>"110000000",
  65251=>"100000000",
  65252=>"000000000",
  65253=>"110111111",
  65254=>"000000000",
  65255=>"101111101",
  65256=>"111111001",
  65257=>"000011011",
  65258=>"111011111",
  65259=>"000011001",
  65260=>"111111111",
  65261=>"111011111",
  65262=>"000000111",
  65263=>"111111111",
  65264=>"000000000",
  65265=>"111001001",
  65266=>"110111111",
  65267=>"000000000",
  65268=>"000000000",
  65269=>"111111100",
  65270=>"111111011",
  65271=>"111111011",
  65272=>"001011010",
  65273=>"100000000",
  65274=>"101111111",
  65275=>"001100100",
  65276=>"111111101",
  65277=>"111011011",
  65278=>"000000110",
  65279=>"111111111",
  65280=>"000000000",
  65281=>"001001001",
  65282=>"111111111",
  65283=>"000000111",
  65284=>"111110000",
  65285=>"110100000",
  65286=>"111110111",
  65287=>"000001000",
  65288=>"100000000",
  65289=>"000000011",
  65290=>"111100100",
  65291=>"100100100",
  65292=>"111001000",
  65293=>"100000000",
  65294=>"111111010",
  65295=>"000000000",
  65296=>"100111111",
  65297=>"111111111",
  65298=>"111111101",
  65299=>"110110101",
  65300=>"010000000",
  65301=>"111000000",
  65302=>"001011101",
  65303=>"011011000",
  65304=>"111111100",
  65305=>"000000000",
  65306=>"000000000",
  65307=>"111111000",
  65308=>"011011111",
  65309=>"111110101",
  65310=>"000000000",
  65311=>"111111111",
  65312=>"110110010",
  65313=>"000000110",
  65314=>"111111111",
  65315=>"000000000",
  65316=>"000110110",
  65317=>"000000000",
  65318=>"011111111",
  65319=>"000110111",
  65320=>"000000000",
  65321=>"011001000",
  65322=>"000000000",
  65323=>"000000000",
  65324=>"111111111",
  65325=>"011111111",
  65326=>"000000000",
  65327=>"100111011",
  65328=>"111111111",
  65329=>"111111111",
  65330=>"001001001",
  65331=>"000000000",
  65332=>"000000111",
  65333=>"111111111",
  65334=>"111111010",
  65335=>"000000000",
  65336=>"000000000",
  65337=>"001011000",
  65338=>"000010000",
  65339=>"111111100",
  65340=>"110111111",
  65341=>"000010010",
  65342=>"100101111",
  65343=>"100100000",
  65344=>"000000000",
  65345=>"001001001",
  65346=>"110110111",
  65347=>"001000000",
  65348=>"001011000",
  65349=>"011000110",
  65350=>"000000000",
  65351=>"111101100",
  65352=>"000000000",
  65353=>"111000000",
  65354=>"000000000",
  65355=>"111110000",
  65356=>"000000000",
  65357=>"111111000",
  65358=>"000010100",
  65359=>"001011110",
  65360=>"000000100",
  65361=>"000000001",
  65362=>"000000000",
  65363=>"111110000",
  65364=>"111110011",
  65365=>"011011011",
  65366=>"000000111",
  65367=>"100111011",
  65368=>"111101111",
  65369=>"111100100",
  65370=>"001000000",
  65371=>"000000111",
  65372=>"110111111",
  65373=>"111111111",
  65374=>"011111111",
  65375=>"111111000",
  65376=>"010000100",
  65377=>"111111111",
  65378=>"111111111",
  65379=>"111100000",
  65380=>"000101100",
  65381=>"000000000",
  65382=>"001011111",
  65383=>"000000000",
  65384=>"011011011",
  65385=>"000000010",
  65386=>"111111011",
  65387=>"100010001",
  65388=>"100000000",
  65389=>"000011111",
  65390=>"000000000",
  65391=>"000000010",
  65392=>"000011011",
  65393=>"000001111",
  65394=>"000000000",
  65395=>"111110110",
  65396=>"000110010",
  65397=>"001000000",
  65398=>"110100000",
  65399=>"111111101",
  65400=>"000000000",
  65401=>"111111111",
  65402=>"100111011",
  65403=>"001000000",
  65404=>"011111000",
  65405=>"011000000",
  65406=>"000100111",
  65407=>"111111111",
  65408=>"111110110",
  65409=>"110011011",
  65410=>"000001000",
  65411=>"111100100",
  65412=>"001000100",
  65413=>"000111111",
  65414=>"000000101",
  65415=>"000000111",
  65416=>"000000000",
  65417=>"001001111",
  65418=>"000000000",
  65419=>"001000011",
  65420=>"000000000",
  65421=>"000000000",
  65422=>"000000000",
  65423=>"111000000",
  65424=>"000000000",
  65425=>"000000000",
  65426=>"110110110",
  65427=>"010000000",
  65428=>"111111000",
  65429=>"000000000",
  65430=>"000100000",
  65431=>"101111110",
  65432=>"111111111",
  65433=>"000000000",
  65434=>"101101000",
  65435=>"011111111",
  65436=>"000000000",
  65437=>"001001101",
  65438=>"000000000",
  65439=>"001011111",
  65440=>"000000000",
  65441=>"011001000",
  65442=>"110011111",
  65443=>"111111111",
  65444=>"000000100",
  65445=>"000000000",
  65446=>"001001000",
  65447=>"111111111",
  65448=>"100000000",
  65449=>"000000000",
  65450=>"111110110",
  65451=>"000000000",
  65452=>"111111000",
  65453=>"100001011",
  65454=>"111111011",
  65455=>"000000000",
  65456=>"000000000",
  65457=>"111111111",
  65458=>"111111111",
  65459=>"000000000",
  65460=>"111111111",
  65461=>"110000001",
  65462=>"111111111",
  65463=>"000000000",
  65464=>"110110110",
  65465=>"010111111",
  65466=>"110110100",
  65467=>"111111101",
  65468=>"011001001",
  65469=>"111111111",
  65470=>"111111001",
  65471=>"001001001",
  65472=>"000000000",
  65473=>"000000000",
  65474=>"000000000",
  65475=>"000100000",
  65476=>"000000000",
  65477=>"000101000",
  65478=>"000000000",
  65479=>"000000001",
  65480=>"111111111",
  65481=>"000000000",
  65482=>"000000000",
  65483=>"000000000",
  65484=>"010010000",
  65485=>"000000000",
  65486=>"001000000",
  65487=>"001110110",
  65488=>"101001000",
  65489=>"100100011",
  65490=>"111111110",
  65491=>"000000000",
  65492=>"000001000",
  65493=>"000000000",
  65494=>"011000110",
  65495=>"011111111",
  65496=>"111010010",
  65497=>"000000000",
  65498=>"001100000",
  65499=>"101101100",
  65500=>"101100111",
  65501=>"000010000",
  65502=>"100100000",
  65503=>"110110100",
  65504=>"011111111",
  65505=>"101111111",
  65506=>"110111100",
  65507=>"110001001",
  65508=>"111111111",
  65509=>"000000000",
  65510=>"111111111",
  65511=>"001111110",
  65512=>"000000000",
  65513=>"111011001",
  65514=>"111000000",
  65515=>"110111111",
  65516=>"111001001",
  65517=>"111111111",
  65518=>"011001011",
  65519=>"000000000",
  65520=>"000000110",
  65521=>"000000000",
  65522=>"111111111",
  65523=>"000000001",
  65524=>"011111110",
  65525=>"000000000",
  65526=>"011011111",
  65527=>"001011111",
  65528=>"111111111",
  65529=>"000000010",
  65530=>"101111111",
  65531=>"001001000",
  65532=>"001001111",
  65533=>"111111111",
  65534=>"000010000",
  65535=>"000000000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;