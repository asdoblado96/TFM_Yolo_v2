LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_1_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(6 DOWNTO 0));
END L7_1_BNROM;

ARCHITECTURE RTL OF L7_1_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"1101110110101010"&"0010001110100000",
  1=>"0000001100011000"&"0010100100001000",
  2=>"1111111010011100"&"0010101101111001",
  3=>"1111010110011001"&"0010000110010110",
  4=>"1111001001000001"&"0010010001010101",
  5=>"1110110111000000"&"0010011101011001",
  6=>"1110111010111111"&"0010010011101011",
  7=>"1110100000101110"&"0010100111110001",
  8=>"1110110000001001"&"0010100001100100",
  9=>"1110001001011111"&"0010010100011100",
  10=>"1111000000010010"&"0010001001011101",
  11=>"1111110110000100"&"0010001100111100",
  12=>"1110100100010101"&"0010001010011101",
  13=>"1111000101100111"&"0010010100011000",
  14=>"1111010011100111"&"0010001100100011",
  15=>"1110011010101001"&"0010101011101100",
  16=>"1110110001100111"&"0010010100010100",
  17=>"1110110010010101"&"0010010101010100",
  18=>"1111000100000011"&"0010010111111000",
  19=>"1111000010110101"&"0010010000100011",
  20=>"1101111111100010"&"0010100001001011",
  21=>"1110000101111010"&"0010010001010111",
  22=>"1111010111000011"&"0010010111011101",
  23=>"1101101110000010"&"0001111111100001",
  24=>"1110000011001011"&"0010011111011001",
  25=>"1111011011100110"&"0010010100100001",
  26=>"1110100110001000"&"0010000100001001",
  27=>"1111010111001001"&"0010010101000110",
  28=>"1110111000011110"&"0010001001010110",
  29=>"1111110010011010"&"0010010111010001",
  30=>"1111001110010100"&"0010010110010110",
  31=>"1110110110111111"&"0010000111001111",
  32=>"1110001101110001"&"0010100010000111",
  33=>"1110111111001111"&"0010010111101101",
  34=>"1111010011100011"&"0010101101001011",
  35=>"1110011110110001"&"0010100100010110",
  36=>"1110101010110101"&"0010111110100000",
  37=>"1110011110010111"&"0010011011100000",
  38=>"1110100001110001"&"0010010010000010",
  39=>"0000000101100000"&"0010010111110010",
  40=>"1110010011101101"&"0010011011110110",
  41=>"1111010101100011"&"0010010011000101",
  42=>"1110001100110101"&"0010100010000100",
  43=>"1111010100001110"&"0010001011100010",
  44=>"1101101010100001"&"0010100001111100",
  45=>"1110110100111111"&"0010010111100010",
  46=>"1110011001100101"&"0010010110011101",
  47=>"1101110001010010"&"0010010110000100",
  48=>"1110111001110100"&"0010101111101100",
  49=>"1111011001000000"&"0010000000010110",
  50=>"1111010111001000"&"0010110001000010",
  51=>"1110100001100111"&"0010010011100001",
  52=>"1111011111000011"&"0010001010011000",
  53=>"1110001001001010"&"0010001100110011",
  54=>"1110101101111011"&"0010010000010001",
  55=>"1110111111110001"&"0010010010000110",
  56=>"1111000101010001"&"0011000110111100",
  57=>"1110010101111111"&"0010011001100000",
  58=>"1110000011000101"&"0010101000100011",
  59=>"1110001111001011"&"0010101100111101",
  60=>"1111000001111101"&"0010010011101101",
  61=>"1110101100000110"&"0010010101111011",
  62=>"1110011010000000"&"0010010000111011",
  63=>"1111000010011100"&"0001111110100000",
  64=>"1110100110001011"&"0010010000000110",
  65=>"1110101100101011"&"0001110010000110",
  66=>"1111110100100011"&"0010010100110000",
  67=>"1111010100111010"&"0010001011001110",
  68=>"0000001110000110"&"0010000000111011",
  69=>"1110011110010101"&"0010100000001001",
  70=>"1101101010100101"&"0010110011001100",
  71=>"1110101010100100"&"0010011110011100",
  72=>"1111100010111110"&"0010001001011000",
  73=>"1111000010111110"&"0010100000001111",
  74=>"1111011110110000"&"0010001111110110",
  75=>"1110100101110101"&"0010100100000110",
  76=>"1110011000011101"&"0010001010110101",
  77=>"1101100011110010"&"0010101011111001",
  78=>"1111001011110011"&"0010001011100011",
  79=>"1111001011001000"&"0010001111011011",
  80=>"1110100000001110"&"0010101000001001",
  81=>"1101111011100010"&"0010001111101100",
  82=>"1111010011101100"&"0010101000100111",
  83=>"1111000011001001"&"0010100001011100",
  84=>"1111010001001111"&"0010001011010101",
  85=>"1110110101111101"&"0010110110110000",
  86=>"0000010111101001"&"0010010011001100",
  87=>"1111000110001010"&"0010010011011011",
  88=>"1111011100111111"&"0010010100011100",
  89=>"1110110101101000"&"0010011011000011",
  90=>"1110011010111011"&"0010010011111001",
  91=>"1111001000101101"&"0010000001101010",
  92=>"1110111011010111"&"0010011110101001",
  93=>"1110001100101011"&"0010100010000100",
  94=>"1110111111111010"&"0010011010111011",
  95=>"1110011100011110"&"0010101110101011",
  96=>"1101010111001101"&"0010010011101100",
  97=>"1111010001000110"&"0010000101100011",
  98=>"1110101101111000"&"0010010111101101",
  99=>"1111000010001100"&"0010001001100100",
  100=>"1110110001001011"&"0010000011000101",
  101=>"1111001111110001"&"0010100111101011",
  102=>"0000001001001111"&"0010010001101001",
  103=>"1111010010010010"&"0010000010001101",
  104=>"1110110110110010"&"0010001101100110",
  105=>"1101000001011011"&"0010100001011000",
  106=>"1111100011101100"&"0010010000100010",
  107=>"1111011110001011"&"0010000010111011",
  108=>"1111000100010111"&"0010011000000000",
  109=>"1110111001000000"&"0010010000011110",
  110=>"1110001000111111"&"0010000111011111",
  111=>"1101100110111110"&"0010101010100110",
  112=>"1111100110011101"&"0010111110111100",
  113=>"1111110110001110"&"0010000001001100",
  114=>"1110000000001101"&"0010110001001100",
  115=>"1101011001100110"&"0010110101001111",
  116=>"1110111000110100"&"0010011110010111",
  117=>"1111001101101001"&"0010010100110101",
  118=>"1111011111000001"&"0010101100101010",
  119=>"1111010100111001"&"0010011101010110",
  120=>"1110101010001101"&"0010001001100011",
  121=>"1111001000011011"&"0010010000011110",
  122=>"1111110101111000"&"0010010100010001",
  123=>"1111100000011000"&"0010011100001010",
  124=>"1110001110011111"&"0010001010100010",
  125=>"1110100001001100"&"0010100010011001",
  126=>"1110110110111001"&"0010010110001110",
  127=>"1110100111100001"&"0010010010000100");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;