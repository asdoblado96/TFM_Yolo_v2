LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_4_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_4_BNROM;

ARCHITECTURE RTL OF L8_4_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0010010101111000"&"0010001001011010",
  1=>"0000111111101111"&"0001101011010011",
  2=>"0001100001101100"&"0010000101101111",
  3=>"0001110111001101"&"0010001010001010",
  4=>"0001011010001011"&"0010000100011000",
  5=>"0001100011101110"&"0010010101000000",
  6=>"0001000110111001"&"0010011001011100",
  7=>"0010010001000101"&"0010010001010111",
  8=>"0000000011100110"&"0010000011011111",
  9=>"0010110001100010"&"0010001100101100",
  10=>"0000010111001111"&"0001111000100111",
  11=>"1110111000010000"&"0010000100111111",
  12=>"0001101111110000"&"0010010111000011",
  13=>"0001010001001000"&"0010000011111011",
  14=>"0001001111011001"&"0001111000110001",
  15=>"1111011010010100"&"0010010010100110",
  16=>"0010011000101110"&"0010001111101100",
  17=>"0001110001000011"&"0010011110100000",
  18=>"0010001100010111"&"0001100111111100",
  19=>"0001011101001000"&"0010010000010011",
  20=>"0001011100010011"&"0001100001111001",
  21=>"0000110001001100"&"0010011100100001",
  22=>"0001110010101010"&"0001111101111110",
  23=>"0010001011010000"&"0010001110110101",
  24=>"0000100001010100"&"0010001111111011",
  25=>"0001011011111000"&"0001111110100010",
  26=>"0010011100000110"&"0010000011100000",
  27=>"0010000010100011"&"0010011111110100",
  28=>"0001101100101010"&"0010010110001001",
  29=>"0001100111111001"&"0010011011111010",
  30=>"0001111001101101"&"0010011001000001",
  31=>"0001001101010010"&"0010010011101100",
  32=>"0001111001010001"&"0010000001100001",
  33=>"0001010111101100"&"0010011010000011",
  34=>"0000011110111101"&"0010001110011110",
  35=>"0010011101111101"&"0010000111111011",
  36=>"0001000010100101"&"0010001000001011",
  37=>"0000001111110110"&"0010011001100010",
  38=>"0001101011010000"&"0010010100101011",
  39=>"0000001101110011"&"0010011000001000",
  40=>"0001101010000111"&"0001100100100110",
  41=>"0000010101101000"&"0010010100100010",
  42=>"0001100111101001"&"0010001111100000",
  43=>"0001000010010011"&"0001101001001011",
  44=>"0010010010000000"&"0001100011100100",
  45=>"0000110101100001"&"0010001101111010",
  46=>"0001001011010011"&"0010010011010010",
  47=>"0010011111000101"&"0001101000001011",
  48=>"0000000101100101"&"0010100001000100",
  49=>"0000000111010000"&"0010011100011110",
  50=>"0001101101000000"&"0010010101000101",
  51=>"0001000000000110"&"0010000110000100",
  52=>"0010011111110111"&"0010010010001011",
  53=>"0001101010001010"&"0010001111111001",
  54=>"0001101101110000"&"0001111101100011",
  55=>"0010000001111111"&"0010010010110101",
  56=>"0000000000011000"&"0010001001100011",
  57=>"0001011010100000"&"0001111000101011",
  58=>"0000011101100001"&"0010010100100100",
  59=>"0001111101100101"&"0001111011010110",
  60=>"0001011100001101"&"0010001111001100",
  61=>"0001011100101010"&"0010000001010101",
  62=>"0001010001110011"&"0001111110001010",
  63=>"0000011011011001"&"0001111101010011");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;