LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L4_2_WROM IS
    PORT (
        weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        address : IN unsigned(weightsbitsAddress(4)-1 DOWNTO 0));
END L4_2_WROM;

ARCHITECTURE RTL OF L4_2_WROM IS

    TYPE ROM_mem IS ARRAY (0 TO 4095) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem := (0=>"100100000",
    1=>"110111001",
    2=>"110110111",
    3=>"111001001",
    4=>"000000000",
    5=>"000100110",
    6=>"100110110",
    7=>"001101101",
    8=>"111011101",
    9=>"000110000",
    10=>"000100000",
    11=>"101011001",
    12=>"110111111",
    13=>"111111111",
    14=>"000100110",
    15=>"100110001",
    16=>"010110100",
    17=>"111110010",
    18=>"000001101",
    19=>"000000101",
    20=>"111001101",
    21=>"000000000",
    22=>"100100100",
    23=>"000001010",
    24=>"111000101",
    25=>"000110000",
    26=>"001101011",
    27=>"110110100",
    28=>"000001000",
    29=>"001001111",
    30=>"100000110",
    31=>"000010000",
    32=>"000000010",
    33=>"001100100",
    34=>"111010000",
    35=>"110100000",
    36=>"000000000",
    37=>"000110101",
    38=>"000010110",
    39=>"110111111",
    40=>"110111111",
    41=>"000110111",
    42=>"000100110",
    43=>"010000001",
    44=>"101001101",
    45=>"001101101",
    46=>"010000000",
    47=>"110110100",
    48=>"111111111",
    49=>"000010000",
    50=>"110111001",
    51=>"111101111",
    52=>"111011001",
    53=>"110000001",
    54=>"000010000",
    55=>"000110010",
    56=>"101110001",
    57=>"110011011",
    58=>"000101111",
    59=>"001011011",
    60=>"100000000",
    61=>"000010111",
    62=>"000111101",
    63=>"110111111",
    64=>"010010100",
    65=>"000100011",
    66=>"110111001",
    67=>"111111100",
    68=>"100100110",
    69=>"100101001",
    70=>"111111110",
    71=>"011001110",
    72=>"111100010",
    73=>"101101000",
    74=>"001001111",
    75=>"000010011",
    76=>"101001111",
    77=>"000000000",
    78=>"000010010",
    79=>"111000101",
    80=>"000111111",
    81=>"101100101",
    82=>"111111011",
    83=>"000000000",
    84=>"100011001",
    85=>"000000100",
    86=>"000111111",
    87=>"000111100",
    88=>"000100010",
    89=>"000000111",
    90=>"001101100",
    91=>"011010000",
    92=>"000101111",
    93=>"111101001",
    94=>"100111011",
    95=>"000011010",
    96=>"010010010",
    97=>"011011001",
    98=>"000011000",
    99=>"001010110",
    100=>"001111011",
    101=>"110000011",
    102=>"110110100",
    103=>"000000000",
    104=>"111011010",
    105=>"000000000",
    106=>"100010010",
    107=>"001111111",
    108=>"010010011",
    109=>"001010110",
    110=>"111001101",
    111=>"000010000",
    112=>"001000000",
    113=>"000000111",
    114=>"101100011",
    115=>"011000000",
    116=>"111110000",
    117=>"111110110",
    118=>"000010000",
    119=>"000010011",
    120=>"000010110",
    121=>"100010110",
    122=>"111111110",
    123=>"001011110",
    124=>"000101101",
    125=>"100000001",
    126=>"000000000",
    127=>"000010111",
    128=>"000101111",
    129=>"111111000",
    130=>"100111111",
    131=>"011010111",
    132=>"000110111",
    133=>"101111111",
    134=>"110100001",
    135=>"000100111",
    136=>"101100000",
    137=>"111110000",
    138=>"011110111",
    139=>"000000011",
    140=>"011000111",
    141=>"101000000",
    142=>"111001001",
    143=>"111000000",
    144=>"100000011",
    145=>"111000000",
    146=>"001011100",
    147=>"111011001",
    148=>"001000010",
    149=>"111000000",
    150=>"000111111",
    151=>"111110000",
    152=>"000010111",
    153=>"111000000",
    154=>"101011111",
    155=>"110000001",
    156=>"111100010",
    157=>"111000111",
    158=>"111111000",
    159=>"111010000",
    160=>"000001111",
    161=>"111001000",
    162=>"100000000",
    163=>"000000111",
    164=>"111010010",
    165=>"000000111",
    166=>"111001000",
    167=>"111111101",
    168=>"000001111",
    169=>"111110000",
    170=>"111011000",
    171=>"111000011",
    172=>"001101111",
    173=>"110000111",
    174=>"000001111",
    175=>"001101000",
    176=>"111000000",
    177=>"111000000",
    178=>"000000111",
    179=>"001001000",
    180=>"111110000",
    181=>"000000001",
    182=>"000110110",
    183=>"000100111",
    184=>"111011000",
    185=>"001011111",
    186=>"100010001",
    187=>"110011111",
    188=>"000001111",
    189=>"000001111",
    190=>"111111001",
    191=>"111000010",
    192=>"000111001",
    193=>"111010010",
    194=>"011111001",
    195=>"100001111",
    196=>"011011100",
    197=>"000110110",
    198=>"111011110",
    199=>"110101001",
    200=>"111011000",
    201=>"101101001",
    202=>"110100000",
    203=>"101110100",
    204=>"111111010",
    205=>"010010000",
    206=>"001101100",
    207=>"001001101",
    208=>"110010110",
    209=>"110000010",
    210=>"011110100",
    211=>"010000001",
    212=>"111000000",
    213=>"010010000",
    214=>"110000111",
    215=>"010010011",
    216=>"010010010",
    217=>"010010010",
    218=>"100011011",
    219=>"110111010",
    220=>"000010010",
    221=>"001101111",
    222=>"011111010",
    223=>"000000000",
    224=>"111111000",
    225=>"001110110",
    226=>"000000110",
    227=>"000000111",
    228=>"000000000",
    229=>"001100100",
    230=>"010011011",
    231=>"000000000",
    232=>"111111100",
    233=>"101111000",
    234=>"001101110",
    235=>"010000011",
    236=>"001111100",
    237=>"111111001",
    238=>"111101101",
    239=>"000000000",
    240=>"111111110",
    241=>"111011000",
    242=>"011001000",
    243=>"111111110",
    244=>"000000000",
    245=>"100111001",
    246=>"000001001",
    247=>"000111010",
    248=>"110010011",
    249=>"111101001",
    250=>"110111001",
    251=>"100111000",
    252=>"111110111",
    253=>"011001000",
    254=>"000000000",
    255=>"000000000",
    256=>"000001000",
    257=>"110110011",
    258=>"100010001",
    259=>"001110011",
    260=>"111011000",
    261=>"100110111",
    262=>"001010000",
    263=>"011111001",
    264=>"011001001",
    265=>"011010100",
    266=>"001001011",
    267=>"000110011",
    268=>"111011111",
    269=>"110011000",
    270=>"010001100",
    271=>"110100011",
    272=>"000000000",
    273=>"111110001",
    274=>"111001101",
    275=>"111100000",
    276=>"011001100",
    277=>"001100100",
    278=>"011111100",
    279=>"101001001",
    280=>"111000100",
    281=>"101001110",
    282=>"111000011",
    283=>"011001101",
    284=>"100100001",
    285=>"100011100",
    286=>"000000110",
    287=>"001011100",
    288=>"011100110",
    289=>"000100110",
    290=>"000110110",
    291=>"111100000",
    292=>"100011111",
    293=>"001100110",
    294=>"111110100",
    295=>"001000110",
    296=>"001010100",
    297=>"101001101",
    298=>"101001000",
    299=>"000001100",
    300=>"101100101",
    301=>"000110000",
    302=>"011110110",
    303=>"101001101",
    304=>"001011010",
    305=>"001011011",
    306=>"111110111",
    307=>"000100110",
    308=>"001110001",
    309=>"110100000",
    310=>"101100010",
    311=>"001100101",
    312=>"110001011",
    313=>"011001110",
    314=>"101111011",
    315=>"000110100",
    316=>"100100010",
    317=>"000000001",
    318=>"110100101",
    319=>"001100100",
    320=>"001111011",
    321=>"101100011",
    322=>"011111010",
    323=>"011011001",
    324=>"111111110",
    325=>"010011110",
    326=>"111111011",
    327=>"100000000",
    328=>"111111110",
    329=>"111111110",
    330=>"000000000",
    331=>"001101101",
    332=>"111111110",
    333=>"110010010",
    334=>"110101100",
    335=>"010011111",
    336=>"111111011",
    337=>"011111111",
    338=>"001101111",
    339=>"110110110",
    340=>"011011111",
    341=>"100100100",
    342=>"000010111",
    343=>"110100011",
    344=>"101101101",
    345=>"100100100",
    346=>"110011010",
    347=>"101000100",
    348=>"010000011",
    349=>"000010110",
    350=>"011011111",
    351=>"001000001",
    352=>"001001011",
    353=>"000000000",
    354=>"000100100",
    355=>"000000000",
    356=>"111111110",
    357=>"000000100",
    358=>"110111111",
    359=>"100101111",
    360=>"000001000",
    361=>"110111111",
    362=>"101001101",
    363=>"000000000",
    364=>"101101101",
    365=>"000000001",
    366=>"000110010",
    367=>"000001001",
    368=>"000101101",
    369=>"000100100",
    370=>"011010011",
    371=>"000101011",
    372=>"000011011",
    373=>"111111111",
    374=>"101100100",
    375=>"100000100",
    376=>"101001111",
    377=>"100101101",
    378=>"100111001",
    379=>"100000000",
    380=>"000000010",
    381=>"000000000",
    382=>"111100101",
    383=>"100000000",
    384=>"000000000",
    385=>"111000000",
    386=>"000100000",
    387=>"000011000",
    388=>"011011000",
    389=>"010111000",
    390=>"110111011",
    391=>"110111000",
    392=>"000100100",
    393=>"111111111",
    394=>"111111110",
    395=>"111111001",
    396=>"010110010",
    397=>"111111111",
    398=>"000111110",
    399=>"111101000",
    400=>"000010101",
    401=>"110010110",
    402=>"010100100",
    403=>"000111000",
    404=>"110111111",
    405=>"010111010",
    406=>"011011011",
    407=>"110000111",
    408=>"000110101",
    409=>"000000110",
    410=>"000011001",
    411=>"010110001",
    412=>"111101111",
    413=>"000111000",
    414=>"101111010",
    415=>"000101111",
    416=>"110011000",
    417=>"100110110",
    418=>"001000000",
    419=>"000010000",
    420=>"111011100",
    421=>"111111100",
    422=>"000111010",
    423=>"000001100",
    424=>"000010110",
    425=>"100100000",
    426=>"101011010",
    427=>"111100111",
    428=>"000010000",
    429=>"000000000",
    430=>"010010010",
    431=>"011100000",
    432=>"000000000",
    433=>"010011001",
    434=>"000111000",
    435=>"000000100",
    436=>"100111111",
    437=>"100110100",
    438=>"110111011",
    439=>"110110000",
    440=>"000100000",
    441=>"011111100",
    442=>"010010110",
    443=>"000111000",
    444=>"000010000",
    445=>"011001110",
    446=>"110110010",
    447=>"111111111",
    448=>"101001000",
    449=>"000100110",
    450=>"111111001",
    451=>"111010000",
    452=>"111111000",
    453=>"001000101",
    454=>"000000111",
    455=>"111111000",
    456=>"111000000",
    457=>"010000111",
    458=>"111010000",
    459=>"001000110",
    460=>"111000000",
    461=>"010100010",
    462=>"010100011",
    463=>"111101000",
    464=>"000000111",
    465=>"000000111",
    466=>"000101000",
    467=>"011000001",
    468=>"011110111",
    469=>"000000111",
    470=>"000000111",
    471=>"000111111",
    472=>"111110110",
    473=>"000001111",
    474=>"100000111",
    475=>"000000111",
    476=>"000101111",
    477=>"111111000",
    478=>"000000111",
    479=>"000000111",
    480=>"111111000",
    481=>"000110110",
    482=>"011110101",
    483=>"111111000",
    484=>"000101111",
    485=>"111111000",
    486=>"000001011",
    487=>"111011101",
    488=>"111111001",
    489=>"000100111",
    490=>"000011111",
    491=>"000000100",
    492=>"100101000",
    493=>"000000111",
    494=>"111111000",
    495=>"000100111",
    496=>"000010110",
    497=>"000111111",
    498=>"001101000",
    499=>"001001111",
    500=>"000000111",
    501=>"111101000",
    502=>"000100001",
    503=>"111111000",
    504=>"000000111",
    505=>"111011110",
    506=>"000100000",
    507=>"111111000",
    508=>"110000010",
    509=>"111101000",
    510=>"110110000",
    511=>"000011000",
    512=>"100111011",
    513=>"110111011",
    514=>"000000000",
    515=>"010111011",
    516=>"000000011",
    517=>"000000000",
    518=>"111111111",
    519=>"111111111",
    520=>"000000000",
    521=>"010110101",
    522=>"111110101",
    523=>"100000000",
    524=>"010111000",
    525=>"101011010",
    526=>"100000000",
    527=>"000110000",
    528=>"111011100",
    529=>"011110000",
    530=>"000000000",
    531=>"101101000",
    532=>"000000101",
    533=>"000000000",
    534=>"001001011",
    535=>"110100110",
    536=>"001011011",
    537=>"011100000",
    538=>"111111111",
    539=>"110110110",
    540=>"100101110",
    541=>"000000000",
    542=>"000000000",
    543=>"100100001",
    544=>"110100011",
    545=>"010110000",
    546=>"100100101",
    547=>"101011101",
    548=>"010111001",
    549=>"000000000",
    550=>"111111000",
    551=>"000000000",
    552=>"111111111",
    553=>"010010000",
    554=>"000100010",
    555=>"001000101",
    556=>"100000010",
    557=>"110111011",
    558=>"100100100",
    559=>"111111100",
    560=>"100100100",
    561=>"110110000",
    562=>"000000001",
    563=>"001011100",
    564=>"000111001",
    565=>"010101001",
    566=>"000110110",
    567=>"100000001",
    568=>"011110000",
    569=>"110100000",
    570=>"100100100",
    571=>"110110111",
    572=>"001000010",
    573=>"000000000",
    574=>"110111111",
    575=>"011000001",
    576=>"100000100",
    577=>"000000010",
    578=>"011101111",
    579=>"000111111",
    580=>"000110110",
    581=>"000000100",
    582=>"111111111",
    583=>"100000110",
    584=>"111110110",
    585=>"010010010",
    586=>"110011011",
    587=>"101111101",
    588=>"110111111",
    589=>"010000100",
    590=>"011011101",
    591=>"000111101",
    592=>"001110111",
    593=>"000101101",
    594=>"000100011",
    595=>"110101110",
    596=>"001000000",
    597=>"011111011",
    598=>"101101000",
    599=>"010010100",
    600=>"001000000",
    601=>"111110100",
    602=>"001000100",
    603=>"111010010",
    604=>"111110010",
    605=>"100000000",
    606=>"011111100",
    607=>"011011000",
    608=>"101001111",
    609=>"010001000",
    610=>"001001100",
    611=>"100000100",
    612=>"000000000",
    613=>"100100011",
    614=>"100100000",
    615=>"000101011",
    616=>"111110111",
    617=>"011010010",
    618=>"011001001",
    619=>"001000000",
    620=>"100000001",
    621=>"011110011",
    622=>"100000011",
    623=>"110100100",
    624=>"001111000",
    625=>"000000010",
    626=>"001000101",
    627=>"111110110",
    628=>"010011000",
    629=>"111001001",
    630=>"111111111",
    631=>"100000100",
    632=>"000110100",
    633=>"110111001",
    634=>"001101111",
    635=>"110110100",
    636=>"101101101",
    637=>"000000001",
    638=>"001101101",
    639=>"100100000",
    640=>"111010000",
    641=>"110111111",
    642=>"110110111",
    643=>"110111111",
    644=>"111101110",
    645=>"101100110",
    646=>"111111011",
    647=>"001000101",
    648=>"110110001",
    649=>"011000100",
    650=>"011001111",
    651=>"000000000",
    652=>"101101101",
    653=>"111100010",
    654=>"111111011",
    655=>"011001001",
    656=>"000100110",
    657=>"000000000",
    658=>"000110010",
    659=>"100001110",
    660=>"111100010",
    661=>"000000110",
    662=>"000100101",
    663=>"111111111",
    664=>"001100110",
    665=>"001101101",
    666=>"010101111",
    667=>"111000101",
    668=>"000110111",
    669=>"110100000",
    670=>"110010001",
    671=>"100100001",
    672=>"000100111",
    673=>"111000111",
    674=>"011100110",
    675=>"001100100",
    676=>"111111110",
    677=>"111110010",
    678=>"101000110",
    679=>"110111111",
    680=>"111111110",
    681=>"111011000",
    682=>"100100111",
    683=>"011101101",
    684=>"111000001",
    685=>"000000111",
    686=>"000100111",
    687=>"110110010",
    688=>"111111001",
    689=>"100101001",
    690=>"000111101",
    691=>"100010110",
    692=>"111001000",
    693=>"110110110",
    694=>"111001000",
    695=>"000000100",
    696=>"000000000",
    697=>"100100111",
    698=>"010010100",
    699=>"111101000",
    700=>"100101111",
    701=>"000000011",
    702=>"110011101",
    703=>"111101000",
    704=>"110110111",
    705=>"011000011",
    706=>"010000001",
    707=>"100000000",
    708=>"001011010",
    709=>"111111111",
    710=>"111011001",
    711=>"111011111",
    712=>"000011000",
    713=>"000000000",
    714=>"000110000",
    715=>"111111100",
    716=>"000111010",
    717=>"110010010",
    718=>"110111011",
    719=>"000000000",
    720=>"111111111",
    721=>"000000100",
    722=>"111111111",
    723=>"111111101",
    724=>"110110111",
    725=>"111011010",
    726=>"111111111",
    727=>"011011110",
    728=>"111111111",
    729=>"001000111",
    730=>"111111111",
    731=>"111110100",
    732=>"111111111",
    733=>"101101001",
    734=>"111111110",
    735=>"111000000",
    736=>"111111111",
    737=>"000010011",
    738=>"111111111",
    739=>"000000011",
    740=>"111111111",
    741=>"111111111",
    742=>"000011110",
    743=>"111111011",
    744=>"111111111",
    745=>"000000000",
    746=>"011001011",
    747=>"111111000",
    748=>"111111111",
    749=>"111110101",
    750=>"110100111",
    751=>"111011111",
    752=>"000000110",
    753=>"010011100",
    754=>"111111111",
    755=>"111111101",
    756=>"000110111",
    757=>"111111011",
    758=>"111110110",
    759=>"100111110",
    760=>"110110101",
    761=>"110111100",
    762=>"111111110",
    763=>"111110111",
    764=>"111111111",
    765=>"000000001",
    766=>"111110111",
    767=>"111110010",
    768=>"111101111",
    769=>"000010010",
    770=>"000110010",
    771=>"010010010",
    772=>"111111111",
    773=>"010000100",
    774=>"011100011",
    775=>"110111101",
    776=>"111111111",
    777=>"100100111",
    778=>"111111111",
    779=>"011001100",
    780=>"111111110",
    781=>"000000011",
    782=>"000000011",
    783=>"101001001",
    784=>"111100110",
    785=>"111101000",
    786=>"011001100",
    787=>"110001011",
    788=>"111111111",
    789=>"000000111",
    790=>"000000000",
    791=>"110110010",
    792=>"101111111",
    793=>"111001011",
    794=>"110000001",
    795=>"100000001",
    796=>"100000000",
    797=>"111000101",
    798=>"001000110",
    799=>"011001000",
    800=>"000111101",
    801=>"000000000",
    802=>"000000000",
    803=>"010111101",
    804=>"111111111",
    805=>"001000110",
    806=>"000000000",
    807=>"000000010",
    808=>"000010011",
    809=>"000001111",
    810=>"011000111",
    811=>"111010010",
    812=>"001101111",
    813=>"111100001",
    814=>"000000000",
    815=>"111111111",
    816=>"111111000",
    817=>"111111111",
    818=>"111001000",
    819=>"010001110",
    820=>"110110010",
    821=>"100001100",
    822=>"000100111",
    823=>"000111000",
    824=>"110000000",
    825=>"000100011",
    826=>"110110101",
    827=>"100101010",
    828=>"101000000",
    829=>"001110001",
    830=>"000001000",
    831=>"000000111",
    832=>"100100000",
    833=>"110110110",
    834=>"011011010",
    835=>"000110110",
    836=>"001110110",
    837=>"000101101",
    838=>"110110111",
    839=>"100000000",
    840=>"011011111",
    841=>"001011010",
    842=>"100110110",
    843=>"011011011",
    844=>"110111111",
    845=>"000010000",
    846=>"100100000",
    847=>"000000010",
    848=>"100111111",
    849=>"000000000",
    850=>"010100110",
    851=>"010111110",
    852=>"111001001",
    853=>"000000110",
    854=>"101001001",
    855=>"000000110",
    856=>"111001000",
    857=>"110110000",
    858=>"001001001",
    859=>"000011011",
    860=>"101000000",
    861=>"001011000",
    862=>"000111010",
    863=>"110111111",
    864=>"111001001",
    865=>"100111110",
    866=>"111101101",
    867=>"110000011",
    868=>"000000000",
    869=>"111000111",
    870=>"110111111",
    871=>"010110111",
    872=>"100111111",
    873=>"010111110",
    874=>"011111001",
    875=>"001000101",
    876=>"001011000",
    877=>"010110000",
    878=>"101001001",
    879=>"110110001",
    880=>"011111111",
    881=>"110101101",
    882=>"011000000",
    883=>"100010000",
    884=>"000111110",
    885=>"011110010",
    886=>"001011111",
    887=>"000000000",
    888=>"010000001",
    889=>"000000110",
    890=>"010001111",
    891=>"001000000",
    892=>"110000101",
    893=>"110000000",
    894=>"100111111",
    895=>"110111001",
    896=>"100101011",
    897=>"010111111",
    898=>"110011010",
    899=>"000111111",
    900=>"111110000",
    901=>"000001101",
    902=>"000000001",
    903=>"110100111",
    904=>"111000000",
    905=>"111111000",
    906=>"111110000",
    907=>"001111111",
    908=>"111110000",
    909=>"010000000",
    910=>"111011001",
    911=>"101111111",
    912=>"000000000",
    913=>"101001111",
    914=>"001100111",
    915=>"100000000",
    916=>"001000100",
    917=>"101111011",
    918=>"111101111",
    919=>"110010000",
    920=>"000100000",
    921=>"111001111",
    922=>"111001101",
    923=>"000000110",
    924=>"111000000",
    925=>"101000111",
    926=>"000000000",
    927=>"111101101",
    928=>"111011011",
    929=>"000011111",
    930=>"000000011",
    931=>"101100100",
    932=>"111111111",
    933=>"101100100",
    934=>"000011111",
    935=>"101111100",
    936=>"010001000",
    937=>"000000000",
    938=>"110110110",
    939=>"111000001",
    940=>"000001101",
    941=>"110000001",
    942=>"111100111",
    943=>"111000001",
    944=>"111100000",
    945=>"111000100",
    946=>"101000100",
    947=>"000111111",
    948=>"000010111",
    949=>"001001101",
    950=>"100110111",
    951=>"000111000",
    952=>"011011111",
    953=>"000001011",
    954=>"111000000",
    955=>"100000001",
    956=>"000000011",
    957=>"101001001",
    958=>"101010000",
    959=>"101001111",
    960=>"110100100",
    961=>"011101110",
    962=>"100101001",
    963=>"111111111",
    964=>"001101100",
    965=>"110011011",
    966=>"101011011",
    967=>"111001000",
    968=>"011111111",
    969=>"110000000",
    970=>"100101011",
    971=>"000000000",
    972=>"111110111",
    973=>"010011000",
    974=>"000000000",
    975=>"010010111",
    976=>"000110010",
    977=>"000000111",
    978=>"110110110",
    979=>"000100111",
    980=>"001000100",
    981=>"101101111",
    982=>"000000101",
    983=>"000000000",
    984=>"000001101",
    985=>"110100000",
    986=>"001111110",
    987=>"101000001",
    988=>"000000111",
    989=>"100000000",
    990=>"111111111",
    991=>"101000101",
    992=>"001001110",
    993=>"001000101",
    994=>"000011101",
    995=>"001100100",
    996=>"000010100",
    997=>"111010011",
    998=>"001100001",
    999=>"001110111",
    1000=>"111111011",
    1001=>"111111010",
    1002=>"100000100",
    1003=>"000000000",
    1004=>"001011100",
    1005=>"000000001",
    1006=>"000000101",
    1007=>"011111101",
    1008=>"111111111",
    1009=>"010001110",
    1010=>"000010100",
    1011=>"111111010",
    1012=>"111111111",
    1013=>"000000101",
    1014=>"111111111",
    1015=>"000000100",
    1016=>"000000000",
    1017=>"101000101",
    1018=>"111011011",
    1019=>"000000000",
    1020=>"000101111",
    1021=>"000000001",
    1022=>"110111111",
    1023=>"100000101",
    1024=>"001000000",
    1025=>"111111111",
    1026=>"000000000",
    1027=>"010111010",
    1028=>"110000001",
    1029=>"111101111",
    1030=>"011111111",
    1031=>"000000000",
    1032=>"111111111",
    1033=>"000111110",
    1034=>"101111111",
    1035=>"100000111",
    1036=>"010111110",
    1037=>"000111101",
    1038=>"001000001",
    1039=>"001001000",
    1040=>"110110111",
    1041=>"111001101",
    1042=>"000000001",
    1043=>"110101111",
    1044=>"100111000",
    1045=>"000101001",
    1046=>"011000000",
    1047=>"110111111",
    1048=>"101000100",
    1049=>"001000101",
    1050=>"001101111",
    1051=>"000101101",
    1052=>"111000111",
    1053=>"111000111",
    1054=>"110111111",
    1055=>"101000000",
    1056=>"111111111",
    1057=>"110111111",
    1058=>"111111111",
    1059=>"101000100",
    1060=>"111101101",
    1061=>"001000000",
    1062=>"111111110",
    1063=>"000000000",
    1064=>"000000000",
    1065=>"000000000",
    1066=>"100111111",
    1067=>"010110111",
    1068=>"000001001",
    1069=>"001001110",
    1070=>"111111111",
    1071=>"100110101",
    1072=>"110100100",
    1073=>"000111101",
    1074=>"001001111",
    1075=>"000000011",
    1076=>"011111110",
    1077=>"001000000",
    1078=>"000000000",
    1079=>"101100000",
    1080=>"111111111",
    1081=>"000000000",
    1082=>"100001001",
    1083=>"001000000",
    1084=>"001000000",
    1085=>"101000101",
    1086=>"000000000",
    1087=>"110111000",
    1088=>"111111111",
    1089=>"000000000",
    1090=>"000000110",
    1091=>"011011011",
    1092=>"111011011",
    1093=>"000000001",
    1094=>"000000000",
    1095=>"011111111",
    1096=>"000000000",
    1097=>"111010110",
    1098=>"111111110",
    1099=>"000000000",
    1100=>"000110110",
    1101=>"000000010",
    1102=>"101000001",
    1103=>"011111010",
    1104=>"000000000",
    1105=>"111111111",
    1106=>"000000000",
    1107=>"110000001",
    1108=>"000000000",
    1109=>"000000000",
    1110=>"000100111",
    1111=>"111000011",
    1112=>"000000111",
    1113=>"111110100",
    1114=>"000000110",
    1115=>"111111111",
    1116=>"111100100",
    1117=>"011010110",
    1118=>"000000000",
    1119=>"100100110",
    1120=>"100000001",
    1121=>"100000000",
    1122=>"000000000",
    1123=>"111111110",
    1124=>"000001000",
    1125=>"111100100",
    1126=>"111111111",
    1127=>"000000000",
    1128=>"011111111",
    1129=>"011111011",
    1130=>"000000100",
    1131=>"110100100",
    1132=>"111111011",
    1133=>"111111111",
    1134=>"001011111",
    1135=>"000000000",
    1136=>"011000000",
    1137=>"101000001",
    1138=>"111111011",
    1139=>"111111110",
    1140=>"110111110",
    1141=>"111111111",
    1142=>"111111111",
    1143=>"110100001",
    1144=>"100100001",
    1145=>"110100101",
    1146=>"110101101",
    1147=>"111111011",
    1148=>"110111111",
    1149=>"000000000",
    1150=>"111111111",
    1151=>"101101001",
    1152=>"111001100",
    1153=>"001111000",
    1154=>"000000101",
    1155=>"000000101",
    1156=>"100110110",
    1157=>"100011001",
    1158=>"110111100",
    1159=>"011100100",
    1160=>"111101011",
    1161=>"010000000",
    1162=>"001101101",
    1163=>"110111011",
    1164=>"000111010",
    1165=>"001001001",
    1166=>"100110011",
    1167=>"011001100",
    1168=>"000000001",
    1169=>"001000101",
    1170=>"100110011",
    1171=>"001001001",
    1172=>"110110010",
    1173=>"000000000",
    1174=>"000110111",
    1175=>"001111111",
    1176=>"000000110",
    1177=>"000000000",
    1178=>"001001111",
    1179=>"100111100",
    1180=>"010110111",
    1181=>"000000001",
    1182=>"111111111",
    1183=>"111111111",
    1184=>"100100101",
    1185=>"111111110",
    1186=>"000111000",
    1187=>"000100101",
    1188=>"000100000",
    1189=>"111011011",
    1190=>"111111100",
    1191=>"100001101",
    1192=>"111111000",
    1193=>"111101000",
    1194=>"000110010",
    1195=>"000110111",
    1196=>"111111011",
    1197=>"111111100",
    1198=>"000110010",
    1199=>"100101010",
    1200=>"110111110",
    1201=>"011001011",
    1202=>"000000011",
    1203=>"110111110",
    1204=>"110110110",
    1205=>"110111001",
    1206=>"101100111",
    1207=>"001001111",
    1208=>"000111011",
    1209=>"000010110",
    1210=>"011111100",
    1211=>"011100100",
    1212=>"011001111",
    1213=>"001000101",
    1214=>"001000011",
    1215=>"001000110",
    1216=>"101000011",
    1217=>"010110011",
    1218=>"011100011",
    1219=>"110110000",
    1220=>"001101011",
    1221=>"001100101",
    1222=>"000111000",
    1223=>"101011111",
    1224=>"011001100",
    1225=>"000001111",
    1226=>"001010110",
    1227=>"010101111",
    1228=>"111111111",
    1229=>"110110000",
    1230=>"011101000",
    1231=>"111000010",
    1232=>"000110110",
    1233=>"011011111",
    1234=>"000001110",
    1235=>"000000110",
    1236=>"110100100",
    1237=>"101000000",
    1238=>"001101111",
    1239=>"000000110",
    1240=>"001011111",
    1241=>"011101011",
    1242=>"001011111",
    1243=>"011011011",
    1244=>"000001011",
    1245=>"001001110",
    1246=>"100000100",
    1247=>"110110000",
    1248=>"000010011",
    1249=>"011100110",
    1250=>"000000010",
    1251=>"001001101",
    1252=>"111100000",
    1253=>"011111100",
    1254=>"100101111",
    1255=>"011110110",
    1256=>"111011001",
    1257=>"110001000",
    1258=>"010001110",
    1259=>"111110000",
    1260=>"001001001",
    1261=>"001000010",
    1262=>"001001110",
    1263=>"110111010",
    1264=>"001001011",
    1265=>"001001111",
    1266=>"011001111",
    1267=>"000000101",
    1268=>"100110110",
    1269=>"001001010",
    1270=>"110010000",
    1271=>"000000000",
    1272=>"100000111",
    1273=>"001101011",
    1274=>"000001001",
    1275=>"001011001",
    1276=>"001001111",
    1277=>"001011111",
    1278=>"101110001",
    1279=>"110110000",
    1280=>"110110101",
    1281=>"000011100",
    1282=>"000000000",
    1283=>"110110100",
    1284=>"000000000",
    1285=>"111000000",
    1286=>"110111111",
    1287=>"000000000",
    1288=>"100000100",
    1289=>"100001001",
    1290=>"111111111",
    1291=>"000000100",
    1292=>"111111011",
    1293=>"011001000",
    1294=>"001101000",
    1295=>"111010011",
    1296=>"111110110",
    1297=>"000000001",
    1298=>"011100100",
    1299=>"001000011",
    1300=>"000100100",
    1301=>"011001001",
    1302=>"110000001",
    1303=>"000100011",
    1304=>"000001001",
    1305=>"001001101",
    1306=>"000010000",
    1307=>"111000001",
    1308=>"001100011",
    1309=>"011011010",
    1310=>"111111110",
    1311=>"100100100",
    1312=>"100110100",
    1313=>"111111111",
    1314=>"011101011",
    1315=>"011001001",
    1316=>"111111111",
    1317=>"000110000",
    1318=>"000000000",
    1319=>"011011111",
    1320=>"111111110",
    1321=>"000100000",
    1322=>"011001100",
    1323=>"111000111",
    1324=>"101101101",
    1325=>"111101101",
    1326=>"100110010",
    1327=>"111111101",
    1328=>"110110110",
    1329=>"000000001",
    1330=>"011000001",
    1331=>"111111110",
    1332=>"010110010",
    1333=>"000000000",
    1334=>"001101000",
    1335=>"101100000",
    1336=>"010110111",
    1337=>"100100000",
    1338=>"110111111",
    1339=>"110111111",
    1340=>"110010011",
    1341=>"000010000",
    1342=>"001001001",
    1343=>"001001000",
    1344=>"000000000",
    1345=>"000000000",
    1346=>"100010001",
    1347=>"001001111",
    1348=>"000000000",
    1349=>"111000111",
    1350=>"111111111",
    1351=>"100001011",
    1352=>"111001010",
    1353=>"000000000",
    1354=>"000000000",
    1355=>"101000000",
    1356=>"101101111",
    1357=>"101111111",
    1358=>"000101100",
    1359=>"100110110",
    1360=>"011110110",
    1361=>"111001000",
    1362=>"000100100",
    1363=>"100100111",
    1364=>"100000000",
    1365=>"111111111",
    1366=>"001000000",
    1367=>"111011101",
    1368=>"111011011",
    1369=>"000000000",
    1370=>"110000011",
    1371=>"101111000",
    1372=>"000101000",
    1373=>"111000100",
    1374=>"111111111",
    1375=>"000100111",
    1376=>"000111111",
    1377=>"000000000",
    1378=>"001000000",
    1379=>"000000000",
    1380=>"111001101",
    1381=>"001100100",
    1382=>"000000000",
    1383=>"100010010",
    1384=>"000001000",
    1385=>"000100000",
    1386=>"011101110",
    1387=>"000000000",
    1388=>"000000000",
    1389=>"111000111",
    1390=>"000000000",
    1391=>"111111110",
    1392=>"111100100",
    1393=>"000000000",
    1394=>"111011000",
    1395=>"111011111",
    1396=>"100111101",
    1397=>"000000000",
    1398=>"000000000",
    1399=>"100111111",
    1400=>"001100001",
    1401=>"111001001",
    1402=>"101010000",
    1403=>"100001000",
    1404=>"000011010",
    1405=>"000010010",
    1406=>"110111111",
    1407=>"000000000",
    1408=>"111011101",
    1409=>"011110111",
    1410=>"010000111",
    1411=>"101101101",
    1412=>"011111101",
    1413=>"110110100",
    1414=>"111011011",
    1415=>"011001001",
    1416=>"111100101",
    1417=>"001001111",
    1418=>"001011111",
    1419=>"111100100",
    1420=>"110000111",
    1421=>"011010011",
    1422=>"101100100",
    1423=>"011001001",
    1424=>"010110110",
    1425=>"110100000",
    1426=>"000001001",
    1427=>"011011011",
    1428=>"000110100",
    1429=>"000000000",
    1430=>"100111111",
    1431=>"000111111",
    1432=>"100110110",
    1433=>"110110010",
    1434=>"011011011",
    1435=>"001011010",
    1436=>"110010110",
    1437=>"000100111",
    1438=>"100100100",
    1439=>"101000010",
    1440=>"011001001",
    1441=>"110101100",
    1442=>"100110110",
    1443=>"001010001",
    1444=>"100100100",
    1445=>"100100111",
    1446=>"011011011",
    1447=>"111001001",
    1448=>"000000110",
    1449=>"100100000",
    1450=>"101100011",
    1451=>"100000010",
    1452=>"101100000",
    1453=>"100001001",
    1454=>"001001101",
    1455=>"000000011",
    1456=>"010010110",
    1457=>"010010111",
    1458=>"100100000",
    1459=>"111100100",
    1460=>"110011111",
    1461=>"001001000",
    1462=>"111001000",
    1463=>"110000000",
    1464=>"000011011",
    1465=>"101101001",
    1466=>"101101100",
    1467=>"101001001",
    1468=>"110111000",
    1469=>"110100100",
    1470=>"111000100",
    1471=>"001101111",
    1472=>"100111011",
    1473=>"111111011",
    1474=>"111101110",
    1475=>"011001111",
    1476=>"001110110",
    1477=>"000110110",
    1478=>"010101101",
    1479=>"110100101",
    1480=>"011000110",
    1481=>"101001000",
    1482=>"100011011",
    1483=>"001110100",
    1484=>"000101111",
    1485=>"011011000",
    1486=>"001111100",
    1487=>"100000100",
    1488=>"010000111",
    1489=>"010000110",
    1490=>"001100100",
    1491=>"110010001",
    1492=>"000000000",
    1493=>"010010000",
    1494=>"011010111",
    1495=>"011000001",
    1496=>"000000000",
    1497=>"010000000",
    1498=>"100000001",
    1499=>"100000101",
    1500=>"111111000",
    1501=>"101100111",
    1502=>"010111111",
    1503=>"000011000",
    1504=>"000000101",
    1505=>"111001001",
    1506=>"001010010",
    1507=>"000000101",
    1508=>"000000000",
    1509=>"000110110",
    1510=>"111111110",
    1511=>"011111101",
    1512=>"101000011",
    1513=>"000000010",
    1514=>"011000010",
    1515=>"000011011",
    1516=>"110111100",
    1517=>"100011001",
    1518=>"100100100",
    1519=>"110110000",
    1520=>"000010001",
    1521=>"011000000",
    1522=>"011001000",
    1523=>"110110010",
    1524=>"110101000",
    1525=>"100001001",
    1526=>"001011100",
    1527=>"000001000",
    1528=>"110010011",
    1529=>"110111001",
    1530=>"110011111",
    1531=>"110110001",
    1532=>"000010111",
    1533=>"000000100",
    1534=>"110111111",
    1535=>"010111000",
    1536=>"001101000",
    1537=>"011100010",
    1538=>"001000110",
    1539=>"101101100",
    1540=>"100110110",
    1541=>"001000001",
    1542=>"000100110",
    1543=>"111001101",
    1544=>"000000010",
    1545=>"011001011",
    1546=>"000100110",
    1547=>"000100100",
    1548=>"111111000",
    1549=>"011101110",
    1550=>"100110011",
    1551=>"011011010",
    1552=>"000100011",
    1553=>"011001001",
    1554=>"100110000",
    1555=>"000110111",
    1556=>"000001000",
    1557=>"100100110",
    1558=>"011011011",
    1559=>"100110011",
    1560=>"001001001",
    1561=>"011001011",
    1562=>"001001101",
    1563=>"100010110",
    1564=>"100111001",
    1565=>"011011001",
    1566=>"011001110",
    1567=>"001001011",
    1568=>"100100100",
    1569=>"000100100",
    1570=>"110110011",
    1571=>"001001100",
    1572=>"110011001",
    1573=>"101000010",
    1574=>"000001000",
    1575=>"000100110",
    1576=>"000110100",
    1577=>"000000011",
    1578=>"111110011",
    1579=>"011000001",
    1580=>"101010011",
    1581=>"100110110",
    1582=>"110111100",
    1583=>"000000110",
    1584=>"110011011",
    1585=>"100100000",
    1586=>"000100010",
    1587=>"100001000",
    1588=>"110001001",
    1589=>"000000100",
    1590=>"110110011",
    1591=>"100100110",
    1592=>"001100110",
    1593=>"100001100",
    1594=>"100110010",
    1595=>"101001011",
    1596=>"111010011",
    1597=>"010001011",
    1598=>"110101101",
    1599=>"000100100",
    1600=>"000001100",
    1601=>"111011110",
    1602=>"011000001",
    1603=>"011001011",
    1604=>"001011011",
    1605=>"001001001",
    1606=>"110110110",
    1607=>"000110110",
    1608=>"001001001",
    1609=>"011001001",
    1610=>"100100110",
    1611=>"001001001",
    1612=>"111000011",
    1613=>"111010010",
    1614=>"000001001",
    1615=>"100100101",
    1616=>"011011011",
    1617=>"000110011",
    1618=>"000000001",
    1619=>"110110110",
    1620=>"100001000",
    1621=>"000000111",
    1622=>"111111111",
    1623=>"110110100",
    1624=>"111010010",
    1625=>"111110110",
    1626=>"110110110",
    1627=>"110110101",
    1628=>"001111000",
    1629=>"111001001",
    1630=>"001011011",
    1631=>"000001010",
    1632=>"001100100",
    1633=>"001011111",
    1634=>"011011001",
    1635=>"101110110",
    1636=>"000001000",
    1637=>"100001001",
    1638=>"111110110",
    1639=>"000000000",
    1640=>"000000101",
    1641=>"100100101",
    1642=>"011011001",
    1643=>"010010010",
    1644=>"011110100",
    1645=>"100100110",
    1646=>"101100000",
    1647=>"001000110",
    1648=>"100100110",
    1649=>"000110110",
    1650=>"001011011",
    1651=>"010010000",
    1652=>"001010111",
    1653=>"000000101",
    1654=>"000000001",
    1655=>"100010011",
    1656=>"100110101",
    1657=>"100100101",
    1658=>"000000010",
    1659=>"100100100",
    1660=>"000100111",
    1661=>"000001011",
    1662=>"000101100",
    1663=>"000010001",
    1664=>"011010010",
    1665=>"111011011",
    1666=>"100100100",
    1667=>"101101001",
    1668=>"110100100",
    1669=>"001001101",
    1670=>"110100111",
    1671=>"010110100",
    1672=>"101100011",
    1673=>"111111000",
    1674=>"100100100",
    1675=>"010010110",
    1676=>"101000101",
    1677=>"110100111",
    1678=>"110010110",
    1679=>"100100100",
    1680=>"000000100",
    1681=>"001001001",
    1682=>"001001000",
    1683=>"000100001",
    1684=>"011011011",
    1685=>"011010010",
    1686=>"011011011",
    1687=>"001011010",
    1688=>"001011000",
    1689=>"010010010",
    1690=>"100110010",
    1691=>"110110110",
    1692=>"100100110",
    1693=>"001001011",
    1694=>"011000110",
    1695=>"011110000",
    1696=>"100100100",
    1697=>"000011110",
    1698=>"011010011",
    1699=>"000000111",
    1700=>"001001001",
    1701=>"001100000",
    1702=>"111001011",
    1703=>"100000111",
    1704=>"010010100",
    1705=>"011000000",
    1706=>"101010010",
    1707=>"011011011",
    1708=>"011010010",
    1709=>"111100000",
    1710=>"100100100",
    1711=>"010000100",
    1712=>"111011011",
    1713=>"000011110",
    1714=>"101110110",
    1715=>"110101110",
    1716=>"110110100",
    1717=>"010110111",
    1718=>"111110110",
    1719=>"011011111",
    1720=>"011001011",
    1721=>"010110000",
    1722=>"011010110",
    1723=>"010110100",
    1724=>"100100101",
    1725=>"001001001",
    1726=>"111110100",
    1727=>"110000100",
    1728=>"111001000",
    1729=>"011110110",
    1730=>"111110110",
    1731=>"001111111",
    1732=>"101111001",
    1733=>"000110111",
    1734=>"111111110",
    1735=>"011101001",
    1736=>"100011101",
    1737=>"011000110",
    1738=>"101011000",
    1739=>"011101110",
    1740=>"111111111",
    1741=>"011000000",
    1742=>"000010000",
    1743=>"110011000",
    1744=>"111110110",
    1745=>"001000111",
    1746=>"110010100",
    1747=>"111000000",
    1748=>"011000100",
    1749=>"101111001",
    1750=>"000000000",
    1751=>"111011111",
    1752=>"010000101",
    1753=>"000100000",
    1754=>"110010111",
    1755=>"110100111",
    1756=>"000000000",
    1757=>"011111010",
    1758=>"110111111",
    1759=>"000000110",
    1760=>"110111000",
    1761=>"011001000",
    1762=>"010011000",
    1763=>"100000100",
    1764=>"111111101",
    1765=>"001111110",
    1766=>"110000001",
    1767=>"001100110",
    1768=>"110111111",
    1769=>"011111000",
    1770=>"001001011",
    1771=>"100000000",
    1772=>"110110000",
    1773=>"111111111",
    1774=>"111000111",
    1775=>"110010000",
    1776=>"000101111",
    1777=>"000000000",
    1778=>"101000111",
    1779=>"101010001",
    1780=>"011010000",
    1781=>"100101100",
    1782=>"001001100",
    1783=>"000011000",
    1784=>"000000000",
    1785=>"111100001",
    1786=>"011011010",
    1787=>"000000000",
    1788=>"000001011",
    1789=>"010000001",
    1790=>"100011001",
    1791=>"010010000",
    1792=>"101000111",
    1793=>"101101001",
    1794=>"000001011",
    1795=>"111111111",
    1796=>"101101001",
    1797=>"011000100",
    1798=>"111001010",
    1799=>"001000001",
    1800=>"001000011",
    1801=>"011000000",
    1802=>"001001111",
    1803=>"000000000",
    1804=>"101100101",
    1805=>"000101111",
    1806=>"111111111",
    1807=>"110100100",
    1808=>"000101110",
    1809=>"111100100",
    1810=>"100111111",
    1811=>"011011011",
    1812=>"000000001",
    1813=>"000000000",
    1814=>"100100100",
    1815=>"000000000",
    1816=>"100100111",
    1817=>"100100100",
    1818=>"000000111",
    1819=>"000000000",
    1820=>"110110100",
    1821=>"101101110",
    1822=>"001001010",
    1823=>"000001011",
    1824=>"100110001",
    1825=>"001001000",
    1826=>"000100111",
    1827=>"111111100",
    1828=>"000110000",
    1829=>"000110000",
    1830=>"101100101",
    1831=>"010111111",
    1832=>"111110111",
    1833=>"011011111",
    1834=>"100000100",
    1835=>"100000000",
    1836=>"011011111",
    1837=>"110110110",
    1838=>"100100100",
    1839=>"100111110",
    1840=>"111111111",
    1841=>"000100000",
    1842=>"110100100",
    1843=>"000010000",
    1844=>"001001011",
    1845=>"000001101",
    1846=>"010101011",
    1847=>"000100001",
    1848=>"011011111",
    1849=>"111111111",
    1850=>"011101011",
    1851=>"000000000",
    1852=>"000001111",
    1853=>"110100000",
    1854=>"001000010",
    1855=>"101111110",
    1856=>"001000100",
    1857=>"100100000",
    1858=>"111111011",
    1859=>"111011000",
    1860=>"111011111",
    1861=>"110001000",
    1862=>"001100100",
    1863=>"000000000",
    1864=>"111001001",
    1865=>"111100110",
    1866=>"000000110",
    1867=>"101111011",
    1868=>"111011101",
    1869=>"111100101",
    1870=>"111011101",
    1871=>"000000101",
    1872=>"111100110",
    1873=>"110011000",
    1874=>"101111001",
    1875=>"000000100",
    1876=>"001111100",
    1877=>"001000101",
    1878=>"111011001",
    1879=>"100100100",
    1880=>"101101111",
    1881=>"001001000",
    1882=>"100000000",
    1883=>"001000100",
    1884=>"110111101",
    1885=>"110011001",
    1886=>"111111110",
    1887=>"011001100",
    1888=>"001100110",
    1889=>"111011011",
    1890=>"111110110",
    1891=>"000110011",
    1892=>"110011100",
    1893=>"000001001",
    1894=>"000100100",
    1895=>"001001111",
    1896=>"001100011",
    1897=>"000000100",
    1898=>"111011101",
    1899=>"111100100",
    1900=>"001100111",
    1901=>"001100100",
    1902=>"010011011",
    1903=>"001101111",
    1904=>"111011101",
    1905=>"100100100",
    1906=>"100110011",
    1907=>"011101101",
    1908=>"111100100",
    1909=>"001000100",
    1910=>"001100111",
    1911=>"000000100",
    1912=>"000100100",
    1913=>"100100001",
    1914=>"000000000",
    1915=>"001000100",
    1916=>"000000000",
    1917=>"000000000",
    1918=>"000000000",
    1919=>"001101111",
    1920=>"101100100",
    1921=>"011011110",
    1922=>"100100100",
    1923=>"011011111",
    1924=>"000001101",
    1925=>"011001011",
    1926=>"110110100",
    1927=>"100100100",
    1928=>"011011001",
    1929=>"100100100",
    1930=>"000100111",
    1931=>"100110100",
    1932=>"001100001",
    1933=>"101100101",
    1934=>"100100100",
    1935=>"011011011",
    1936=>"110000100",
    1937=>"011011011",
    1938=>"000010000",
    1939=>"111001110",
    1940=>"110111100",
    1941=>"100000100",
    1942=>"111111111",
    1943=>"010011011",
    1944=>"100100100",
    1945=>"000000000",
    1946=>"010011010",
    1947=>"100010100",
    1948=>"001101101",
    1949=>"111110000",
    1950=>"111011110",
    1951=>"100100100",
    1952=>"001000001",
    1953=>"000001111",
    1954=>"011011000",
    1955=>"001001001",
    1956=>"010010010",
    1957=>"100100100",
    1958=>"010011010",
    1959=>"000011001",
    1960=>"100100100",
    1961=>"001001000",
    1962=>"010110110",
    1963=>"011010010",
    1964=>"100100100",
    1965=>"001100100",
    1966=>"101100100",
    1967=>"100111100",
    1968=>"010110110",
    1969=>"011010010",
    1970=>"010010100",
    1971=>"111111111",
    1972=>"000100100",
    1973=>"100100100",
    1974=>"100000100",
    1975=>"011011010",
    1976=>"011011010",
    1977=>"101101110",
    1978=>"000001001",
    1979=>"100111100",
    1980=>"010011011",
    1981=>"011011011",
    1982=>"000001000",
    1983=>"000000100",
    1984=>"011011100",
    1985=>"111001101",
    1986=>"110100001",
    1987=>"111111000",
    1988=>"111111011",
    1989=>"010000111",
    1990=>"111111111",
    1991=>"111010000",
    1992=>"000000101",
    1993=>"100101111",
    1994=>"111111010",
    1995=>"100101001",
    1996=>"111101101",
    1997=>"111100111",
    1998=>"001000000",
    1999=>"100001010",
    2000=>"111000000",
    2001=>"101000111",
    2002=>"111111101",
    2003=>"000000000",
    2004=>"111111101",
    2005=>"111010000",
    2006=>"111100101",
    2007=>"110010000",
    2008=>"011010000",
    2009=>"101011010",
    2010=>"100000011",
    2011=>"001001001",
    2012=>"000000000",
    2013=>"001000111",
    2014=>"011111111",
    2015=>"111101011",
    2016=>"111110000",
    2017=>"110011111",
    2018=>"000000000",
    2019=>"000000000",
    2020=>"010110101",
    2021=>"111100000",
    2022=>"000110111",
    2023=>"000000000",
    2024=>"011111011",
    2025=>"000000010",
    2026=>"100111110",
    2027=>"111110110",
    2028=>"001001000",
    2029=>"001011010",
    2030=>"111111000",
    2031=>"011111000",
    2032=>"110100001",
    2033=>"000000000",
    2034=>"111001101",
    2035=>"000000001",
    2036=>"000111111",
    2037=>"111100010",
    2038=>"010010001",
    2039=>"011011011",
    2040=>"000100100",
    2041=>"000111111",
    2042=>"011111011",
    2043=>"001011011",
    2044=>"010010100",
    2045=>"001010000",
    2046=>"000000000",
    2047=>"011010000",
    2048=>"000001101",
    2049=>"011111011",
    2050=>"110111110",
    2051=>"100110110",
    2052=>"100100110",
    2053=>"011111111",
    2054=>"110100100",
    2055=>"111101000",
    2056=>"110110110",
    2057=>"110100100",
    2058=>"100110100",
    2059=>"000100100",
    2060=>"001001101",
    2061=>"011100011",
    2062=>"110000100",
    2063=>"110110100",
    2064=>"101101010",
    2065=>"011011011",
    2066=>"000000100",
    2067=>"110000100",
    2068=>"000000100",
    2069=>"010001000",
    2070=>"001011011",
    2071=>"111101111",
    2072=>"001001001",
    2073=>"001011011",
    2074=>"011011000",
    2075=>"100101001",
    2076=>"011111011",
    2077=>"001101101",
    2078=>"011110111",
    2079=>"110100110",
    2080=>"110100100",
    2081=>"110110100",
    2082=>"000010001",
    2083=>"111000001",
    2084=>"110010100",
    2085=>"100110111",
    2086=>"100100100",
    2087=>"011000000",
    2088=>"010011011",
    2089=>"000110000",
    2090=>"011100101",
    2091=>"001001001",
    2092=>"001101101",
    2093=>"100000011",
    2094=>"110100110",
    2095=>"111100100",
    2096=>"100101001",
    2097=>"110000110",
    2098=>"000011011",
    2099=>"000111001",
    2100=>"101100100",
    2101=>"000000101",
    2102=>"100001101",
    2103=>"011010001",
    2104=>"111011011",
    2105=>"100101100",
    2106=>"100110111",
    2107=>"100100100",
    2108=>"011011011",
    2109=>"001001011",
    2110=>"011110110",
    2111=>"110100001",
    2112=>"100100100",
    2113=>"001011101",
    2114=>"111111111",
    2115=>"011111000",
    2116=>"111111111",
    2117=>"001001100",
    2118=>"001000001",
    2119=>"110111111",
    2120=>"111111111",
    2121=>"001011011",
    2122=>"011000001",
    2123=>"111111111",
    2124=>"011111011",
    2125=>"000111110",
    2126=>"110110110",
    2127=>"000111010",
    2128=>"111111010",
    2129=>"111110100",
    2130=>"101111110",
    2131=>"100000000",
    2132=>"000111111",
    2133=>"000110110",
    2134=>"111001000",
    2135=>"000000001",
    2136=>"000000000",
    2137=>"110100100",
    2138=>"110111111",
    2139=>"000001000",
    2140=>"000110110",
    2141=>"010110100",
    2142=>"010111111",
    2143=>"111111011",
    2144=>"001011011",
    2145=>"110110111",
    2146=>"000100110",
    2147=>"111001100",
    2148=>"110101110",
    2149=>"000000001",
    2150=>"001001000",
    2151=>"111111111",
    2152=>"000100110",
    2153=>"000000000",
    2154=>"001110111",
    2155=>"000000000",
    2156=>"000100010",
    2157=>"000000000",
    2158=>"011011011",
    2159=>"100100011",
    2160=>"000110110",
    2161=>"001000001",
    2162=>"000000000",
    2163=>"100000000",
    2164=>"011111011",
    2165=>"100000100",
    2166=>"100110110",
    2167=>"001001001",
    2168=>"001001001",
    2169=>"000111011",
    2170=>"000000000",
    2171=>"100000000",
    2172=>"110110110",
    2173=>"000000000",
    2174=>"000000001",
    2175=>"001111100",
    2176=>"100000000",
    2177=>"111111111",
    2178=>"011111111",
    2179=>"111011010",
    2180=>"000100011",
    2181=>"000000001",
    2182=>"000000000",
    2183=>"011110110",
    2184=>"011111111",
    2185=>"110110000",
    2186=>"000111111",
    2187=>"001000111",
    2188=>"111011011",
    2189=>"101110010",
    2190=>"101011110",
    2191=>"001011000",
    2192=>"000111011",
    2193=>"111111000",
    2194=>"000000000",
    2195=>"101111110",
    2196=>"000000000",
    2197=>"000000000",
    2198=>"000000011",
    2199=>"110101011",
    2200=>"000001111",
    2201=>"110000010",
    2202=>"100000000",
    2203=>"010001000",
    2204=>"001000010",
    2205=>"000000000",
    2206=>"001100100",
    2207=>"000000000",
    2208=>"000000000",
    2209=>"111111000",
    2210=>"111111111",
    2211=>"000000000",
    2212=>"000000000",
    2213=>"001101011",
    2214=>"111111010",
    2215=>"110111111",
    2216=>"001101110",
    2217=>"110110110",
    2218=>"100100100",
    2219=>"000000000",
    2220=>"111011001",
    2221=>"100000000",
    2222=>"000000111",
    2223=>"000000000",
    2224=>"111111010",
    2225=>"100110111",
    2226=>"101001011",
    2227=>"111111111",
    2228=>"011111010",
    2229=>"000000001",
    2230=>"100100100",
    2231=>"101000000",
    2232=>"111111010",
    2233=>"000001111",
    2234=>"000000001",
    2235=>"111101011",
    2236=>"000001110",
    2237=>"000000000",
    2238=>"111111111",
    2239=>"000000000",
    2240=>"111111111",
    2241=>"000001111",
    2242=>"110010111",
    2243=>"110111010",
    2244=>"101000000",
    2245=>"000110000",
    2246=>"111000010",
    2247=>"100000100",
    2248=>"010011110",
    2249=>"000000011",
    2250=>"000010110",
    2251=>"100000110",
    2252=>"110110111",
    2253=>"010111111",
    2254=>"101011011",
    2255=>"000000000",
    2256=>"000110010",
    2257=>"110110100",
    2258=>"101000000",
    2259=>"110111011",
    2260=>"110110001",
    2261=>"111111000",
    2262=>"101100101",
    2263=>"000110000",
    2264=>"000000000",
    2265=>"001001011",
    2266=>"010110000",
    2267=>"001011111",
    2268=>"000000000",
    2269=>"100000000",
    2270=>"000000110",
    2271=>"000000000",
    2272=>"110110110",
    2273=>"000010000",
    2274=>"111111110",
    2275=>"000000000",
    2276=>"110111110",
    2277=>"001000000",
    2278=>"000010000",
    2279=>"111111111",
    2280=>"000001101",
    2281=>"000000101",
    2282=>"100100110",
    2283=>"001000000",
    2284=>"111110111",
    2285=>"000000000",
    2286=>"111000000",
    2287=>"001001101",
    2288=>"000000000",
    2289=>"000111111",
    2290=>"111011011",
    2291=>"011111111",
    2292=>"101000101",
    2293=>"010100000",
    2294=>"111111110",
    2295=>"000000010",
    2296=>"111111111",
    2297=>"000111111",
    2298=>"101111110",
    2299=>"011111111",
    2300=>"011110000",
    2301=>"100000001",
    2302=>"111111111",
    2303=>"111111110",
    2304=>"101001110",
    2305=>"000100111",
    2306=>"111110010",
    2307=>"111010000",
    2308=>"010000111",
    2309=>"100110111",
    2310=>"000001111",
    2311=>"111001000",
    2312=>"111100111",
    2313=>"111011000",
    2314=>"010010011",
    2315=>"100110110",
    2316=>"111100000",
    2317=>"011010000",
    2318=>"001000100",
    2319=>"111111000",
    2320=>"000110111",
    2321=>"011000000",
    2322=>"000100110",
    2323=>"100000100",
    2324=>"000100111",
    2325=>"001000000",
    2326=>"000101111",
    2327=>"100000100",
    2328=>"000110110",
    2329=>"111010000",
    2330=>"000011111",
    2331=>"001001011",
    2332=>"000010010",
    2333=>"111011000",
    2334=>"000110111",
    2335=>"000100111",
    2336=>"000100111",
    2337=>"110010111",
    2338=>"000000000",
    2339=>"001011000",
    2340=>"010100111",
    2341=>"111110000",
    2342=>"001001111",
    2343=>"000100111",
    2344=>"101111111",
    2345=>"111110000",
    2346=>"110110010",
    2347=>"000000111",
    2348=>"110010001",
    2349=>"000101011",
    2350=>"101110100",
    2351=>"010000001",
    2352=>"100000111",
    2353=>"010000000",
    2354=>"000100111",
    2355=>"000010010",
    2356=>"000000111",
    2357=>"000000010",
    2358=>"001001100",
    2359=>"000100111",
    2360=>"000011111",
    2361=>"110000011",
    2362=>"100001111",
    2363=>"100001111",
    2364=>"000100111",
    2365=>"100111100",
    2366=>"000101111",
    2367=>"101001111",
    2368=>"101111110",
    2369=>"111111111",
    2370=>"110111111",
    2371=>"000110110",
    2372=>"111111011",
    2373=>"011110110",
    2374=>"000000010",
    2375=>"111111111",
    2376=>"101111011",
    2377=>"111111111",
    2378=>"110111110",
    2379=>"001001010",
    2380=>"010111111",
    2381=>"010001011",
    2382=>"111100101",
    2383=>"000110010",
    2384=>"001000111",
    2385=>"111111010",
    2386=>"110111101",
    2387=>"111111110",
    2388=>"111101100",
    2389=>"001001000",
    2390=>"100000111",
    2391=>"110100111",
    2392=>"111110100",
    2393=>"111111010",
    2394=>"110111111",
    2395=>"001001111",
    2396=>"111111111",
    2397=>"010111010",
    2398=>"010010111",
    2399=>"100100111",
    2400=>"101001001",
    2401=>"111111011",
    2402=>"111111111",
    2403=>"100001111",
    2404=>"111111111",
    2405=>"111111111",
    2406=>"111111011",
    2407=>"111111111",
    2408=>"101101100",
    2409=>"000000000",
    2410=>"011000100",
    2411=>"111110111",
    2412=>"101101001",
    2413=>"111111011",
    2414=>"000111110",
    2415=>"000000001",
    2416=>"010111111",
    2417=>"111101001",
    2418=>"111111111",
    2419=>"000010001",
    2420=>"000000001",
    2421=>"001101111",
    2422=>"001001011",
    2423=>"000000000",
    2424=>"101000000",
    2425=>"100100001",
    2426=>"100101101",
    2427=>"111101001",
    2428=>"110000110",
    2429=>"011011111",
    2430=>"111111011",
    2431=>"111001001",
    2432=>"101100100",
    2433=>"000000000",
    2434=>"111111111",
    2435=>"110110110",
    2436=>"111111111",
    2437=>"001001111",
    2438=>"000000000",
    2439=>"110111110",
    2440=>"111111111",
    2441=>"110000000",
    2442=>"000000000",
    2443=>"111111111",
    2444=>"000100111",
    2445=>"111010011",
    2446=>"111111111",
    2447=>"111111011",
    2448=>"001000000",
    2449=>"111011101",
    2450=>"111101100",
    2451=>"001000000",
    2452=>"111101100",
    2453=>"111111000",
    2454=>"000000111",
    2455=>"001000100",
    2456=>"100110111",
    2457=>"110010011",
    2458=>"110010000",
    2459=>"001000000",
    2460=>"111111011",
    2461=>"110111111",
    2462=>"000000000",
    2463=>"010011010",
    2464=>"001100100",
    2465=>"111111111",
    2466=>"000001100",
    2467=>"000000110",
    2468=>"000000000",
    2469=>"111111111",
    2470=>"000000000",
    2471=>"111111111",
    2472=>"010001001",
    2473=>"111111110",
    2474=>"011001101",
    2475=>"001000000",
    2476=>"111111111",
    2477=>"000000000",
    2478=>"100110111",
    2479=>"001000000",
    2480=>"111111010",
    2481=>"111011000",
    2482=>"000000100",
    2483=>"011010101",
    2484=>"111110100",
    2485=>"000000000",
    2486=>"111111111",
    2487=>"011001001",
    2488=>"001001000",
    2489=>"100110011",
    2490=>"000000000",
    2491=>"000000000",
    2492=>"111111111",
    2493=>"111111111",
    2494=>"000000000",
    2495=>"001100100",
    2496=>"010010100",
    2497=>"000001000",
    2498=>"000010011",
    2499=>"000011111",
    2500=>"001100111",
    2501=>"111001110",
    2502=>"000111111",
    2503=>"110110110",
    2504=>"001001011",
    2505=>"000000010",
    2506=>"000001111",
    2507=>"011010110",
    2508=>"110000111",
    2509=>"000000010",
    2510=>"110111001",
    2511=>"001001111",
    2512=>"011111111",
    2513=>"000111000",
    2514=>"100001001",
    2515=>"001010110",
    2516=>"111000000",
    2517=>"000000000",
    2518=>"111101000",
    2519=>"010110110",
    2520=>"111000000",
    2521=>"000111111",
    2522=>"111100110",
    2523=>"000110010",
    2524=>"110111111",
    2525=>"000111111",
    2526=>"000111011",
    2527=>"000111111",
    2528=>"111101000",
    2529=>"011001110",
    2530=>"100111110",
    2531=>"010101000",
    2532=>"000000000",
    2533=>"100001001",
    2534=>"111000111",
    2535=>"000000110",
    2536=>"000110110",
    2537=>"000000111",
    2538=>"010110100",
    2539=>"110111111",
    2540=>"000000000",
    2541=>"100001000",
    2542=>"111101000",
    2543=>"011110110",
    2544=>"000011111",
    2545=>"000111111",
    2546=>"111001001",
    2547=>"111111110",
    2548=>"000000111",
    2549=>"011011111",
    2550=>"100000111",
    2551=>"111000000",
    2552=>"100001000",
    2553=>"110000011",
    2554=>"010111110",
    2555=>"010110111",
    2556=>"111011000",
    2557=>"101000000",
    2558=>"000000000",
    2559=>"110111100",
    2560=>"100000010",
    2561=>"001111101",
    2562=>"111111111",
    2563=>"110000100",
    2564=>"000000111",
    2565=>"000000000",
    2566=>"111111111",
    2567=>"000000000",
    2568=>"010000000",
    2569=>"110010010",
    2570=>"111111111",
    2571=>"101011010",
    2572=>"111101111",
    2573=>"111110111",
    2574=>"010101001",
    2575=>"000000000",
    2576=>"100001000",
    2577=>"000001100",
    2578=>"111111111",
    2579=>"111111111",
    2580=>"111100101",
    2581=>"000000000",
    2582=>"001101101",
    2583=>"011100100",
    2584=>"011111110",
    2585=>"001111100",
    2586=>"101111101",
    2587=>"100110111",
    2588=>"000111110",
    2589=>"111000010",
    2590=>"000000000",
    2591=>"000001111",
    2592=>"111000011",
    2593=>"001000000",
    2594=>"000000100",
    2595=>"001000100",
    2596=>"000000000",
    2597=>"111010011",
    2598=>"001111111",
    2599=>"111110111",
    2600=>"110010010",
    2601=>"000000000",
    2602=>"001110010",
    2603=>"011101101",
    2604=>"110111111",
    2605=>"111001010",
    2606=>"111000011",
    2607=>"010001011",
    2608=>"000101111",
    2609=>"010110001",
    2610=>"001000011",
    2611=>"010110111",
    2612=>"000101101",
    2613=>"000000101",
    2614=>"010000000",
    2615=>"111100100",
    2616=>"000111101",
    2617=>"111010111",
    2618=>"000000000",
    2619=>"111000100",
    2620=>"000001000",
    2621=>"100000000",
    2622=>"000000000",
    2623=>"000010100",
    2624=>"001001011",
    2625=>"111111111",
    2626=>"000000000",
    2627=>"110110100",
    2628=>"000000000",
    2629=>"011000110",
    2630=>"110110000",
    2631=>"000111001",
    2632=>"010010000",
    2633=>"001001111",
    2634=>"000000000",
    2635=>"001000101",
    2636=>"111101100",
    2637=>"110100101",
    2638=>"001001101",
    2639=>"000100000",
    2640=>"000000000",
    2641=>"110110110",
    2642=>"001101101",
    2643=>"100011111",
    2644=>"110100111",
    2645=>"000000111",
    2646=>"011011111",
    2647=>"001000111",
    2648=>"111110000",
    2649=>"000001001",
    2650=>"000000000",
    2651=>"001001111",
    2652=>"000100111",
    2653=>"111111110",
    2654=>"010001001",
    2655=>"000000001",
    2656=>"000000000",
    2657=>"000000000",
    2658=>"000100101",
    2659=>"111110000",
    2660=>"001111111",
    2661=>"000010000",
    2662=>"100000001",
    2663=>"111111111",
    2664=>"000000000",
    2665=>"110100100",
    2666=>"110100111",
    2667=>"111111111",
    2668=>"101001111",
    2669=>"000001001",
    2670=>"000000001",
    2671=>"001001011",
    2672=>"111011111",
    2673=>"100001111",
    2674=>"100000100",
    2675=>"101101011",
    2676=>"101000001",
    2677=>"001001011",
    2678=>"000000000",
    2679=>"111110000",
    2680=>"101001111",
    2681=>"001101011",
    2682=>"000001010",
    2683=>"000001010",
    2684=>"000100000",
    2685=>"110111010",
    2686=>"111111011",
    2687=>"000001001",
    2688=>"100100100",
    2689=>"100100100",
    2690=>"110100110",
    2691=>"000001111",
    2692=>"101101101",
    2693=>"001001001",
    2694=>"001010100",
    2695=>"001001000",
    2696=>"010011001",
    2697=>"111011000",
    2698=>"111000101",
    2699=>"111111111",
    2700=>"111110111",
    2701=>"101001100",
    2702=>"000000000",
    2703=>"001010010",
    2704=>"001001001",
    2705=>"101011001",
    2706=>"111001001",
    2707=>"111011111",
    2708=>"100000011",
    2709=>"001001011",
    2710=>"000001111",
    2711=>"011111111",
    2712=>"100000011",
    2713=>"110100100",
    2714=>"011011101",
    2715=>"100000000",
    2716=>"001001011",
    2717=>"010011011",
    2718=>"000101011",
    2719=>"100001011",
    2720=>"001001011",
    2721=>"001101001",
    2722=>"001101111",
    2723=>"100101111",
    2724=>"000000101",
    2725=>"100000010",
    2726=>"110011111",
    2727=>"110110100",
    2728=>"010010110",
    2729=>"111110100",
    2730=>"001000000",
    2731=>"000000100",
    2732=>"111110101",
    2733=>"001001001",
    2734=>"001001111",
    2735=>"001001011",
    2736=>"110110100",
    2737=>"000000000",
    2738=>"000001011",
    2739=>"000001100",
    2740=>"010100111",
    2741=>"110100111",
    2742=>"111110110",
    2743=>"100100000",
    2744=>"100000000",
    2745=>"111111111",
    2746=>"101000000",
    2747=>"111110111",
    2748=>"000001011",
    2749=>"100000001",
    2750=>"011110110",
    2751=>"110100100",
    2752=>"001100110",
    2753=>"111011101",
    2754=>"000000111",
    2755=>"111011000",
    2756=>"001001011",
    2757=>"000101001",
    2758=>"000000111",
    2759=>"111100111",
    2760=>"001001111",
    2761=>"111000000",
    2762=>"100100111",
    2763=>"000001011",
    2764=>"111101101",
    2765=>"000011000",
    2766=>"000000111",
    2767=>"010000100",
    2768=>"000010010",
    2769=>"011111000",
    2770=>"001001111",
    2771=>"010010010",
    2772=>"000011011",
    2773=>"000000111",
    2774=>"011111100",
    2775=>"011110000",
    2776=>"101101101",
    2777=>"100000010",
    2778=>"011111100",
    2779=>"100000111",
    2780=>"101000011",
    2781=>"111111000",
    2782=>"000000101",
    2783=>"000010111",
    2784=>"001001011",
    2785=>"000001011",
    2786=>"111011001",
    2787=>"000000100",
    2788=>"101111000",
    2789=>"100100011",
    2790=>"011110100",
    2791=>"000011111",
    2792=>"000000111",
    2793=>"000000011",
    2794=>"001011011",
    2795=>"110111000",
    2796=>"100000011",
    2797=>"000110111",
    2798=>"011101101",
    2799=>"010110111",
    2800=>"111000001",
    2801=>"000000101",
    2802=>"010011111",
    2803=>"000110111",
    2804=>"000010111",
    2805=>"000100111",
    2806=>"000001011",
    2807=>"001101000",
    2808=>"011010100",
    2809=>"000110110",
    2810=>"000010111",
    2811=>"000110111",
    2812=>"011111001",
    2813=>"110000000",
    2814=>"000000011",
    2815=>"010010010",
    2816=>"111111111",
    2817=>"000000000",
    2818=>"111111011",
    2819=>"010110010",
    2820=>"111111110",
    2821=>"000000000",
    2822=>"000100010",
    2823=>"110001011",
    2824=>"100000001",
    2825=>"000000000",
    2826=>"111011110",
    2827=>"111111111",
    2828=>"111110110",
    2829=>"000000000",
    2830=>"111110111",
    2831=>"100100110",
    2832=>"000000001",
    2833=>"011001000",
    2834=>"111101110",
    2835=>"000000100",
    2836=>"011011001",
    2837=>"110110011",
    2838=>"111111111",
    2839=>"101000000",
    2840=>"000000000",
    2841=>"111111010",
    2842=>"000000000",
    2843=>"011000010",
    2844=>"000010000",
    2845=>"111111000",
    2846=>"000000000",
    2847=>"100000111",
    2848=>"000000000",
    2849=>"000100000",
    2850=>"000000000",
    2851=>"000100111",
    2852=>"000000000",
    2853=>"111111111",
    2854=>"001001000",
    2855=>"111111111",
    2856=>"111111111",
    2857=>"000000000",
    2858=>"010000000",
    2859=>"100000000",
    2860=>"111111011",
    2861=>"010110111",
    2862=>"000000000",
    2863=>"110001101",
    2864=>"011011011",
    2865=>"000000000",
    2866=>"001001010",
    2867=>"000001000",
    2868=>"010110110",
    2869=>"111111111",
    2870=>"111111111",
    2871=>"010000011",
    2872=>"000000101",
    2873=>"010111111",
    2874=>"110101100",
    2875=>"111111111",
    2876=>"111111111",
    2877=>"100001101",
    2878=>"111011111",
    2879=>"100100100",
    2880=>"110111111",
    2881=>"000000100",
    2882=>"000000000",
    2883=>"111001111",
    2884=>"000000100",
    2885=>"011011000",
    2886=>"000000000",
    2887=>"111111011",
    2888=>"000000000",
    2889=>"000101111",
    2890=>"000000000",
    2891=>"101100110",
    2892=>"111100110",
    2893=>"111010111",
    2894=>"001000111",
    2895=>"111010001",
    2896=>"101101011",
    2897=>"111011000",
    2898=>"110101110",
    2899=>"101000001",
    2900=>"111111111",
    2901=>"000100100",
    2902=>"111111100",
    2903=>"101101110",
    2904=>"010111110",
    2905=>"000001111",
    2906=>"111111100",
    2907=>"000011011",
    2908=>"000111001",
    2909=>"111001001",
    2910=>"000000000",
    2911=>"000110000",
    2912=>"111100000",
    2913=>"000000100",
    2914=>"101101110",
    2915=>"111110000",
    2916=>"011111100",
    2917=>"011000010",
    2918=>"100000001",
    2919=>"000000000",
    2920=>"000000000",
    2921=>"111001101",
    2922=>"000110000",
    2923=>"111101111",
    2924=>"100100110",
    2925=>"100111111",
    2926=>"111111111",
    2927=>"001111111",
    2928=>"000000000",
    2929=>"000111110",
    2930=>"110111110",
    2931=>"000010010",
    2932=>"000000001",
    2933=>"000001110",
    2934=>"110110010",
    2935=>"111001111",
    2936=>"101001100",
    2937=>"111101110",
    2938=>"100101000",
    2939=>"010010010",
    2940=>"111000000",
    2941=>"001101000",
    2942=>"000000100",
    2943=>"001101111",
    2944=>"010110110",
    2945=>"000011110",
    2946=>"110110000",
    2947=>"100100111",
    2948=>"001100111",
    2949=>"100110111",
    2950=>"101111011",
    2951=>"100000100",
    2952=>"111110110",
    2953=>"011010100",
    2954=>"111101001",
    2955=>"001001100",
    2956=>"111110110",
    2957=>"011100110",
    2958=>"001010000",
    2959=>"000000011",
    2960=>"000101011",
    2961=>"100100000",
    2962=>"100100111",
    2963=>"110111000",
    2964=>"101000000",
    2965=>"010010000",
    2966=>"010011010",
    2967=>"000011011",
    2968=>"100100100",
    2969=>"111010000",
    2970=>"100101101",
    2971=>"100110111",
    2972=>"101111111",
    2973=>"100100111",
    2974=>"110110110",
    2975=>"000010000",
    2976=>"100000001",
    2977=>"110111111",
    2978=>"100100011",
    2979=>"100000001",
    2980=>"000111110",
    2981=>"110000001",
    2982=>"001011011",
    2983=>"111011001",
    2984=>"100101100",
    2985=>"000000000",
    2986=>"001001000",
    2987=>"000100111",
    2988=>"101101000",
    2989=>"011100001",
    2990=>"100010011",
    2991=>"010000110",
    2992=>"110100111",
    2993=>"111000000",
    2994=>"101100000",
    2995=>"000011011",
    2996=>"110110100",
    2997=>"100100111",
    2998=>"101001111",
    2999=>"001000000",
    3000=>"010010000",
    3001=>"110100000",
    3002=>"000001000",
    3003=>"110011100",
    3004=>"000000011",
    3005=>"100000000",
    3006=>"011110110",
    3007=>"100100111",
    3008=>"000000001",
    3009=>"001011001",
    3010=>"110111111",
    3011=>"101111101",
    3012=>"100111101",
    3013=>"001111000",
    3014=>"011001011",
    3015=>"110110101",
    3016=>"110111001",
    3017=>"000000111",
    3018=>"100100100",
    3019=>"000111011",
    3020=>"100100101",
    3021=>"000000001",
    3022=>"100111100",
    3023=>"000100000",
    3024=>"000001001",
    3025=>"101101101",
    3026=>"001100010",
    3027=>"011000011",
    3028=>"000110010",
    3029=>"001001001",
    3030=>"101101111",
    3031=>"001001001",
    3032=>"000001110",
    3033=>"111101100",
    3034=>"001001000",
    3035=>"111001100",
    3036=>"001001001",
    3037=>"100110110",
    3038=>"011011011",
    3039=>"001001001",
    3040=>"110100000",
    3041=>"001000111",
    3042=>"001001110",
    3043=>"100100110",
    3044=>"000110101",
    3045=>"100110111",
    3046=>"011010000",
    3047=>"001010110",
    3048=>"011010001",
    3049=>"001001000",
    3050=>"001001100",
    3051=>"110001000",
    3052=>"111011001",
    3053=>"001001000",
    3054=>"110110110",
    3055=>"111011001",
    3056=>"111100000",
    3057=>"001001001",
    3058=>"000001000",
    3059=>"011011001",
    3060=>"011001001",
    3061=>"111100000",
    3062=>"000000000",
    3063=>"100110011",
    3064=>"011001001",
    3065=>"110111001",
    3066=>"011001001",
    3067=>"110001001",
    3068=>"110100110",
    3069=>"110000000",
    3070=>"011110000",
    3071=>"001001001",
    3072=>"000000000",
    3073=>"000000111",
    3074=>"000001010",
    3075=>"011001001",
    3076=>"011111110",
    3077=>"001000010",
    3078=>"011111111",
    3079=>"000100000",
    3080=>"011111111",
    3081=>"010000011",
    3082=>"110111011",
    3083=>"001001100",
    3084=>"111101001",
    3085=>"101010111",
    3086=>"001001100",
    3087=>"100000101",
    3088=>"000000000",
    3089=>"111111101",
    3090=>"001001000",
    3091=>"111111111",
    3092=>"001001110",
    3093=>"111111110",
    3094=>"111111111",
    3095=>"110010111",
    3096=>"000000000",
    3097=>"111100000",
    3098=>"000000000",
    3099=>"100100001",
    3100=>"001001101",
    3101=>"011011101",
    3102=>"001111110",
    3103=>"101101111",
    3104=>"000000110",
    3105=>"111111111",
    3106=>"011000110",
    3107=>"001000000",
    3108=>"111111111",
    3109=>"000000000",
    3110=>"110110011",
    3111=>"111011111",
    3112=>"000010100",
    3113=>"000000000",
    3114=>"001011111",
    3115=>"110100001",
    3116=>"000000000",
    3117=>"100100011",
    3118=>"001000110",
    3119=>"101100011",
    3120=>"111111101",
    3121=>"111110010",
    3122=>"000000000",
    3123=>"111111111",
    3124=>"000000100",
    3125=>"110111111",
    3126=>"100011111",
    3127=>"101111111",
    3128=>"111101111",
    3129=>"001100100",
    3130=>"100100100",
    3131=>"100100010",
    3132=>"101111111",
    3133=>"000100000",
    3134=>"111110111",
    3135=>"111000000",
    3136=>"100110110",
    3137=>"100010000",
    3138=>"000111001",
    3139=>"000111111",
    3140=>"010011001",
    3141=>"011000110",
    3142=>"011011100",
    3143=>"100111011",
    3144=>"011001000",
    3145=>"100011000",
    3146=>"100100000",
    3147=>"010011000",
    3148=>"110111111",
    3149=>"001000000",
    3150=>"010011100",
    3151=>"011111101",
    3152=>"111011000",
    3153=>"111001100",
    3154=>"100111111",
    3155=>"000000100",
    3156=>"001110010",
    3157=>"000111000",
    3158=>"111000000",
    3159=>"110011000",
    3160=>"110110011",
    3161=>"100100110",
    3162=>"110100101",
    3163=>"111000000",
    3164=>"111001001",
    3165=>"001000111",
    3166=>"110011110",
    3167=>"010001001",
    3168=>"000111011",
    3169=>"110000000",
    3170=>"110110000",
    3171=>"000000100",
    3172=>"000100111",
    3173=>"000111101",
    3174=>"101100100",
    3175=>"000000010",
    3176=>"100111111",
    3177=>"010000000",
    3178=>"111110000",
    3179=>"100110110",
    3180=>"001101110",
    3181=>"100110000",
    3182=>"001001001",
    3183=>"100000000",
    3184=>"111011000",
    3185=>"001100000",
    3186=>"011001000",
    3187=>"111011010",
    3188=>"111011000",
    3189=>"000111111",
    3190=>"111011001",
    3191=>"000110111",
    3192=>"111111000",
    3193=>"101011000",
    3194=>"000110110",
    3195=>"000110011",
    3196=>"110100111",
    3197=>"000000011",
    3198=>"000000000",
    3199=>"000100010",
    3200=>"110001110",
    3201=>"000101000",
    3202=>"111101010",
    3203=>"101001001",
    3204=>"100000100",
    3205=>"000000001",
    3206=>"000000100",
    3207=>"011010110",
    3208=>"001101000",
    3209=>"010110110",
    3210=>"000011000",
    3211=>"111101111",
    3212=>"010000111",
    3213=>"101111101",
    3214=>"100111010",
    3215=>"001001001",
    3216=>"001001000",
    3217=>"101101001",
    3218=>"100101111",
    3219=>"101101000",
    3220=>"111101000",
    3221=>"000100110",
    3222=>"001001001",
    3223=>"001000000",
    3224=>"111000111",
    3225=>"001000101",
    3226=>"000000101",
    3227=>"010111011",
    3228=>"010001010",
    3229=>"100000101",
    3230=>"001001101",
    3231=>"110111111",
    3232=>"110111110",
    3233=>"011001001",
    3234=>"101001101",
    3235=>"101001001",
    3236=>"011000001",
    3237=>"110010011",
    3238=>"101000000",
    3239=>"100101100",
    3240=>"111111111",
    3241=>"000000100",
    3242=>"000011110",
    3243=>"001101101",
    3244=>"111011011",
    3245=>"110111101",
    3246=>"111010110",
    3247=>"111011010",
    3248=>"000001111",
    3249=>"001011000",
    3250=>"101101110",
    3251=>"011010010",
    3252=>"000000000",
    3253=>"010100100",
    3254=>"100100100",
    3255=>"000000000",
    3256=>"000000001",
    3257=>"110110110",
    3258=>"001111111",
    3259=>"011011101",
    3260=>"001001001",
    3261=>"011101100",
    3262=>"011000001",
    3263=>"000000000",
    3264=>"111101001",
    3265=>"000000000",
    3266=>"000000000",
    3267=>"000100110",
    3268=>"110100110",
    3269=>"111100111",
    3270=>"100011010",
    3271=>"111111001",
    3272=>"000000000",
    3273=>"011111010",
    3274=>"111011011",
    3275=>"001100100",
    3276=>"000000000",
    3277=>"111111101",
    3278=>"111001000",
    3279=>"100011110",
    3280=>"111101111",
    3281=>"001111011",
    3282=>"111111111",
    3283=>"110001011",
    3284=>"111111111",
    3285=>"011101010",
    3286=>"110100101",
    3287=>"001000101",
    3288=>"000000000",
    3289=>"111111010",
    3290=>"110101011",
    3291=>"001011111",
    3292=>"111011011",
    3293=>"111111000",
    3294=>"000000000",
    3295=>"001110111",
    3296=>"010100001",
    3297=>"101100110",
    3298=>"100110100",
    3299=>"110001010",
    3300=>"111111111",
    3301=>"111111100",
    3302=>"010111111",
    3303=>"000000000",
    3304=>"000000000",
    3305=>"001010000",
    3306=>"001000000",
    3307=>"111111111",
    3308=>"100110001",
    3309=>"110000001",
    3310=>"000100001",
    3311=>"011111111",
    3312=>"010111011",
    3313=>"101000000",
    3314=>"011101101",
    3315=>"001000101",
    3316=>"100101111",
    3317=>"111111111",
    3318=>"111101110",
    3319=>"000000000",
    3320=>"100001010",
    3321=>"100101111",
    3322=>"111110111",
    3323=>"000000001",
    3324=>"000000000",
    3325=>"110000001",
    3326=>"000000000",
    3327=>"001000001",
    3328=>"001100000",
    3329=>"111101111",
    3330=>"111101111",
    3331=>"101101001",
    3332=>"001100010",
    3333=>"111101000",
    3334=>"111111111",
    3335=>"001000000",
    3336=>"110111111",
    3337=>"000000000",
    3338=>"000011011",
    3339=>"111001000",
    3340=>"111101111",
    3341=>"111000110",
    3342=>"100110111",
    3343=>"111110101",
    3344=>"111110010",
    3345=>"001000000",
    3346=>"111111011",
    3347=>"111000101",
    3348=>"100001000",
    3349=>"100000000",
    3350=>"111101111",
    3351=>"111011011",
    3352=>"111111111",
    3353=>"000000000",
    3354=>"001100001",
    3355=>"101010000",
    3356=>"000000101",
    3357=>"000000000",
    3358=>"101111111",
    3359=>"000000000",
    3360=>"111111111",
    3361=>"010011000",
    3362=>"001010000",
    3363=>"000000000",
    3364=>"000000000",
    3365=>"000000000",
    3366=>"011010000",
    3367=>"111101111",
    3368=>"111011111",
    3369=>"111111111",
    3370=>"001111110",
    3371=>"011000000",
    3372=>"111101101",
    3373=>"111110111",
    3374=>"111111111",
    3375=>"111110111",
    3376=>"000011000",
    3377=>"001000000",
    3378=>"101101101",
    3379=>"000000000",
    3380=>"101111100",
    3381=>"001001001",
    3382=>"000001000",
    3383=>"111111111",
    3384=>"110011111",
    3385=>"111001100",
    3386=>"001010000",
    3387=>"101101110",
    3388=>"111111111",
    3389=>"000000000",
    3390=>"111111111",
    3391=>"111000101",
    3392=>"000000010",
    3393=>"110000110",
    3394=>"000011001",
    3395=>"111111111",
    3396=>"010011001",
    3397=>"111011000",
    3398=>"011110011",
    3399=>"111111111",
    3400=>"111010001",
    3401=>"000100101",
    3402=>"000110100",
    3403=>"011011001",
    3404=>"000010110",
    3405=>"000000010",
    3406=>"010011001",
    3407=>"111111111",
    3408=>"110111111",
    3409=>"111111100",
    3410=>"110011001",
    3411=>"011111100",
    3412=>"011001001",
    3413=>"000000000",
    3414=>"000111000",
    3415=>"111111000",
    3416=>"101111111",
    3417=>"111000000",
    3418=>"111111110",
    3419=>"100110000",
    3420=>"011110010",
    3421=>"101001111",
    3422=>"111011000",
    3423=>"111110000",
    3424=>"010011111",
    3425=>"000011011",
    3426=>"011001010",
    3427=>"001001111",
    3428=>"110111111",
    3429=>"011111111",
    3430=>"011110110",
    3431=>"000010011",
    3432=>"000000111",
    3433=>"111000000",
    3434=>"011111001",
    3435=>"111111101",
    3436=>"000000000",
    3437=>"100100100",
    3438=>"000101001",
    3439=>"000000100",
    3440=>"111000000",
    3441=>"111100000",
    3442=>"111111111",
    3443=>"000000010",
    3444=>"000000111",
    3445=>"000100000",
    3446=>"000000000",
    3447=>"000011111",
    3448=>"110111000",
    3449=>"110101000",
    3450=>"011110111",
    3451=>"000100100",
    3452=>"111111000",
    3453=>"111010101",
    3454=>"000100110",
    3455=>"110110010",
    3456=>"000011111",
    3457=>"111111000",
    3458=>"000101111",
    3459=>"011111111",
    3460=>"000100110",
    3461=>"111001100",
    3462=>"011111100",
    3463=>"000000111",
    3464=>"011011000",
    3465=>"101001101",
    3466=>"000111101",
    3467=>"000001110",
    3468=>"111111111",
    3469=>"100111001",
    3470=>"010000101",
    3471=>"000000111",
    3472=>"101111111",
    3473=>"111000000",
    3474=>"111011011",
    3475=>"000000111",
    3476=>"000000001",
    3477=>"110000000",
    3478=>"111111000",
    3479=>"111111000",
    3480=>"010111010",
    3481=>"010000000",
    3482=>"111100011",
    3483=>"101111000",
    3484=>"000010111",
    3485=>"111000000",
    3486=>"111111000",
    3487=>"000111011",
    3488=>"000000111",
    3489=>"111000000",
    3490=>"011000011",
    3491=>"100000111",
    3492=>"111000111",
    3493=>"000000111",
    3494=>"111100000",
    3495=>"000100111",
    3496=>"000111010",
    3497=>"000000101",
    3498=>"001000110",
    3499=>"010000110",
    3500=>"000111110",
    3501=>"000000010",
    3502=>"000000111",
    3503=>"110111000",
    3504=>"000111110",
    3505=>"000001000",
    3506=>"011101111",
    3507=>"101001100",
    3508=>"011111000",
    3509=>"000010011",
    3510=>"000000011",
    3511=>"010000101",
    3512=>"111101000",
    3513=>"000001111",
    3514=>"000000100",
    3515=>"000000111",
    3516=>"010000000",
    3517=>"111100100",
    3518=>"000010100",
    3519=>"110010000",
    3520=>"000000010",
    3521=>"100100000",
    3522=>"000001010",
    3523=>"110011001",
    3524=>"000011011",
    3525=>"000011111",
    3526=>"011110000",
    3527=>"111101000",
    3528=>"000011111",
    3529=>"001000111",
    3530=>"111110000",
    3531=>"000000111",
    3532=>"110011111",
    3533=>"100000000",
    3534=>"001000111",
    3535=>"010000000",
    3536=>"001100001",
    3537=>"110110000",
    3538=>"111111110",
    3539=>"011111100",
    3540=>"001011010",
    3541=>"000010100",
    3542=>"111100110",
    3543=>"011110000",
    3544=>"000001111",
    3545=>"011110001",
    3546=>"111100000",
    3547=>"111110000",
    3548=>"010100001",
    3549=>"000001111",
    3550=>"000011111",
    3551=>"001110100",
    3552=>"111011110",
    3553=>"001011000",
    3554=>"111000001",
    3555=>"100000001",
    3556=>"011100000",
    3557=>"000001111",
    3558=>"110100000",
    3559=>"111011110",
    3560=>"000100000",
    3561=>"001110000",
    3562=>"000011110",
    3563=>"001010100",
    3564=>"000110100",
    3565=>"011110000",
    3566=>"100001111",
    3567=>"001100000",
    3568=>"110110000",
    3569=>"010100001",
    3570=>"000001111",
    3571=>"111110000",
    3572=>"111100000",
    3573=>"011100000",
    3574=>"011100100",
    3575=>"100001111",
    3576=>"011110000",
    3577=>"001000000",
    3578=>"011010100",
    3579=>"011110100",
    3580=>"111111000",
    3581=>"000001011",
    3582=>"011000000",
    3583=>"111100000",
    3584=>"100100011",
    3585=>"010110001",
    3586=>"010010111",
    3587=>"111011000",
    3588=>"111101111",
    3589=>"100000111",
    3590=>"010010000",
    3591=>"100110110",
    3592=>"000000000",
    3593=>"110100001",
    3594=>"110010111",
    3595=>"111111111",
    3596=>"111000111",
    3597=>"010110111",
    3598=>"000000000",
    3599=>"010111011",
    3600=>"000100110",
    3601=>"010000100",
    3602=>"011100111",
    3603=>"110000001",
    3604=>"010000100",
    3605=>"111100000",
    3606=>"100110111",
    3607=>"000000000",
    3608=>"000000100",
    3609=>"001000001",
    3610=>"101000111",
    3611=>"100000100",
    3612=>"111011000",
    3613=>"000000000",
    3614=>"000010000",
    3615=>"000110111",
    3616=>"110100110",
    3617=>"011001100",
    3618=>"011111111",
    3619=>"000000100",
    3620=>"001000110",
    3621=>"010010010",
    3622=>"010000000",
    3623=>"001110000",
    3624=>"100011111",
    3625=>"111110000",
    3626=>"111001100",
    3627=>"010100011",
    3628=>"110001010",
    3629=>"111011100",
    3630=>"100110111",
    3631=>"011011010",
    3632=>"111111001",
    3633=>"110100110",
    3634=>"111001001",
    3635=>"111110010",
    3636=>"000100111",
    3637=>"000001110",
    3638=>"011010100",
    3639=>"000000110",
    3640=>"111111111",
    3641=>"110000000",
    3642=>"010000000",
    3643=>"000010011",
    3644=>"101000011",
    3645=>"110010000",
    3646=>"010011000",
    3647=>"000110111",
    3648=>"000001001",
    3649=>"001000010",
    3650=>"011111111",
    3651=>"000001110",
    3652=>"000110010",
    3653=>"111000000",
    3654=>"101000110",
    3655=>"000111111",
    3656=>"000111111",
    3657=>"000000101",
    3658=>"000111110",
    3659=>"001111110",
    3660=>"000111111",
    3661=>"011001111",
    3662=>"000000111",
    3663=>"000111111",
    3664=>"111000000",
    3665=>"111100000",
    3666=>"001001000",
    3667=>"111100100",
    3668=>"111100011",
    3669=>"111010000",
    3670=>"111000000",
    3671=>"111000000",
    3672=>"110000000",
    3673=>"111000010",
    3674=>"110000000",
    3675=>"110000000",
    3676=>"111000101",
    3677=>"000111111",
    3678=>"001000010",
    3679=>"001000000",
    3680=>"000111111",
    3681=>"111010000",
    3682=>"111000000",
    3683=>"000111111",
    3684=>"101000000",
    3685=>"000111111",
    3686=>"111110000",
    3687=>"000000001",
    3688=>"111111111",
    3689=>"000000111",
    3690=>"111000000",
    3691=>"111110001",
    3692=>"000000100",
    3693=>"110000100",
    3694=>"000111111",
    3695=>"011010010",
    3696=>"111000011",
    3697=>"111000000",
    3698=>"101001010",
    3699=>"110110110",
    3700=>"111010000",
    3701=>"000000100",
    3702=>"100111111",
    3703=>"000110111",
    3704=>"111000000",
    3705=>"000101111",
    3706=>"100101110",
    3707=>"000001111",
    3708=>"010110010",
    3709=>"000111101",
    3710=>"000011111",
    3711=>"111000000",
    3712=>"111111111",
    3713=>"110111101",
    3714=>"000000010",
    3715=>"101001010",
    3716=>"111011011",
    3717=>"111011100",
    3718=>"000000000",
    3719=>"011000111",
    3720=>"111011000",
    3721=>"111010010",
    3722=>"001010110",
    3723=>"000111000",
    3724=>"111100111",
    3725=>"110111111",
    3726=>"011001011",
    3727=>"001000000",
    3728=>"001100111",
    3729=>"100111001",
    3730=>"000000000",
    3731=>"000000000",
    3732=>"011000101",
    3733=>"000000000",
    3734=>"100101101",
    3735=>"001000000",
    3736=>"010111011",
    3737=>"110111000",
    3738=>"100000000",
    3739=>"001101100",
    3740=>"001011000",
    3741=>"100000000",
    3742=>"111111111",
    3743=>"110000101",
    3744=>"000000111",
    3745=>"110111111",
    3746=>"111111111",
    3747=>"001000111",
    3748=>"111000111",
    3749=>"000000000",
    3750=>"000000010",
    3751=>"000000000",
    3752=>"011010111",
    3753=>"101000100",
    3754=>"101101101",
    3755=>"010101001",
    3756=>"000000010",
    3757=>"111010110",
    3758=>"011000111",
    3759=>"001000000",
    3760=>"000111101",
    3761=>"000011100",
    3762=>"000110001",
    3763=>"011011110",
    3764=>"001001111",
    3765=>"011111111",
    3766=>"011010110",
    3767=>"111001111",
    3768=>"101111010",
    3769=>"001010110",
    3770=>"111101111",
    3771=>"111000111",
    3772=>"000000000",
    3773=>"100100000",
    3774=>"111111111",
    3775=>"000111011",
    3776=>"101001011",
    3777=>"111111111",
    3778=>"000000000",
    3779=>"100111000",
    3780=>"000110110",
    3781=>"110111001",
    3782=>"101110110",
    3783=>"000001001",
    3784=>"001000100",
    3785=>"000000001",
    3786=>"010000001",
    3787=>"110000011",
    3788=>"111101000",
    3789=>"010001000",
    3790=>"010000000",
    3791=>"000000110",
    3792=>"000001011",
    3793=>"000111111",
    3794=>"111000100",
    3795=>"000010110",
    3796=>"101100111",
    3797=>"110110111",
    3798=>"111111111",
    3799=>"111111011",
    3800=>"000010101",
    3801=>"010110000",
    3802=>"001010100",
    3803=>"011001111",
    3804=>"111111000",
    3805=>"000000001",
    3806=>"111011011",
    3807=>"111101000",
    3808=>"000000001",
    3809=>"011111011",
    3810=>"000000101",
    3811=>"000100000",
    3812=>"100101111",
    3813=>"001000100",
    3814=>"111010110",
    3815=>"010000100",
    3816=>"000000000",
    3817=>"010000000",
    3818=>"010100000",
    3819=>"111111100",
    3820=>"111100111",
    3821=>"111001010",
    3822=>"000000000",
    3823=>"100111110",
    3824=>"000111010",
    3825=>"000101111",
    3826=>"000000110",
    3827=>"111111010",
    3828=>"111111111",
    3829=>"111001111",
    3830=>"011111011",
    3831=>"000000000",
    3832=>"110111111",
    3833=>"000001011",
    3834=>"010000001",
    3835=>"000000101",
    3836=>"110111111",
    3837=>"000000011",
    3838=>"000000000",
    3839=>"000011111",
    3840=>"110110110",
    3841=>"100110110",
    3842=>"011011011",
    3843=>"101001001",
    3844=>"011011011",
    3845=>"101101101",
    3846=>"101000011",
    3847=>"001001001",
    3848=>"111011111",
    3849=>"010011001",
    3850=>"011011011",
    3851=>"010010011",
    3852=>"111111111",
    3853=>"011011011",
    3854=>"110010011",
    3855=>"000001001",
    3856=>"000000011",
    3857=>"101101100",
    3858=>"100110010",
    3859=>"100110011",
    3860=>"000010010",
    3861=>"000010110",
    3862=>"111110110",
    3863=>"100100100",
    3864=>"000100100",
    3865=>"000000011",
    3866=>"101100100",
    3867=>"101100110",
    3868=>"000010011",
    3869=>"000011101",
    3870=>"111101110",
    3871=>"110010010",
    3872=>"010010000",
    3873=>"011010001",
    3874=>"111100100",
    3875=>"001000000",
    3876=>"101101100",
    3877=>"010011001",
    3878=>"100100110",
    3879=>"100110010",
    3880=>"010000001",
    3881=>"100000000",
    3882=>"110100110",
    3883=>"100100100",
    3884=>"110111010",
    3885=>"010110010",
    3886=>"011011011",
    3887=>"011111011",
    3888=>"101110110",
    3889=>"000110111",
    3890=>"000000000",
    3891=>"000001011",
    3892=>"001001001",
    3893=>"111011011",
    3894=>"011011011",
    3895=>"100100100",
    3896=>"101100100",
    3897=>"110011111",
    3898=>"001100000",
    3899=>"010010010",
    3900=>"001100100",
    3901=>"000101101",
    3902=>"011011011",
    3903=>"100100010",
    3904=>"100000011",
    3905=>"000000011",
    3906=>"111110000",
    3907=>"000000111",
    3908=>"000001111",
    3909=>"100000110",
    3910=>"101111011",
    3911=>"011000001",
    3912=>"000000010",
    3913=>"111110000",
    3914=>"100000111",
    3915=>"111011000",
    3916=>"111000111",
    3917=>"000101011",
    3918=>"111001100",
    3919=>"001000000",
    3920=>"111101101",
    3921=>"001100111",
    3922=>"000110111",
    3923=>"001100110",
    3924=>"000001000",
    3925=>"000000000",
    3926=>"000101111",
    3927=>"101000010",
    3928=>"110000000",
    3929=>"001110110",
    3930=>"001010011",
    3931=>"101010000",
    3932=>"000000010",
    3933=>"100001000",
    3934=>"001011010",
    3935=>"100111010",
    3936=>"111000000",
    3937=>"011011010",
    3938=>"001010000",
    3939=>"100000000",
    3940=>"001001111",
    3941=>"110011100",
    3942=>"000011010",
    3943=>"000111011",
    3944=>"010011000",
    3945=>"111010000",
    3946=>"001010110",
    3947=>"000000110",
    3948=>"011001100",
    3949=>"101110111",
    3950=>"111111000",
    3951=>"110101100",
    3952=>"001000111",
    3953=>"001000000",
    3954=>"100101001",
    3955=>"001110111",
    3956=>"010000111",
    3957=>"000100001",
    3958=>"110111001",
    3959=>"000000100",
    3960=>"001110010",
    3961=>"010000101",
    3962=>"001001100",
    3963=>"010010111",
    3964=>"000001111",
    3965=>"101000000",
    3966=>"011011001",
    3967=>"110000000",
    3968=>"100101000",
    3969=>"000000010",
    3970=>"000010000",
    3971=>"111100111",
    3972=>"001110100",
    3973=>"001000000",
    3974=>"111000111",
    3975=>"100100000",
    3976=>"011011000",
    3977=>"100000010",
    3978=>"100100001",
    3979=>"001111001",
    3980=>"101101111",
    3981=>"011111010",
    3982=>"011111100",
    3983=>"000010111",
    3984=>"101000000",
    3985=>"111010000",
    3986=>"010101100",
    3987=>"111011101",
    3988=>"111001101",
    3989=>"000100111",
    3990=>"110110111",
    3991=>"110000011",
    3992=>"001001001",
    3993=>"011101000",
    3994=>"110000000",
    3995=>"100001000",
    3996=>"111111000",
    3997=>"011111000",
    3998=>"011100111",
    3999=>"010000100",
    4000=>"111000001",
    4001=>"011010010",
    4002=>"101110111",
    4003=>"010000001",
    4004=>"111001111",
    4005=>"000001000",
    4006=>"110010010",
    4007=>"111101101",
    4008=>"000101000",
    4009=>"000000000",
    4010=>"010001101",
    4011=>"000000100",
    4012=>"000101100",
    4013=>"111100100",
    4014=>"100111101",
    4015=>"101100000",
    4016=>"111110000",
    4017=>"111000000",
    4018=>"011000000",
    4019=>"001000000",
    4020=>"000011010",
    4021=>"000011111",
    4022=>"000000110",
    4023=>"110100100",
    4024=>"110010011",
    4025=>"001100100",
    4026=>"110110000",
    4027=>"110111001",
    4028=>"111000100",
    4029=>"100000000",
    4030=>"110001001",
    4031=>"111000101",
    4032=>"010110111",
    4033=>"100101101",
    4034=>"010000010",
    4035=>"001000101",
    4036=>"010000000",
    4037=>"100001001",
    4038=>"011010110",
    4039=>"001010010",
    4040=>"110011011",
    4041=>"010010010",
    4042=>"011010111",
    4043=>"000010100",
    4044=>"111111111",
    4045=>"110101001",
    4046=>"001010000",
    4047=>"000010010",
    4048=>"001001100",
    4049=>"100101001",
    4050=>"110100111",
    4051=>"011000000",
    4052=>"111010011",
    4053=>"000010010",
    4054=>"100101111",
    4055=>"011010110",
    4056=>"100101001",
    4057=>"101010100",
    4058=>"001001000",
    4059=>"011110110",
    4060=>"000011111",
    4061=>"100101001",
    4062=>"111111111",
    4063=>"011010110",
    4064=>"011010000",
    4065=>"010110110",
    4066=>"110101001",
    4067=>"000000000",
    4068=>"110111100",
    4069=>"100000001",
    4070=>"010110110",
    4071=>"110000000",
    4072=>"001010110",
    4073=>"000000000",
    4074=>"010011001",
    4075=>"000001000",
    4076=>"101011111",
    4077=>"011010100",
    4078=>"110111010",
    4079=>"110110110",
    4080=>"100100100",
    4081=>"000001001",
    4082=>"110100001",
    4083=>"011110111",
    4084=>"010111100",
    4085=>"010111100",
    4086=>"011010110",
    4087=>"100000000",
    4088=>"110001011",
    4089=>"011100110",
    4090=>"011010010",
    4091=>"011010100",
    4092=>"100001001",
    4093=>"100001001",
    4094=>"011010110",
    4095=>"010100110");

BEGIN
    weight <= ROM_content(to_integer(address));
END RTL;