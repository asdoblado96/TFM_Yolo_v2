LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_6_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_6_WROM;

ARCHITECTURE RTL OF L8_6_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"000110001",
  1=>"101011100",
  2=>"001110101",
  3=>"100100000",
  4=>"000001111",
  5=>"000010001",
  6=>"010010001",
  7=>"100001011",
  8=>"101111001",
  9=>"100001100",
  10=>"011010011",
  11=>"100101001",
  12=>"000001011",
  13=>"010110111",
  14=>"101010111",
  15=>"100111011",
  16=>"111100011",
  17=>"000010000",
  18=>"100111110",
  19=>"111111001",
  20=>"010001001",
  21=>"011101001",
  22=>"110110101",
  23=>"000100000",
  24=>"011100011",
  25=>"001011111",
  26=>"101100000",
  27=>"011010101",
  28=>"011001101",
  29=>"110010001",
  30=>"001101011",
  31=>"110110010",
  32=>"110000011",
  33=>"011001010",
  34=>"101000011",
  35=>"011110001",
  36=>"101111011",
  37=>"011010110",
  38=>"100110001",
  39=>"111110110",
  40=>"111111000",
  41=>"110101100",
  42=>"011100101",
  43=>"011010000",
  44=>"110000011",
  45=>"110011110",
  46=>"010010101",
  47=>"000111000",
  48=>"001011011",
  49=>"101110010",
  50=>"111011000",
  51=>"010001000",
  52=>"001100010",
  53=>"101011000",
  54=>"110011001",
  55=>"001000000",
  56=>"010011011",
  57=>"101010101",
  58=>"110011000",
  59=>"000000110",
  60=>"011111001",
  61=>"001010010",
  62=>"110100011",
  63=>"000101101",
  64=>"001000011",
  65=>"111101101",
  66=>"001111010",
  67=>"010100001",
  68=>"000000011",
  69=>"011010110",
  70=>"111110011",
  71=>"110000110",
  72=>"001101001",
  73=>"001011011",
  74=>"110110001",
  75=>"001001011",
  76=>"000110010",
  77=>"111001100",
  78=>"101011110",
  79=>"100001110",
  80=>"101101110",
  81=>"000001010",
  82=>"101011000",
  83=>"111010010",
  84=>"111110000",
  85=>"101101101",
  86=>"100100101",
  87=>"101000100",
  88=>"100000101",
  89=>"111010001",
  90=>"000011010",
  91=>"011110111",
  92=>"001111100",
  93=>"100011111",
  94=>"000001010",
  95=>"100000000",
  96=>"110100110",
  97=>"001000110",
  98=>"101010001",
  99=>"000001110",
  100=>"001011000",
  101=>"001110110",
  102=>"111101111",
  103=>"101100010",
  104=>"010000000",
  105=>"011111000",
  106=>"100110000",
  107=>"010010111",
  108=>"101001000",
  109=>"101000001",
  110=>"011011000",
  111=>"110110111",
  112=>"011101111",
  113=>"011001000",
  114=>"110110101",
  115=>"010100011",
  116=>"101110111",
  117=>"110110101",
  118=>"110010100",
  119=>"111100101",
  120=>"101111110",
  121=>"001110011",
  122=>"011010001",
  123=>"110110011",
  124=>"010010110",
  125=>"110000000",
  126=>"100110110",
  127=>"011010100",
  128=>"001001110",
  129=>"001110110",
  130=>"100010100",
  131=>"011101110",
  132=>"010000010",
  133=>"011010111",
  134=>"001111001",
  135=>"000010000",
  136=>"010010001",
  137=>"001010010",
  138=>"100101110",
  139=>"001000011",
  140=>"110111000",
  141=>"101100010",
  142=>"111011101",
  143=>"110100010",
  144=>"110000000",
  145=>"001100100",
  146=>"000001100",
  147=>"100100101",
  148=>"001100010",
  149=>"011111011",
  150=>"000010001",
  151=>"101101110",
  152=>"101111000",
  153=>"000001011",
  154=>"100011111",
  155=>"101011010",
  156=>"101001000",
  157=>"101001101",
  158=>"100110000",
  159=>"001111010",
  160=>"001101001",
  161=>"110110110",
  162=>"010100010",
  163=>"101100000",
  164=>"000000010",
  165=>"111100111",
  166=>"000011000",
  167=>"010011111",
  168=>"001000010",
  169=>"110011010",
  170=>"111000010",
  171=>"011001110",
  172=>"110011101",
  173=>"000100101",
  174=>"100001111",
  175=>"110000000",
  176=>"010100011",
  177=>"110000001",
  178=>"010001101",
  179=>"000011100",
  180=>"011100101",
  181=>"010100100",
  182=>"110001011",
  183=>"000010010",
  184=>"111011001",
  185=>"111001110",
  186=>"101010010",
  187=>"101110101",
  188=>"111001000",
  189=>"011000001",
  190=>"111101101",
  191=>"100111001",
  192=>"000010000",
  193=>"001111110",
  194=>"100111100",
  195=>"011000111",
  196=>"111010010",
  197=>"111001111",
  198=>"010110000",
  199=>"101010000",
  200=>"001000000",
  201=>"010101011",
  202=>"000000001",
  203=>"111000110",
  204=>"100000010",
  205=>"010101111",
  206=>"110100100",
  207=>"100000000",
  208=>"100000000",
  209=>"101100111",
  210=>"100001111",
  211=>"101010011",
  212=>"010011001",
  213=>"001000001",
  214=>"010110110",
  215=>"111101011",
  216=>"010100100",
  217=>"111111100",
  218=>"001011011",
  219=>"101100100",
  220=>"010010001",
  221=>"000111111",
  222=>"001001111",
  223=>"010101001",
  224=>"001010101",
  225=>"010110001",
  226=>"100101110",
  227=>"110001000",
  228=>"101010100",
  229=>"010010111",
  230=>"000100010",
  231=>"111111011",
  232=>"001010100",
  233=>"000111010",
  234=>"011011100",
  235=>"101000110",
  236=>"000011111",
  237=>"110001101",
  238=>"101101100",
  239=>"000100110",
  240=>"111010111",
  241=>"111001001",
  242=>"100000011",
  243=>"111100011",
  244=>"011000110",
  245=>"010011010",
  246=>"100011010",
  247=>"000001000",
  248=>"010001001",
  249=>"111101111",
  250=>"111001011",
  251=>"001111100",
  252=>"101000111",
  253=>"110001010",
  254=>"011101011",
  255=>"001110000",
  256=>"010010001",
  257=>"000000110",
  258=>"111111001",
  259=>"101111110",
  260=>"101110100",
  261=>"000101000",
  262=>"111101111",
  263=>"010111001",
  264=>"100110000",
  265=>"101001111",
  266=>"011101010",
  267=>"111001001",
  268=>"001101111",
  269=>"001001001",
  270=>"101010110",
  271=>"100010111",
  272=>"110100000",
  273=>"100010111",
  274=>"111111111",
  275=>"011111001",
  276=>"010100000",
  277=>"000100101",
  278=>"100000001",
  279=>"011111001",
  280=>"000100011",
  281=>"011101100",
  282=>"111110011",
  283=>"111001101",
  284=>"001100111",
  285=>"011110001",
  286=>"110011010",
  287=>"000000101",
  288=>"000110110",
  289=>"000110001",
  290=>"010011010",
  291=>"110011111",
  292=>"011111011",
  293=>"010111010",
  294=>"000001001",
  295=>"001100111",
  296=>"011100001",
  297=>"101000010",
  298=>"001101100",
  299=>"110100000",
  300=>"000011000",
  301=>"001110011",
  302=>"111010010",
  303=>"001111101",
  304=>"101111110",
  305=>"111011011",
  306=>"110100110",
  307=>"100001110",
  308=>"111010100",
  309=>"111001001",
  310=>"100101101",
  311=>"001111010",
  312=>"001010010",
  313=>"001101010",
  314=>"010100110",
  315=>"001100010",
  316=>"100100000",
  317=>"010010100",
  318=>"100011101",
  319=>"111000001",
  320=>"011110101",
  321=>"000000001",
  322=>"010111010",
  323=>"110001011",
  324=>"110110000",
  325=>"010010011",
  326=>"010110101",
  327=>"100100110",
  328=>"011001110",
  329=>"000000101",
  330=>"010011100",
  331=>"001101010",
  332=>"110010011",
  333=>"111011111",
  334=>"011011000",
  335=>"011001010",
  336=>"110101110",
  337=>"101010110",
  338=>"100101110",
  339=>"001111110",
  340=>"100111010",
  341=>"111100000",
  342=>"000000011",
  343=>"000010010",
  344=>"101110111",
  345=>"100000010",
  346=>"000100000",
  347=>"100100110",
  348=>"001000101",
  349=>"101001001",
  350=>"010101110",
  351=>"011000100",
  352=>"010010101",
  353=>"101000110",
  354=>"110110110",
  355=>"000101100",
  356=>"010111100",
  357=>"010111100",
  358=>"010000010",
  359=>"110000101",
  360=>"011011000",
  361=>"000110100",
  362=>"100001000",
  363=>"010001111",
  364=>"100111000",
  365=>"000101101",
  366=>"000000011",
  367=>"011001001",
  368=>"101000010",
  369=>"110111001",
  370=>"111100001",
  371=>"010111110",
  372=>"101110001",
  373=>"000011110",
  374=>"110010111",
  375=>"001001001",
  376=>"101001111",
  377=>"010110001",
  378=>"010001111",
  379=>"111010110",
  380=>"100110011",
  381=>"010101010",
  382=>"011101100",
  383=>"101100100",
  384=>"001001000",
  385=>"011010011",
  386=>"110011000",
  387=>"101101100",
  388=>"011011011",
  389=>"100001100",
  390=>"111101011",
  391=>"010101100",
  392=>"010000110",
  393=>"011110000",
  394=>"110101101",
  395=>"011001101",
  396=>"110000001",
  397=>"010100000",
  398=>"111101110",
  399=>"100100010",
  400=>"011000111",
  401=>"100000000",
  402=>"110001000",
  403=>"001111111",
  404=>"100101011",
  405=>"111110110",
  406=>"100110011",
  407=>"101001111",
  408=>"100000101",
  409=>"110000100",
  410=>"101101011",
  411=>"001111000",
  412=>"000010101",
  413=>"011000100",
  414=>"110111011",
  415=>"110100000",
  416=>"110011010",
  417=>"111011001",
  418=>"010100000",
  419=>"000010011",
  420=>"011001111",
  421=>"000001110",
  422=>"000111010",
  423=>"101001010",
  424=>"101111110",
  425=>"100111110",
  426=>"000111000",
  427=>"101111111",
  428=>"000011001",
  429=>"100101000",
  430=>"100101001",
  431=>"010100111",
  432=>"010010101",
  433=>"000101111",
  434=>"100011101",
  435=>"001010110",
  436=>"000001011",
  437=>"111110111",
  438=>"001110011",
  439=>"001000110",
  440=>"110000011",
  441=>"000111000",
  442=>"100011000",
  443=>"001111100",
  444=>"101100010",
  445=>"100011000",
  446=>"001111111",
  447=>"011011000",
  448=>"001100100",
  449=>"100111101",
  450=>"011011100",
  451=>"101111101",
  452=>"101011010",
  453=>"100111111",
  454=>"010111000",
  455=>"001001001",
  456=>"000001101",
  457=>"110100101",
  458=>"110110010",
  459=>"010000111",
  460=>"001101000",
  461=>"111000000",
  462=>"111111100",
  463=>"011001001",
  464=>"011101010",
  465=>"010100010",
  466=>"010000001",
  467=>"110111111",
  468=>"010100110",
  469=>"100101001",
  470=>"000001000",
  471=>"110101000",
  472=>"011110110",
  473=>"110101101",
  474=>"111011001",
  475=>"001011000",
  476=>"001011111",
  477=>"010001011",
  478=>"101100100",
  479=>"001111001",
  480=>"110101000",
  481=>"001111011",
  482=>"100100010",
  483=>"100000110",
  484=>"000110000",
  485=>"101101110",
  486=>"011000010",
  487=>"010101111",
  488=>"001010010",
  489=>"100001000",
  490=>"010100110",
  491=>"000010110",
  492=>"001111101",
  493=>"000101000",
  494=>"010000000",
  495=>"100110000",
  496=>"001011010",
  497=>"011011101",
  498=>"111001100",
  499=>"001101111",
  500=>"011110000",
  501=>"110010101",
  502=>"101011000",
  503=>"011010110",
  504=>"010100011",
  505=>"010110011",
  506=>"100100111",
  507=>"101110101",
  508=>"100101100",
  509=>"011000000",
  510=>"001000001",
  511=>"011011000",
  512=>"000010011",
  513=>"011100111",
  514=>"111001001",
  515=>"000010101",
  516=>"001110001",
  517=>"110100011",
  518=>"011101100",
  519=>"001001101",
  520=>"101101001",
  521=>"100011011",
  522=>"010010111",
  523=>"111111111",
  524=>"001000100",
  525=>"110011001",
  526=>"110111110",
  527=>"100000001",
  528=>"111000001",
  529=>"011011001",
  530=>"000100001",
  531=>"110001011",
  532=>"000001001",
  533=>"011100001",
  534=>"110111110",
  535=>"111101110",
  536=>"111000000",
  537=>"101000011",
  538=>"000000111",
  539=>"110111001",
  540=>"101100111",
  541=>"110011111",
  542=>"011101100",
  543=>"111111110",
  544=>"100010000",
  545=>"101101100",
  546=>"011100011",
  547=>"001011100",
  548=>"101100101",
  549=>"010100110",
  550=>"110100001",
  551=>"111000000",
  552=>"001110011",
  553=>"100100100",
  554=>"000100110",
  555=>"011101010",
  556=>"100011010",
  557=>"110111010",
  558=>"001100101",
  559=>"101011111",
  560=>"001110111",
  561=>"001010001",
  562=>"111000001",
  563=>"001001001",
  564=>"111101000",
  565=>"010100110",
  566=>"100101100",
  567=>"110010110",
  568=>"011000101",
  569=>"110110001",
  570=>"110110011",
  571=>"100010110",
  572=>"010010101",
  573=>"000110111",
  574=>"000110010",
  575=>"010001100",
  576=>"110010010",
  577=>"111011011",
  578=>"111001011",
  579=>"000001001",
  580=>"110111111",
  581=>"110010011",
  582=>"000001110",
  583=>"000110011",
  584=>"011010010",
  585=>"111100010",
  586=>"010000100",
  587=>"001011111",
  588=>"100000000",
  589=>"001101101",
  590=>"011000000",
  591=>"100001110",
  592=>"110011011",
  593=>"110010010",
  594=>"110011000",
  595=>"000011101",
  596=>"000101000",
  597=>"000100001",
  598=>"111001101",
  599=>"000000000",
  600=>"000100000",
  601=>"111000010",
  602=>"001011011",
  603=>"100110110",
  604=>"011000111",
  605=>"001000000",
  606=>"100111100",
  607=>"001101110",
  608=>"000100110",
  609=>"011101101",
  610=>"001110100",
  611=>"111110111",
  612=>"110000011",
  613=>"110010011",
  614=>"000110110",
  615=>"100001111",
  616=>"100010000",
  617=>"000000100",
  618=>"101111100",
  619=>"110110000",
  620=>"100101010",
  621=>"001100000",
  622=>"000010101",
  623=>"110101010",
  624=>"001110000",
  625=>"011110001",
  626=>"110110110",
  627=>"010000011",
  628=>"100010000",
  629=>"010000110",
  630=>"011001111",
  631=>"101111000",
  632=>"011101010",
  633=>"000101010",
  634=>"101100100",
  635=>"111010010",
  636=>"101011010",
  637=>"110010111",
  638=>"100101001",
  639=>"110111111",
  640=>"100101101",
  641=>"111011110",
  642=>"001011010",
  643=>"110010010",
  644=>"010100111",
  645=>"001111111",
  646=>"110011011",
  647=>"000000011",
  648=>"110111001",
  649=>"100001100",
  650=>"000110111",
  651=>"001111101",
  652=>"001000110",
  653=>"011110101",
  654=>"101100011",
  655=>"110001010",
  656=>"100011011",
  657=>"001000101",
  658=>"011101011",
  659=>"111011000",
  660=>"100101111",
  661=>"101000101",
  662=>"001001001",
  663=>"001001010",
  664=>"101110100",
  665=>"001110010",
  666=>"101100111",
  667=>"101111011",
  668=>"000100001",
  669=>"000100011",
  670=>"110010100",
  671=>"100110101",
  672=>"011101010",
  673=>"101011000",
  674=>"101000011",
  675=>"100001101",
  676=>"101111001",
  677=>"010010010",
  678=>"001110011",
  679=>"100111100",
  680=>"011010001",
  681=>"100110100",
  682=>"001000001",
  683=>"100011111",
  684=>"001110011",
  685=>"100111011",
  686=>"111110110",
  687=>"001010111",
  688=>"010101000",
  689=>"101001010",
  690=>"101110110",
  691=>"110110011",
  692=>"111000110",
  693=>"100111010",
  694=>"100101011",
  695=>"111011011",
  696=>"111101011",
  697=>"100100001",
  698=>"111100011",
  699=>"101110100",
  700=>"111000100",
  701=>"000100011",
  702=>"100101010",
  703=>"011000110",
  704=>"100011111",
  705=>"110000000",
  706=>"100110101",
  707=>"101010101",
  708=>"110011101",
  709=>"001110011",
  710=>"010000110",
  711=>"111100110",
  712=>"000001011",
  713=>"100110010",
  714=>"000000100",
  715=>"011100011",
  716=>"111101010",
  717=>"010001010",
  718=>"001100100",
  719=>"100001101",
  720=>"001111110",
  721=>"101111000",
  722=>"101011000",
  723=>"000001000",
  724=>"010000101",
  725=>"110010110",
  726=>"111101110",
  727=>"000100101",
  728=>"100100101",
  729=>"011000101",
  730=>"111101101",
  731=>"010010000",
  732=>"101001111",
  733=>"111001110",
  734=>"010000000",
  735=>"111011111",
  736=>"001000111",
  737=>"100100010",
  738=>"111011110",
  739=>"110111011",
  740=>"010100001",
  741=>"010100000",
  742=>"101011000",
  743=>"100010000",
  744=>"101010100",
  745=>"001000000",
  746=>"011111001",
  747=>"001101111",
  748=>"111010000",
  749=>"111100011",
  750=>"111010111",
  751=>"100001011",
  752=>"010000100",
  753=>"001101101",
  754=>"100001111",
  755=>"011010101",
  756=>"101001010",
  757=>"110001111",
  758=>"010001101",
  759=>"011110110",
  760=>"000011001",
  761=>"101011111",
  762=>"000010011",
  763=>"001011011",
  764=>"111100110",
  765=>"000111110",
  766=>"111100000",
  767=>"011010001",
  768=>"000111110",
  769=>"001101000",
  770=>"110100101",
  771=>"000100011",
  772=>"110111100",
  773=>"110111111",
  774=>"100000111",
  775=>"000011000",
  776=>"001011010",
  777=>"011011010",
  778=>"010110011",
  779=>"100000100",
  780=>"111111110",
  781=>"000011011",
  782=>"110011011",
  783=>"111101100",
  784=>"011011100",
  785=>"001100001",
  786=>"010001000",
  787=>"110001111",
  788=>"001110000",
  789=>"001010011",
  790=>"000010100",
  791=>"010000111",
  792=>"000011011",
  793=>"010011111",
  794=>"101011011",
  795=>"101001010",
  796=>"100010110",
  797=>"101001101",
  798=>"000001110",
  799=>"110010111",
  800=>"111100000",
  801=>"011101000",
  802=>"101001110",
  803=>"010001100",
  804=>"010010100",
  805=>"111001110",
  806=>"110011001",
  807=>"000001110",
  808=>"111000111",
  809=>"000000000",
  810=>"010000010",
  811=>"101000111",
  812=>"000111001",
  813=>"110110100",
  814=>"101100110",
  815=>"011010001",
  816=>"001011001",
  817=>"111110101",
  818=>"100001000",
  819=>"010010011",
  820=>"101011010",
  821=>"101001010",
  822=>"011101010",
  823=>"100010010",
  824=>"011000110",
  825=>"011101000",
  826=>"101011001",
  827=>"100110011",
  828=>"110110110",
  829=>"001001001",
  830=>"010001110",
  831=>"000011111",
  832=>"101001110",
  833=>"100001001",
  834=>"011010111",
  835=>"000000001",
  836=>"000011000",
  837=>"010000101",
  838=>"101110101",
  839=>"000101011",
  840=>"011001111",
  841=>"100001010",
  842=>"010001001",
  843=>"000100011",
  844=>"000010101",
  845=>"001111011",
  846=>"101100011",
  847=>"100010000",
  848=>"110101010",
  849=>"000010110",
  850=>"010001110",
  851=>"000000010",
  852=>"000010010",
  853=>"111011100",
  854=>"011100000",
  855=>"000101110",
  856=>"001000010",
  857=>"001111001",
  858=>"100110010",
  859=>"110100111",
  860=>"000101010",
  861=>"000111110",
  862=>"100001011",
  863=>"111011110",
  864=>"011010111",
  865=>"000101101",
  866=>"101101000",
  867=>"110001101",
  868=>"001111000",
  869=>"011000010",
  870=>"111011010",
  871=>"011011111",
  872=>"101101100",
  873=>"111001011",
  874=>"011010110",
  875=>"110001011",
  876=>"100000010",
  877=>"101101010",
  878=>"110011110",
  879=>"000001101",
  880=>"101001110",
  881=>"000101010",
  882=>"010010001",
  883=>"101101000",
  884=>"000111111",
  885=>"110101001",
  886=>"100000010",
  887=>"001000011",
  888=>"111001101",
  889=>"101000100",
  890=>"101111010",
  891=>"010011110",
  892=>"010001011",
  893=>"001100111",
  894=>"010100011",
  895=>"110000000",
  896=>"110010011",
  897=>"100010111",
  898=>"110000010",
  899=>"011010100",
  900=>"101110111",
  901=>"001100011",
  902=>"010100010",
  903=>"100010010",
  904=>"000000101",
  905=>"001101011",
  906=>"001000001",
  907=>"010001001",
  908=>"100110011",
  909=>"110101010",
  910=>"011000100",
  911=>"110101110",
  912=>"001100010",
  913=>"100011100",
  914=>"000110100",
  915=>"010101011",
  916=>"111010111",
  917=>"100100001",
  918=>"000111011",
  919=>"001010000",
  920=>"001110101",
  921=>"011110100",
  922=>"111101111",
  923=>"100100000",
  924=>"101000001",
  925=>"000011011",
  926=>"000101100",
  927=>"001010010",
  928=>"000000100",
  929=>"100001100",
  930=>"101011101",
  931=>"011010100",
  932=>"010101010",
  933=>"010111010",
  934=>"010111000",
  935=>"110100000",
  936=>"111010011",
  937=>"100100001",
  938=>"101001110",
  939=>"100110110",
  940=>"001001101",
  941=>"000000000",
  942=>"100010000",
  943=>"100101001",
  944=>"111110111",
  945=>"011101101",
  946=>"101000000",
  947=>"111101000",
  948=>"100000011",
  949=>"101000010",
  950=>"011110111",
  951=>"000110110",
  952=>"101011101",
  953=>"000110011",
  954=>"100111110",
  955=>"100100010",
  956=>"001011101",
  957=>"110111000",
  958=>"100111010",
  959=>"111100000",
  960=>"001111000",
  961=>"000000101",
  962=>"101101111",
  963=>"000000000",
  964=>"110011001",
  965=>"100110010",
  966=>"101001101",
  967=>"010011001",
  968=>"011011001",
  969=>"110000111",
  970=>"000001000",
  971=>"011100101",
  972=>"011100100",
  973=>"011100100",
  974=>"001110000",
  975=>"001110100",
  976=>"101111101",
  977=>"101010001",
  978=>"101000101",
  979=>"010111111",
  980=>"100011010",
  981=>"000001000",
  982=>"010010110",
  983=>"001111001",
  984=>"100011010",
  985=>"001000110",
  986=>"100011010",
  987=>"010111000",
  988=>"110110001",
  989=>"011000111",
  990=>"010011110",
  991=>"010011111",
  992=>"000001110",
  993=>"111000110",
  994=>"101011000",
  995=>"010000001",
  996=>"000000000",
  997=>"100111100",
  998=>"110011010",
  999=>"000000110",
  1000=>"010100100",
  1001=>"000011010",
  1002=>"010000101",
  1003=>"000110100",
  1004=>"101111000",
  1005=>"100011100",
  1006=>"001010101",
  1007=>"101011110",
  1008=>"010111101",
  1009=>"110101101",
  1010=>"111110010",
  1011=>"001000100",
  1012=>"100110010",
  1013=>"111000001",
  1014=>"010010101",
  1015=>"000010110",
  1016=>"111000010",
  1017=>"111101100",
  1018=>"000110000",
  1019=>"010001000",
  1020=>"001111111",
  1021=>"000001100",
  1022=>"000101110",
  1023=>"011001111",
  1024=>"000000110",
  1025=>"011011100",
  1026=>"111011101",
  1027=>"101100101",
  1028=>"001100001",
  1029=>"010011011",
  1030=>"111010101",
  1031=>"011101010",
  1032=>"100100111",
  1033=>"111000010",
  1034=>"010110010",
  1035=>"101110001",
  1036=>"100110001",
  1037=>"101111011",
  1038=>"000010010",
  1039=>"011001000",
  1040=>"101101101",
  1041=>"010110111",
  1042=>"011100111",
  1043=>"010011101",
  1044=>"000001010",
  1045=>"110000100",
  1046=>"011001000",
  1047=>"011001010",
  1048=>"010010000",
  1049=>"001000010",
  1050=>"001001000",
  1051=>"011011100",
  1052=>"100010101",
  1053=>"010111111",
  1054=>"000000111",
  1055=>"001000101",
  1056=>"101101111",
  1057=>"001010110",
  1058=>"100010001",
  1059=>"010010000",
  1060=>"111001000",
  1061=>"000111001",
  1062=>"110100111",
  1063=>"111011101",
  1064=>"101111001",
  1065=>"001001011",
  1066=>"010111101",
  1067=>"011000101",
  1068=>"111111011",
  1069=>"111110010",
  1070=>"100111010",
  1071=>"110111100",
  1072=>"100101011",
  1073=>"111110001",
  1074=>"011010101",
  1075=>"001110100",
  1076=>"110000101",
  1077=>"010010101",
  1078=>"011000011",
  1079=>"110101100",
  1080=>"100001111",
  1081=>"101010001",
  1082=>"101110110",
  1083=>"001100011",
  1084=>"010100110",
  1085=>"000011101",
  1086=>"101010100",
  1087=>"101101001",
  1088=>"011001101",
  1089=>"001111110",
  1090=>"111011100",
  1091=>"001010101",
  1092=>"110100100",
  1093=>"010111010",
  1094=>"011000001",
  1095=>"100101100",
  1096=>"010000010",
  1097=>"011001111",
  1098=>"010101011",
  1099=>"111010100",
  1100=>"101111011",
  1101=>"110010110",
  1102=>"010011001",
  1103=>"110101100",
  1104=>"010000111",
  1105=>"111111111",
  1106=>"001110100",
  1107=>"011100111",
  1108=>"000000101",
  1109=>"101110001",
  1110=>"000110110",
  1111=>"100110011",
  1112=>"001010111",
  1113=>"100110110",
  1114=>"101000011",
  1115=>"100001111",
  1116=>"011111100",
  1117=>"000000110",
  1118=>"010110010",
  1119=>"110011011",
  1120=>"101010100",
  1121=>"101000000",
  1122=>"001101001",
  1123=>"001100110",
  1124=>"111001110",
  1125=>"010000000",
  1126=>"001010001",
  1127=>"100001100",
  1128=>"011001101",
  1129=>"011111111",
  1130=>"011110010",
  1131=>"000100110",
  1132=>"011110110",
  1133=>"101111101",
  1134=>"010000101",
  1135=>"110111011",
  1136=>"100011010",
  1137=>"111011000",
  1138=>"111100110",
  1139=>"001000001",
  1140=>"011100001",
  1141=>"011110010",
  1142=>"000001000",
  1143=>"111000111",
  1144=>"001010010",
  1145=>"111000111",
  1146=>"100010100",
  1147=>"000011010",
  1148=>"000100110",
  1149=>"110001001",
  1150=>"110000001",
  1151=>"110101110",
  1152=>"101000110",
  1153=>"011111011",
  1154=>"001001101",
  1155=>"000111010",
  1156=>"101101100",
  1157=>"101010000",
  1158=>"111101101",
  1159=>"100110011",
  1160=>"101100110",
  1161=>"100111100",
  1162=>"000111010",
  1163=>"011010101",
  1164=>"001001101",
  1165=>"010100110",
  1166=>"001101100",
  1167=>"000100110",
  1168=>"111010110",
  1169=>"110100011",
  1170=>"011110111",
  1171=>"011100110",
  1172=>"001010100",
  1173=>"110000010",
  1174=>"000011101",
  1175=>"001001100",
  1176=>"011101101",
  1177=>"010011010",
  1178=>"010010110",
  1179=>"011011001",
  1180=>"100100010",
  1181=>"101100001",
  1182=>"001111110",
  1183=>"001010011",
  1184=>"111101000",
  1185=>"101110000",
  1186=>"001101001",
  1187=>"110001100",
  1188=>"111001001",
  1189=>"111111001",
  1190=>"111000000",
  1191=>"001100011",
  1192=>"110010010",
  1193=>"010111110",
  1194=>"111100011",
  1195=>"011110000",
  1196=>"011011111",
  1197=>"101100101",
  1198=>"111110001",
  1199=>"101111100",
  1200=>"010010110",
  1201=>"101001110",
  1202=>"100111010",
  1203=>"000010001",
  1204=>"100010101",
  1205=>"010011101",
  1206=>"000111000",
  1207=>"011000001",
  1208=>"111011110",
  1209=>"100111101",
  1210=>"011000101",
  1211=>"011111101",
  1212=>"111111101",
  1213=>"000110010",
  1214=>"110110011",
  1215=>"111001110",
  1216=>"101101101",
  1217=>"011011101",
  1218=>"110000010",
  1219=>"001010101",
  1220=>"101100110",
  1221=>"001101000",
  1222=>"111110100",
  1223=>"101001010",
  1224=>"101110000",
  1225=>"011110010",
  1226=>"001011101",
  1227=>"111100011",
  1228=>"100101011",
  1229=>"110100000",
  1230=>"000011010",
  1231=>"001011001",
  1232=>"000010010",
  1233=>"101100000",
  1234=>"001011010",
  1235=>"101110011",
  1236=>"010001101",
  1237=>"000010111",
  1238=>"101010111",
  1239=>"101111000",
  1240=>"100101100",
  1241=>"100100000",
  1242=>"110110000",
  1243=>"111101011",
  1244=>"100101001",
  1245=>"011101110",
  1246=>"001100011",
  1247=>"101010111",
  1248=>"010101110",
  1249=>"100000101",
  1250=>"000000000",
  1251=>"111000001",
  1252=>"000011010",
  1253=>"111000110",
  1254=>"111111100",
  1255=>"011111111",
  1256=>"100000111",
  1257=>"101010100",
  1258=>"111010111",
  1259=>"101000100",
  1260=>"001101101",
  1261=>"100000000",
  1262=>"001000001",
  1263=>"001000110",
  1264=>"100000010",
  1265=>"111100000",
  1266=>"101001011",
  1267=>"001111000",
  1268=>"101010110",
  1269=>"101111101",
  1270=>"101110011",
  1271=>"111000100",
  1272=>"111011001",
  1273=>"111000010",
  1274=>"011110110",
  1275=>"001001011",
  1276=>"011110111",
  1277=>"100001100",
  1278=>"010110001",
  1279=>"100001100",
  1280=>"010110010",
  1281=>"011110100",
  1282=>"000101110",
  1283=>"100010010",
  1284=>"100000111",
  1285=>"010111110",
  1286=>"001110000",
  1287=>"110000100",
  1288=>"110101110",
  1289=>"000001001",
  1290=>"101000010",
  1291=>"101101101",
  1292=>"100111100",
  1293=>"000000001",
  1294=>"110001100",
  1295=>"100011110",
  1296=>"100111000",
  1297=>"101000100",
  1298=>"101101100",
  1299=>"110110110",
  1300=>"110000110",
  1301=>"011101000",
  1302=>"100110100",
  1303=>"111101111",
  1304=>"011100010",
  1305=>"000100111",
  1306=>"000011010",
  1307=>"110001010",
  1308=>"001110000",
  1309=>"111001010",
  1310=>"010111101",
  1311=>"101100100",
  1312=>"101111110",
  1313=>"000010000",
  1314=>"001011010",
  1315=>"000100011",
  1316=>"011100001",
  1317=>"010110000",
  1318=>"001000110",
  1319=>"100111111",
  1320=>"110101011",
  1321=>"110011111",
  1322=>"101000001",
  1323=>"011011011",
  1324=>"101010111",
  1325=>"110000011",
  1326=>"001001101",
  1327=>"110010000",
  1328=>"000101101",
  1329=>"000001101",
  1330=>"101010000",
  1331=>"100011010",
  1332=>"010100001",
  1333=>"100011011",
  1334=>"100000001",
  1335=>"001011111",
  1336=>"000011100",
  1337=>"110111110",
  1338=>"000101101",
  1339=>"010001010",
  1340=>"110010101",
  1341=>"010111011",
  1342=>"100000111",
  1343=>"001110001",
  1344=>"011101000",
  1345=>"001000010",
  1346=>"100000100",
  1347=>"000000000",
  1348=>"110111101",
  1349=>"010000111",
  1350=>"001110010",
  1351=>"011000100",
  1352=>"000100110",
  1353=>"101100101",
  1354=>"101010111",
  1355=>"011100010",
  1356=>"001100011",
  1357=>"100000000",
  1358=>"000001011",
  1359=>"000000010",
  1360=>"000011001",
  1361=>"001011100",
  1362=>"000100110",
  1363=>"010000100",
  1364=>"100101001",
  1365=>"000000001",
  1366=>"001100111",
  1367=>"100100110",
  1368=>"100101101",
  1369=>"000010101",
  1370=>"101011000",
  1371=>"100110110",
  1372=>"011010111",
  1373=>"001100011",
  1374=>"100110100",
  1375=>"101010000",
  1376=>"011110100",
  1377=>"010000010",
  1378=>"000001011",
  1379=>"011110110",
  1380=>"101001001",
  1381=>"111111010",
  1382=>"111001110",
  1383=>"000110011",
  1384=>"100011101",
  1385=>"100100110",
  1386=>"001110100",
  1387=>"000011100",
  1388=>"001010110",
  1389=>"101111110",
  1390=>"001011111",
  1391=>"101010101",
  1392=>"110011010",
  1393=>"111110001",
  1394=>"011111110",
  1395=>"100100101",
  1396=>"100111110",
  1397=>"100100001",
  1398=>"000001101",
  1399=>"000110110",
  1400=>"100000101",
  1401=>"100101110",
  1402=>"010010001",
  1403=>"101001000",
  1404=>"110111101",
  1405=>"111100010",
  1406=>"111000100",
  1407=>"111100001",
  1408=>"100111110",
  1409=>"011010001",
  1410=>"011101000",
  1411=>"000010011",
  1412=>"001100010",
  1413=>"110000010",
  1414=>"010001011",
  1415=>"000001011",
  1416=>"000000100",
  1417=>"111110111",
  1418=>"101111111",
  1419=>"111100010",
  1420=>"111010100",
  1421=>"100011100",
  1422=>"100011110",
  1423=>"010001100",
  1424=>"000110100",
  1425=>"101111111",
  1426=>"010110100",
  1427=>"111001111",
  1428=>"010111010",
  1429=>"010000111",
  1430=>"110100110",
  1431=>"100110011",
  1432=>"100000110",
  1433=>"000011110",
  1434=>"110100000",
  1435=>"101011101",
  1436=>"011000111",
  1437=>"000100100",
  1438=>"001011101",
  1439=>"001100101",
  1440=>"110101011",
  1441=>"001111111",
  1442=>"011101011",
  1443=>"000001110",
  1444=>"000011011",
  1445=>"111100011",
  1446=>"101010011",
  1447=>"011111100",
  1448=>"101001101",
  1449=>"001001111",
  1450=>"001010110",
  1451=>"110001011",
  1452=>"011010001",
  1453=>"101001011",
  1454=>"011000010",
  1455=>"001100000",
  1456=>"100100011",
  1457=>"000000100",
  1458=>"110010111",
  1459=>"001000011",
  1460=>"101101101",
  1461=>"010110010",
  1462=>"111000111",
  1463=>"110010111",
  1464=>"001001101",
  1465=>"100100101",
  1466=>"101001101",
  1467=>"100000011",
  1468=>"000001001",
  1469=>"110010000",
  1470=>"111110110",
  1471=>"001000010",
  1472=>"110000110",
  1473=>"010010001",
  1474=>"001111011",
  1475=>"010110001",
  1476=>"101100010",
  1477=>"011000111",
  1478=>"100010100",
  1479=>"111101010",
  1480=>"001111011",
  1481=>"000111111",
  1482=>"100001111",
  1483=>"111100111",
  1484=>"000100001",
  1485=>"000101101",
  1486=>"111100011",
  1487=>"101000001",
  1488=>"111110011",
  1489=>"110101011",
  1490=>"011001100",
  1491=>"010101111",
  1492=>"000101010",
  1493=>"110010111",
  1494=>"111011111",
  1495=>"101001001",
  1496=>"011011000",
  1497=>"100001111",
  1498=>"110101110",
  1499=>"010001001",
  1500=>"110010010",
  1501=>"101000001",
  1502=>"110000010",
  1503=>"001010001",
  1504=>"000001100",
  1505=>"010110011",
  1506=>"101101011",
  1507=>"011001100",
  1508=>"000110001",
  1509=>"110000111",
  1510=>"000010111",
  1511=>"100111000",
  1512=>"011001011",
  1513=>"001011101",
  1514=>"011011111",
  1515=>"000111110",
  1516=>"011100110",
  1517=>"010000101",
  1518=>"011101100",
  1519=>"110110111",
  1520=>"101100100",
  1521=>"101101100",
  1522=>"000111111",
  1523=>"001101000",
  1524=>"100010111",
  1525=>"101110101",
  1526=>"111010101",
  1527=>"101011001",
  1528=>"000011000",
  1529=>"000110100",
  1530=>"110111111",
  1531=>"001011110",
  1532=>"110011010",
  1533=>"111111000",
  1534=>"111011101",
  1535=>"010000111",
  1536=>"010111111",
  1537=>"011001001",
  1538=>"011111000",
  1539=>"101101000",
  1540=>"010111001",
  1541=>"000100110",
  1542=>"010001101",
  1543=>"101001010",
  1544=>"111111010",
  1545=>"010010100",
  1546=>"000011011",
  1547=>"111000101",
  1548=>"101010011",
  1549=>"011111001",
  1550=>"100110001",
  1551=>"001000101",
  1552=>"000110100",
  1553=>"110010100",
  1554=>"100011011",
  1555=>"011110011",
  1556=>"010101110",
  1557=>"110001010",
  1558=>"110001011",
  1559=>"001110101",
  1560=>"111110111",
  1561=>"100100010",
  1562=>"010110001",
  1563=>"100010000",
  1564=>"000101001",
  1565=>"000100111",
  1566=>"000101011",
  1567=>"010101101",
  1568=>"001011001",
  1569=>"111110000",
  1570=>"100001011",
  1571=>"011110011",
  1572=>"001110111",
  1573=>"011110111",
  1574=>"010011110",
  1575=>"110000110",
  1576=>"111111101",
  1577=>"001101101",
  1578=>"100000010",
  1579=>"000100110",
  1580=>"010110101",
  1581=>"100010100",
  1582=>"101110000",
  1583=>"010010111",
  1584=>"010001011",
  1585=>"111101110",
  1586=>"110100000",
  1587=>"001000000",
  1588=>"000101010",
  1589=>"011001110",
  1590=>"111111110",
  1591=>"001000100",
  1592=>"001101110",
  1593=>"111100000",
  1594=>"011000111",
  1595=>"101110101",
  1596=>"011101010",
  1597=>"000000001",
  1598=>"100011001",
  1599=>"000101010",
  1600=>"110101011",
  1601=>"010011110",
  1602=>"111001000",
  1603=>"011111100",
  1604=>"101111110",
  1605=>"000001010",
  1606=>"110101101",
  1607=>"100111000",
  1608=>"010000010",
  1609=>"011001101",
  1610=>"111000011",
  1611=>"001000110",
  1612=>"101011101",
  1613=>"111101111",
  1614=>"101001110",
  1615=>"000100110",
  1616=>"000101110",
  1617=>"010100010",
  1618=>"001010001",
  1619=>"110111101",
  1620=>"100000101",
  1621=>"100101110",
  1622=>"000111011",
  1623=>"010011111",
  1624=>"101100011",
  1625=>"010010110",
  1626=>"101111110",
  1627=>"000000010",
  1628=>"000100010",
  1629=>"111100111",
  1630=>"000000110",
  1631=>"010100001",
  1632=>"001010010",
  1633=>"111010100",
  1634=>"110001011",
  1635=>"111000110",
  1636=>"001000000",
  1637=>"010110111",
  1638=>"010000011",
  1639=>"000110110",
  1640=>"101101010",
  1641=>"001011100",
  1642=>"001110000",
  1643=>"010000010",
  1644=>"100111101",
  1645=>"111110111",
  1646=>"011000111",
  1647=>"111001101",
  1648=>"100011001",
  1649=>"011001011",
  1650=>"100010101",
  1651=>"111111110",
  1652=>"101010011",
  1653=>"100010100",
  1654=>"010110101",
  1655=>"011100011",
  1656=>"111101111",
  1657=>"101101100",
  1658=>"100110100",
  1659=>"110111001",
  1660=>"110111110",
  1661=>"100011100",
  1662=>"011100110",
  1663=>"000111001",
  1664=>"010010001",
  1665=>"010100011",
  1666=>"101101001",
  1667=>"110010111",
  1668=>"101111010",
  1669=>"101001001",
  1670=>"100101010",
  1671=>"000001000",
  1672=>"000010110",
  1673=>"010110011",
  1674=>"110110011",
  1675=>"101101000",
  1676=>"000111111",
  1677=>"011101100",
  1678=>"010100001",
  1679=>"011010011",
  1680=>"001100101",
  1681=>"000101000",
  1682=>"111010101",
  1683=>"111100001",
  1684=>"010100001",
  1685=>"110001111",
  1686=>"110101100",
  1687=>"100101100",
  1688=>"000000000",
  1689=>"000110101",
  1690=>"110110100",
  1691=>"001111110",
  1692=>"111001010",
  1693=>"101101111",
  1694=>"000111010",
  1695=>"001001101",
  1696=>"001110100",
  1697=>"101010001",
  1698=>"101010000",
  1699=>"110101100",
  1700=>"101111011",
  1701=>"001010010",
  1702=>"110010111",
  1703=>"000100101",
  1704=>"111001110",
  1705=>"000100101",
  1706=>"001100000",
  1707=>"010101010",
  1708=>"111110000",
  1709=>"011001110",
  1710=>"011101110",
  1711=>"101011011",
  1712=>"010100101",
  1713=>"000100100",
  1714=>"000010100",
  1715=>"001101001",
  1716=>"111100011",
  1717=>"101111011",
  1718=>"111111110",
  1719=>"010100100",
  1720=>"101010011",
  1721=>"101010110",
  1722=>"101111011",
  1723=>"000000010",
  1724=>"100111110",
  1725=>"111110001",
  1726=>"111111100",
  1727=>"000000101",
  1728=>"111001110",
  1729=>"111010100",
  1730=>"101100000",
  1731=>"001000001",
  1732=>"010110000",
  1733=>"000001100",
  1734=>"000000010",
  1735=>"000000100",
  1736=>"011010110",
  1737=>"010110101",
  1738=>"000011001",
  1739=>"110100111",
  1740=>"100100011",
  1741=>"011010101",
  1742=>"001111010",
  1743=>"001000001",
  1744=>"100110111",
  1745=>"111111111",
  1746=>"011000100",
  1747=>"001111000",
  1748=>"110001010",
  1749=>"000100010",
  1750=>"011111111",
  1751=>"110100101",
  1752=>"000101101",
  1753=>"111010010",
  1754=>"011101111",
  1755=>"010101011",
  1756=>"010101011",
  1757=>"110111111",
  1758=>"011111111",
  1759=>"011001000",
  1760=>"111011111",
  1761=>"010000111",
  1762=>"000000010",
  1763=>"110111100",
  1764=>"010001000",
  1765=>"110001100",
  1766=>"111100000",
  1767=>"110000000",
  1768=>"000011101",
  1769=>"100111111",
  1770=>"011011010",
  1771=>"001000000",
  1772=>"100001010",
  1773=>"101101110",
  1774=>"000110111",
  1775=>"100111001",
  1776=>"110101000",
  1777=>"110000010",
  1778=>"110000001",
  1779=>"111000011",
  1780=>"000111110",
  1781=>"000001000",
  1782=>"010001001",
  1783=>"111111111",
  1784=>"110110001",
  1785=>"100110100",
  1786=>"010000001",
  1787=>"011110001",
  1788=>"111100001",
  1789=>"000011100",
  1790=>"100000011",
  1791=>"000111101",
  1792=>"110110111",
  1793=>"101100000",
  1794=>"010110010",
  1795=>"001000010",
  1796=>"110111111",
  1797=>"110010011",
  1798=>"100010100",
  1799=>"110000101",
  1800=>"110010110",
  1801=>"100100001",
  1802=>"011110111",
  1803=>"001101000",
  1804=>"011100110",
  1805=>"101001010",
  1806=>"010011011",
  1807=>"100110000",
  1808=>"110100011",
  1809=>"100000001",
  1810=>"001101010",
  1811=>"011101100",
  1812=>"011011111",
  1813=>"110100011",
  1814=>"001000010",
  1815=>"110101111",
  1816=>"000110100",
  1817=>"010110101",
  1818=>"000100001",
  1819=>"001110101",
  1820=>"001011100",
  1821=>"011100000",
  1822=>"100101110",
  1823=>"001111100",
  1824=>"110110001",
  1825=>"101111010",
  1826=>"011010010",
  1827=>"000001110",
  1828=>"011110111",
  1829=>"111111101",
  1830=>"010010101",
  1831=>"010101011",
  1832=>"010000101",
  1833=>"000111101",
  1834=>"001111001",
  1835=>"101111011",
  1836=>"111101001",
  1837=>"001100100",
  1838=>"100100001",
  1839=>"100100100",
  1840=>"111010011",
  1841=>"110100111",
  1842=>"101010011",
  1843=>"001101000",
  1844=>"111100111",
  1845=>"110100000",
  1846=>"101110000",
  1847=>"000010110",
  1848=>"100001010",
  1849=>"010011010",
  1850=>"111111101",
  1851=>"110110010",
  1852=>"001011100",
  1853=>"100100010",
  1854=>"000110010",
  1855=>"010110100",
  1856=>"100111011",
  1857=>"101100001",
  1858=>"101111101",
  1859=>"101110100",
  1860=>"110100011",
  1861=>"001010111",
  1862=>"110100111",
  1863=>"000111111",
  1864=>"011110100",
  1865=>"111101111",
  1866=>"110010100",
  1867=>"111011011",
  1868=>"001001011",
  1869=>"111010100",
  1870=>"000110110",
  1871=>"101010100",
  1872=>"110010101",
  1873=>"010000111",
  1874=>"011011111",
  1875=>"011100101",
  1876=>"101101110",
  1877=>"101101010",
  1878=>"100010011",
  1879=>"011010000",
  1880=>"001000011",
  1881=>"111100011",
  1882=>"011100110",
  1883=>"111011011",
  1884=>"110101100",
  1885=>"001101000",
  1886=>"111111000",
  1887=>"100000111",
  1888=>"111011010",
  1889=>"010010011",
  1890=>"110011000",
  1891=>"001100011",
  1892=>"110110000",
  1893=>"001001000",
  1894=>"101110111",
  1895=>"010010110",
  1896=>"110100001",
  1897=>"001110011",
  1898=>"111111010",
  1899=>"111001101",
  1900=>"001110000",
  1901=>"000000100",
  1902=>"010101110",
  1903=>"110011000",
  1904=>"010101000",
  1905=>"001111001",
  1906=>"111100001",
  1907=>"100111001",
  1908=>"000010101",
  1909=>"000001101",
  1910=>"100110111",
  1911=>"111010010",
  1912=>"011000000",
  1913=>"101101111",
  1914=>"000000100",
  1915=>"001101001",
  1916=>"000100001",
  1917=>"100101111",
  1918=>"010010011",
  1919=>"101110010",
  1920=>"101011100",
  1921=>"011010100",
  1922=>"001100111",
  1923=>"110000010",
  1924=>"100011111",
  1925=>"001000000",
  1926=>"011011010",
  1927=>"111110111",
  1928=>"111100001",
  1929=>"110001001",
  1930=>"000100101",
  1931=>"101111001",
  1932=>"110111000",
  1933=>"000100111",
  1934=>"110100000",
  1935=>"011110110",
  1936=>"110101011",
  1937=>"000001000",
  1938=>"011010001",
  1939=>"000100000",
  1940=>"011000101",
  1941=>"110101100",
  1942=>"001110000",
  1943=>"011100100",
  1944=>"010011010",
  1945=>"111101101",
  1946=>"001110100",
  1947=>"001011010",
  1948=>"011011101",
  1949=>"001011011",
  1950=>"010100100",
  1951=>"011110010",
  1952=>"011100010",
  1953=>"011111000",
  1954=>"000111001",
  1955=>"110000110",
  1956=>"101100100",
  1957=>"001110101",
  1958=>"101101101",
  1959=>"100010110",
  1960=>"010101010",
  1961=>"010010000",
  1962=>"100001100",
  1963=>"100101101",
  1964=>"011100011",
  1965=>"111101011",
  1966=>"010100011",
  1967=>"001010011",
  1968=>"000010100",
  1969=>"110101101",
  1970=>"101110000",
  1971=>"111110010",
  1972=>"011110011",
  1973=>"101100010",
  1974=>"001100101",
  1975=>"111111111",
  1976=>"010111011",
  1977=>"001110000",
  1978=>"011010011",
  1979=>"101000111",
  1980=>"001011000",
  1981=>"011100100",
  1982=>"111101010",
  1983=>"001100000",
  1984=>"101011010",
  1985=>"011110001",
  1986=>"010001010",
  1987=>"011110111",
  1988=>"011101010",
  1989=>"000101111",
  1990=>"011000010",
  1991=>"000011000",
  1992=>"001100110",
  1993=>"110100010",
  1994=>"010010110",
  1995=>"011101110",
  1996=>"110011100",
  1997=>"101100110",
  1998=>"000101010",
  1999=>"100010001",
  2000=>"011000001",
  2001=>"010100110",
  2002=>"111100010",
  2003=>"000000000",
  2004=>"111101111",
  2005=>"001000000",
  2006=>"101111010",
  2007=>"011110010",
  2008=>"010001111",
  2009=>"101101110",
  2010=>"110001011",
  2011=>"110100001",
  2012=>"111010010",
  2013=>"000100110",
  2014=>"101111111",
  2015=>"010010101",
  2016=>"101010000",
  2017=>"010110100",
  2018=>"001011010",
  2019=>"000101010",
  2020=>"110100111",
  2021=>"000010001",
  2022=>"011110111",
  2023=>"100111010",
  2024=>"010100110",
  2025=>"111100110",
  2026=>"110001001",
  2027=>"001010000",
  2028=>"111111010",
  2029=>"001000100",
  2030=>"111000111",
  2031=>"011111011",
  2032=>"101101011",
  2033=>"010101111",
  2034=>"000000000",
  2035=>"111111100",
  2036=>"001001001",
  2037=>"011000000",
  2038=>"111110100",
  2039=>"010100000",
  2040=>"010011100",
  2041=>"110110001",
  2042=>"111101111",
  2043=>"001000010",
  2044=>"000101110",
  2045=>"001111100",
  2046=>"010000101",
  2047=>"110101111",
  2048=>"111000011",
  2049=>"101011000",
  2050=>"010011110",
  2051=>"000000000",
  2052=>"001100100",
  2053=>"100011101",
  2054=>"000011101",
  2055=>"000010001",
  2056=>"110100100",
  2057=>"111111101",
  2058=>"010101110",
  2059=>"001000010",
  2060=>"110011101",
  2061=>"001011101",
  2062=>"111111111",
  2063=>"101000001",
  2064=>"101110001",
  2065=>"110100100",
  2066=>"100010101",
  2067=>"010010001",
  2068=>"011000101",
  2069=>"000010000",
  2070=>"110000001",
  2071=>"001010001",
  2072=>"101101001",
  2073=>"001000101",
  2074=>"110101011",
  2075=>"001000100",
  2076=>"100010100",
  2077=>"110010100",
  2078=>"000110111",
  2079=>"110110000",
  2080=>"000110111",
  2081=>"100010000",
  2082=>"110111101",
  2083=>"011001010",
  2084=>"010111110",
  2085=>"100000011",
  2086=>"000111100",
  2087=>"011000100",
  2088=>"011110010",
  2089=>"101111111",
  2090=>"111110100",
  2091=>"011001110",
  2092=>"011010000",
  2093=>"110010011",
  2094=>"100101100",
  2095=>"001101110",
  2096=>"110100010",
  2097=>"011001000",
  2098=>"011001010",
  2099=>"101010111",
  2100=>"110100000",
  2101=>"010110000",
  2102=>"101001100",
  2103=>"111111100",
  2104=>"001110111",
  2105=>"011010011",
  2106=>"101001111",
  2107=>"010001111",
  2108=>"111001011",
  2109=>"111010011",
  2110=>"111100100",
  2111=>"001110001",
  2112=>"111101000",
  2113=>"000000011",
  2114=>"011111101",
  2115=>"101100001",
  2116=>"000101000",
  2117=>"001100000",
  2118=>"000000011",
  2119=>"001011000",
  2120=>"010010011",
  2121=>"111100001",
  2122=>"000111010",
  2123=>"011000010",
  2124=>"111000111",
  2125=>"111011001",
  2126=>"111110010",
  2127=>"100111001",
  2128=>"110000101",
  2129=>"110100001",
  2130=>"111011011",
  2131=>"101110000",
  2132=>"001000010",
  2133=>"100010001",
  2134=>"100100010",
  2135=>"000000100",
  2136=>"101100010",
  2137=>"010011001",
  2138=>"001000100",
  2139=>"110000001",
  2140=>"000110010",
  2141=>"000010101",
  2142=>"100011000",
  2143=>"000100000",
  2144=>"010100111",
  2145=>"110100000",
  2146=>"000000001",
  2147=>"000011011",
  2148=>"111001001",
  2149=>"000010111",
  2150=>"100100011",
  2151=>"111000111",
  2152=>"110111100",
  2153=>"111111011",
  2154=>"011001000",
  2155=>"110111111",
  2156=>"111101101",
  2157=>"100110000",
  2158=>"011011000",
  2159=>"100011101",
  2160=>"111011010",
  2161=>"001110111",
  2162=>"010011010",
  2163=>"101110111",
  2164=>"100011000",
  2165=>"010011101",
  2166=>"000110000",
  2167=>"101011111",
  2168=>"011101100",
  2169=>"111101010",
  2170=>"101010001",
  2171=>"111000000",
  2172=>"010111000",
  2173=>"101010000",
  2174=>"111100010",
  2175=>"101010000",
  2176=>"010011001",
  2177=>"010111100",
  2178=>"011010111",
  2179=>"000000110",
  2180=>"100100000",
  2181=>"001101010",
  2182=>"111111011",
  2183=>"000100000",
  2184=>"110111111",
  2185=>"001010110",
  2186=>"011001000",
  2187=>"111100100",
  2188=>"000011100",
  2189=>"010011110",
  2190=>"110001101",
  2191=>"001011011",
  2192=>"111111110",
  2193=>"010110011",
  2194=>"010011000",
  2195=>"100001111",
  2196=>"001010110",
  2197=>"101100000",
  2198=>"000101001",
  2199=>"000110101",
  2200=>"101111110",
  2201=>"011110100",
  2202=>"011111111",
  2203=>"000000100",
  2204=>"110010101",
  2205=>"100000100",
  2206=>"101100010",
  2207=>"000101101",
  2208=>"110010111",
  2209=>"111111000",
  2210=>"001110100",
  2211=>"110110111",
  2212=>"001100110",
  2213=>"100111110",
  2214=>"101100011",
  2215=>"001110111",
  2216=>"100001010",
  2217=>"010100010",
  2218=>"110010010",
  2219=>"001100000",
  2220=>"110001011",
  2221=>"111011001",
  2222=>"100111101",
  2223=>"110001001",
  2224=>"101111000",
  2225=>"001111011",
  2226=>"101100001",
  2227=>"111110000",
  2228=>"010001110",
  2229=>"000111111",
  2230=>"010111110",
  2231=>"001010100",
  2232=>"010100000",
  2233=>"110010111",
  2234=>"001000111",
  2235=>"001111011",
  2236=>"101111101",
  2237=>"010011101",
  2238=>"010111111",
  2239=>"111001010",
  2240=>"011110000",
  2241=>"011110011",
  2242=>"100001101",
  2243=>"111101101",
  2244=>"111010010",
  2245=>"010111001",
  2246=>"100110000",
  2247=>"010111101",
  2248=>"101011101",
  2249=>"001000011",
  2250=>"111111001",
  2251=>"010111100",
  2252=>"110001101",
  2253=>"000111010",
  2254=>"011111011",
  2255=>"101011011",
  2256=>"111110010",
  2257=>"101011110",
  2258=>"000010000",
  2259=>"010101111",
  2260=>"001010001",
  2261=>"111011011",
  2262=>"101000001",
  2263=>"101001011",
  2264=>"010011100",
  2265=>"110000011",
  2266=>"001001110",
  2267=>"111011110",
  2268=>"010000001",
  2269=>"010100101",
  2270=>"001110000",
  2271=>"011100010",
  2272=>"001100111",
  2273=>"000000010",
  2274=>"110010100",
  2275=>"000100110",
  2276=>"010110000",
  2277=>"000111101",
  2278=>"011100100",
  2279=>"000100000",
  2280=>"000100010",
  2281=>"100010011",
  2282=>"011110010",
  2283=>"011000100",
  2284=>"100010101",
  2285=>"111000000",
  2286=>"001111101",
  2287=>"011110110",
  2288=>"010000110",
  2289=>"000011100",
  2290=>"110011000",
  2291=>"000001110",
  2292=>"110010001",
  2293=>"000001001",
  2294=>"011000001",
  2295=>"001110101",
  2296=>"001011110",
  2297=>"110001000",
  2298=>"000010110",
  2299=>"110111001",
  2300=>"011000000",
  2301=>"000011110",
  2302=>"010011111",
  2303=>"111110001",
  2304=>"011010101",
  2305=>"001101010",
  2306=>"110100001",
  2307=>"001000000",
  2308=>"011001111",
  2309=>"010000101",
  2310=>"111100010",
  2311=>"011111011",
  2312=>"010100011",
  2313=>"110001000",
  2314=>"111111000",
  2315=>"100000000",
  2316=>"010011100",
  2317=>"011010000",
  2318=>"110011001",
  2319=>"000010111",
  2320=>"111110001",
  2321=>"110100001",
  2322=>"000111100",
  2323=>"110100001",
  2324=>"110111101",
  2325=>"110011110",
  2326=>"011011101",
  2327=>"100110100",
  2328=>"101110100",
  2329=>"100011100",
  2330=>"000001111",
  2331=>"111001011",
  2332=>"100011010",
  2333=>"110010000",
  2334=>"010101100",
  2335=>"001001101",
  2336=>"000101001",
  2337=>"001010001",
  2338=>"110001100",
  2339=>"100010101",
  2340=>"111110001",
  2341=>"011110011",
  2342=>"011000011",
  2343=>"111111000",
  2344=>"111011010",
  2345=>"110010001",
  2346=>"000001000",
  2347=>"101100110",
  2348=>"101000110",
  2349=>"101011111",
  2350=>"000001101",
  2351=>"101011111",
  2352=>"000001111",
  2353=>"110100001",
  2354=>"000001100",
  2355=>"010111000",
  2356=>"100000001",
  2357=>"000000111",
  2358=>"100010000",
  2359=>"011010000",
  2360=>"000000010",
  2361=>"110001110",
  2362=>"111011000",
  2363=>"010010010",
  2364=>"110001100",
  2365=>"110110100",
  2366=>"000101011",
  2367=>"001100100",
  2368=>"010100101",
  2369=>"011000010",
  2370=>"001110110",
  2371=>"110111000",
  2372=>"000011111",
  2373=>"001100000",
  2374=>"010101101",
  2375=>"000001101",
  2376=>"100000001",
  2377=>"011000011",
  2378=>"011001111",
  2379=>"110000111",
  2380=>"001111000",
  2381=>"110011001",
  2382=>"101110100",
  2383=>"010111011",
  2384=>"001110100",
  2385=>"101111001",
  2386=>"101101001",
  2387=>"100111110",
  2388=>"000101000",
  2389=>"110001101",
  2390=>"000101101",
  2391=>"000101111",
  2392=>"001100011",
  2393=>"011111011",
  2394=>"001110000",
  2395=>"010000110",
  2396=>"001111101",
  2397=>"000011100",
  2398=>"011011101",
  2399=>"111010111",
  2400=>"010000001",
  2401=>"000100100",
  2402=>"010001101",
  2403=>"001111111",
  2404=>"000000001",
  2405=>"111010101",
  2406=>"111011011",
  2407=>"011111100",
  2408=>"010000110",
  2409=>"010000110",
  2410=>"101000000",
  2411=>"111000100",
  2412=>"100101010",
  2413=>"011010100",
  2414=>"110100001",
  2415=>"001010111",
  2416=>"010110110",
  2417=>"110101010",
  2418=>"010100000",
  2419=>"101010110",
  2420=>"010001101",
  2421=>"001011101",
  2422=>"010111011",
  2423=>"110010000",
  2424=>"011101000",
  2425=>"101011100",
  2426=>"010001011",
  2427=>"011111011",
  2428=>"000101010",
  2429=>"001100101",
  2430=>"100101001",
  2431=>"011101001",
  2432=>"011110010",
  2433=>"010100111",
  2434=>"100111000",
  2435=>"111100010",
  2436=>"011001111",
  2437=>"011010001",
  2438=>"111001101",
  2439=>"110010000",
  2440=>"110010010",
  2441=>"101100101",
  2442=>"111010111",
  2443=>"100011001",
  2444=>"011011100",
  2445=>"100101111",
  2446=>"101101111",
  2447=>"111101010",
  2448=>"011010000",
  2449=>"001011111",
  2450=>"000110100",
  2451=>"000101111",
  2452=>"110100101",
  2453=>"110101000",
  2454=>"001111101",
  2455=>"111101100",
  2456=>"010110011",
  2457=>"110110001",
  2458=>"001010011",
  2459=>"011000000",
  2460=>"110101101",
  2461=>"110010100",
  2462=>"011111000",
  2463=>"110100001",
  2464=>"011011001",
  2465=>"101000000",
  2466=>"111101000",
  2467=>"111000000",
  2468=>"100000111",
  2469=>"011001100",
  2470=>"111000111",
  2471=>"011010010",
  2472=>"101010101",
  2473=>"001010111",
  2474=>"000111111",
  2475=>"100001110",
  2476=>"001100101",
  2477=>"101010011",
  2478=>"000111111",
  2479=>"111001011",
  2480=>"001000111",
  2481=>"001101001",
  2482=>"001011011",
  2483=>"011001100",
  2484=>"101100000",
  2485=>"011011100",
  2486=>"000010000",
  2487=>"011011011",
  2488=>"100011101",
  2489=>"101010010",
  2490=>"001001110",
  2491=>"100110110",
  2492=>"011100101",
  2493=>"010011100",
  2494=>"001110100",
  2495=>"110011111",
  2496=>"100011000",
  2497=>"000101000",
  2498=>"001010000",
  2499=>"100111011",
  2500=>"111001100",
  2501=>"111111001",
  2502=>"101100100",
  2503=>"100000110",
  2504=>"110110100",
  2505=>"010101001",
  2506=>"011101000",
  2507=>"001111011",
  2508=>"000110011",
  2509=>"111101011",
  2510=>"001101001",
  2511=>"001011110",
  2512=>"111011001",
  2513=>"011111010",
  2514=>"000111011",
  2515=>"000100110",
  2516=>"111111101",
  2517=>"001101100",
  2518=>"101000100",
  2519=>"011001100",
  2520=>"110010111",
  2521=>"101000001",
  2522=>"001100110",
  2523=>"001001000",
  2524=>"100100101",
  2525=>"101010100",
  2526=>"010011001",
  2527=>"100100101",
  2528=>"011100111",
  2529=>"001000010",
  2530=>"110001000",
  2531=>"100011000",
  2532=>"010001101",
  2533=>"011110010",
  2534=>"100001100",
  2535=>"111100001",
  2536=>"100101000",
  2537=>"100100101",
  2538=>"100110001",
  2539=>"111000000",
  2540=>"011111101",
  2541=>"000110111",
  2542=>"110001010",
  2543=>"001111111",
  2544=>"001100101",
  2545=>"001100110",
  2546=>"110001000",
  2547=>"101010010",
  2548=>"011011101",
  2549=>"000100100",
  2550=>"000101010",
  2551=>"010101100",
  2552=>"111000110",
  2553=>"111010001",
  2554=>"011100101",
  2555=>"000101111",
  2556=>"011110011",
  2557=>"100000101",
  2558=>"001111110",
  2559=>"001100111",
  2560=>"100100010",
  2561=>"001101111",
  2562=>"100010101",
  2563=>"101010100",
  2564=>"101110010",
  2565=>"111101111",
  2566=>"010000111",
  2567=>"100101111",
  2568=>"111001111",
  2569=>"010100000",
  2570=>"010010101",
  2571=>"010000010",
  2572=>"110001001",
  2573=>"001101100",
  2574=>"010010101",
  2575=>"111001011",
  2576=>"001000010",
  2577=>"111010111",
  2578=>"101101110",
  2579=>"000000010",
  2580=>"010010010",
  2581=>"000110110",
  2582=>"000010010",
  2583=>"110010100",
  2584=>"111110110",
  2585=>"011110111",
  2586=>"111110110",
  2587=>"001010010",
  2588=>"000001001",
  2589=>"000000110",
  2590=>"010010000",
  2591=>"100000011",
  2592=>"011101110",
  2593=>"010011101",
  2594=>"010010110",
  2595=>"100100011",
  2596=>"010011110",
  2597=>"111010100",
  2598=>"110010100",
  2599=>"010110100",
  2600=>"001010101",
  2601=>"010011010",
  2602=>"111110000",
  2603=>"101111111",
  2604=>"011001000",
  2605=>"001011011",
  2606=>"001110111",
  2607=>"111011101",
  2608=>"110111110",
  2609=>"010111100",
  2610=>"100011001",
  2611=>"101100111",
  2612=>"001111000",
  2613=>"111001011",
  2614=>"011111100",
  2615=>"000001000",
  2616=>"101010110",
  2617=>"101001000",
  2618=>"001001110",
  2619=>"000000110",
  2620=>"010100010",
  2621=>"001001000",
  2622=>"011110110",
  2623=>"110101111",
  2624=>"001111001",
  2625=>"001011100",
  2626=>"100010010",
  2627=>"111010001",
  2628=>"111010011",
  2629=>"000000101",
  2630=>"101010101",
  2631=>"000101011",
  2632=>"100101000",
  2633=>"100101101",
  2634=>"100100110",
  2635=>"000100011",
  2636=>"010010100",
  2637=>"011011010",
  2638=>"101010111",
  2639=>"110011001",
  2640=>"101111111",
  2641=>"010000000",
  2642=>"111010010",
  2643=>"001001110",
  2644=>"101011001",
  2645=>"000000010",
  2646=>"101011100",
  2647=>"110000011",
  2648=>"101100111",
  2649=>"011000000",
  2650=>"000100101",
  2651=>"000111100",
  2652=>"011010100",
  2653=>"000001001",
  2654=>"000100010",
  2655=>"110001000",
  2656=>"101101000",
  2657=>"001111111",
  2658=>"011010110",
  2659=>"101001110",
  2660=>"100011101",
  2661=>"100000111",
  2662=>"001010100",
  2663=>"111110010",
  2664=>"000110001",
  2665=>"010010100",
  2666=>"000010011",
  2667=>"001101111",
  2668=>"001011110",
  2669=>"011111011",
  2670=>"101011100",
  2671=>"110111100",
  2672=>"000000001",
  2673=>"001101010",
  2674=>"011001110",
  2675=>"000101110",
  2676=>"100101000",
  2677=>"101010101",
  2678=>"010101111",
  2679=>"101001100",
  2680=>"010001001",
  2681=>"101101001",
  2682=>"101111010",
  2683=>"000010010",
  2684=>"001111110",
  2685=>"010000100",
  2686=>"111101010",
  2687=>"001000001",
  2688=>"000011110",
  2689=>"101100110",
  2690=>"111111100",
  2691=>"010101100",
  2692=>"100000001",
  2693=>"100110000",
  2694=>"011000100",
  2695=>"000111100",
  2696=>"110001110",
  2697=>"001011011",
  2698=>"000110110",
  2699=>"110001000",
  2700=>"100001011",
  2701=>"111100111",
  2702=>"001111000",
  2703=>"000001000",
  2704=>"011101111",
  2705=>"111101111",
  2706=>"101100110",
  2707=>"000101100",
  2708=>"011011101",
  2709=>"111111010",
  2710=>"100111000",
  2711=>"000000011",
  2712=>"101101011",
  2713=>"000111110",
  2714=>"111101100",
  2715=>"001000010",
  2716=>"111001111",
  2717=>"010101010",
  2718=>"010101101",
  2719=>"000000011",
  2720=>"111110111",
  2721=>"101100000",
  2722=>"111011110",
  2723=>"011110010",
  2724=>"000101011",
  2725=>"101011101",
  2726=>"101101111",
  2727=>"111000001",
  2728=>"110111110",
  2729=>"011101101",
  2730=>"001101101",
  2731=>"011101010",
  2732=>"101011100",
  2733=>"101001001",
  2734=>"100001011",
  2735=>"111110010",
  2736=>"010001010",
  2737=>"110100010",
  2738=>"100110110",
  2739=>"011011100",
  2740=>"001111111",
  2741=>"011011001",
  2742=>"100001001",
  2743=>"111101011",
  2744=>"011001100",
  2745=>"101001101",
  2746=>"100000011",
  2747=>"000110111",
  2748=>"000000000",
  2749=>"110110000",
  2750=>"001100001",
  2751=>"010001011",
  2752=>"010110011",
  2753=>"111000101",
  2754=>"001101001",
  2755=>"011000010",
  2756=>"011001011",
  2757=>"010011001",
  2758=>"111110000",
  2759=>"001000011",
  2760=>"111110100",
  2761=>"011110101",
  2762=>"000011100",
  2763=>"111000110",
  2764=>"011001100",
  2765=>"101010000",
  2766=>"110101101",
  2767=>"101101101",
  2768=>"011101111",
  2769=>"111011011",
  2770=>"100010010",
  2771=>"011010011",
  2772=>"001100000",
  2773=>"000000110",
  2774=>"110101011",
  2775=>"110111011",
  2776=>"111000001",
  2777=>"110111100",
  2778=>"101001110",
  2779=>"111111111",
  2780=>"001011010",
  2781=>"011101011",
  2782=>"010110010",
  2783=>"100000000",
  2784=>"110001110",
  2785=>"000001111",
  2786=>"010011001",
  2787=>"100010010",
  2788=>"100011000",
  2789=>"101101011",
  2790=>"110110011",
  2791=>"010011110",
  2792=>"101111100",
  2793=>"001001100",
  2794=>"100000000",
  2795=>"001001001",
  2796=>"000000001",
  2797=>"000010101",
  2798=>"010011001",
  2799=>"011110000",
  2800=>"101101101",
  2801=>"111001100",
  2802=>"001010100",
  2803=>"100101010",
  2804=>"100000000",
  2805=>"011010001",
  2806=>"010111101",
  2807=>"011010100",
  2808=>"110011101",
  2809=>"011111110",
  2810=>"101000111",
  2811=>"110000010",
  2812=>"111010111",
  2813=>"110010101",
  2814=>"001010001",
  2815=>"111000101",
  2816=>"101110111",
  2817=>"010110101",
  2818=>"101100100",
  2819=>"001001110",
  2820=>"110100100",
  2821=>"110000010",
  2822=>"011100000",
  2823=>"010110000",
  2824=>"000010101",
  2825=>"001001001",
  2826=>"110010111",
  2827=>"110010001",
  2828=>"000000011",
  2829=>"100111100",
  2830=>"111111111",
  2831=>"101101110",
  2832=>"011111111",
  2833=>"111100111",
  2834=>"011101010",
  2835=>"010010000",
  2836=>"001110110",
  2837=>"110111101",
  2838=>"111100011",
  2839=>"010001111",
  2840=>"011111101",
  2841=>"011001001",
  2842=>"000001111",
  2843=>"000001100",
  2844=>"110001111",
  2845=>"110100010",
  2846=>"101000011",
  2847=>"111101001",
  2848=>"101111100",
  2849=>"111010000",
  2850=>"100101000",
  2851=>"101101111",
  2852=>"011000001",
  2853=>"001010101",
  2854=>"100101011",
  2855=>"101011001",
  2856=>"101011001",
  2857=>"111101001",
  2858=>"001000011",
  2859=>"000110001",
  2860=>"011101100",
  2861=>"010001011",
  2862=>"111101111",
  2863=>"101111111",
  2864=>"011101111",
  2865=>"010010100",
  2866=>"111010000",
  2867=>"101011001",
  2868=>"100001111",
  2869=>"110001110",
  2870=>"111001010",
  2871=>"111001100",
  2872=>"110111010",
  2873=>"111011001",
  2874=>"101000111",
  2875=>"100001011",
  2876=>"110010100",
  2877=>"000001101",
  2878=>"000000001",
  2879=>"001101001",
  2880=>"101110110",
  2881=>"111110100",
  2882=>"010011111",
  2883=>"110010101",
  2884=>"111000110",
  2885=>"111000011",
  2886=>"000110011",
  2887=>"111011011",
  2888=>"111110011",
  2889=>"100001101",
  2890=>"000010001",
  2891=>"110110011",
  2892=>"000011111",
  2893=>"011100010",
  2894=>"011110100",
  2895=>"001011100",
  2896=>"011101111",
  2897=>"100001101",
  2898=>"111101111",
  2899=>"011100011",
  2900=>"111000001",
  2901=>"010111110",
  2902=>"000110111",
  2903=>"110001000",
  2904=>"010010010",
  2905=>"001101001",
  2906=>"110011001",
  2907=>"010011011",
  2908=>"100010100",
  2909=>"101000000",
  2910=>"011000000",
  2911=>"000010011",
  2912=>"111101010",
  2913=>"110011100",
  2914=>"000010101",
  2915=>"111010001",
  2916=>"011110100",
  2917=>"110111000",
  2918=>"010000101",
  2919=>"000001001",
  2920=>"111000000",
  2921=>"001101111",
  2922=>"001011011",
  2923=>"000101010",
  2924=>"111101010",
  2925=>"010010110",
  2926=>"000010001",
  2927=>"011100000",
  2928=>"000001111",
  2929=>"101010001",
  2930=>"110011011",
  2931=>"011110011",
  2932=>"010111100",
  2933=>"000100010",
  2934=>"111101011",
  2935=>"110101111",
  2936=>"010111100",
  2937=>"011111001",
  2938=>"011111101",
  2939=>"111100100",
  2940=>"000001010",
  2941=>"111110010",
  2942=>"000100111",
  2943=>"101011000",
  2944=>"011011001",
  2945=>"010011101",
  2946=>"111011011",
  2947=>"000001000",
  2948=>"111000110",
  2949=>"111001110",
  2950=>"000001011",
  2951=>"101011000",
  2952=>"101000100",
  2953=>"101011110",
  2954=>"010110010",
  2955=>"011000101",
  2956=>"100001010",
  2957=>"001000001",
  2958=>"111110011",
  2959=>"000001111",
  2960=>"011011100",
  2961=>"010111010",
  2962=>"000001100",
  2963=>"010011101",
  2964=>"100111011",
  2965=>"110001011",
  2966=>"001111101",
  2967=>"101011001",
  2968=>"000100001",
  2969=>"111001011",
  2970=>"101101001",
  2971=>"001110010",
  2972=>"111011111",
  2973=>"001000110",
  2974=>"101000001",
  2975=>"001100111",
  2976=>"011000100",
  2977=>"000100011",
  2978=>"011001100",
  2979=>"100100110",
  2980=>"001010101",
  2981=>"010110011",
  2982=>"000100101",
  2983=>"110001111",
  2984=>"000101100",
  2985=>"010100111",
  2986=>"011111111",
  2987=>"110111110",
  2988=>"010111110",
  2989=>"010111111",
  2990=>"010110000",
  2991=>"111101000",
  2992=>"110000010",
  2993=>"001100001",
  2994=>"001011011",
  2995=>"110010100",
  2996=>"101010100",
  2997=>"010100000",
  2998=>"010000010",
  2999=>"000000010",
  3000=>"001011101",
  3001=>"010010101",
  3002=>"100101110",
  3003=>"111110101",
  3004=>"110010101",
  3005=>"001110111",
  3006=>"111100100",
  3007=>"001110100",
  3008=>"101111101",
  3009=>"011000001",
  3010=>"001100100",
  3011=>"000000110",
  3012=>"110010101",
  3013=>"010110101",
  3014=>"000001111",
  3015=>"111001111",
  3016=>"001011010",
  3017=>"011010100",
  3018=>"110001110",
  3019=>"011011011",
  3020=>"100110010",
  3021=>"110110010",
  3022=>"110001101",
  3023=>"001001100",
  3024=>"111010110",
  3025=>"000000000",
  3026=>"000011101",
  3027=>"110110110",
  3028=>"010110101",
  3029=>"101010100",
  3030=>"000011101",
  3031=>"001100110",
  3032=>"010001001",
  3033=>"011000011",
  3034=>"011000000",
  3035=>"000010011",
  3036=>"010101100",
  3037=>"111000001",
  3038=>"110011000",
  3039=>"000010010",
  3040=>"010010100",
  3041=>"110100110",
  3042=>"010100111",
  3043=>"001001100",
  3044=>"001100011",
  3045=>"010101010",
  3046=>"001011110",
  3047=>"110101000",
  3048=>"001001011",
  3049=>"000001001",
  3050=>"101000001",
  3051=>"000011100",
  3052=>"000010000",
  3053=>"010011110",
  3054=>"010001001",
  3055=>"001010010",
  3056=>"001111111",
  3057=>"100111010",
  3058=>"110100001",
  3059=>"011101000",
  3060=>"011000011",
  3061=>"000000110",
  3062=>"011011101",
  3063=>"000101111",
  3064=>"001000110",
  3065=>"111011010",
  3066=>"000000001",
  3067=>"011000001",
  3068=>"010011000",
  3069=>"101010011",
  3070=>"100100100",
  3071=>"001101010",
  3072=>"111011010",
  3073=>"101010110",
  3074=>"011111010",
  3075=>"011001110",
  3076=>"010000010",
  3077=>"101100010",
  3078=>"100000111",
  3079=>"101010001",
  3080=>"010010010",
  3081=>"110010111",
  3082=>"001000101",
  3083=>"001111010",
  3084=>"010101110",
  3085=>"011100110",
  3086=>"001101100",
  3087=>"001101100",
  3088=>"100100101",
  3089=>"110010110",
  3090=>"110100111",
  3091=>"010000101",
  3092=>"101101101",
  3093=>"110000110",
  3094=>"000110111",
  3095=>"000000000",
  3096=>"111001100",
  3097=>"101000000",
  3098=>"101001110",
  3099=>"110011101",
  3100=>"110111111",
  3101=>"001001001",
  3102=>"111111110",
  3103=>"110110001",
  3104=>"010000000",
  3105=>"010100000",
  3106=>"001111100",
  3107=>"000010111",
  3108=>"001000101",
  3109=>"100100011",
  3110=>"110110010",
  3111=>"111110111",
  3112=>"110101101",
  3113=>"001001001",
  3114=>"100010101",
  3115=>"111111011",
  3116=>"101100101",
  3117=>"110100000",
  3118=>"001001011",
  3119=>"101000010",
  3120=>"111110011",
  3121=>"100111111",
  3122=>"001011101",
  3123=>"001100000",
  3124=>"001011010",
  3125=>"110000000",
  3126=>"110111000",
  3127=>"010001000",
  3128=>"010111101",
  3129=>"001101111",
  3130=>"100100000",
  3131=>"111111000",
  3132=>"100111100",
  3133=>"101010100",
  3134=>"110001101",
  3135=>"000001110",
  3136=>"110110000",
  3137=>"001010011",
  3138=>"011011010",
  3139=>"101000000",
  3140=>"100111101",
  3141=>"111111000",
  3142=>"011010011",
  3143=>"100110000",
  3144=>"000101000",
  3145=>"110011110",
  3146=>"010100000",
  3147=>"110111011",
  3148=>"100001001",
  3149=>"001111101",
  3150=>"000011111",
  3151=>"100100100",
  3152=>"101011100",
  3153=>"000001011",
  3154=>"011001010",
  3155=>"010101010",
  3156=>"001001111",
  3157=>"101100000",
  3158=>"010110010",
  3159=>"001000011",
  3160=>"011011101",
  3161=>"100010101",
  3162=>"100001001",
  3163=>"000000111",
  3164=>"000100011",
  3165=>"011101100",
  3166=>"011011110",
  3167=>"101101110",
  3168=>"010000100",
  3169=>"011011100",
  3170=>"010110000",
  3171=>"110010010",
  3172=>"000001111",
  3173=>"111001000",
  3174=>"010100110",
  3175=>"010000010",
  3176=>"000001110",
  3177=>"001000000",
  3178=>"110000000",
  3179=>"110101100",
  3180=>"111000101",
  3181=>"001001100",
  3182=>"011011101",
  3183=>"001101110",
  3184=>"111110000",
  3185=>"001001010",
  3186=>"000110100",
  3187=>"001010111",
  3188=>"100001010",
  3189=>"010011110",
  3190=>"100001111",
  3191=>"011101010",
  3192=>"100101110",
  3193=>"000000111",
  3194=>"000101000",
  3195=>"000000000",
  3196=>"010101011",
  3197=>"000011000",
  3198=>"010010010",
  3199=>"110011101",
  3200=>"100110011",
  3201=>"001000111",
  3202=>"101010011",
  3203=>"101000001",
  3204=>"101000011",
  3205=>"000101000",
  3206=>"110010010",
  3207=>"100001110",
  3208=>"111110111",
  3209=>"101111100",
  3210=>"100010011",
  3211=>"110011101",
  3212=>"011001011",
  3213=>"100101111",
  3214=>"010010011",
  3215=>"111111011",
  3216=>"011010000",
  3217=>"010000000",
  3218=>"101101111",
  3219=>"100000011",
  3220=>"000111111",
  3221=>"000000000",
  3222=>"100000010",
  3223=>"000000010",
  3224=>"010010001",
  3225=>"100000011",
  3226=>"101101101",
  3227=>"011001011",
  3228=>"011101001",
  3229=>"011101000",
  3230=>"101111100",
  3231=>"011110111",
  3232=>"011001010",
  3233=>"100011111",
  3234=>"001000001",
  3235=>"111001011",
  3236=>"110110010",
  3237=>"001110111",
  3238=>"000110100",
  3239=>"101000110",
  3240=>"001000011",
  3241=>"001001001",
  3242=>"100101111",
  3243=>"111111100",
  3244=>"000100101",
  3245=>"001110010",
  3246=>"101110001",
  3247=>"001000000",
  3248=>"101010101",
  3249=>"100011001",
  3250=>"011010011",
  3251=>"110000011",
  3252=>"011100000",
  3253=>"011100101",
  3254=>"010001001",
  3255=>"000101000",
  3256=>"111010110",
  3257=>"001010111",
  3258=>"111000001",
  3259=>"000001000",
  3260=>"010100111",
  3261=>"001100101",
  3262=>"111110100",
  3263=>"000110111",
  3264=>"010111000",
  3265=>"010110000",
  3266=>"110001101",
  3267=>"010110011",
  3268=>"001001100",
  3269=>"111000011",
  3270=>"011111011",
  3271=>"010011010",
  3272=>"110010011",
  3273=>"000001111",
  3274=>"101010111",
  3275=>"011010100",
  3276=>"101111111",
  3277=>"111100001",
  3278=>"000111101",
  3279=>"001001111",
  3280=>"111110001",
  3281=>"101001100",
  3282=>"001011110",
  3283=>"101100011",
  3284=>"110100010",
  3285=>"110000101",
  3286=>"100100110",
  3287=>"011010101",
  3288=>"101000100",
  3289=>"111111010",
  3290=>"011000100",
  3291=>"001010100",
  3292=>"110010011",
  3293=>"011001101",
  3294=>"001001000",
  3295=>"011001001",
  3296=>"100111110",
  3297=>"100011100",
  3298=>"001100010",
  3299=>"000111110",
  3300=>"100111010",
  3301=>"100010100",
  3302=>"100010101",
  3303=>"001111110",
  3304=>"000001101",
  3305=>"101001000",
  3306=>"111001111",
  3307=>"111001011",
  3308=>"010100110",
  3309=>"010100110",
  3310=>"111001101",
  3311=>"111010010",
  3312=>"101111000",
  3313=>"101111011",
  3314=>"010001111",
  3315=>"010111010",
  3316=>"001011101",
  3317=>"010000001",
  3318=>"101000101",
  3319=>"001000000",
  3320=>"100110110",
  3321=>"110110001",
  3322=>"010010000",
  3323=>"101001101",
  3324=>"000010101",
  3325=>"010111001",
  3326=>"001111001",
  3327=>"010100000",
  3328=>"001011010",
  3329=>"010101000",
  3330=>"000010110",
  3331=>"011000011",
  3332=>"110100111",
  3333=>"000001011",
  3334=>"110010110",
  3335=>"100110010",
  3336=>"000011100",
  3337=>"000001000",
  3338=>"110010101",
  3339=>"001011100",
  3340=>"110101101",
  3341=>"101101111",
  3342=>"010011101",
  3343=>"011100001",
  3344=>"000110110",
  3345=>"100111110",
  3346=>"100011110",
  3347=>"011010011",
  3348=>"011111101",
  3349=>"010111001",
  3350=>"000101001",
  3351=>"010001110",
  3352=>"010000001",
  3353=>"101011000",
  3354=>"111010111",
  3355=>"000000100",
  3356=>"101000011",
  3357=>"010011001",
  3358=>"110011100",
  3359=>"010000011",
  3360=>"100110000",
  3361=>"111110110",
  3362=>"110110001",
  3363=>"111111111",
  3364=>"111001111",
  3365=>"111110110",
  3366=>"111111110",
  3367=>"011110011",
  3368=>"100100101",
  3369=>"111100110",
  3370=>"111010000",
  3371=>"011010010",
  3372=>"101000111",
  3373=>"100100111",
  3374=>"011100000",
  3375=>"010110100",
  3376=>"100001110",
  3377=>"111101011",
  3378=>"011001010",
  3379=>"100001110",
  3380=>"100100010",
  3381=>"010001010",
  3382=>"101000100",
  3383=>"101100011",
  3384=>"010000110",
  3385=>"011010011",
  3386=>"110100100",
  3387=>"001100110",
  3388=>"101010010",
  3389=>"101111100",
  3390=>"100100101",
  3391=>"101111110",
  3392=>"110100101",
  3393=>"100101101",
  3394=>"101001111",
  3395=>"000110111",
  3396=>"111101010",
  3397=>"110001001",
  3398=>"111001111",
  3399=>"111010100",
  3400=>"101100011",
  3401=>"111011001",
  3402=>"101100000",
  3403=>"000000001",
  3404=>"001110001",
  3405=>"001000100",
  3406=>"000011100",
  3407=>"000000110",
  3408=>"101100101",
  3409=>"101010110",
  3410=>"101101111",
  3411=>"010111000",
  3412=>"101011010",
  3413=>"011000011",
  3414=>"110000001",
  3415=>"110010000",
  3416=>"010001000",
  3417=>"000011000",
  3418=>"001000000",
  3419=>"111000001",
  3420=>"110101010",
  3421=>"110011101",
  3422=>"011000111",
  3423=>"000101000",
  3424=>"111100001",
  3425=>"110111100",
  3426=>"101001100",
  3427=>"001110001",
  3428=>"011111001",
  3429=>"011111000",
  3430=>"010100011",
  3431=>"110001101",
  3432=>"101010000",
  3433=>"000000010",
  3434=>"101011110",
  3435=>"010001001",
  3436=>"101100001",
  3437=>"011011000",
  3438=>"111000010",
  3439=>"011110100",
  3440=>"001011100",
  3441=>"010110111",
  3442=>"010100010",
  3443=>"101110101",
  3444=>"110111000",
  3445=>"000100100",
  3446=>"011000110",
  3447=>"110101010",
  3448=>"011100101",
  3449=>"101100110",
  3450=>"110101001",
  3451=>"101000101",
  3452=>"110100001",
  3453=>"011011000",
  3454=>"000001100",
  3455=>"011110001",
  3456=>"001001010",
  3457=>"100111111",
  3458=>"011101001",
  3459=>"000111100",
  3460=>"110100000",
  3461=>"010001000",
  3462=>"000101001",
  3463=>"111101101",
  3464=>"000001011",
  3465=>"111110111",
  3466=>"110111010",
  3467=>"110100011",
  3468=>"100110100",
  3469=>"000110001",
  3470=>"101001010",
  3471=>"101000100",
  3472=>"010101101",
  3473=>"011010110",
  3474=>"101100111",
  3475=>"110001110",
  3476=>"111010101",
  3477=>"010000001",
  3478=>"010100100",
  3479=>"101010110",
  3480=>"110010101",
  3481=>"001010111",
  3482=>"110010110",
  3483=>"101001000",
  3484=>"001110110",
  3485=>"011001100",
  3486=>"001100000",
  3487=>"101101111",
  3488=>"100100100",
  3489=>"100110110",
  3490=>"100011000",
  3491=>"011001100",
  3492=>"101011010",
  3493=>"110111010",
  3494=>"100100111",
  3495=>"111100110",
  3496=>"100111000",
  3497=>"101100000",
  3498=>"000100101",
  3499=>"110000000",
  3500=>"101000110",
  3501=>"100100100",
  3502=>"110110010",
  3503=>"110011110",
  3504=>"000100111",
  3505=>"100000111",
  3506=>"000010101",
  3507=>"000101010",
  3508=>"011100010",
  3509=>"111011100",
  3510=>"100101111",
  3511=>"000001000",
  3512=>"010101010",
  3513=>"111000110",
  3514=>"010100011",
  3515=>"011101111",
  3516=>"001110000",
  3517=>"011000010",
  3518=>"100001010",
  3519=>"110110100",
  3520=>"010011101",
  3521=>"001010101",
  3522=>"100101110",
  3523=>"000001011",
  3524=>"010010000",
  3525=>"011100000",
  3526=>"000001111",
  3527=>"010000111",
  3528=>"001011010",
  3529=>"001101110",
  3530=>"011001111",
  3531=>"110011001",
  3532=>"011001010",
  3533=>"000011010",
  3534=>"001100000",
  3535=>"011010101",
  3536=>"111111110",
  3537=>"100000000",
  3538=>"011011011",
  3539=>"111100011",
  3540=>"111011011",
  3541=>"110101111",
  3542=>"010101001",
  3543=>"011101000",
  3544=>"011000001",
  3545=>"000110101",
  3546=>"100111110",
  3547=>"101001000",
  3548=>"110011100",
  3549=>"001011111",
  3550=>"100010111",
  3551=>"000000010",
  3552=>"000111001",
  3553=>"010111010",
  3554=>"110011101",
  3555=>"101110001",
  3556=>"100000101",
  3557=>"001110001",
  3558=>"110100001",
  3559=>"001010001",
  3560=>"111000000",
  3561=>"011000101",
  3562=>"101111000",
  3563=>"011111111",
  3564=>"111000101",
  3565=>"111010100",
  3566=>"110001110",
  3567=>"110011011",
  3568=>"100011001",
  3569=>"111100111",
  3570=>"110100101",
  3571=>"110010100",
  3572=>"100010011",
  3573=>"111101001",
  3574=>"000100011",
  3575=>"010110001",
  3576=>"000101000",
  3577=>"011001001",
  3578=>"101111101",
  3579=>"001110111",
  3580=>"000100000",
  3581=>"010011001",
  3582=>"100101101",
  3583=>"110010001",
  3584=>"101000111",
  3585=>"110110101",
  3586=>"011101110",
  3587=>"000100011",
  3588=>"100000101",
  3589=>"010101110",
  3590=>"010010101",
  3591=>"111100010",
  3592=>"110010011",
  3593=>"011001011",
  3594=>"110001000",
  3595=>"101111010",
  3596=>"011100000",
  3597=>"010110101",
  3598=>"101110000",
  3599=>"000001111",
  3600=>"000110100",
  3601=>"000011001",
  3602=>"000101101",
  3603=>"111110011",
  3604=>"000010100",
  3605=>"100001111",
  3606=>"111111110",
  3607=>"111100110",
  3608=>"111101111",
  3609=>"101000000",
  3610=>"010110001",
  3611=>"011011111",
  3612=>"000001100",
  3613=>"010100000",
  3614=>"110111000",
  3615=>"101111001",
  3616=>"010000100",
  3617=>"011110101",
  3618=>"001001101",
  3619=>"111111001",
  3620=>"001111000",
  3621=>"011000001",
  3622=>"110110000",
  3623=>"100110110",
  3624=>"010100001",
  3625=>"010010111",
  3626=>"110110000",
  3627=>"100100011",
  3628=>"100000111",
  3629=>"110000101",
  3630=>"010100100",
  3631=>"000101110",
  3632=>"101110001",
  3633=>"010011000",
  3634=>"000000101",
  3635=>"010010000",
  3636=>"110101100",
  3637=>"010100101",
  3638=>"001111001",
  3639=>"000100010",
  3640=>"010100110",
  3641=>"111110111",
  3642=>"111010110",
  3643=>"011000000",
  3644=>"010111101",
  3645=>"100000101",
  3646=>"011111101",
  3647=>"000111111",
  3648=>"100000100",
  3649=>"101111100",
  3650=>"000101111",
  3651=>"100110101",
  3652=>"011010000",
  3653=>"010011111",
  3654=>"000000100",
  3655=>"110010111",
  3656=>"010010101",
  3657=>"010100001",
  3658=>"101110110",
  3659=>"111101111",
  3660=>"001000101",
  3661=>"100000000",
  3662=>"110010000",
  3663=>"101100000",
  3664=>"101000111",
  3665=>"111010011",
  3666=>"001010010",
  3667=>"110110100",
  3668=>"011100011",
  3669=>"011001011",
  3670=>"000000000",
  3671=>"000110001",
  3672=>"100110000",
  3673=>"100100001",
  3674=>"001000011",
  3675=>"111010111",
  3676=>"101000010",
  3677=>"010101101",
  3678=>"111011110",
  3679=>"100110110",
  3680=>"100001111",
  3681=>"010000001",
  3682=>"100111100",
  3683=>"010011011",
  3684=>"011010000",
  3685=>"100000000",
  3686=>"100000111",
  3687=>"000000110",
  3688=>"010101101",
  3689=>"101001110",
  3690=>"111100001",
  3691=>"110000100",
  3692=>"011011010",
  3693=>"000001011",
  3694=>"000110010",
  3695=>"010000010",
  3696=>"111100010",
  3697=>"111101101",
  3698=>"101000011",
  3699=>"100100000",
  3700=>"000100111",
  3701=>"110000001",
  3702=>"111010010",
  3703=>"000000010",
  3704=>"110011000",
  3705=>"101111010",
  3706=>"110110000",
  3707=>"010100011",
  3708=>"101000010",
  3709=>"110000000",
  3710=>"101110111",
  3711=>"111101101",
  3712=>"111100110",
  3713=>"111101101",
  3714=>"101100001",
  3715=>"000011101",
  3716=>"101110010",
  3717=>"011111000",
  3718=>"101001011",
  3719=>"111111111",
  3720=>"111001010",
  3721=>"011110011",
  3722=>"010011011",
  3723=>"000000000",
  3724=>"110011100",
  3725=>"110001101",
  3726=>"111001111",
  3727=>"110011111",
  3728=>"001101011",
  3729=>"000000110",
  3730=>"100101011",
  3731=>"100101101",
  3732=>"001010010",
  3733=>"110001001",
  3734=>"011101101",
  3735=>"000010000",
  3736=>"111111010",
  3737=>"111110000",
  3738=>"101100101",
  3739=>"011001001",
  3740=>"110100111",
  3741=>"000000111",
  3742=>"000010111",
  3743=>"110100000",
  3744=>"001010111",
  3745=>"001111001",
  3746=>"010010011",
  3747=>"110001010",
  3748=>"100100100",
  3749=>"000011100",
  3750=>"101111101",
  3751=>"000000110",
  3752=>"011100010",
  3753=>"000001011",
  3754=>"111000110",
  3755=>"011110101",
  3756=>"111010001",
  3757=>"001110000",
  3758=>"010000010",
  3759=>"100000011",
  3760=>"001111001",
  3761=>"110000010",
  3762=>"001100101",
  3763=>"100111010",
  3764=>"001010010",
  3765=>"010001010",
  3766=>"100001110",
  3767=>"101100001",
  3768=>"111010101",
  3769=>"110010000",
  3770=>"100111011",
  3771=>"000001101",
  3772=>"100010011",
  3773=>"000000101",
  3774=>"011111111",
  3775=>"110011100",
  3776=>"100101111",
  3777=>"100101001",
  3778=>"001100111",
  3779=>"101011000",
  3780=>"000111001",
  3781=>"101110111",
  3782=>"110010010",
  3783=>"000011100",
  3784=>"111001000",
  3785=>"011011000",
  3786=>"111100011",
  3787=>"010001110",
  3788=>"010000001",
  3789=>"010100100",
  3790=>"010011010",
  3791=>"001000111",
  3792=>"100100000",
  3793=>"001100100",
  3794=>"111011000",
  3795=>"001010110",
  3796=>"110011011",
  3797=>"000110100",
  3798=>"100110110",
  3799=>"100100111",
  3800=>"000011110",
  3801=>"110101011",
  3802=>"110001100",
  3803=>"000010101",
  3804=>"010101000",
  3805=>"100111111",
  3806=>"100111110",
  3807=>"011110111",
  3808=>"111001011",
  3809=>"011101000",
  3810=>"110011111",
  3811=>"110001000",
  3812=>"011100000",
  3813=>"011101010",
  3814=>"000111001",
  3815=>"010001100",
  3816=>"010001110",
  3817=>"011101101",
  3818=>"000011010",
  3819=>"110011011",
  3820=>"111011111",
  3821=>"101100111",
  3822=>"111100110",
  3823=>"110111000",
  3824=>"000000011",
  3825=>"010011100",
  3826=>"100100011",
  3827=>"100000111",
  3828=>"110100101",
  3829=>"111010010",
  3830=>"010010000",
  3831=>"011110101",
  3832=>"111101111",
  3833=>"110010011",
  3834=>"111000101",
  3835=>"011111100",
  3836=>"011100000",
  3837=>"011111110",
  3838=>"110110111",
  3839=>"000111100",
  3840=>"100010000",
  3841=>"011010110",
  3842=>"000011010",
  3843=>"011010111",
  3844=>"011011001",
  3845=>"100001000",
  3846=>"001001010",
  3847=>"011110100",
  3848=>"101001101",
  3849=>"010111101",
  3850=>"000110100",
  3851=>"000001101",
  3852=>"101111111",
  3853=>"110001110",
  3854=>"111011001",
  3855=>"110101100",
  3856=>"011111101",
  3857=>"010010010",
  3858=>"100100011",
  3859=>"101101111",
  3860=>"011101111",
  3861=>"110001101",
  3862=>"100100101",
  3863=>"010110110",
  3864=>"000010011",
  3865=>"001000001",
  3866=>"111001101",
  3867=>"111110101",
  3868=>"110001000",
  3869=>"010101110",
  3870=>"000100100",
  3871=>"010100011",
  3872=>"011001011",
  3873=>"000010010",
  3874=>"011000101",
  3875=>"100000010",
  3876=>"110101100",
  3877=>"110110100",
  3878=>"111011110",
  3879=>"001111100",
  3880=>"110000111",
  3881=>"101000000",
  3882=>"110110100",
  3883=>"101110001",
  3884=>"010001011",
  3885=>"110011010",
  3886=>"010111010",
  3887=>"111000110",
  3888=>"001000000",
  3889=>"100001101",
  3890=>"000010101",
  3891=>"111111101",
  3892=>"101000010",
  3893=>"111101101",
  3894=>"000110010",
  3895=>"100101101",
  3896=>"000101011",
  3897=>"110111000",
  3898=>"010110011",
  3899=>"101001100",
  3900=>"101101010",
  3901=>"100010111",
  3902=>"011111000",
  3903=>"001101110",
  3904=>"111011101",
  3905=>"110100011",
  3906=>"010111000",
  3907=>"010010110",
  3908=>"100100010",
  3909=>"110011100",
  3910=>"010011110",
  3911=>"110111000",
  3912=>"001010110",
  3913=>"001000110",
  3914=>"000111000",
  3915=>"011110000",
  3916=>"101101100",
  3917=>"011000000",
  3918=>"011100010",
  3919=>"110000101",
  3920=>"110001010",
  3921=>"101111011",
  3922=>"000000100",
  3923=>"101011011",
  3924=>"110010111",
  3925=>"000001111",
  3926=>"011010011",
  3927=>"111011000",
  3928=>"100011010",
  3929=>"011000011",
  3930=>"011011101",
  3931=>"111001110",
  3932=>"000000011",
  3933=>"011011110",
  3934=>"111000101",
  3935=>"010100001",
  3936=>"000011011",
  3937=>"100011010",
  3938=>"011001011",
  3939=>"111000001",
  3940=>"010111101",
  3941=>"101010101",
  3942=>"000110101",
  3943=>"101001101",
  3944=>"110010001",
  3945=>"011100010",
  3946=>"010100001",
  3947=>"000110001",
  3948=>"001001101",
  3949=>"011010001",
  3950=>"110100110",
  3951=>"111101100",
  3952=>"000001000",
  3953=>"001111011",
  3954=>"101000011",
  3955=>"000010101",
  3956=>"000110010",
  3957=>"111000111",
  3958=>"000101001",
  3959=>"011011100",
  3960=>"010100000",
  3961=>"110000101",
  3962=>"101000010",
  3963=>"001111100",
  3964=>"100000110",
  3965=>"100010101",
  3966=>"100100111",
  3967=>"110110101",
  3968=>"110111011",
  3969=>"011000110",
  3970=>"100101001",
  3971=>"011110010",
  3972=>"111101101",
  3973=>"101001011",
  3974=>"001101111",
  3975=>"110110110",
  3976=>"101111011",
  3977=>"111101100",
  3978=>"110010111",
  3979=>"100011100",
  3980=>"110111111",
  3981=>"001110101",
  3982=>"100101001",
  3983=>"110001101",
  3984=>"100100110",
  3985=>"110011110",
  3986=>"011010001",
  3987=>"111110000",
  3988=>"110001001",
  3989=>"110100100",
  3990=>"100011110",
  3991=>"111011011",
  3992=>"110111011",
  3993=>"010111110",
  3994=>"110000001",
  3995=>"010101001",
  3996=>"100110001",
  3997=>"100001010",
  3998=>"011011111",
  3999=>"000001011",
  4000=>"001010001",
  4001=>"100110111",
  4002=>"001011101",
  4003=>"001011101",
  4004=>"010110110",
  4005=>"100111100",
  4006=>"010001011",
  4007=>"001101011",
  4008=>"010101001",
  4009=>"101011101",
  4010=>"000001100",
  4011=>"100111110",
  4012=>"110001011",
  4013=>"101100011",
  4014=>"111000011",
  4015=>"001001101",
  4016=>"000001001",
  4017=>"001001100",
  4018=>"101101011",
  4019=>"101110001",
  4020=>"111101000",
  4021=>"010011000",
  4022=>"111000000",
  4023=>"010011111",
  4024=>"101111011",
  4025=>"101110101",
  4026=>"100110011",
  4027=>"010000001",
  4028=>"111011101",
  4029=>"011011011",
  4030=>"100010111",
  4031=>"001000101",
  4032=>"001111111",
  4033=>"011001010",
  4034=>"100111111",
  4035=>"000100101",
  4036=>"100110011",
  4037=>"000001101",
  4038=>"101011111",
  4039=>"100100011",
  4040=>"010000100",
  4041=>"000011010",
  4042=>"100111111",
  4043=>"110000100",
  4044=>"001001110",
  4045=>"000110100",
  4046=>"101011011",
  4047=>"110010111",
  4048=>"110001001",
  4049=>"100010011",
  4050=>"101010010",
  4051=>"110101000",
  4052=>"110000001",
  4053=>"100111110",
  4054=>"001100101",
  4055=>"111101101",
  4056=>"000000101",
  4057=>"001101110",
  4058=>"011100011",
  4059=>"111100111",
  4060=>"001011010",
  4061=>"110010100",
  4062=>"000000001",
  4063=>"101010010",
  4064=>"010010110",
  4065=>"010111100",
  4066=>"000101100",
  4067=>"001010011",
  4068=>"110000110",
  4069=>"111110010",
  4070=>"011010110",
  4071=>"001000000",
  4072=>"000011111",
  4073=>"000000110",
  4074=>"011110000",
  4075=>"101011001",
  4076=>"101001001",
  4077=>"000001001",
  4078=>"000110111",
  4079=>"001001101",
  4080=>"110000001",
  4081=>"101110101",
  4082=>"001010010",
  4083=>"110000011",
  4084=>"111010001",
  4085=>"000000110",
  4086=>"100011101",
  4087=>"010100101",
  4088=>"110110111",
  4089=>"011111111",
  4090=>"001011100",
  4091=>"110010011",
  4092=>"100100000",
  4093=>"110011000",
  4094=>"010010111",
  4095=>"100001010",
  4096=>"100111110",
  4097=>"011010010",
  4098=>"011011111",
  4099=>"011011011",
  4100=>"000101100",
  4101=>"010001000",
  4102=>"001000100",
  4103=>"101000000",
  4104=>"011110111",
  4105=>"010110010",
  4106=>"110100111",
  4107=>"101001011",
  4108=>"100110100",
  4109=>"001110111",
  4110=>"000101101",
  4111=>"111100001",
  4112=>"101110000",
  4113=>"001000110",
  4114=>"011010010",
  4115=>"100011001",
  4116=>"111100100",
  4117=>"100011011",
  4118=>"110101010",
  4119=>"001110100",
  4120=>"001001110",
  4121=>"111010001",
  4122=>"110101110",
  4123=>"110111100",
  4124=>"001011110",
  4125=>"001011111",
  4126=>"000010110",
  4127=>"100110110",
  4128=>"011001001",
  4129=>"000111110",
  4130=>"110111110",
  4131=>"100110100",
  4132=>"101110111",
  4133=>"100110010",
  4134=>"111010001",
  4135=>"001110101",
  4136=>"100110010",
  4137=>"111101000",
  4138=>"010001011",
  4139=>"001101011",
  4140=>"010101110",
  4141=>"000011010",
  4142=>"111000011",
  4143=>"110110100",
  4144=>"110011000",
  4145=>"001001001",
  4146=>"001001110",
  4147=>"111010010",
  4148=>"100101101",
  4149=>"110100101",
  4150=>"111111010",
  4151=>"010110111",
  4152=>"110001110",
  4153=>"011100111",
  4154=>"000000000",
  4155=>"101010000",
  4156=>"100100100",
  4157=>"111111000",
  4158=>"110101100",
  4159=>"101001101",
  4160=>"111100111",
  4161=>"000101011",
  4162=>"101010110",
  4163=>"000000001",
  4164=>"010000100",
  4165=>"010011011",
  4166=>"000011010",
  4167=>"100110100",
  4168=>"011101110",
  4169=>"001110001",
  4170=>"011010101",
  4171=>"101001111",
  4172=>"110110001",
  4173=>"110101010",
  4174=>"000110101",
  4175=>"011000011",
  4176=>"101110101",
  4177=>"001100100",
  4178=>"110100001",
  4179=>"011011101",
  4180=>"011011000",
  4181=>"110110000",
  4182=>"001111000",
  4183=>"100000000",
  4184=>"110000100",
  4185=>"101010101",
  4186=>"110000110",
  4187=>"110100010",
  4188=>"101001100",
  4189=>"100100101",
  4190=>"100000101",
  4191=>"111100010",
  4192=>"101000110",
  4193=>"110001100",
  4194=>"011110100",
  4195=>"111000000",
  4196=>"000011110",
  4197=>"111100010",
  4198=>"100101000",
  4199=>"111011000",
  4200=>"010001100",
  4201=>"011000101",
  4202=>"010101011",
  4203=>"001101110",
  4204=>"100101000",
  4205=>"100010111",
  4206=>"001101111",
  4207=>"100100011",
  4208=>"000010100",
  4209=>"001101000",
  4210=>"101110100",
  4211=>"001001011",
  4212=>"000111011",
  4213=>"010010101",
  4214=>"001000011",
  4215=>"010101011",
  4216=>"000011011",
  4217=>"011111100",
  4218=>"100100110",
  4219=>"100011010",
  4220=>"101000000",
  4221=>"100010110",
  4222=>"000111110",
  4223=>"010010000",
  4224=>"001000100",
  4225=>"101000010",
  4226=>"100010001",
  4227=>"000110101",
  4228=>"111011100",
  4229=>"001010111",
  4230=>"110100111",
  4231=>"110011010",
  4232=>"011011101",
  4233=>"101111111",
  4234=>"111101000",
  4235=>"101000010",
  4236=>"011001111",
  4237=>"110101101",
  4238=>"000000111",
  4239=>"001011010",
  4240=>"110001010",
  4241=>"001010011",
  4242=>"110100111",
  4243=>"010100110",
  4244=>"000101111",
  4245=>"011001111",
  4246=>"001000100",
  4247=>"011000111",
  4248=>"101011110",
  4249=>"010011111",
  4250=>"100111010",
  4251=>"000010010",
  4252=>"110100100",
  4253=>"111110111",
  4254=>"001110100",
  4255=>"001011011",
  4256=>"110000100",
  4257=>"101110101",
  4258=>"101100110",
  4259=>"011010110",
  4260=>"111010011",
  4261=>"000001011",
  4262=>"011001100",
  4263=>"000100101",
  4264=>"100101101",
  4265=>"001010111",
  4266=>"110110010",
  4267=>"000111000",
  4268=>"011111101",
  4269=>"000110100",
  4270=>"011111010",
  4271=>"110100010",
  4272=>"001101000",
  4273=>"001100011",
  4274=>"110010000",
  4275=>"100011100",
  4276=>"000010100",
  4277=>"100100111",
  4278=>"010011010",
  4279=>"001000010",
  4280=>"111110110",
  4281=>"100101110",
  4282=>"100101100",
  4283=>"111101111",
  4284=>"001100110",
  4285=>"110100100",
  4286=>"010101110",
  4287=>"001111101",
  4288=>"101101111",
  4289=>"100111000",
  4290=>"000010111",
  4291=>"000001011",
  4292=>"010000011",
  4293=>"001000100",
  4294=>"010000101",
  4295=>"101000010",
  4296=>"000010010",
  4297=>"100010010",
  4298=>"100011010",
  4299=>"000011010",
  4300=>"101110111",
  4301=>"110101111",
  4302=>"000101110",
  4303=>"000000011",
  4304=>"011000101",
  4305=>"011101011",
  4306=>"110010010",
  4307=>"010011110",
  4308=>"011111001",
  4309=>"111111001",
  4310=>"110001001",
  4311=>"101000101",
  4312=>"010010101",
  4313=>"110011010",
  4314=>"010101111",
  4315=>"101100001",
  4316=>"000111111",
  4317=>"110100010",
  4318=>"100100111",
  4319=>"010010011",
  4320=>"110011111",
  4321=>"000101111",
  4322=>"011110100",
  4323=>"001010110",
  4324=>"011111011",
  4325=>"001011100",
  4326=>"100011111",
  4327=>"101110101",
  4328=>"110111010",
  4329=>"011000101",
  4330=>"100111010",
  4331=>"100011000",
  4332=>"100001100",
  4333=>"001101011",
  4334=>"100000110",
  4335=>"111011101",
  4336=>"001101011",
  4337=>"001101100",
  4338=>"010100000",
  4339=>"011101001",
  4340=>"101111001",
  4341=>"111101111",
  4342=>"011010011",
  4343=>"100100010",
  4344=>"101010011",
  4345=>"110111011",
  4346=>"101011101",
  4347=>"100010100",
  4348=>"010001010",
  4349=>"010000110",
  4350=>"010100110",
  4351=>"111110111",
  4352=>"101101100",
  4353=>"001000001",
  4354=>"110011001",
  4355=>"111101000",
  4356=>"001101001",
  4357=>"110011110",
  4358=>"011010101",
  4359=>"111111101",
  4360=>"010101010",
  4361=>"110001101",
  4362=>"101110110",
  4363=>"001000001",
  4364=>"001000010",
  4365=>"001101110",
  4366=>"100000111",
  4367=>"111000000",
  4368=>"010100001",
  4369=>"011011000",
  4370=>"101001011",
  4371=>"010100101",
  4372=>"011011000",
  4373=>"001101000",
  4374=>"011110011",
  4375=>"010101101",
  4376=>"010101010",
  4377=>"111100100",
  4378=>"000011010",
  4379=>"101110110",
  4380=>"111111110",
  4381=>"110110101",
  4382=>"011110011",
  4383=>"000100100",
  4384=>"110010100",
  4385=>"101111010",
  4386=>"111010101",
  4387=>"101010000",
  4388=>"110011101",
  4389=>"110101111",
  4390=>"000100000",
  4391=>"100000001",
  4392=>"001011010",
  4393=>"111011011",
  4394=>"000011001",
  4395=>"011000001",
  4396=>"111100000",
  4397=>"110110100",
  4398=>"001110110",
  4399=>"110111110",
  4400=>"010110010",
  4401=>"011110011",
  4402=>"011001101",
  4403=>"100101001",
  4404=>"001010000",
  4405=>"100111110",
  4406=>"001111010",
  4407=>"011101110",
  4408=>"100111100",
  4409=>"110101101",
  4410=>"000100101",
  4411=>"110000100",
  4412=>"101011111",
  4413=>"010100111",
  4414=>"011100000",
  4415=>"001111010",
  4416=>"101101101",
  4417=>"110100011",
  4418=>"110100100",
  4419=>"000100011",
  4420=>"111111101",
  4421=>"001111011",
  4422=>"001110100",
  4423=>"110110001",
  4424=>"111110010",
  4425=>"110100100",
  4426=>"101001010",
  4427=>"101110011",
  4428=>"001000101",
  4429=>"011111011",
  4430=>"000110000",
  4431=>"000011101",
  4432=>"011110101",
  4433=>"100011101",
  4434=>"101011000",
  4435=>"110111010",
  4436=>"100000101",
  4437=>"101001100",
  4438=>"110110100",
  4439=>"110001111",
  4440=>"010000110",
  4441=>"111010110",
  4442=>"100100100",
  4443=>"110110101",
  4444=>"000001001",
  4445=>"110010001",
  4446=>"001111000",
  4447=>"110101010",
  4448=>"110010011",
  4449=>"100010010",
  4450=>"000110100",
  4451=>"000010101",
  4452=>"001101111",
  4453=>"001100111",
  4454=>"001101011",
  4455=>"011110000",
  4456=>"000100011",
  4457=>"111001100",
  4458=>"101000010",
  4459=>"001000111",
  4460=>"100100010",
  4461=>"110111011",
  4462=>"001001110",
  4463=>"000000111",
  4464=>"110011010",
  4465=>"100010111",
  4466=>"110111101",
  4467=>"000110111",
  4468=>"100001100",
  4469=>"100100100",
  4470=>"011001110",
  4471=>"010000111",
  4472=>"100111001",
  4473=>"010100110",
  4474=>"010111000",
  4475=>"110111100",
  4476=>"100010111",
  4477=>"000110010",
  4478=>"100010001",
  4479=>"011000010",
  4480=>"011100010",
  4481=>"010010110",
  4482=>"101111010",
  4483=>"010011001",
  4484=>"111001010",
  4485=>"100011000",
  4486=>"101011011",
  4487=>"011000011",
  4488=>"110010100",
  4489=>"001000010",
  4490=>"001100111",
  4491=>"010110110",
  4492=>"000001100",
  4493=>"011101110",
  4494=>"110101001",
  4495=>"011001100",
  4496=>"101110110",
  4497=>"100110110",
  4498=>"110000000",
  4499=>"101110011",
  4500=>"111000010",
  4501=>"111111001",
  4502=>"110101100",
  4503=>"000000100",
  4504=>"000101100",
  4505=>"101000100",
  4506=>"000111000",
  4507=>"000111101",
  4508=>"010100111",
  4509=>"111000010",
  4510=>"101101010",
  4511=>"101111111",
  4512=>"000100100",
  4513=>"111100000",
  4514=>"100000101",
  4515=>"101011000",
  4516=>"010000101",
  4517=>"001100110",
  4518=>"011100001",
  4519=>"011001010",
  4520=>"101000101",
  4521=>"000110100",
  4522=>"110111010",
  4523=>"001110001",
  4524=>"000101010",
  4525=>"011100101",
  4526=>"011000011",
  4527=>"010000010",
  4528=>"100111000",
  4529=>"011001111",
  4530=>"101111111",
  4531=>"010101100",
  4532=>"101101111",
  4533=>"111000001",
  4534=>"101001101",
  4535=>"101000111",
  4536=>"010001111",
  4537=>"110100010",
  4538=>"100101101",
  4539=>"101000000",
  4540=>"110101001",
  4541=>"111111000",
  4542=>"000000011",
  4543=>"000111101",
  4544=>"110101010",
  4545=>"101001010",
  4546=>"111101001",
  4547=>"101110000",
  4548=>"000000001",
  4549=>"011110110",
  4550=>"111001010",
  4551=>"111110110",
  4552=>"111101001",
  4553=>"100101010",
  4554=>"110001011",
  4555=>"000101001",
  4556=>"000111101",
  4557=>"110110110",
  4558=>"101001011",
  4559=>"001001110",
  4560=>"111000101",
  4561=>"111111110",
  4562=>"111100000",
  4563=>"010111010",
  4564=>"100100011",
  4565=>"001001001",
  4566=>"000101100",
  4567=>"100001011",
  4568=>"111100011",
  4569=>"011001011",
  4570=>"001100000",
  4571=>"011111110",
  4572=>"111001101",
  4573=>"110011100",
  4574=>"011111111",
  4575=>"101100101",
  4576=>"001010010",
  4577=>"010101011",
  4578=>"010100110",
  4579=>"011111110",
  4580=>"100110000",
  4581=>"000101110",
  4582=>"110011111",
  4583=>"111101001",
  4584=>"001101011",
  4585=>"011110110",
  4586=>"011111010",
  4587=>"110010011",
  4588=>"101111000",
  4589=>"011100000",
  4590=>"111110000",
  4591=>"111110001",
  4592=>"001011011",
  4593=>"001110011",
  4594=>"010001110",
  4595=>"100001100",
  4596=>"110110000",
  4597=>"011111110",
  4598=>"010101000",
  4599=>"111110110",
  4600=>"001110100",
  4601=>"010010110",
  4602=>"011010011",
  4603=>"001111000",
  4604=>"111110001",
  4605=>"010010100",
  4606=>"101110001",
  4607=>"010101011",
  4608=>"111111001",
  4609=>"001000001",
  4610=>"010100000",
  4611=>"100000010",
  4612=>"110001011",
  4613=>"000010110",
  4614=>"111010000",
  4615=>"000101101",
  4616=>"010000111",
  4617=>"010000011",
  4618=>"011100111",
  4619=>"010001100",
  4620=>"110011111",
  4621=>"011010100",
  4622=>"100100110",
  4623=>"110100010",
  4624=>"110101001",
  4625=>"001101001",
  4626=>"000010111",
  4627=>"111110000",
  4628=>"100100001",
  4629=>"001101001",
  4630=>"001001011",
  4631=>"101000110",
  4632=>"010100101",
  4633=>"100100000",
  4634=>"110110000",
  4635=>"110111010",
  4636=>"110100110",
  4637=>"010000101",
  4638=>"101011010",
  4639=>"010101001",
  4640=>"001000110",
  4641=>"110101111",
  4642=>"011110111",
  4643=>"001011100",
  4644=>"110111100",
  4645=>"110011010",
  4646=>"101010111",
  4647=>"111001000",
  4648=>"011101101",
  4649=>"110110111",
  4650=>"101111110",
  4651=>"000100111",
  4652=>"010100101",
  4653=>"011010100",
  4654=>"010111101",
  4655=>"011100101",
  4656=>"111000001",
  4657=>"010100110",
  4658=>"101101101",
  4659=>"000111100",
  4660=>"000010000",
  4661=>"010111000",
  4662=>"000100100",
  4663=>"111011001",
  4664=>"001111101",
  4665=>"110110010",
  4666=>"111010011",
  4667=>"101011000",
  4668=>"011110100",
  4669=>"111000100",
  4670=>"010100100",
  4671=>"110110100",
  4672=>"110111001",
  4673=>"101001011",
  4674=>"000111011",
  4675=>"101111001",
  4676=>"111111100",
  4677=>"001011001",
  4678=>"000100100",
  4679=>"110010010",
  4680=>"010010111",
  4681=>"110001000",
  4682=>"111000101",
  4683=>"000001000",
  4684=>"100110011",
  4685=>"010110110",
  4686=>"101011100",
  4687=>"000001011",
  4688=>"101001011",
  4689=>"101110001",
  4690=>"010100110",
  4691=>"000110111",
  4692=>"100010100",
  4693=>"100101000",
  4694=>"110100010",
  4695=>"101010011",
  4696=>"110111100",
  4697=>"100111110",
  4698=>"011000001",
  4699=>"111000100",
  4700=>"010101100",
  4701=>"101100100",
  4702=>"110100111",
  4703=>"001011100",
  4704=>"000000000",
  4705=>"011010101",
  4706=>"011111101",
  4707=>"010111111",
  4708=>"010111101",
  4709=>"010001111",
  4710=>"011001111",
  4711=>"011011011",
  4712=>"001000000",
  4713=>"001110111",
  4714=>"011111101",
  4715=>"010100001",
  4716=>"110000100",
  4717=>"111101010",
  4718=>"101011001",
  4719=>"110010001",
  4720=>"011011000",
  4721=>"101100101",
  4722=>"010000010",
  4723=>"101000111",
  4724=>"110101101",
  4725=>"000000000",
  4726=>"111100000",
  4727=>"100000011",
  4728=>"010010100",
  4729=>"101110110",
  4730=>"101010100",
  4731=>"111100110",
  4732=>"100010110",
  4733=>"011100111",
  4734=>"000101100",
  4735=>"111011001",
  4736=>"100101100",
  4737=>"111110101",
  4738=>"101101000",
  4739=>"000110101",
  4740=>"101111111",
  4741=>"111000100",
  4742=>"010011100",
  4743=>"010110110",
  4744=>"100011011",
  4745=>"100001100",
  4746=>"000000101",
  4747=>"000110101",
  4748=>"000011010",
  4749=>"100111010",
  4750=>"000110000",
  4751=>"100011111",
  4752=>"001001100",
  4753=>"000101100",
  4754=>"001011110",
  4755=>"101011111",
  4756=>"011110101",
  4757=>"001101011",
  4758=>"100110011",
  4759=>"101011010",
  4760=>"010100011",
  4761=>"110000010",
  4762=>"011001111",
  4763=>"010101101",
  4764=>"100000101",
  4765=>"001010000",
  4766=>"010100110",
  4767=>"100001010",
  4768=>"000101100",
  4769=>"101011111",
  4770=>"011101110",
  4771=>"111100000",
  4772=>"111100010",
  4773=>"101110101",
  4774=>"100110110",
  4775=>"110111100",
  4776=>"100100001",
  4777=>"110010110",
  4778=>"001100100",
  4779=>"000011010",
  4780=>"011000010",
  4781=>"011101010",
  4782=>"101101001",
  4783=>"001011011",
  4784=>"010001110",
  4785=>"100101111",
  4786=>"000110101",
  4787=>"000000101",
  4788=>"101011001",
  4789=>"011010011",
  4790=>"101000110",
  4791=>"001100001",
  4792=>"010011011",
  4793=>"000110111",
  4794=>"110011011",
  4795=>"001110010",
  4796=>"010100001",
  4797=>"010010000",
  4798=>"000100100",
  4799=>"011011101",
  4800=>"101001001",
  4801=>"001100101",
  4802=>"010011010",
  4803=>"001000011",
  4804=>"111100101",
  4805=>"100101111",
  4806=>"100011010",
  4807=>"011111100",
  4808=>"000010111",
  4809=>"110001110",
  4810=>"110101110",
  4811=>"011011101",
  4812=>"101010101",
  4813=>"100011010",
  4814=>"001101111",
  4815=>"110110011",
  4816=>"010000100",
  4817=>"001010001",
  4818=>"010111101",
  4819=>"000111001",
  4820=>"100111000",
  4821=>"011111010",
  4822=>"100001101",
  4823=>"000000001",
  4824=>"001110010",
  4825=>"011100011",
  4826=>"110101001",
  4827=>"010000011",
  4828=>"110101010",
  4829=>"010111101",
  4830=>"000010010",
  4831=>"011000011",
  4832=>"000100101",
  4833=>"110100101",
  4834=>"001011001",
  4835=>"011110010",
  4836=>"100100101",
  4837=>"001101110",
  4838=>"000110110",
  4839=>"101010101",
  4840=>"110111111",
  4841=>"110011101",
  4842=>"100101100",
  4843=>"101101000",
  4844=>"010000011",
  4845=>"000101001",
  4846=>"010010000",
  4847=>"101011110",
  4848=>"000001001",
  4849=>"010111011",
  4850=>"011001010",
  4851=>"010110001",
  4852=>"100100100",
  4853=>"100011000",
  4854=>"101010001",
  4855=>"000000010",
  4856=>"011001111",
  4857=>"111111110",
  4858=>"011101001",
  4859=>"001100100",
  4860=>"011111010",
  4861=>"010111011",
  4862=>"010100111",
  4863=>"001111011",
  4864=>"001011100",
  4865=>"001000001",
  4866=>"100101110",
  4867=>"100000111",
  4868=>"101010101",
  4869=>"110110111",
  4870=>"001101111",
  4871=>"100011000",
  4872=>"101011110",
  4873=>"001100010",
  4874=>"111001111",
  4875=>"100010101",
  4876=>"010101111",
  4877=>"001111101",
  4878=>"111111110",
  4879=>"111001110",
  4880=>"000011011",
  4881=>"101111000",
  4882=>"010110010",
  4883=>"101011011",
  4884=>"110010000",
  4885=>"100010001",
  4886=>"100111110",
  4887=>"100100011",
  4888=>"111100100",
  4889=>"110000000",
  4890=>"110000001",
  4891=>"000000010",
  4892=>"010110101",
  4893=>"100101110",
  4894=>"100011110",
  4895=>"011001110",
  4896=>"110000011",
  4897=>"000110001",
  4898=>"111101111",
  4899=>"101110100",
  4900=>"010100000",
  4901=>"000010110",
  4902=>"011001111",
  4903=>"001101100",
  4904=>"100010110",
  4905=>"110101001",
  4906=>"110001010",
  4907=>"000101111",
  4908=>"011000100",
  4909=>"101110100",
  4910=>"110110101",
  4911=>"100000111",
  4912=>"101011111",
  4913=>"101001011",
  4914=>"110101100",
  4915=>"111011110",
  4916=>"001000000",
  4917=>"110000011",
  4918=>"010000011",
  4919=>"100001111",
  4920=>"011100011",
  4921=>"010110100",
  4922=>"001000101",
  4923=>"101000001",
  4924=>"100001111",
  4925=>"100000010",
  4926=>"100010010",
  4927=>"011011011",
  4928=>"011110010",
  4929=>"001011111",
  4930=>"111001000",
  4931=>"111110110",
  4932=>"100000111",
  4933=>"111011000",
  4934=>"101100100",
  4935=>"000000000",
  4936=>"001000011",
  4937=>"010001000",
  4938=>"101001001",
  4939=>"000110100",
  4940=>"100111101",
  4941=>"100100011",
  4942=>"010100010",
  4943=>"100001010",
  4944=>"111101101",
  4945=>"000100100",
  4946=>"001110010",
  4947=>"000110001",
  4948=>"100111010",
  4949=>"010001011",
  4950=>"001001110",
  4951=>"110110011",
  4952=>"011000100",
  4953=>"100101101",
  4954=>"111111011",
  4955=>"010011101",
  4956=>"000011101",
  4957=>"101101000",
  4958=>"111011000",
  4959=>"110011100",
  4960=>"010111100",
  4961=>"001100110",
  4962=>"000010110",
  4963=>"111111000",
  4964=>"101000101",
  4965=>"010101000",
  4966=>"100111010",
  4967=>"111111001",
  4968=>"010100000",
  4969=>"111000010",
  4970=>"001111010",
  4971=>"010000101",
  4972=>"100101101",
  4973=>"100011101",
  4974=>"010100011",
  4975=>"101110111",
  4976=>"001000100",
  4977=>"111000100",
  4978=>"001101101",
  4979=>"010100000",
  4980=>"110100001",
  4981=>"100101101",
  4982=>"011010001",
  4983=>"100110010",
  4984=>"101110000",
  4985=>"110000011",
  4986=>"101101111",
  4987=>"000100100",
  4988=>"100110010",
  4989=>"000010101",
  4990=>"000101111",
  4991=>"011011110",
  4992=>"010101101",
  4993=>"001010100",
  4994=>"110011110",
  4995=>"110010100",
  4996=>"100110111",
  4997=>"101011011",
  4998=>"111011110",
  4999=>"010101100",
  5000=>"010111111",
  5001=>"001001110",
  5002=>"000010111",
  5003=>"101000100",
  5004=>"111000100",
  5005=>"101101010",
  5006=>"001000101",
  5007=>"011010001",
  5008=>"110110101",
  5009=>"000111101",
  5010=>"110000010",
  5011=>"101011000",
  5012=>"010101010",
  5013=>"100100001",
  5014=>"101011100",
  5015=>"000010110",
  5016=>"110100010",
  5017=>"101010011",
  5018=>"110011110",
  5019=>"101000001",
  5020=>"101001001",
  5021=>"111000101",
  5022=>"011111010",
  5023=>"100111101",
  5024=>"110011010",
  5025=>"110010001",
  5026=>"100001001",
  5027=>"010100011",
  5028=>"100110101",
  5029=>"010001101",
  5030=>"111001100",
  5031=>"100000010",
  5032=>"011010001",
  5033=>"000111001",
  5034=>"111010001",
  5035=>"001100010",
  5036=>"010110100",
  5037=>"111110111",
  5038=>"001110000",
  5039=>"100001111",
  5040=>"010010101",
  5041=>"101101110",
  5042=>"100000101",
  5043=>"010010101",
  5044=>"110110001",
  5045=>"110001001",
  5046=>"111011111",
  5047=>"101110111",
  5048=>"111000100",
  5049=>"010101100",
  5050=>"010110100",
  5051=>"111011001",
  5052=>"000110100",
  5053=>"100010010",
  5054=>"001111100",
  5055=>"100110001",
  5056=>"000100001",
  5057=>"011010100",
  5058=>"010111110",
  5059=>"101100001",
  5060=>"001011110",
  5061=>"010000010",
  5062=>"001000111",
  5063=>"111100001",
  5064=>"100100000",
  5065=>"110110000",
  5066=>"110000000",
  5067=>"010011111",
  5068=>"100010000",
  5069=>"100010101",
  5070=>"000000100",
  5071=>"010010110",
  5072=>"111101001",
  5073=>"011111000",
  5074=>"010100110",
  5075=>"101001100",
  5076=>"001000100",
  5077=>"110100000",
  5078=>"100101101",
  5079=>"111100001",
  5080=>"100111111",
  5081=>"001111111",
  5082=>"010100111",
  5083=>"101111101",
  5084=>"100100010",
  5085=>"010010010",
  5086=>"000100100",
  5087=>"000011011",
  5088=>"011100100",
  5089=>"100011010",
  5090=>"101111011",
  5091=>"100001001",
  5092=>"000100100",
  5093=>"000100011",
  5094=>"001111101",
  5095=>"110110110",
  5096=>"000111000",
  5097=>"011000111",
  5098=>"000010000",
  5099=>"101110101",
  5100=>"110111000",
  5101=>"111100100",
  5102=>"011101100",
  5103=>"110101111",
  5104=>"001001001",
  5105=>"010000010",
  5106=>"100001110",
  5107=>"101011100",
  5108=>"011010110",
  5109=>"100101010",
  5110=>"001010110",
  5111=>"100010101",
  5112=>"110011010",
  5113=>"111111011",
  5114=>"110011110",
  5115=>"001010000",
  5116=>"010010101",
  5117=>"001001001",
  5118=>"111001111",
  5119=>"001010010",
  5120=>"010001011",
  5121=>"011010001",
  5122=>"000110000",
  5123=>"100101000",
  5124=>"110001011",
  5125=>"111001111",
  5126=>"001011000",
  5127=>"001001001",
  5128=>"010100100",
  5129=>"011111011",
  5130=>"011010100",
  5131=>"011001000",
  5132=>"010101000",
  5133=>"010110110",
  5134=>"110000110",
  5135=>"010100101",
  5136=>"010111011",
  5137=>"011001111",
  5138=>"100000100",
  5139=>"111101101",
  5140=>"000011100",
  5141=>"000001100",
  5142=>"110011100",
  5143=>"001011001",
  5144=>"000010110",
  5145=>"101101111",
  5146=>"101110011",
  5147=>"000010001",
  5148=>"001110010",
  5149=>"101011011",
  5150=>"011000000",
  5151=>"000111011",
  5152=>"100110110",
  5153=>"011001000",
  5154=>"000010110",
  5155=>"110000100",
  5156=>"110001110",
  5157=>"110111000",
  5158=>"101010101",
  5159=>"111100101",
  5160=>"100101001",
  5161=>"110110110",
  5162=>"101010011",
  5163=>"100001011",
  5164=>"000111010",
  5165=>"101010100",
  5166=>"001110110",
  5167=>"101100101",
  5168=>"000100100",
  5169=>"111101010",
  5170=>"110100111",
  5171=>"111010111",
  5172=>"001101011",
  5173=>"000010000",
  5174=>"100111101",
  5175=>"100111111",
  5176=>"000111101",
  5177=>"110010101",
  5178=>"010010101",
  5179=>"010111000",
  5180=>"001110001",
  5181=>"010000001",
  5182=>"110011001",
  5183=>"111011110",
  5184=>"101110010",
  5185=>"001110011",
  5186=>"011001000",
  5187=>"000100111",
  5188=>"110000110",
  5189=>"101110000",
  5190=>"100000111",
  5191=>"000110000",
  5192=>"110111011",
  5193=>"101001011",
  5194=>"101101001",
  5195=>"100101001",
  5196=>"110100000",
  5197=>"100011011",
  5198=>"011000000",
  5199=>"000001110",
  5200=>"000111110",
  5201=>"001111010",
  5202=>"101100010",
  5203=>"000000000",
  5204=>"001000000",
  5205=>"001011010",
  5206=>"011101110",
  5207=>"110111011",
  5208=>"001001100",
  5209=>"100010100",
  5210=>"101110101",
  5211=>"000000000",
  5212=>"000100001",
  5213=>"000010110",
  5214=>"001010110",
  5215=>"011000000",
  5216=>"000111111",
  5217=>"010001111",
  5218=>"000001101",
  5219=>"100000001",
  5220=>"101111111",
  5221=>"100000110",
  5222=>"000001011",
  5223=>"110111110",
  5224=>"011101001",
  5225=>"100111110",
  5226=>"001011101",
  5227=>"010001001",
  5228=>"100010101",
  5229=>"101101110",
  5230=>"101101111",
  5231=>"001010001",
  5232=>"010000101",
  5233=>"010100011",
  5234=>"000111100",
  5235=>"011001010",
  5236=>"110001010",
  5237=>"000001101",
  5238=>"011110011",
  5239=>"100010110",
  5240=>"101001010",
  5241=>"100000011",
  5242=>"011001101",
  5243=>"111111111",
  5244=>"110110101",
  5245=>"101111111",
  5246=>"100111111",
  5247=>"100010000",
  5248=>"000101101",
  5249=>"111110011",
  5250=>"110001100",
  5251=>"101000110",
  5252=>"000000001",
  5253=>"011010110",
  5254=>"010100000",
  5255=>"111010101",
  5256=>"110110011",
  5257=>"100011000",
  5258=>"011011011",
  5259=>"111000010",
  5260=>"100011100",
  5261=>"101001100",
  5262=>"110001001",
  5263=>"111100100",
  5264=>"000110110",
  5265=>"101000001",
  5266=>"110001011",
  5267=>"010010110",
  5268=>"111111111",
  5269=>"000011001",
  5270=>"001111010",
  5271=>"001011010",
  5272=>"110110101",
  5273=>"000100100",
  5274=>"010000010",
  5275=>"001110100",
  5276=>"111110011",
  5277=>"111111000",
  5278=>"010011001",
  5279=>"111011110",
  5280=>"110011001",
  5281=>"111000100",
  5282=>"010100100",
  5283=>"110010111",
  5284=>"101011001",
  5285=>"110101001",
  5286=>"000111110",
  5287=>"100010001",
  5288=>"100111000",
  5289=>"110110100",
  5290=>"011110000",
  5291=>"111011001",
  5292=>"010101010",
  5293=>"000110010",
  5294=>"111100011",
  5295=>"000001100",
  5296=>"101110000",
  5297=>"001000011",
  5298=>"001001110",
  5299=>"100100100",
  5300=>"100111100",
  5301=>"000000101",
  5302=>"010100100",
  5303=>"100111011",
  5304=>"010001000",
  5305=>"101010011",
  5306=>"110010110",
  5307=>"111110101",
  5308=>"100100000",
  5309=>"111110110",
  5310=>"101110100",
  5311=>"010101101",
  5312=>"000000011",
  5313=>"000101010",
  5314=>"111011110",
  5315=>"110001111",
  5316=>"101010000",
  5317=>"110001011",
  5318=>"110100010",
  5319=>"101110110",
  5320=>"100001010",
  5321=>"111011111",
  5322=>"100100001",
  5323=>"101110011",
  5324=>"111010011",
  5325=>"000011010",
  5326=>"011111100",
  5327=>"100010000",
  5328=>"000011111",
  5329=>"010100010",
  5330=>"010111001",
  5331=>"001111101",
  5332=>"010100111",
  5333=>"010000101",
  5334=>"110010100",
  5335=>"110010101",
  5336=>"011111000",
  5337=>"000011011",
  5338=>"101101000",
  5339=>"100101000",
  5340=>"100110000",
  5341=>"001100101",
  5342=>"111010000",
  5343=>"011001101",
  5344=>"011010000",
  5345=>"011100101",
  5346=>"110011101",
  5347=>"101000011",
  5348=>"001110011",
  5349=>"110000011",
  5350=>"100100011",
  5351=>"011011001",
  5352=>"000011100",
  5353=>"000001111",
  5354=>"001110100",
  5355=>"010000110",
  5356=>"000111100",
  5357=>"010000110",
  5358=>"111100111",
  5359=>"100100110",
  5360=>"100100010",
  5361=>"000100000",
  5362=>"111101010",
  5363=>"010111010",
  5364=>"010100011",
  5365=>"001110110",
  5366=>"000011100",
  5367=>"000111111",
  5368=>"011101110",
  5369=>"101111001",
  5370=>"100011111",
  5371=>"000010000",
  5372=>"110011000",
  5373=>"011010101",
  5374=>"010100001",
  5375=>"100000101",
  5376=>"010001010",
  5377=>"000100000",
  5378=>"010001101",
  5379=>"111010101",
  5380=>"010110111",
  5381=>"100011000",
  5382=>"011110110",
  5383=>"000101110",
  5384=>"011010110",
  5385=>"011110011",
  5386=>"101101010",
  5387=>"001000000",
  5388=>"011000000",
  5389=>"000001011",
  5390=>"101001111",
  5391=>"000010011",
  5392=>"011000010",
  5393=>"110111011",
  5394=>"110101010",
  5395=>"111011110",
  5396=>"011101111",
  5397=>"000110011",
  5398=>"110000101",
  5399=>"110111110",
  5400=>"010110010",
  5401=>"010011100",
  5402=>"010111000",
  5403=>"011111111",
  5404=>"110000000",
  5405=>"010000111",
  5406=>"111110001",
  5407=>"011111101",
  5408=>"000000010",
  5409=>"010011101",
  5410=>"010110011",
  5411=>"011000111",
  5412=>"101011011",
  5413=>"011011001",
  5414=>"010011000",
  5415=>"011000101",
  5416=>"010111110",
  5417=>"101001111",
  5418=>"011010011",
  5419=>"010111000",
  5420=>"010000001",
  5421=>"010111011",
  5422=>"011111000",
  5423=>"101000111",
  5424=>"001101011",
  5425=>"000100101",
  5426=>"000000111",
  5427=>"101101101",
  5428=>"111110011",
  5429=>"110111111",
  5430=>"010000111",
  5431=>"110001000",
  5432=>"000001000",
  5433=>"001111111",
  5434=>"001100101",
  5435=>"110101101",
  5436=>"000110111",
  5437=>"011010110",
  5438=>"001001011",
  5439=>"110100010",
  5440=>"101000110",
  5441=>"011101001",
  5442=>"011110011",
  5443=>"010001011",
  5444=>"110111100",
  5445=>"001110000",
  5446=>"001111000",
  5447=>"110001000",
  5448=>"000011100",
  5449=>"001010011",
  5450=>"010111011",
  5451=>"001111111",
  5452=>"101110111",
  5453=>"100000101",
  5454=>"010111000",
  5455=>"011100001",
  5456=>"010000001",
  5457=>"110011111",
  5458=>"111101100",
  5459=>"011100001",
  5460=>"011100110",
  5461=>"110100100",
  5462=>"001000110",
  5463=>"011001100",
  5464=>"000101110",
  5465=>"101101111",
  5466=>"111110001",
  5467=>"010000000",
  5468=>"111011110",
  5469=>"001001011",
  5470=>"001001001",
  5471=>"001101011",
  5472=>"001111100",
  5473=>"001110110",
  5474=>"101110101",
  5475=>"010000111",
  5476=>"101100101",
  5477=>"101000111",
  5478=>"100011011",
  5479=>"111101110",
  5480=>"100101100",
  5481=>"100110110",
  5482=>"010011011",
  5483=>"001011110",
  5484=>"101001010",
  5485=>"010000001",
  5486=>"110110000",
  5487=>"101111000",
  5488=>"100111111",
  5489=>"000100111",
  5490=>"100100100",
  5491=>"110101101",
  5492=>"100000100",
  5493=>"110111110",
  5494=>"101010001",
  5495=>"110001110",
  5496=>"010101101",
  5497=>"010111000",
  5498=>"110001011",
  5499=>"111110101",
  5500=>"111111101",
  5501=>"001110011",
  5502=>"101101010",
  5503=>"011111100",
  5504=>"000011110",
  5505=>"010000110",
  5506=>"101010000",
  5507=>"100111010",
  5508=>"111100001",
  5509=>"001001100",
  5510=>"001100011",
  5511=>"000110000",
  5512=>"011111011",
  5513=>"010111101",
  5514=>"101001100",
  5515=>"110111110",
  5516=>"000011001",
  5517=>"100111001",
  5518=>"011011111",
  5519=>"000101110",
  5520=>"111111000",
  5521=>"011111101",
  5522=>"010010011",
  5523=>"000000000",
  5524=>"111010001",
  5525=>"100011010",
  5526=>"101000111",
  5527=>"001000110",
  5528=>"000101000",
  5529=>"011000100",
  5530=>"101000011",
  5531=>"100101010",
  5532=>"111001001",
  5533=>"011110001",
  5534=>"110001000",
  5535=>"000101110",
  5536=>"000101110",
  5537=>"100010101",
  5538=>"010110111",
  5539=>"010010111",
  5540=>"101010001",
  5541=>"010111111",
  5542=>"110111001",
  5543=>"000001001",
  5544=>"001000010",
  5545=>"010101110",
  5546=>"011001011",
  5547=>"011110100",
  5548=>"001001010",
  5549=>"110001000",
  5550=>"111111111",
  5551=>"001001000",
  5552=>"100001011",
  5553=>"010111111",
  5554=>"001100110",
  5555=>"010110011",
  5556=>"110111111",
  5557=>"011100110",
  5558=>"111100010",
  5559=>"011110111",
  5560=>"000000000",
  5561=>"010111011",
  5562=>"111010110",
  5563=>"101100011",
  5564=>"010100111",
  5565=>"100111001",
  5566=>"111010100",
  5567=>"110101001",
  5568=>"111011101",
  5569=>"110101001",
  5570=>"001101101",
  5571=>"100110010",
  5572=>"001100111",
  5573=>"101110111",
  5574=>"000100010",
  5575=>"010110011",
  5576=>"111011000",
  5577=>"011111010",
  5578=>"101000000",
  5579=>"101111000",
  5580=>"111111111",
  5581=>"011010110",
  5582=>"000001001",
  5583=>"011000001",
  5584=>"110001001",
  5585=>"011011101",
  5586=>"011110111",
  5587=>"100011000",
  5588=>"011010111",
  5589=>"100111110",
  5590=>"100010010",
  5591=>"001000010",
  5592=>"000001010",
  5593=>"001011100",
  5594=>"010001100",
  5595=>"111000101",
  5596=>"110011001",
  5597=>"011111011",
  5598=>"110010000",
  5599=>"011010111",
  5600=>"101011000",
  5601=>"110101001",
  5602=>"000011010",
  5603=>"000010101",
  5604=>"001000001",
  5605=>"001100110",
  5606=>"011000000",
  5607=>"100001010",
  5608=>"110011011",
  5609=>"111111011",
  5610=>"001110000",
  5611=>"010000101",
  5612=>"001010101",
  5613=>"111101101",
  5614=>"001101011",
  5615=>"000000010",
  5616=>"011000101",
  5617=>"111011010",
  5618=>"111100101",
  5619=>"001010000",
  5620=>"101010100",
  5621=>"100000010",
  5622=>"111111000",
  5623=>"011111110",
  5624=>"010111101",
  5625=>"100011001",
  5626=>"101111110",
  5627=>"100000010",
  5628=>"110110010",
  5629=>"001111001",
  5630=>"011110010",
  5631=>"100101000",
  5632=>"000000001",
  5633=>"010100101",
  5634=>"111001000",
  5635=>"000011100",
  5636=>"101001101",
  5637=>"110111011",
  5638=>"000000111",
  5639=>"011010110",
  5640=>"111001110",
  5641=>"010000000",
  5642=>"000001110",
  5643=>"011000011",
  5644=>"100110110",
  5645=>"111000100",
  5646=>"000001111",
  5647=>"111001101",
  5648=>"000100100",
  5649=>"100001010",
  5650=>"101011101",
  5651=>"110111101",
  5652=>"110000111",
  5653=>"100111011",
  5654=>"111111100",
  5655=>"001010000",
  5656=>"010001100",
  5657=>"100000010",
  5658=>"110110010",
  5659=>"010100011",
  5660=>"100010101",
  5661=>"100011100",
  5662=>"100000101",
  5663=>"100111101",
  5664=>"011110011",
  5665=>"100000101",
  5666=>"010110010",
  5667=>"110110010",
  5668=>"101001101",
  5669=>"100101011",
  5670=>"000101011",
  5671=>"101101011",
  5672=>"010001101",
  5673=>"001011101",
  5674=>"011000110",
  5675=>"100101010",
  5676=>"100011010",
  5677=>"001100110",
  5678=>"100000101",
  5679=>"001011101",
  5680=>"000001000",
  5681=>"011111110",
  5682=>"000111011",
  5683=>"011100000",
  5684=>"101011111",
  5685=>"101111110",
  5686=>"011011001",
  5687=>"010100100",
  5688=>"001110000",
  5689=>"001101010",
  5690=>"101010000",
  5691=>"010000100",
  5692=>"110101011",
  5693=>"111011100",
  5694=>"111111010",
  5695=>"010000110",
  5696=>"001011000",
  5697=>"100111101",
  5698=>"101010001",
  5699=>"111101100",
  5700=>"011011000",
  5701=>"010011110",
  5702=>"101010001",
  5703=>"100001001",
  5704=>"000110011",
  5705=>"101101111",
  5706=>"010110010",
  5707=>"001111011",
  5708=>"110010001",
  5709=>"000100101",
  5710=>"000111110",
  5711=>"011101010",
  5712=>"000000000",
  5713=>"101010101",
  5714=>"010001000",
  5715=>"001110010",
  5716=>"101111111",
  5717=>"000010010",
  5718=>"000001010",
  5719=>"110110100",
  5720=>"000111111",
  5721=>"000100111",
  5722=>"000010111",
  5723=>"000110110",
  5724=>"101001100",
  5725=>"000100010",
  5726=>"110111001",
  5727=>"100111101",
  5728=>"111110111",
  5729=>"001000010",
  5730=>"111010111",
  5731=>"101110110",
  5732=>"000100110",
  5733=>"000000000",
  5734=>"110000010",
  5735=>"001100110",
  5736=>"000000110",
  5737=>"000010011",
  5738=>"110001010",
  5739=>"111111100",
  5740=>"010110111",
  5741=>"001110110",
  5742=>"100101001",
  5743=>"011010001",
  5744=>"111101010",
  5745=>"010100101",
  5746=>"110000011",
  5747=>"100010110",
  5748=>"110111011",
  5749=>"010010110",
  5750=>"011000111",
  5751=>"010111111",
  5752=>"011000111",
  5753=>"001111101",
  5754=>"101100010",
  5755=>"001110111",
  5756=>"100100010",
  5757=>"110101011",
  5758=>"001000001",
  5759=>"111110100",
  5760=>"000101011",
  5761=>"111000100",
  5762=>"010101010",
  5763=>"110111010",
  5764=>"111101110",
  5765=>"110110101",
  5766=>"111010110",
  5767=>"001101111",
  5768=>"011001111",
  5769=>"010111010",
  5770=>"001110010",
  5771=>"100011110",
  5772=>"110000001",
  5773=>"011101111",
  5774=>"000111100",
  5775=>"100110101",
  5776=>"111110010",
  5777=>"100110110",
  5778=>"010001100",
  5779=>"000110001",
  5780=>"111010011",
  5781=>"111010101",
  5782=>"010010100",
  5783=>"111111000",
  5784=>"110001100",
  5785=>"001000001",
  5786=>"000000011",
  5787=>"111101100",
  5788=>"100011011",
  5789=>"010000111",
  5790=>"110111100",
  5791=>"010000111",
  5792=>"111001101",
  5793=>"111111101",
  5794=>"111101000",
  5795=>"001011111",
  5796=>"010110011",
  5797=>"110001000",
  5798=>"010111000",
  5799=>"110010000",
  5800=>"001010001",
  5801=>"000001101",
  5802=>"011011010",
  5803=>"100100110",
  5804=>"100100111",
  5805=>"110010010",
  5806=>"111010000",
  5807=>"110110111",
  5808=>"001000001",
  5809=>"111001011",
  5810=>"000001010",
  5811=>"011000100",
  5812=>"111100111",
  5813=>"010000001",
  5814=>"011000001",
  5815=>"001110001",
  5816=>"100110110",
  5817=>"010000110",
  5818=>"001101001",
  5819=>"110111011",
  5820=>"010000101",
  5821=>"011010101",
  5822=>"110011010",
  5823=>"110001100",
  5824=>"000000000",
  5825=>"111101101",
  5826=>"110110010",
  5827=>"010101100",
  5828=>"110000110",
  5829=>"011001101",
  5830=>"001001111",
  5831=>"110011010",
  5832=>"110001000",
  5833=>"100011011",
  5834=>"111101101",
  5835=>"110001011",
  5836=>"000100110",
  5837=>"110101110",
  5838=>"111010110",
  5839=>"111100110",
  5840=>"101000010",
  5841=>"110110001",
  5842=>"110100110",
  5843=>"111110111",
  5844=>"000000101",
  5845=>"001100001",
  5846=>"111100110",
  5847=>"001101010",
  5848=>"010011110",
  5849=>"100111110",
  5850=>"001110001",
  5851=>"000010010",
  5852=>"011000111",
  5853=>"111100111",
  5854=>"001100011",
  5855=>"100101111",
  5856=>"101110011",
  5857=>"000001100",
  5858=>"110001110",
  5859=>"010010100",
  5860=>"001111010",
  5861=>"011110110",
  5862=>"000001000",
  5863=>"100101000",
  5864=>"000110001",
  5865=>"011110100",
  5866=>"001001010",
  5867=>"101010010",
  5868=>"010001111",
  5869=>"111000100",
  5870=>"100011001",
  5871=>"111110110",
  5872=>"110100010",
  5873=>"110010100",
  5874=>"101111110",
  5875=>"110101000",
  5876=>"011101011",
  5877=>"011110100",
  5878=>"011010111",
  5879=>"011000011",
  5880=>"111101000",
  5881=>"011010001",
  5882=>"011110110",
  5883=>"100100111",
  5884=>"010100010",
  5885=>"111100000",
  5886=>"110011111",
  5887=>"010100110",
  5888=>"000001011",
  5889=>"101111010",
  5890=>"000110011",
  5891=>"001101011",
  5892=>"001010001",
  5893=>"111100010",
  5894=>"111000101",
  5895=>"110101101",
  5896=>"100100100",
  5897=>"100101000",
  5898=>"111010101",
  5899=>"101010101",
  5900=>"001100101",
  5901=>"110111110",
  5902=>"011011011",
  5903=>"110101011",
  5904=>"011011100",
  5905=>"110000101",
  5906=>"111000011",
  5907=>"000110101",
  5908=>"000010110",
  5909=>"110101000",
  5910=>"111010110",
  5911=>"101111000",
  5912=>"011011001",
  5913=>"010011011",
  5914=>"101101010",
  5915=>"100100110",
  5916=>"011111100",
  5917=>"110100001",
  5918=>"000101101",
  5919=>"010001111",
  5920=>"111111100",
  5921=>"010011000",
  5922=>"100000111",
  5923=>"100110010",
  5924=>"001000110",
  5925=>"111111010",
  5926=>"011011001",
  5927=>"110101001",
  5928=>"101011110",
  5929=>"110110010",
  5930=>"010111011",
  5931=>"100101000",
  5932=>"110001000",
  5933=>"111111001",
  5934=>"111111101",
  5935=>"101111011",
  5936=>"000011010",
  5937=>"011111001",
  5938=>"100110011",
  5939=>"100000100",
  5940=>"001111110",
  5941=>"010010001",
  5942=>"010011001",
  5943=>"011000001",
  5944=>"110100000",
  5945=>"010000101",
  5946=>"111001110",
  5947=>"010100001",
  5948=>"111001011",
  5949=>"010110110",
  5950=>"110111010",
  5951=>"101010001",
  5952=>"100110011",
  5953=>"000100101",
  5954=>"111001110",
  5955=>"000000101",
  5956=>"100111000",
  5957=>"011010110",
  5958=>"011111000",
  5959=>"011111001",
  5960=>"111011110",
  5961=>"011000010",
  5962=>"110100011",
  5963=>"000111100",
  5964=>"010000100",
  5965=>"001011111",
  5966=>"001011001",
  5967=>"101100011",
  5968=>"001110010",
  5969=>"000100101",
  5970=>"110100001",
  5971=>"000010010",
  5972=>"000101101",
  5973=>"100011111",
  5974=>"100010010",
  5975=>"110110011",
  5976=>"001000011",
  5977=>"001100000",
  5978=>"101100100",
  5979=>"000110101",
  5980=>"110011010",
  5981=>"111001010",
  5982=>"110100111",
  5983=>"010010000",
  5984=>"110001010",
  5985=>"001111101",
  5986=>"001000010",
  5987=>"011110111",
  5988=>"000111100",
  5989=>"011001111",
  5990=>"001000010",
  5991=>"001000000",
  5992=>"100001100",
  5993=>"001111010",
  5994=>"111100100",
  5995=>"010010110",
  5996=>"001110001",
  5997=>"011010011",
  5998=>"100000111",
  5999=>"101000001",
  6000=>"000100001",
  6001=>"110101111",
  6002=>"101101100",
  6003=>"100101101",
  6004=>"111110101",
  6005=>"101000010",
  6006=>"100101000",
  6007=>"110110011",
  6008=>"110000010",
  6009=>"010011110",
  6010=>"010011101",
  6011=>"001100110",
  6012=>"011001010",
  6013=>"110000011",
  6014=>"011110000",
  6015=>"001001000",
  6016=>"110111011",
  6017=>"111010110",
  6018=>"001111001",
  6019=>"010111111",
  6020=>"100101011",
  6021=>"000110101",
  6022=>"111101110",
  6023=>"010011000",
  6024=>"000110011",
  6025=>"001000000",
  6026=>"100010010",
  6027=>"111111111",
  6028=>"010001001",
  6029=>"000000000",
  6030=>"010000100",
  6031=>"111100000",
  6032=>"101110011",
  6033=>"001110101",
  6034=>"000100100",
  6035=>"100000000",
  6036=>"010110000",
  6037=>"100010111",
  6038=>"101100011",
  6039=>"111010011",
  6040=>"010110010",
  6041=>"001010011",
  6042=>"100001110",
  6043=>"110100101",
  6044=>"110000100",
  6045=>"010001001",
  6046=>"110011000",
  6047=>"101100001",
  6048=>"100111100",
  6049=>"011001000",
  6050=>"011001101",
  6051=>"101111100",
  6052=>"011100000",
  6053=>"111111111",
  6054=>"000000011",
  6055=>"001010101",
  6056=>"001010111",
  6057=>"100111010",
  6058=>"100000111",
  6059=>"010110101",
  6060=>"110001110",
  6061=>"000010000",
  6062=>"101100101",
  6063=>"110100010",
  6064=>"000110100",
  6065=>"000001001",
  6066=>"000011010",
  6067=>"110100110",
  6068=>"010011100",
  6069=>"100110110",
  6070=>"000101100",
  6071=>"001001111",
  6072=>"011001101",
  6073=>"010000111",
  6074=>"010010000",
  6075=>"011111001",
  6076=>"010111001",
  6077=>"111001101",
  6078=>"001101100",
  6079=>"111000000",
  6080=>"111111001",
  6081=>"011110100",
  6082=>"000110110",
  6083=>"010011010",
  6084=>"111011010",
  6085=>"110111010",
  6086=>"011011001",
  6087=>"011000100",
  6088=>"000000100",
  6089=>"011111101",
  6090=>"010011110",
  6091=>"011000100",
  6092=>"001110010",
  6093=>"110011011",
  6094=>"101100110",
  6095=>"100110101",
  6096=>"110101000",
  6097=>"110001100",
  6098=>"111110101",
  6099=>"110011111",
  6100=>"110011001",
  6101=>"101011110",
  6102=>"011001010",
  6103=>"010001101",
  6104=>"111111111",
  6105=>"110111110",
  6106=>"001000000",
  6107=>"101010000",
  6108=>"101010001",
  6109=>"011000010",
  6110=>"100101101",
  6111=>"111001101",
  6112=>"111101111",
  6113=>"001001111",
  6114=>"000101100",
  6115=>"101011011",
  6116=>"010011101",
  6117=>"111010100",
  6118=>"111101111",
  6119=>"000010111",
  6120=>"110011100",
  6121=>"101010111",
  6122=>"001011000",
  6123=>"111100111",
  6124=>"000000001",
  6125=>"101010101",
  6126=>"011101111",
  6127=>"111110000",
  6128=>"101100001",
  6129=>"001011011",
  6130=>"101110100",
  6131=>"010111101",
  6132=>"100011001",
  6133=>"100100110",
  6134=>"011101100",
  6135=>"111101111",
  6136=>"101001000",
  6137=>"111001010",
  6138=>"110000111",
  6139=>"010000111",
  6140=>"101101001",
  6141=>"011010110",
  6142=>"100010111",
  6143=>"011111111",
  6144=>"100101000",
  6145=>"000111010",
  6146=>"000010111",
  6147=>"100001110",
  6148=>"001111010",
  6149=>"111101100",
  6150=>"011100010",
  6151=>"000010011",
  6152=>"110001101",
  6153=>"000100110",
  6154=>"101110111",
  6155=>"110001111",
  6156=>"001000110",
  6157=>"011100101",
  6158=>"101010001",
  6159=>"011001011",
  6160=>"000010011",
  6161=>"001011001",
  6162=>"010010101",
  6163=>"000001100",
  6164=>"011100100",
  6165=>"100111011",
  6166=>"011000010",
  6167=>"101011011",
  6168=>"000001100",
  6169=>"001010000",
  6170=>"010111100",
  6171=>"001000111",
  6172=>"100011100",
  6173=>"111011011",
  6174=>"100011110",
  6175=>"111001111",
  6176=>"100011100",
  6177=>"100000001",
  6178=>"011010001",
  6179=>"011101101",
  6180=>"111110010",
  6181=>"011010100",
  6182=>"000000010",
  6183=>"111100000",
  6184=>"100011111",
  6185=>"110000110",
  6186=>"110110100",
  6187=>"011011111",
  6188=>"001001110",
  6189=>"011010101",
  6190=>"111011100",
  6191=>"111001001",
  6192=>"001001011",
  6193=>"001010000",
  6194=>"111101101",
  6195=>"010110101",
  6196=>"111010000",
  6197=>"010000001",
  6198=>"111110110",
  6199=>"010101100",
  6200=>"101011000",
  6201=>"111110000",
  6202=>"010101011",
  6203=>"000100000",
  6204=>"000011011",
  6205=>"101011011",
  6206=>"010101101",
  6207=>"111010000",
  6208=>"111110000",
  6209=>"010100010",
  6210=>"111000000",
  6211=>"111100100",
  6212=>"000000110",
  6213=>"010011101",
  6214=>"010000101",
  6215=>"000100100",
  6216=>"000100101",
  6217=>"001110110",
  6218=>"111111110",
  6219=>"110110001",
  6220=>"010110100",
  6221=>"111011001",
  6222=>"001010011",
  6223=>"010100001",
  6224=>"101100110",
  6225=>"111101111",
  6226=>"111110101",
  6227=>"000100111",
  6228=>"100010110",
  6229=>"111000101",
  6230=>"000101111",
  6231=>"011010110",
  6232=>"000001010",
  6233=>"100100111",
  6234=>"110101001",
  6235=>"100100110",
  6236=>"001011100",
  6237=>"111011010",
  6238=>"101010111",
  6239=>"110011000",
  6240=>"110000111",
  6241=>"001111101",
  6242=>"000010000",
  6243=>"101001010",
  6244=>"110100010",
  6245=>"111001100",
  6246=>"001110000",
  6247=>"011011001",
  6248=>"101100011",
  6249=>"110110010",
  6250=>"100100111",
  6251=>"011111001",
  6252=>"110101010",
  6253=>"100000010",
  6254=>"111011100",
  6255=>"110110011",
  6256=>"000110110",
  6257=>"000011000",
  6258=>"111011110",
  6259=>"110010010",
  6260=>"000111001",
  6261=>"001101000",
  6262=>"111111011",
  6263=>"111110001",
  6264=>"111010110",
  6265=>"010110111",
  6266=>"111000101",
  6267=>"100011011",
  6268=>"010100011",
  6269=>"000010010",
  6270=>"000100011",
  6271=>"111100100",
  6272=>"100010100",
  6273=>"110111111",
  6274=>"110010000",
  6275=>"111110100",
  6276=>"111101101",
  6277=>"010111100",
  6278=>"101011110",
  6279=>"111100110",
  6280=>"111100010",
  6281=>"110011100",
  6282=>"011010100",
  6283=>"100110010",
  6284=>"111101011",
  6285=>"111111100",
  6286=>"001111010",
  6287=>"011010010",
  6288=>"011101010",
  6289=>"011011011",
  6290=>"110010001",
  6291=>"101110100",
  6292=>"010111101",
  6293=>"101100110",
  6294=>"010001000",
  6295=>"100001011",
  6296=>"001000011",
  6297=>"110110011",
  6298=>"110100001",
  6299=>"000110110",
  6300=>"001001100",
  6301=>"101110100",
  6302=>"110001100",
  6303=>"101000010",
  6304=>"100111100",
  6305=>"110110000",
  6306=>"100101101",
  6307=>"010000111",
  6308=>"001111111",
  6309=>"010000100",
  6310=>"001000011",
  6311=>"111011111",
  6312=>"110010001",
  6313=>"011101101",
  6314=>"111101111",
  6315=>"100000101",
  6316=>"001101111",
  6317=>"110010100",
  6318=>"110111011",
  6319=>"011111111",
  6320=>"001010010",
  6321=>"000001000",
  6322=>"101100100",
  6323=>"001010111",
  6324=>"001111100",
  6325=>"000110101",
  6326=>"010001100",
  6327=>"001100110",
  6328=>"010101100",
  6329=>"011010010",
  6330=>"111111111",
  6331=>"111001111",
  6332=>"001011011",
  6333=>"100110111",
  6334=>"111101001",
  6335=>"111110101",
  6336=>"011111101",
  6337=>"110100000",
  6338=>"111000101",
  6339=>"111100011",
  6340=>"000000101",
  6341=>"110111110",
  6342=>"011110111",
  6343=>"001000000",
  6344=>"000111100",
  6345=>"101101000",
  6346=>"111010111",
  6347=>"010111100",
  6348=>"100111110",
  6349=>"110111101",
  6350=>"100101101",
  6351=>"001000001",
  6352=>"110000101",
  6353=>"011101001",
  6354=>"100001011",
  6355=>"001111101",
  6356=>"100001001",
  6357=>"101111000",
  6358=>"000001001",
  6359=>"100101100",
  6360=>"111011001",
  6361=>"011111100",
  6362=>"000100000",
  6363=>"001001101",
  6364=>"111011000",
  6365=>"001010110",
  6366=>"101101010",
  6367=>"011110011",
  6368=>"111010001",
  6369=>"111111001",
  6370=>"101111000",
  6371=>"100101010",
  6372=>"011000001",
  6373=>"001000101",
  6374=>"111000011",
  6375=>"010100001",
  6376=>"000001100",
  6377=>"001110001",
  6378=>"100000111",
  6379=>"000111111",
  6380=>"010011111",
  6381=>"011000110",
  6382=>"100110110",
  6383=>"001111010",
  6384=>"111111000",
  6385=>"001110000",
  6386=>"010001010",
  6387=>"000101010",
  6388=>"001010011",
  6389=>"011111111",
  6390=>"000001001",
  6391=>"011111110",
  6392=>"101011000",
  6393=>"110100011",
  6394=>"010101011",
  6395=>"000000010",
  6396=>"010110100",
  6397=>"011001100",
  6398=>"011110011",
  6399=>"011000001",
  6400=>"100100110",
  6401=>"100111101",
  6402=>"100010111",
  6403=>"110111110",
  6404=>"101100011",
  6405=>"000000100",
  6406=>"111010100",
  6407=>"010111110",
  6408=>"011010111",
  6409=>"001101111",
  6410=>"000110101",
  6411=>"111000100",
  6412=>"110111101",
  6413=>"000000011",
  6414=>"100101010",
  6415=>"101000001",
  6416=>"100111111",
  6417=>"010001001",
  6418=>"101100001",
  6419=>"111011100",
  6420=>"000111010",
  6421=>"100111001",
  6422=>"110110111",
  6423=>"110000011",
  6424=>"011011000",
  6425=>"011101011",
  6426=>"011010010",
  6427=>"000000110",
  6428=>"000100110",
  6429=>"000111111",
  6430=>"110010011",
  6431=>"000010011",
  6432=>"000011000",
  6433=>"000000000",
  6434=>"110111011",
  6435=>"000001011",
  6436=>"000011110",
  6437=>"001000101",
  6438=>"000111011",
  6439=>"100111011",
  6440=>"110000111",
  6441=>"001101101",
  6442=>"001000101",
  6443=>"101101001",
  6444=>"000100001",
  6445=>"000001010",
  6446=>"000100000",
  6447=>"101110111",
  6448=>"001010000",
  6449=>"000010111",
  6450=>"011111101",
  6451=>"100011000",
  6452=>"011100011",
  6453=>"101111000",
  6454=>"011000010",
  6455=>"101100100",
  6456=>"111000001",
  6457=>"110010011",
  6458=>"100110011",
  6459=>"000000111",
  6460=>"111111011",
  6461=>"000110011",
  6462=>"111101001",
  6463=>"010111010",
  6464=>"110010100",
  6465=>"101111000",
  6466=>"111111111",
  6467=>"000111111",
  6468=>"110010110",
  6469=>"111110010",
  6470=>"101001010",
  6471=>"000100011",
  6472=>"000000011",
  6473=>"110010100",
  6474=>"010001011",
  6475=>"110101000",
  6476=>"011111011",
  6477=>"111000101",
  6478=>"110110010",
  6479=>"111111010",
  6480=>"100011001",
  6481=>"100001001",
  6482=>"000101111",
  6483=>"110010000",
  6484=>"000111100",
  6485=>"100001110",
  6486=>"011111111",
  6487=>"100000110",
  6488=>"010001101",
  6489=>"101011110",
  6490=>"101101101",
  6491=>"011011000",
  6492=>"100101101",
  6493=>"001001110",
  6494=>"101100010",
  6495=>"011100110",
  6496=>"101001011",
  6497=>"001011110",
  6498=>"010000001",
  6499=>"000111111",
  6500=>"000000110",
  6501=>"111011011",
  6502=>"101111110",
  6503=>"101010101",
  6504=>"010010010",
  6505=>"111111011",
  6506=>"110000001",
  6507=>"001011001",
  6508=>"000001010",
  6509=>"000110101",
  6510=>"101010010",
  6511=>"000110101",
  6512=>"111110110",
  6513=>"101111101",
  6514=>"111101110",
  6515=>"010111000",
  6516=>"001111011",
  6517=>"101011101",
  6518=>"101001001",
  6519=>"011000010",
  6520=>"101100100",
  6521=>"111110011",
  6522=>"001111111",
  6523=>"001001001",
  6524=>"100000110",
  6525=>"100000000",
  6526=>"001100011",
  6527=>"110100101",
  6528=>"110100011",
  6529=>"000001001",
  6530=>"111000011",
  6531=>"001010000",
  6532=>"000000000",
  6533=>"100100000",
  6534=>"100001001",
  6535=>"000110110",
  6536=>"001010110",
  6537=>"111011011",
  6538=>"100110111",
  6539=>"000110000",
  6540=>"100101000",
  6541=>"011001011",
  6542=>"000010111",
  6543=>"000110110",
  6544=>"101100001",
  6545=>"010001011",
  6546=>"000011011",
  6547=>"100010101",
  6548=>"110001001",
  6549=>"100111000",
  6550=>"110001000",
  6551=>"000010000",
  6552=>"000101101",
  6553=>"001001001",
  6554=>"110000100",
  6555=>"101000100",
  6556=>"001011001",
  6557=>"100001101",
  6558=>"000011101",
  6559=>"110000111",
  6560=>"111011001",
  6561=>"000100110",
  6562=>"010000000",
  6563=>"100011101",
  6564=>"000100111",
  6565=>"100110001",
  6566=>"110101100",
  6567=>"110011110",
  6568=>"110111010",
  6569=>"111101000",
  6570=>"000000010",
  6571=>"001101110",
  6572=>"011101100",
  6573=>"010001001",
  6574=>"010011000",
  6575=>"101011001",
  6576=>"001000010",
  6577=>"001100000",
  6578=>"001001000",
  6579=>"111101001",
  6580=>"100011000",
  6581=>"000011011",
  6582=>"110111000",
  6583=>"100010111",
  6584=>"000001110",
  6585=>"011111111",
  6586=>"111100101",
  6587=>"011010000",
  6588=>"110110001",
  6589=>"110001000",
  6590=>"000111110",
  6591=>"011101010",
  6592=>"101011010",
  6593=>"111111110",
  6594=>"001110110",
  6595=>"110100101",
  6596=>"110010001",
  6597=>"001000101",
  6598=>"011000000",
  6599=>"010001111",
  6600=>"110110011",
  6601=>"010011000",
  6602=>"111100001",
  6603=>"000111010",
  6604=>"101011100",
  6605=>"101110000",
  6606=>"000011010",
  6607=>"100111100",
  6608=>"100010110",
  6609=>"011100001",
  6610=>"100001101",
  6611=>"101100001",
  6612=>"001100011",
  6613=>"011111101",
  6614=>"010101101",
  6615=>"100110001",
  6616=>"000011101",
  6617=>"010001101",
  6618=>"101011011",
  6619=>"110111010",
  6620=>"100110001",
  6621=>"111001001",
  6622=>"111000101",
  6623=>"000000110",
  6624=>"010110111",
  6625=>"110010100",
  6626=>"111101101",
  6627=>"000001110",
  6628=>"111111100",
  6629=>"110000111",
  6630=>"110010001",
  6631=>"111101010",
  6632=>"100010101",
  6633=>"000000010",
  6634=>"000011101",
  6635=>"100000111",
  6636=>"111000001",
  6637=>"011110001",
  6638=>"110010010",
  6639=>"101101011",
  6640=>"011000100",
  6641=>"001100010",
  6642=>"011110100",
  6643=>"111001000",
  6644=>"000101010",
  6645=>"001101000",
  6646=>"110101100",
  6647=>"001100001",
  6648=>"001001011",
  6649=>"001100100",
  6650=>"011101010",
  6651=>"000111000",
  6652=>"001001000",
  6653=>"110001101",
  6654=>"001010101",
  6655=>"001101101",
  6656=>"010010111",
  6657=>"101110011",
  6658=>"000001011",
  6659=>"101100100",
  6660=>"011000010",
  6661=>"100111001",
  6662=>"100101111",
  6663=>"000110101",
  6664=>"011010000",
  6665=>"110111001",
  6666=>"000111000",
  6667=>"110100101",
  6668=>"111001111",
  6669=>"011111011",
  6670=>"111001001",
  6671=>"000011100",
  6672=>"101011111",
  6673=>"110010010",
  6674=>"000100010",
  6675=>"111100101",
  6676=>"000000100",
  6677=>"011001110",
  6678=>"001010000",
  6679=>"001110010",
  6680=>"111111101",
  6681=>"011011000",
  6682=>"001000101",
  6683=>"111000110",
  6684=>"010000000",
  6685=>"100111110",
  6686=>"010010110",
  6687=>"011101001",
  6688=>"011110110",
  6689=>"000000011",
  6690=>"000011100",
  6691=>"011000001",
  6692=>"101111000",
  6693=>"001000000",
  6694=>"001011111",
  6695=>"010111000",
  6696=>"000011111",
  6697=>"101111101",
  6698=>"000000111",
  6699=>"010111011",
  6700=>"010001001",
  6701=>"011101010",
  6702=>"111001101",
  6703=>"010000010",
  6704=>"001000001",
  6705=>"001010001",
  6706=>"101010110",
  6707=>"110011101",
  6708=>"010010110",
  6709=>"000111100",
  6710=>"111100000",
  6711=>"110111101",
  6712=>"110001110",
  6713=>"101010011",
  6714=>"001011101",
  6715=>"111011011",
  6716=>"111001101",
  6717=>"001001101",
  6718=>"000110000",
  6719=>"000101010",
  6720=>"111010010",
  6721=>"100000000",
  6722=>"111110001",
  6723=>"001110110",
  6724=>"000010101",
  6725=>"001100100",
  6726=>"011001111",
  6727=>"000110100",
  6728=>"000101000",
  6729=>"010000101",
  6730=>"110000011",
  6731=>"000110001",
  6732=>"001101000",
  6733=>"000000011",
  6734=>"110001000",
  6735=>"010000001",
  6736=>"111101101",
  6737=>"111011001",
  6738=>"010000001",
  6739=>"001110010",
  6740=>"110110000",
  6741=>"100111110",
  6742=>"000111001",
  6743=>"001110000",
  6744=>"010010101",
  6745=>"111011100",
  6746=>"111101011",
  6747=>"010001000",
  6748=>"010000110",
  6749=>"111011101",
  6750=>"010111111",
  6751=>"011001010",
  6752=>"110111010",
  6753=>"011001111",
  6754=>"000110111",
  6755=>"110100101",
  6756=>"111010001",
  6757=>"001000000",
  6758=>"000111000",
  6759=>"000001001",
  6760=>"100010000",
  6761=>"101111111",
  6762=>"110011001",
  6763=>"001110100",
  6764=>"101000000",
  6765=>"100011111",
  6766=>"001100101",
  6767=>"000011011",
  6768=>"001111111",
  6769=>"111001110",
  6770=>"010010000",
  6771=>"001100101",
  6772=>"100000000",
  6773=>"000111011",
  6774=>"111100010",
  6775=>"111010001",
  6776=>"010100000",
  6777=>"001111101",
  6778=>"011101100",
  6779=>"111110111",
  6780=>"100110111",
  6781=>"010010100",
  6782=>"101101111",
  6783=>"000001001",
  6784=>"010000101",
  6785=>"100111011",
  6786=>"001110110",
  6787=>"011001111",
  6788=>"110101110",
  6789=>"100101010",
  6790=>"010101111",
  6791=>"010100010",
  6792=>"111101010",
  6793=>"111001001",
  6794=>"110111110",
  6795=>"011101111",
  6796=>"000000010",
  6797=>"001000100",
  6798=>"011001000",
  6799=>"110100011",
  6800=>"101001110",
  6801=>"000001010",
  6802=>"110011100",
  6803=>"111100011",
  6804=>"110010010",
  6805=>"010011110",
  6806=>"111100010",
  6807=>"000001100",
  6808=>"101001011",
  6809=>"000101110",
  6810=>"100100100",
  6811=>"000011001",
  6812=>"111001101",
  6813=>"111111101",
  6814=>"010000100",
  6815=>"001001100",
  6816=>"100110110",
  6817=>"010000000",
  6818=>"001110100",
  6819=>"001000110",
  6820=>"101111111",
  6821=>"100010010",
  6822=>"101001100",
  6823=>"101000101",
  6824=>"000001001",
  6825=>"110100001",
  6826=>"000000001",
  6827=>"000110010",
  6828=>"101100100",
  6829=>"010110100",
  6830=>"001101000",
  6831=>"000101011",
  6832=>"000101001",
  6833=>"000000000",
  6834=>"101010111",
  6835=>"101110101",
  6836=>"101111100",
  6837=>"001000010",
  6838=>"001000011",
  6839=>"000011110",
  6840=>"101011101",
  6841=>"010010010",
  6842=>"001101111",
  6843=>"000000111",
  6844=>"000010011",
  6845=>"001001100",
  6846=>"101100110",
  6847=>"011000100",
  6848=>"101110010",
  6849=>"010001100",
  6850=>"110001001",
  6851=>"100110101",
  6852=>"111110011",
  6853=>"000111101",
  6854=>"000010111",
  6855=>"000011010",
  6856=>"001110100",
  6857=>"010111101",
  6858=>"000100110",
  6859=>"110101000",
  6860=>"110001010",
  6861=>"010110110",
  6862=>"010100000",
  6863=>"110100000",
  6864=>"010110110",
  6865=>"111001101",
  6866=>"100111000",
  6867=>"011101111",
  6868=>"000000010",
  6869=>"111111100",
  6870=>"110010010",
  6871=>"010010011",
  6872=>"100000110",
  6873=>"011011111",
  6874=>"111101001",
  6875=>"111111110",
  6876=>"111011110",
  6877=>"110000101",
  6878=>"100110011",
  6879=>"101110111",
  6880=>"001100011",
  6881=>"101000010",
  6882=>"111011010",
  6883=>"010000010",
  6884=>"010000000",
  6885=>"010001111",
  6886=>"010000000",
  6887=>"111001100",
  6888=>"111011100",
  6889=>"001011111",
  6890=>"110110100",
  6891=>"101100011",
  6892=>"001011010",
  6893=>"111100001",
  6894=>"000010011",
  6895=>"000111110",
  6896=>"101001101",
  6897=>"100010000",
  6898=>"000101000",
  6899=>"110110111",
  6900=>"011000011",
  6901=>"110110001",
  6902=>"111101000",
  6903=>"000011110",
  6904=>"000111010",
  6905=>"000011110",
  6906=>"010111010",
  6907=>"111010010",
  6908=>"110100000",
  6909=>"101111010",
  6910=>"010101101",
  6911=>"111000001",
  6912=>"100100101",
  6913=>"001101111",
  6914=>"000000100",
  6915=>"000000011",
  6916=>"000010111",
  6917=>"100010010",
  6918=>"000110000",
  6919=>"100111101",
  6920=>"000101100",
  6921=>"010110010",
  6922=>"010011100",
  6923=>"010100011",
  6924=>"111001110",
  6925=>"011011000",
  6926=>"110100000",
  6927=>"100010010",
  6928=>"101011000",
  6929=>"101101001",
  6930=>"000000110",
  6931=>"010010100",
  6932=>"000111110",
  6933=>"011010010",
  6934=>"100110110",
  6935=>"000110110",
  6936=>"000111001",
  6937=>"000111000",
  6938=>"111010000",
  6939=>"100001110",
  6940=>"101111111",
  6941=>"110111111",
  6942=>"001101010",
  6943=>"101000111",
  6944=>"110101000",
  6945=>"110101010",
  6946=>"111110111",
  6947=>"111110110",
  6948=>"110000111",
  6949=>"111101110",
  6950=>"111010100",
  6951=>"100011100",
  6952=>"110010101",
  6953=>"000000011",
  6954=>"010111110",
  6955=>"000101101",
  6956=>"111100001",
  6957=>"000000010",
  6958=>"111101101",
  6959=>"000010010",
  6960=>"101110100",
  6961=>"000101000",
  6962=>"010111011",
  6963=>"010000111",
  6964=>"101010001",
  6965=>"011011010",
  6966=>"111011011",
  6967=>"010001100",
  6968=>"000010101",
  6969=>"100011110",
  6970=>"110010000",
  6971=>"001010110",
  6972=>"110100101",
  6973=>"000011110",
  6974=>"000010011",
  6975=>"100100111",
  6976=>"011010111",
  6977=>"111110001",
  6978=>"011010111",
  6979=>"101000000",
  6980=>"001011010",
  6981=>"101001000",
  6982=>"101011100",
  6983=>"000011111",
  6984=>"000110101",
  6985=>"000110010",
  6986=>"010010101",
  6987=>"011001111",
  6988=>"101100101",
  6989=>"000001011",
  6990=>"000010000",
  6991=>"011010100",
  6992=>"111110011",
  6993=>"000011101",
  6994=>"111101100",
  6995=>"000001110",
  6996=>"100011110",
  6997=>"111011010",
  6998=>"100011111",
  6999=>"001001010",
  7000=>"101000000",
  7001=>"111001000",
  7002=>"010111111",
  7003=>"101001001",
  7004=>"100001100",
  7005=>"110000011",
  7006=>"111101111",
  7007=>"100101011",
  7008=>"110000110",
  7009=>"010111000",
  7010=>"001100110",
  7011=>"111011100",
  7012=>"000000101",
  7013=>"000100000",
  7014=>"111110100",
  7015=>"111111100",
  7016=>"111101110",
  7017=>"011111000",
  7018=>"000110000",
  7019=>"000000110",
  7020=>"001011100",
  7021=>"111100101",
  7022=>"110011101",
  7023=>"101110110",
  7024=>"001111001",
  7025=>"111010101",
  7026=>"011111111",
  7027=>"010001010",
  7028=>"000010001",
  7029=>"111000000",
  7030=>"101011101",
  7031=>"000110000",
  7032=>"011000011",
  7033=>"101100111",
  7034=>"110000110",
  7035=>"110101111",
  7036=>"101011010",
  7037=>"111111101",
  7038=>"101101001",
  7039=>"111010110",
  7040=>"101110110",
  7041=>"000010011",
  7042=>"000000001",
  7043=>"001001010",
  7044=>"001100110",
  7045=>"000000000",
  7046=>"110000011",
  7047=>"001010000",
  7048=>"101110111",
  7049=>"110011101",
  7050=>"000101110",
  7051=>"100111000",
  7052=>"101001101",
  7053=>"011110111",
  7054=>"001010001",
  7055=>"100011001",
  7056=>"111111011",
  7057=>"000000110",
  7058=>"000011101",
  7059=>"001100101",
  7060=>"111111111",
  7061=>"011111011",
  7062=>"001110000",
  7063=>"000011100",
  7064=>"011010000",
  7065=>"011101101",
  7066=>"010110110",
  7067=>"010000001",
  7068=>"110110110",
  7069=>"000110011",
  7070=>"101110010",
  7071=>"010101101",
  7072=>"000000001",
  7073=>"110101011",
  7074=>"011010001",
  7075=>"110100101",
  7076=>"100010101",
  7077=>"100010000",
  7078=>"100111000",
  7079=>"010100100",
  7080=>"101011100",
  7081=>"110010000",
  7082=>"001000000",
  7083=>"001010101",
  7084=>"110010111",
  7085=>"100100111",
  7086=>"111010001",
  7087=>"011011100",
  7088=>"100110110",
  7089=>"101000000",
  7090=>"011001010",
  7091=>"111011000",
  7092=>"010110100",
  7093=>"001110001",
  7094=>"111000111",
  7095=>"000110101",
  7096=>"001111001",
  7097=>"101000000",
  7098=>"110001001",
  7099=>"101010100",
  7100=>"101011100",
  7101=>"110110101",
  7102=>"100011010",
  7103=>"010011000",
  7104=>"000011011",
  7105=>"101010010",
  7106=>"011011110",
  7107=>"111101011",
  7108=>"101111110",
  7109=>"110110000",
  7110=>"011111011",
  7111=>"100000100",
  7112=>"000010000",
  7113=>"100100010",
  7114=>"001101011",
  7115=>"000111001",
  7116=>"100101111",
  7117=>"011101101",
  7118=>"000010001",
  7119=>"111011110",
  7120=>"010000000",
  7121=>"100100010",
  7122=>"001010100",
  7123=>"101110110",
  7124=>"111011111",
  7125=>"011011001",
  7126=>"001010111",
  7127=>"001001111",
  7128=>"000110010",
  7129=>"100100110",
  7130=>"111100001",
  7131=>"110011010",
  7132=>"101111111",
  7133=>"011110000",
  7134=>"000000000",
  7135=>"010011100",
  7136=>"000011110",
  7137=>"000111110",
  7138=>"111101100",
  7139=>"011100100",
  7140=>"101101100",
  7141=>"001100010",
  7142=>"111111111",
  7143=>"110000110",
  7144=>"000001001",
  7145=>"011001000",
  7146=>"111000110",
  7147=>"111110011",
  7148=>"111011000",
  7149=>"000010001",
  7150=>"110101101",
  7151=>"010101111",
  7152=>"111101011",
  7153=>"111000001",
  7154=>"111010010",
  7155=>"010110110",
  7156=>"111000001",
  7157=>"001001000",
  7158=>"110000000",
  7159=>"111001000",
  7160=>"111100000",
  7161=>"011110011",
  7162=>"000110101",
  7163=>"100101110",
  7164=>"000010111",
  7165=>"001001000",
  7166=>"011011100",
  7167=>"011000110",
  7168=>"110110101",
  7169=>"111001100",
  7170=>"111110101",
  7171=>"010011111",
  7172=>"101011101",
  7173=>"010100010",
  7174=>"100110111",
  7175=>"010101110",
  7176=>"001110001",
  7177=>"000011000",
  7178=>"011010011",
  7179=>"000000111",
  7180=>"011000001",
  7181=>"110101101",
  7182=>"010010000",
  7183=>"000000100",
  7184=>"110111101",
  7185=>"100011110",
  7186=>"011101101",
  7187=>"100101110",
  7188=>"011000010",
  7189=>"001111000",
  7190=>"111111101",
  7191=>"010110101",
  7192=>"100100111",
  7193=>"101111110",
  7194=>"111000100",
  7195=>"110110111",
  7196=>"111001010",
  7197=>"101011100",
  7198=>"100010001",
  7199=>"101100010",
  7200=>"000101001",
  7201=>"011010000",
  7202=>"001001011",
  7203=>"111001011",
  7204=>"001101101",
  7205=>"111100010",
  7206=>"001011110",
  7207=>"001001011",
  7208=>"010111100",
  7209=>"110000011",
  7210=>"001011001",
  7211=>"101100001",
  7212=>"001001001",
  7213=>"010011100",
  7214=>"000011110",
  7215=>"011011101",
  7216=>"100100101",
  7217=>"000000000",
  7218=>"011011101",
  7219=>"101110011",
  7220=>"001001010",
  7221=>"011000010",
  7222=>"011110100",
  7223=>"001101011",
  7224=>"000111000",
  7225=>"111000010",
  7226=>"010010101",
  7227=>"110001111",
  7228=>"001001001",
  7229=>"101100110",
  7230=>"011001010",
  7231=>"000100111",
  7232=>"111010011",
  7233=>"001100101",
  7234=>"110100111",
  7235=>"010100110",
  7236=>"000011101",
  7237=>"001111101",
  7238=>"010001110",
  7239=>"010110011",
  7240=>"111010001",
  7241=>"001111000",
  7242=>"101000010",
  7243=>"000001010",
  7244=>"001100110",
  7245=>"101101100",
  7246=>"011110111",
  7247=>"111001011",
  7248=>"111101010",
  7249=>"111011001",
  7250=>"101011101",
  7251=>"011000100",
  7252=>"100101110",
  7253=>"101001011",
  7254=>"110111000",
  7255=>"010001111",
  7256=>"011101110",
  7257=>"010011001",
  7258=>"101111001",
  7259=>"101100001",
  7260=>"011101110",
  7261=>"000010011",
  7262=>"011100000",
  7263=>"111100011",
  7264=>"000110000",
  7265=>"111010011",
  7266=>"000101011",
  7267=>"100011111",
  7268=>"100011111",
  7269=>"000100111",
  7270=>"101101111",
  7271=>"000000000",
  7272=>"000100011",
  7273=>"111001011",
  7274=>"011110010",
  7275=>"101111001",
  7276=>"001110000",
  7277=>"010111000",
  7278=>"110000101",
  7279=>"001010000",
  7280=>"111110011",
  7281=>"000111111",
  7282=>"011110101",
  7283=>"100010011",
  7284=>"000001000",
  7285=>"110001011",
  7286=>"110111111",
  7287=>"001111010",
  7288=>"010010100",
  7289=>"010101001",
  7290=>"100001110",
  7291=>"001101010",
  7292=>"000011010",
  7293=>"010000000",
  7294=>"000010001",
  7295=>"100011010",
  7296=>"010101000",
  7297=>"111101000",
  7298=>"111010111",
  7299=>"001110110",
  7300=>"111100000",
  7301=>"101010101",
  7302=>"011101001",
  7303=>"110110000",
  7304=>"111101111",
  7305=>"110110000",
  7306=>"010000000",
  7307=>"010101100",
  7308=>"011010110",
  7309=>"101011111",
  7310=>"011000111",
  7311=>"001100110",
  7312=>"001011100",
  7313=>"011110100",
  7314=>"010001000",
  7315=>"110110101",
  7316=>"010110010",
  7317=>"100110101",
  7318=>"101111011",
  7319=>"111101001",
  7320=>"011000100",
  7321=>"000111111",
  7322=>"110001011",
  7323=>"001001110",
  7324=>"000100001",
  7325=>"101110100",
  7326=>"111000000",
  7327=>"100101010",
  7328=>"010011101",
  7329=>"111111101",
  7330=>"101001000",
  7331=>"101001100",
  7332=>"010000110",
  7333=>"000111001",
  7334=>"001000100",
  7335=>"011101001",
  7336=>"101000000",
  7337=>"110000010",
  7338=>"001111110",
  7339=>"011011111",
  7340=>"001010000",
  7341=>"100011000",
  7342=>"111011111",
  7343=>"111011110",
  7344=>"100001010",
  7345=>"010011010",
  7346=>"110001101",
  7347=>"111010000",
  7348=>"010110101",
  7349=>"101011101",
  7350=>"000010111",
  7351=>"010110100",
  7352=>"100110100",
  7353=>"011000001",
  7354=>"001001110",
  7355=>"111110010",
  7356=>"000111101",
  7357=>"100110100",
  7358=>"011110001",
  7359=>"100111011",
  7360=>"011100001",
  7361=>"010111000",
  7362=>"011000000",
  7363=>"110011000",
  7364=>"000010100",
  7365=>"111110101",
  7366=>"010001010",
  7367=>"011100010",
  7368=>"000010010",
  7369=>"000001110",
  7370=>"001110000",
  7371=>"100110000",
  7372=>"101110011",
  7373=>"011010111",
  7374=>"001100011",
  7375=>"001001000",
  7376=>"100001011",
  7377=>"011111100",
  7378=>"000010001",
  7379=>"011100000",
  7380=>"010011100",
  7381=>"101100110",
  7382=>"011100011",
  7383=>"110111010",
  7384=>"111100110",
  7385=>"101000101",
  7386=>"010100000",
  7387=>"100001011",
  7388=>"011010111",
  7389=>"010111010",
  7390=>"110111101",
  7391=>"000010011",
  7392=>"111010011",
  7393=>"000010111",
  7394=>"000110001",
  7395=>"001010100",
  7396=>"110111110",
  7397=>"001000011",
  7398=>"010000000",
  7399=>"100011000",
  7400=>"000000001",
  7401=>"110000001",
  7402=>"110101000",
  7403=>"100011000",
  7404=>"111101010",
  7405=>"001010111",
  7406=>"001010000",
  7407=>"011000000",
  7408=>"101011011",
  7409=>"010010010",
  7410=>"001101010",
  7411=>"010100010",
  7412=>"111000101",
  7413=>"011001111",
  7414=>"000110111",
  7415=>"111111011",
  7416=>"000111111",
  7417=>"010001101",
  7418=>"110111101",
  7419=>"101000101",
  7420=>"111001100",
  7421=>"100000111",
  7422=>"111100101",
  7423=>"111111111",
  7424=>"110000010",
  7425=>"010011111",
  7426=>"101001000",
  7427=>"100111011",
  7428=>"101010011",
  7429=>"111110101",
  7430=>"100110010",
  7431=>"110101011",
  7432=>"010010001",
  7433=>"001010010",
  7434=>"111011101",
  7435=>"111010001",
  7436=>"100111100",
  7437=>"110111000",
  7438=>"111110010",
  7439=>"000001000",
  7440=>"100011011",
  7441=>"011111010",
  7442=>"101100010",
  7443=>"110110100",
  7444=>"101011101",
  7445=>"111101111",
  7446=>"110010010",
  7447=>"000110110",
  7448=>"010001111",
  7449=>"110110010",
  7450=>"111101001",
  7451=>"111110111",
  7452=>"000000101",
  7453=>"011000001",
  7454=>"001100010",
  7455=>"110000101",
  7456=>"000101011",
  7457=>"111010011",
  7458=>"010110100",
  7459=>"000000001",
  7460=>"100100111",
  7461=>"110000101",
  7462=>"010000000",
  7463=>"110111100",
  7464=>"110110100",
  7465=>"001000011",
  7466=>"001101110",
  7467=>"110010000",
  7468=>"000011110",
  7469=>"011000101",
  7470=>"001101010",
  7471=>"001110010",
  7472=>"011001001",
  7473=>"100011101",
  7474=>"111111110",
  7475=>"100111100",
  7476=>"000100000",
  7477=>"100101011",
  7478=>"101001010",
  7479=>"001010010",
  7480=>"100101001",
  7481=>"001101011",
  7482=>"111010001",
  7483=>"000000100",
  7484=>"011000101",
  7485=>"100100010",
  7486=>"110110001",
  7487=>"010001000",
  7488=>"100001101",
  7489=>"111110000",
  7490=>"111110100",
  7491=>"011000010",
  7492=>"011000101",
  7493=>"000011000",
  7494=>"100000010",
  7495=>"001000101",
  7496=>"001101001",
  7497=>"010111011",
  7498=>"110111100",
  7499=>"000101001",
  7500=>"100011110",
  7501=>"000111111",
  7502=>"010011111",
  7503=>"010000010",
  7504=>"001000100",
  7505=>"000001011",
  7506=>"100110110",
  7507=>"000001011",
  7508=>"101100111",
  7509=>"100001011",
  7510=>"011110100",
  7511=>"010100111",
  7512=>"111101110",
  7513=>"111001111",
  7514=>"111010110",
  7515=>"100101010",
  7516=>"110110111",
  7517=>"000100010",
  7518=>"001100111",
  7519=>"101011000",
  7520=>"110110011",
  7521=>"110101001",
  7522=>"110001111",
  7523=>"001000101",
  7524=>"010110011",
  7525=>"011001110",
  7526=>"001001111",
  7527=>"100001101",
  7528=>"101011010",
  7529=>"110101101",
  7530=>"010001010",
  7531=>"100000011",
  7532=>"111000001",
  7533=>"111111010",
  7534=>"010011010",
  7535=>"101101100",
  7536=>"000100001",
  7537=>"001101110",
  7538=>"101111101",
  7539=>"101100011",
  7540=>"001000001",
  7541=>"100010110",
  7542=>"000000001",
  7543=>"001000001",
  7544=>"010010000",
  7545=>"100011111",
  7546=>"000010010",
  7547=>"010000000",
  7548=>"110010010",
  7549=>"010100100",
  7550=>"001011011",
  7551=>"000000101",
  7552=>"001111011",
  7553=>"000011010",
  7554=>"000111011",
  7555=>"000011000",
  7556=>"111110100",
  7557=>"110111010",
  7558=>"101110110",
  7559=>"000000010",
  7560=>"110000111",
  7561=>"001011000",
  7562=>"110100001",
  7563=>"100110000",
  7564=>"000000110",
  7565=>"110110010",
  7566=>"001001011",
  7567=>"101111100",
  7568=>"101111011",
  7569=>"010001001",
  7570=>"111101111",
  7571=>"011111111",
  7572=>"010001011",
  7573=>"101100011",
  7574=>"001000101",
  7575=>"110000100",
  7576=>"010010000",
  7577=>"110100001",
  7578=>"010010001",
  7579=>"111001010",
  7580=>"111001111",
  7581=>"101101100",
  7582=>"011111100",
  7583=>"011110111",
  7584=>"001101111",
  7585=>"000010101",
  7586=>"111100010",
  7587=>"000010100",
  7588=>"000011100",
  7589=>"011010100",
  7590=>"110000010",
  7591=>"010100100",
  7592=>"000000111",
  7593=>"000101110",
  7594=>"000011011",
  7595=>"100011100",
  7596=>"111011101",
  7597=>"101110100",
  7598=>"110001111",
  7599=>"011100101",
  7600=>"100111110",
  7601=>"100001010",
  7602=>"101010000",
  7603=>"100000011",
  7604=>"001001100",
  7605=>"011001001",
  7606=>"111010000",
  7607=>"111011001",
  7608=>"010001101",
  7609=>"000111101",
  7610=>"100100110",
  7611=>"110010010",
  7612=>"111100010",
  7613=>"110111111",
  7614=>"101111000",
  7615=>"110011101",
  7616=>"111001011",
  7617=>"000001101",
  7618=>"011100001",
  7619=>"000010000",
  7620=>"001100011",
  7621=>"101110111",
  7622=>"110100100",
  7623=>"000000001",
  7624=>"100001010",
  7625=>"101001011",
  7626=>"011010101",
  7627=>"111100110",
  7628=>"010100010",
  7629=>"100000011",
  7630=>"110011000",
  7631=>"001110101",
  7632=>"110010111",
  7633=>"101100001",
  7634=>"111101110",
  7635=>"101000100",
  7636=>"100111011",
  7637=>"110110010",
  7638=>"001111000",
  7639=>"110011110",
  7640=>"110111001",
  7641=>"010100010",
  7642=>"000000101",
  7643=>"001100000",
  7644=>"000110110",
  7645=>"110101011",
  7646=>"010000111",
  7647=>"001000110",
  7648=>"101001101",
  7649=>"101110110",
  7650=>"010110100",
  7651=>"110110101",
  7652=>"011001101",
  7653=>"010000101",
  7654=>"010110011",
  7655=>"100011000",
  7656=>"000110100",
  7657=>"100110101",
  7658=>"101111000",
  7659=>"101110101",
  7660=>"001101010",
  7661=>"011010010",
  7662=>"010001000",
  7663=>"000001011",
  7664=>"011100100",
  7665=>"110101010",
  7666=>"010111101",
  7667=>"110010000",
  7668=>"101010011",
  7669=>"000111100",
  7670=>"000100001",
  7671=>"000100000",
  7672=>"110010001",
  7673=>"101000101",
  7674=>"111110000",
  7675=>"001101100",
  7676=>"101101100",
  7677=>"111110011",
  7678=>"000101001",
  7679=>"110111011",
  7680=>"001001110",
  7681=>"110100011",
  7682=>"011001001",
  7683=>"110010100",
  7684=>"100101111",
  7685=>"100000010",
  7686=>"101010000",
  7687=>"100000010",
  7688=>"010011110",
  7689=>"100010110",
  7690=>"001000100",
  7691=>"110010000",
  7692=>"010100111",
  7693=>"011010000",
  7694=>"111100110",
  7695=>"110110111",
  7696=>"100100101",
  7697=>"000111011",
  7698=>"111100110",
  7699=>"111111111",
  7700=>"000001010",
  7701=>"100011111",
  7702=>"101010110",
  7703=>"010101010",
  7704=>"100010111",
  7705=>"111101110",
  7706=>"101111001",
  7707=>"010011100",
  7708=>"101010011",
  7709=>"000111110",
  7710=>"001100000",
  7711=>"100000110",
  7712=>"001000111",
  7713=>"001000101",
  7714=>"011010111",
  7715=>"110010001",
  7716=>"011011100",
  7717=>"010101011",
  7718=>"100010100",
  7719=>"000001111",
  7720=>"001001101",
  7721=>"110001100",
  7722=>"111101000",
  7723=>"111100001",
  7724=>"010011001",
  7725=>"000000010",
  7726=>"001000011",
  7727=>"101101101",
  7728=>"000000010",
  7729=>"100000110",
  7730=>"000010001",
  7731=>"000100110",
  7732=>"000000101",
  7733=>"000011111",
  7734=>"100000101",
  7735=>"010001101",
  7736=>"101000111",
  7737=>"101001011",
  7738=>"011111001",
  7739=>"110011001",
  7740=>"010011001",
  7741=>"110110101",
  7742=>"101100001",
  7743=>"011001000",
  7744=>"100000101",
  7745=>"100101010",
  7746=>"011000010",
  7747=>"101010101",
  7748=>"110001101",
  7749=>"001010001",
  7750=>"001101111",
  7751=>"100101010",
  7752=>"100000000",
  7753=>"101100000",
  7754=>"110101101",
  7755=>"000100110",
  7756=>"011101010",
  7757=>"000101111",
  7758=>"001100010",
  7759=>"101111000",
  7760=>"100010000",
  7761=>"010101101",
  7762=>"101101111",
  7763=>"001000001",
  7764=>"111001010",
  7765=>"110101001",
  7766=>"110001011",
  7767=>"000101000",
  7768=>"010001101",
  7769=>"001101010",
  7770=>"000101000",
  7771=>"011000011",
  7772=>"101100100",
  7773=>"101000000",
  7774=>"000011111",
  7775=>"100001011",
  7776=>"011100001",
  7777=>"111110100",
  7778=>"110100000",
  7779=>"111110001",
  7780=>"101011010",
  7781=>"001000101",
  7782=>"100101011",
  7783=>"001111111",
  7784=>"001101010",
  7785=>"101001000",
  7786=>"101010001",
  7787=>"101101011",
  7788=>"010111010",
  7789=>"010011000",
  7790=>"000000000",
  7791=>"011001110",
  7792=>"101001101",
  7793=>"011000100",
  7794=>"011010100",
  7795=>"010110010",
  7796=>"011110001",
  7797=>"110111110",
  7798=>"110000011",
  7799=>"011010000",
  7800=>"110001001",
  7801=>"011010110",
  7802=>"111011001",
  7803=>"100100100",
  7804=>"111010100",
  7805=>"011000000",
  7806=>"001101010",
  7807=>"010100010",
  7808=>"100100110",
  7809=>"001111011",
  7810=>"011011111",
  7811=>"110001110",
  7812=>"000101000",
  7813=>"001000001",
  7814=>"110011010",
  7815=>"101100101",
  7816=>"111101010",
  7817=>"111000000",
  7818=>"010100101",
  7819=>"100110000",
  7820=>"000000110",
  7821=>"101000001",
  7822=>"111110100",
  7823=>"101010111",
  7824=>"110010111",
  7825=>"110011011",
  7826=>"111110011",
  7827=>"001101010",
  7828=>"000010001",
  7829=>"001011110",
  7830=>"011000010",
  7831=>"111101011",
  7832=>"101100111",
  7833=>"011110000",
  7834=>"000110011",
  7835=>"000111111",
  7836=>"100001111",
  7837=>"111001011",
  7838=>"001001001",
  7839=>"110110001",
  7840=>"110010010",
  7841=>"001011110",
  7842=>"000000011",
  7843=>"111110100",
  7844=>"100110111",
  7845=>"101101001",
  7846=>"010010000",
  7847=>"010001000",
  7848=>"100100010",
  7849=>"001111110",
  7850=>"100000010",
  7851=>"011110000",
  7852=>"000001000",
  7853=>"101100001",
  7854=>"010110111",
  7855=>"110000011",
  7856=>"110100100",
  7857=>"011110010",
  7858=>"001000011",
  7859=>"110100001",
  7860=>"100001111",
  7861=>"100100011",
  7862=>"000111000",
  7863=>"011011010",
  7864=>"001100001",
  7865=>"010110110",
  7866=>"110001100",
  7867=>"110011111",
  7868=>"001000000",
  7869=>"000100101",
  7870=>"110001010",
  7871=>"101111011",
  7872=>"100110011",
  7873=>"111101110",
  7874=>"101000010",
  7875=>"001100101",
  7876=>"000101110",
  7877=>"000000111",
  7878=>"110101111",
  7879=>"101011101",
  7880=>"110001011",
  7881=>"000110010",
  7882=>"101111000",
  7883=>"100010111",
  7884=>"010001000",
  7885=>"001101011",
  7886=>"110100110",
  7887=>"111101010",
  7888=>"010100111",
  7889=>"000001000",
  7890=>"010110101",
  7891=>"001010110",
  7892=>"001110101",
  7893=>"100011111",
  7894=>"101010011",
  7895=>"011011001",
  7896=>"001000110",
  7897=>"001001110",
  7898=>"000000101",
  7899=>"110001010",
  7900=>"001111010",
  7901=>"011011100",
  7902=>"101110001",
  7903=>"010010101",
  7904=>"110111100",
  7905=>"101100000",
  7906=>"100100010",
  7907=>"010000100",
  7908=>"010101100",
  7909=>"010010111",
  7910=>"100111000",
  7911=>"110100001",
  7912=>"000001000",
  7913=>"100001100",
  7914=>"111110000",
  7915=>"111111111",
  7916=>"000000011",
  7917=>"010100001",
  7918=>"010101010",
  7919=>"100010111",
  7920=>"011000001",
  7921=>"110001010",
  7922=>"001010001",
  7923=>"111011000",
  7924=>"111110010",
  7925=>"100100110",
  7926=>"001010100",
  7927=>"010011100",
  7928=>"010101000",
  7929=>"100100000",
  7930=>"001001110",
  7931=>"111000111",
  7932=>"001010010",
  7933=>"111001110",
  7934=>"000010010",
  7935=>"000110100",
  7936=>"111111010",
  7937=>"001111011",
  7938=>"001100111",
  7939=>"110111100",
  7940=>"101110001",
  7941=>"001011100",
  7942=>"101111100",
  7943=>"100111110",
  7944=>"001010011",
  7945=>"000000001",
  7946=>"111101101",
  7947=>"001111010",
  7948=>"010010001",
  7949=>"101111010",
  7950=>"110001010",
  7951=>"101010010",
  7952=>"100011001",
  7953=>"000000010",
  7954=>"010001110",
  7955=>"010101010",
  7956=>"101101001",
  7957=>"011110111",
  7958=>"010001110",
  7959=>"011011100",
  7960=>"110101000",
  7961=>"110000100",
  7962=>"001111101",
  7963=>"100010010",
  7964=>"011110101",
  7965=>"011011111",
  7966=>"111001111",
  7967=>"110111101",
  7968=>"000001000",
  7969=>"100011100",
  7970=>"011010100",
  7971=>"101100111",
  7972=>"101000000",
  7973=>"010000100",
  7974=>"010010011",
  7975=>"000100100",
  7976=>"111010001",
  7977=>"111100001",
  7978=>"110111011",
  7979=>"000000101",
  7980=>"011001101",
  7981=>"000001010",
  7982=>"110101111",
  7983=>"101100111",
  7984=>"100111100",
  7985=>"100100110",
  7986=>"000101000",
  7987=>"110011101",
  7988=>"000101111",
  7989=>"000010101",
  7990=>"101111000",
  7991=>"111001011",
  7992=>"110011110",
  7993=>"110101001",
  7994=>"001101011",
  7995=>"001100011",
  7996=>"001000010",
  7997=>"000101101",
  7998=>"010111011",
  7999=>"000001111",
  8000=>"101111100",
  8001=>"001000100",
  8002=>"101010110",
  8003=>"111010111",
  8004=>"010110000",
  8005=>"100111100",
  8006=>"110011011",
  8007=>"101111011",
  8008=>"011101001",
  8009=>"101111100",
  8010=>"001111101",
  8011=>"100010100",
  8012=>"101001111",
  8013=>"110110000",
  8014=>"011110001",
  8015=>"000111100",
  8016=>"101110100",
  8017=>"010010110",
  8018=>"010101001",
  8019=>"111100101",
  8020=>"010001000",
  8021=>"111010101",
  8022=>"011011011",
  8023=>"000011000",
  8024=>"011100011",
  8025=>"100011110",
  8026=>"001000100",
  8027=>"111010011",
  8028=>"010110110",
  8029=>"010100010",
  8030=>"111101111",
  8031=>"100000000",
  8032=>"000001000",
  8033=>"010100001",
  8034=>"100001111",
  8035=>"010011010",
  8036=>"000000110",
  8037=>"000001110",
  8038=>"010011101",
  8039=>"001111000",
  8040=>"101100000",
  8041=>"000011001",
  8042=>"111100000",
  8043=>"001011010",
  8044=>"011110000",
  8045=>"110110101",
  8046=>"011001100",
  8047=>"111001001",
  8048=>"001101101",
  8049=>"010011101",
  8050=>"100110110",
  8051=>"010101110",
  8052=>"010001001",
  8053=>"001101001",
  8054=>"010110010",
  8055=>"010000010",
  8056=>"101001100",
  8057=>"110111001",
  8058=>"011111011",
  8059=>"010111010",
  8060=>"010101001",
  8061=>"100011010",
  8062=>"100111001",
  8063=>"100100001",
  8064=>"001110100",
  8065=>"111111001",
  8066=>"101001100",
  8067=>"110110110",
  8068=>"111100101",
  8069=>"101000101",
  8070=>"100110110",
  8071=>"001000011",
  8072=>"100010011",
  8073=>"111111000",
  8074=>"001100000",
  8075=>"101110110",
  8076=>"101011110",
  8077=>"101011111",
  8078=>"100001111",
  8079=>"010000110",
  8080=>"001101001",
  8081=>"100100101",
  8082=>"100000111",
  8083=>"100111111",
  8084=>"100000001",
  8085=>"101001010",
  8086=>"110101001",
  8087=>"101111011",
  8088=>"101011100",
  8089=>"010111100",
  8090=>"101001000",
  8091=>"100011011",
  8092=>"111000111",
  8093=>"111101000",
  8094=>"110000010",
  8095=>"010110000",
  8096=>"010000100",
  8097=>"101110001",
  8098=>"110110110",
  8099=>"000010100",
  8100=>"110010110",
  8101=>"011101000",
  8102=>"001000101",
  8103=>"101011101",
  8104=>"010010111",
  8105=>"011001010",
  8106=>"001101111",
  8107=>"101011111",
  8108=>"100000110",
  8109=>"111000101",
  8110=>"110111010",
  8111=>"010000111",
  8112=>"111101101",
  8113=>"101011101",
  8114=>"010100100",
  8115=>"111000000",
  8116=>"101101111",
  8117=>"010111010",
  8118=>"000110101",
  8119=>"101010111",
  8120=>"111001001",
  8121=>"011001111",
  8122=>"101000110",
  8123=>"011101011",
  8124=>"110101001",
  8125=>"000100110",
  8126=>"100101000",
  8127=>"001101001",
  8128=>"101110000",
  8129=>"001110111",
  8130=>"100101001",
  8131=>"101000011",
  8132=>"010100111",
  8133=>"000100011",
  8134=>"111110100",
  8135=>"111101011",
  8136=>"111010000",
  8137=>"111001000",
  8138=>"111110110",
  8139=>"010111010",
  8140=>"100101110",
  8141=>"001010011",
  8142=>"000100011",
  8143=>"001111110",
  8144=>"001101001",
  8145=>"000011011",
  8146=>"101001101",
  8147=>"110101001",
  8148=>"110001001",
  8149=>"010110001",
  8150=>"011111010",
  8151=>"101111011",
  8152=>"100101011",
  8153=>"001011110",
  8154=>"010010001",
  8155=>"111011101",
  8156=>"001110011",
  8157=>"111100110",
  8158=>"110110001",
  8159=>"010101110",
  8160=>"100100010",
  8161=>"000001011",
  8162=>"010010010",
  8163=>"100000111",
  8164=>"011100000",
  8165=>"111011111",
  8166=>"000001111",
  8167=>"010011110",
  8168=>"101110100",
  8169=>"010110001",
  8170=>"101000110",
  8171=>"101101111",
  8172=>"101110100",
  8173=>"001100111",
  8174=>"100110110",
  8175=>"011111000",
  8176=>"000101001",
  8177=>"110010010",
  8178=>"001001000",
  8179=>"111010110",
  8180=>"101111100",
  8181=>"010110101",
  8182=>"001100100",
  8183=>"101110100",
  8184=>"011100111",
  8185=>"000101110",
  8186=>"111010000",
  8187=>"010010111",
  8188=>"010010110",
  8189=>"000001101",
  8190=>"011001101",
  8191=>"001110010",
  8192=>"011000000",
  8193=>"010001011",
  8194=>"010011110",
  8195=>"011001101",
  8196=>"010100100",
  8197=>"011001000",
  8198=>"011011011",
  8199=>"000110000",
  8200=>"001011010",
  8201=>"101000111",
  8202=>"101001001",
  8203=>"001100111",
  8204=>"101111101",
  8205=>"101101010",
  8206=>"100011000",
  8207=>"101011111",
  8208=>"001001110",
  8209=>"100100001",
  8210=>"010001110",
  8211=>"101010010",
  8212=>"010000110",
  8213=>"011010010",
  8214=>"111000011",
  8215=>"001110100",
  8216=>"001101000",
  8217=>"101010000",
  8218=>"000011111",
  8219=>"011111010",
  8220=>"111011101",
  8221=>"010100100",
  8222=>"001100110",
  8223=>"100011100",
  8224=>"100101111",
  8225=>"011000000",
  8226=>"110000000",
  8227=>"011111101",
  8228=>"111000110",
  8229=>"111110001",
  8230=>"100111000",
  8231=>"111101011",
  8232=>"100000110",
  8233=>"110101001",
  8234=>"001000010",
  8235=>"101011111",
  8236=>"010011000",
  8237=>"010111111",
  8238=>"111001011",
  8239=>"010111110",
  8240=>"101110000",
  8241=>"100100011",
  8242=>"001000101",
  8243=>"101010111",
  8244=>"111000101",
  8245=>"011011100",
  8246=>"001011100",
  8247=>"110111101",
  8248=>"101101011",
  8249=>"011111011",
  8250=>"111001111",
  8251=>"010110111",
  8252=>"011000010",
  8253=>"010110100",
  8254=>"100011010",
  8255=>"010000100",
  8256=>"001011000",
  8257=>"000000110",
  8258=>"001001101",
  8259=>"100101110",
  8260=>"001110100",
  8261=>"111101100",
  8262=>"001111000",
  8263=>"010000001",
  8264=>"110101001",
  8265=>"110100110",
  8266=>"111111001",
  8267=>"110001000",
  8268=>"001000010",
  8269=>"000011111",
  8270=>"010101111",
  8271=>"100001011",
  8272=>"100001011",
  8273=>"001000001",
  8274=>"100110101",
  8275=>"001111000",
  8276=>"101111010",
  8277=>"110010100",
  8278=>"000000000",
  8279=>"100101110",
  8280=>"010001010",
  8281=>"101111110",
  8282=>"100011001",
  8283=>"111010011",
  8284=>"011101110",
  8285=>"111110011",
  8286=>"110111000",
  8287=>"100111011",
  8288=>"000011010",
  8289=>"111011000",
  8290=>"111011001",
  8291=>"010000010",
  8292=>"000010001",
  8293=>"110000111",
  8294=>"100001110",
  8295=>"100001111",
  8296=>"110001110",
  8297=>"100100010",
  8298=>"010101001",
  8299=>"110111100",
  8300=>"011110010",
  8301=>"011110001",
  8302=>"010110101",
  8303=>"101111011",
  8304=>"110100100",
  8305=>"101011100",
  8306=>"100011000",
  8307=>"110001101",
  8308=>"001111001",
  8309=>"110010101",
  8310=>"110111110",
  8311=>"111101111",
  8312=>"001000000",
  8313=>"110101100",
  8314=>"100000110",
  8315=>"110010000",
  8316=>"001101011",
  8317=>"110010010",
  8318=>"000101000",
  8319=>"111000110",
  8320=>"000001000",
  8321=>"111000010",
  8322=>"101101010",
  8323=>"000010000",
  8324=>"010001110",
  8325=>"001000010",
  8326=>"011110001",
  8327=>"100100101",
  8328=>"111110101",
  8329=>"000010101",
  8330=>"010100111",
  8331=>"000000001",
  8332=>"111000101",
  8333=>"100101101",
  8334=>"010110000",
  8335=>"101011100",
  8336=>"011001001",
  8337=>"111010010",
  8338=>"000011010",
  8339=>"110110010",
  8340=>"010110101",
  8341=>"101001010",
  8342=>"000011111",
  8343=>"110000101",
  8344=>"110110011",
  8345=>"011111111",
  8346=>"111001110",
  8347=>"000101011",
  8348=>"010000111",
  8349=>"000100110",
  8350=>"000101111",
  8351=>"010000110",
  8352=>"111100110",
  8353=>"110101110",
  8354=>"001110100",
  8355=>"111010100",
  8356=>"010011100",
  8357=>"001010110",
  8358=>"110101100",
  8359=>"101000110",
  8360=>"000011011",
  8361=>"101100111",
  8362=>"100001110",
  8363=>"000011000",
  8364=>"010010100",
  8365=>"100111100",
  8366=>"111111001",
  8367=>"100100101",
  8368=>"000110010",
  8369=>"111100100",
  8370=>"100001110",
  8371=>"110100110",
  8372=>"001010111",
  8373=>"010111111",
  8374=>"010000100",
  8375=>"110110100",
  8376=>"000101110",
  8377=>"010100101",
  8378=>"011001001",
  8379=>"101101100",
  8380=>"110000100",
  8381=>"110010001",
  8382=>"100100110",
  8383=>"110100011",
  8384=>"001101011",
  8385=>"111101101",
  8386=>"010101000",
  8387=>"100000001",
  8388=>"100110101",
  8389=>"001111101",
  8390=>"000100101",
  8391=>"101001011",
  8392=>"110011000",
  8393=>"101111110",
  8394=>"110111011",
  8395=>"001010100",
  8396=>"101111000",
  8397=>"111010100",
  8398=>"010100101",
  8399=>"010100001",
  8400=>"110001011",
  8401=>"101100000",
  8402=>"001010011",
  8403=>"100001100",
  8404=>"011100001",
  8405=>"100001110",
  8406=>"000010100",
  8407=>"011000011",
  8408=>"101001100",
  8409=>"000000011",
  8410=>"000101100",
  8411=>"000100101",
  8412=>"100100010",
  8413=>"100111110",
  8414=>"100111101",
  8415=>"111100100",
  8416=>"110000111",
  8417=>"000001000",
  8418=>"111111000",
  8419=>"011110111",
  8420=>"000110011",
  8421=>"011110111",
  8422=>"011111000",
  8423=>"100011001",
  8424=>"010010100",
  8425=>"011111110",
  8426=>"111110010",
  8427=>"101000100",
  8428=>"010100010",
  8429=>"110000111",
  8430=>"001001111",
  8431=>"101111001",
  8432=>"001001100",
  8433=>"101100111",
  8434=>"000000010",
  8435=>"100100000",
  8436=>"001011101",
  8437=>"001111111",
  8438=>"011011010",
  8439=>"101000111",
  8440=>"101111001",
  8441=>"010000001",
  8442=>"111101101",
  8443=>"100011010",
  8444=>"000000110",
  8445=>"111111011",
  8446=>"101111100",
  8447=>"011111000",
  8448=>"100101001",
  8449=>"110001110",
  8450=>"111101111",
  8451=>"100000110",
  8452=>"011011100",
  8453=>"010101000",
  8454=>"100000100",
  8455=>"111001101",
  8456=>"111101111",
  8457=>"000100110",
  8458=>"001100010",
  8459=>"011101111",
  8460=>"011100100",
  8461=>"001000110",
  8462=>"000100000",
  8463=>"010001110",
  8464=>"111101101",
  8465=>"101101000",
  8466=>"110110010",
  8467=>"010100000",
  8468=>"111101100",
  8469=>"100111111",
  8470=>"000101100",
  8471=>"000000011",
  8472=>"110010100",
  8473=>"100011100",
  8474=>"000000110",
  8475=>"010111101",
  8476=>"010111010",
  8477=>"101100101",
  8478=>"110000110",
  8479=>"010010001",
  8480=>"001011001",
  8481=>"001101001",
  8482=>"010001011",
  8483=>"101000100",
  8484=>"111011010",
  8485=>"010100011",
  8486=>"011111111",
  8487=>"111011100",
  8488=>"101001001",
  8489=>"110110011",
  8490=>"101011000",
  8491=>"001100100",
  8492=>"111000001",
  8493=>"000010000",
  8494=>"101001001",
  8495=>"101111010",
  8496=>"000111010",
  8497=>"111111000",
  8498=>"000111110",
  8499=>"001011110",
  8500=>"010110001",
  8501=>"111010011",
  8502=>"010011100",
  8503=>"111101001",
  8504=>"000100101",
  8505=>"111110000",
  8506=>"010110001",
  8507=>"111111000",
  8508=>"011000100",
  8509=>"110110011",
  8510=>"110011110",
  8511=>"111010001",
  8512=>"111011001",
  8513=>"010101111",
  8514=>"111100100",
  8515=>"100010010",
  8516=>"100101100",
  8517=>"101010111",
  8518=>"000110100",
  8519=>"110110001",
  8520=>"011100111",
  8521=>"110110110",
  8522=>"011110101",
  8523=>"001100111",
  8524=>"100110110",
  8525=>"001110001",
  8526=>"111101101",
  8527=>"010010100",
  8528=>"001010101",
  8529=>"000000110",
  8530=>"100010011",
  8531=>"110110111",
  8532=>"010100000",
  8533=>"001110111",
  8534=>"000110111",
  8535=>"000110110",
  8536=>"010010000",
  8537=>"001000101",
  8538=>"110001110",
  8539=>"001010100",
  8540=>"111101100",
  8541=>"100010100",
  8542=>"100001010",
  8543=>"111010100",
  8544=>"101011001",
  8545=>"001110010",
  8546=>"000011011",
  8547=>"101100001",
  8548=>"010000100",
  8549=>"111111101",
  8550=>"001110110",
  8551=>"111111111",
  8552=>"011010101",
  8553=>"001100111",
  8554=>"100001000",
  8555=>"101010010",
  8556=>"111011010",
  8557=>"000111101",
  8558=>"101011000",
  8559=>"100111011",
  8560=>"000001101",
  8561=>"101100110",
  8562=>"110100000",
  8563=>"010110001",
  8564=>"111110101",
  8565=>"000000100",
  8566=>"011110110",
  8567=>"110111010",
  8568=>"000011100",
  8569=>"001100010",
  8570=>"011001010",
  8571=>"000110011",
  8572=>"110110101",
  8573=>"111111111",
  8574=>"011110101",
  8575=>"000100010",
  8576=>"111010001",
  8577=>"001110000",
  8578=>"001000100",
  8579=>"100011100",
  8580=>"101111000",
  8581=>"111101101",
  8582=>"110001000",
  8583=>"000000011",
  8584=>"000011111",
  8585=>"001000001",
  8586=>"100110101",
  8587=>"001001011",
  8588=>"100001001",
  8589=>"001010011",
  8590=>"100000011",
  8591=>"010111100",
  8592=>"001010100",
  8593=>"001000001",
  8594=>"110110001",
  8595=>"000011010",
  8596=>"111110010",
  8597=>"010001001",
  8598=>"010010110",
  8599=>"111000111",
  8600=>"100001010",
  8601=>"011100010",
  8602=>"001100011",
  8603=>"010110010",
  8604=>"111001010",
  8605=>"101110101",
  8606=>"110001101",
  8607=>"000000000",
  8608=>"100010001",
  8609=>"111010000",
  8610=>"010100110",
  8611=>"111110100",
  8612=>"001010111",
  8613=>"010011110",
  8614=>"101001011",
  8615=>"010011100",
  8616=>"011011011",
  8617=>"000001100",
  8618=>"000110100",
  8619=>"000001001",
  8620=>"110110110",
  8621=>"011110010",
  8622=>"100110110",
  8623=>"101100101",
  8624=>"100010000",
  8625=>"010001110",
  8626=>"111100011",
  8627=>"111000011",
  8628=>"110111100",
  8629=>"111111010",
  8630=>"101111111",
  8631=>"111110100",
  8632=>"101011010",
  8633=>"100100111",
  8634=>"000000111",
  8635=>"011111011",
  8636=>"100011011",
  8637=>"001011011",
  8638=>"011001100",
  8639=>"110011110",
  8640=>"011000100",
  8641=>"000011010",
  8642=>"110010101",
  8643=>"010000000",
  8644=>"110001110",
  8645=>"110100011",
  8646=>"001001010",
  8647=>"101111111",
  8648=>"100010010",
  8649=>"000010011",
  8650=>"000010100",
  8651=>"001011011",
  8652=>"001111110",
  8653=>"001111010",
  8654=>"111111110",
  8655=>"100110010",
  8656=>"111000010",
  8657=>"000111011",
  8658=>"000101111",
  8659=>"011011011",
  8660=>"001101110",
  8661=>"011100010",
  8662=>"010010001",
  8663=>"101011000",
  8664=>"111101101",
  8665=>"011110000",
  8666=>"001001011",
  8667=>"010000000",
  8668=>"100001000",
  8669=>"001010110",
  8670=>"101000011",
  8671=>"001101110",
  8672=>"011100001",
  8673=>"011101000",
  8674=>"111110001",
  8675=>"010100010",
  8676=>"001110000",
  8677=>"001011100",
  8678=>"001111011",
  8679=>"101000100",
  8680=>"010110011",
  8681=>"000010001",
  8682=>"101111110",
  8683=>"010111100",
  8684=>"111110101",
  8685=>"011100101",
  8686=>"001010100",
  8687=>"100110110",
  8688=>"000001000",
  8689=>"011001010",
  8690=>"100101010",
  8691=>"110000001",
  8692=>"001100011",
  8693=>"011001101",
  8694=>"011101101",
  8695=>"011000100",
  8696=>"001010111",
  8697=>"011000100",
  8698=>"000001000",
  8699=>"001110111",
  8700=>"000110010",
  8701=>"110000001",
  8702=>"101111001",
  8703=>"101001101",
  8704=>"110111110",
  8705=>"100011011",
  8706=>"001111000",
  8707=>"010101100",
  8708=>"110111001",
  8709=>"000001101",
  8710=>"111110011",
  8711=>"101001100",
  8712=>"100001100",
  8713=>"011100010",
  8714=>"011110101",
  8715=>"011100010",
  8716=>"001010000",
  8717=>"001101010",
  8718=>"110010111",
  8719=>"111011100",
  8720=>"001111100",
  8721=>"001010110",
  8722=>"011010111",
  8723=>"111010001",
  8724=>"011001001",
  8725=>"111110111",
  8726=>"100101100",
  8727=>"111011101",
  8728=>"101110011",
  8729=>"000100111",
  8730=>"101010100",
  8731=>"000101110",
  8732=>"110000111",
  8733=>"110011011",
  8734=>"111100111",
  8735=>"010110110",
  8736=>"000000101",
  8737=>"011101101",
  8738=>"101000101",
  8739=>"101011001",
  8740=>"110111110",
  8741=>"010010111",
  8742=>"001010101",
  8743=>"001001111",
  8744=>"000111110",
  8745=>"010010000",
  8746=>"010000010",
  8747=>"110001110",
  8748=>"010101101",
  8749=>"000000110",
  8750=>"110001111",
  8751=>"001110110",
  8752=>"010101010",
  8753=>"111110111",
  8754=>"000011100",
  8755=>"110000110",
  8756=>"000011000",
  8757=>"000110011",
  8758=>"100000000",
  8759=>"110100011",
  8760=>"110001100",
  8761=>"101110110",
  8762=>"101001011",
  8763=>"101010001",
  8764=>"001100111",
  8765=>"111100110",
  8766=>"000000110",
  8767=>"010001100",
  8768=>"010001000",
  8769=>"010101000",
  8770=>"100101000",
  8771=>"011010011",
  8772=>"010101110",
  8773=>"001101110",
  8774=>"100000101",
  8775=>"001100100",
  8776=>"010111001",
  8777=>"001001001",
  8778=>"001001010",
  8779=>"000101011",
  8780=>"110010010",
  8781=>"101111001",
  8782=>"100101001",
  8783=>"101001110",
  8784=>"110000101",
  8785=>"101000101",
  8786=>"100101010",
  8787=>"100000000",
  8788=>"000011011",
  8789=>"110100000",
  8790=>"011111011",
  8791=>"010101010",
  8792=>"110001001",
  8793=>"110000011",
  8794=>"011001111",
  8795=>"110000101",
  8796=>"110111100",
  8797=>"101001000",
  8798=>"001001101",
  8799=>"001001010",
  8800=>"011001000",
  8801=>"010010110",
  8802=>"000001010",
  8803=>"011101010",
  8804=>"010111101",
  8805=>"100010101",
  8806=>"000010001",
  8807=>"010001101",
  8808=>"111001000",
  8809=>"000011100",
  8810=>"011010010",
  8811=>"010101100",
  8812=>"000010101",
  8813=>"111000000",
  8814=>"110111101",
  8815=>"110011010",
  8816=>"000010001",
  8817=>"000110000",
  8818=>"101110111",
  8819=>"001101111",
  8820=>"010100100",
  8821=>"011100000",
  8822=>"100010110",
  8823=>"110111110",
  8824=>"110011010",
  8825=>"111101111",
  8826=>"101001111",
  8827=>"000101001",
  8828=>"010000110",
  8829=>"011000010",
  8830=>"010111001",
  8831=>"110110001",
  8832=>"000100010",
  8833=>"100001110",
  8834=>"011110010",
  8835=>"110001111",
  8836=>"100001101",
  8837=>"010010111",
  8838=>"001010111",
  8839=>"010111011",
  8840=>"100110110",
  8841=>"001011101",
  8842=>"111100111",
  8843=>"101100010",
  8844=>"010011011",
  8845=>"001101011",
  8846=>"011010100",
  8847=>"110000111",
  8848=>"011100111",
  8849=>"111101110",
  8850=>"101001101",
  8851=>"110100100",
  8852=>"010100100",
  8853=>"011100010",
  8854=>"001111010",
  8855=>"100100111",
  8856=>"111010000",
  8857=>"110110111",
  8858=>"110100110",
  8859=>"110011010",
  8860=>"010100000",
  8861=>"001010001",
  8862=>"111010101",
  8863=>"101001100",
  8864=>"000010111",
  8865=>"000100011",
  8866=>"110100001",
  8867=>"100111000",
  8868=>"110101100",
  8869=>"111100101",
  8870=>"000100000",
  8871=>"100010100",
  8872=>"111010001",
  8873=>"001000000",
  8874=>"001000111",
  8875=>"101001000",
  8876=>"100010000",
  8877=>"111010000",
  8878=>"010111100",
  8879=>"111111011",
  8880=>"011011000",
  8881=>"000110010",
  8882=>"100001111",
  8883=>"000011100",
  8884=>"001101000",
  8885=>"000101111",
  8886=>"001001000",
  8887=>"000011000",
  8888=>"010101111",
  8889=>"011100000",
  8890=>"000100010",
  8891=>"101100010",
  8892=>"110101101",
  8893=>"110010101",
  8894=>"011100001",
  8895=>"111111111",
  8896=>"101110101",
  8897=>"000011111",
  8898=>"010011001",
  8899=>"100010111",
  8900=>"000010011",
  8901=>"110010001",
  8902=>"101011111",
  8903=>"010101001",
  8904=>"011000100",
  8905=>"100001010",
  8906=>"001001111",
  8907=>"000011001",
  8908=>"110110010",
  8909=>"101100110",
  8910=>"101010110",
  8911=>"001010011",
  8912=>"000111110",
  8913=>"101000011",
  8914=>"101111011",
  8915=>"010000111",
  8916=>"001100110",
  8917=>"010000100",
  8918=>"011100100",
  8919=>"010011101",
  8920=>"010101101",
  8921=>"101111111",
  8922=>"110011111",
  8923=>"010110000",
  8924=>"101101100",
  8925=>"111110101",
  8926=>"110101010",
  8927=>"010011100",
  8928=>"010110110",
  8929=>"100100100",
  8930=>"100000110",
  8931=>"010000001",
  8932=>"110001100",
  8933=>"100011101",
  8934=>"011000111",
  8935=>"011001110",
  8936=>"000100010",
  8937=>"111110100",
  8938=>"101101101",
  8939=>"000111100",
  8940=>"001000110",
  8941=>"101000110",
  8942=>"110110101",
  8943=>"100110100",
  8944=>"001101100",
  8945=>"101001010",
  8946=>"011000000",
  8947=>"111001101",
  8948=>"111111101",
  8949=>"000010000",
  8950=>"100100001",
  8951=>"001111011",
  8952=>"001001111",
  8953=>"111010110",
  8954=>"011110110",
  8955=>"101011111",
  8956=>"111101110",
  8957=>"101000100",
  8958=>"011000101",
  8959=>"100100010",
  8960=>"111110010",
  8961=>"000110110",
  8962=>"110011101",
  8963=>"100011000",
  8964=>"001000100",
  8965=>"101011100",
  8966=>"000001100",
  8967=>"101011000",
  8968=>"011011001",
  8969=>"010110000",
  8970=>"110011110",
  8971=>"110000010",
  8972=>"000101010",
  8973=>"011101010",
  8974=>"011100011",
  8975=>"000010110",
  8976=>"100001101",
  8977=>"100101100",
  8978=>"001101010",
  8979=>"110000001",
  8980=>"101110011",
  8981=>"101100100",
  8982=>"000101101",
  8983=>"110100110",
  8984=>"111100010",
  8985=>"001010100",
  8986=>"001001011",
  8987=>"101100110",
  8988=>"101000001",
  8989=>"111000001",
  8990=>"110001001",
  8991=>"101100011",
  8992=>"000000110",
  8993=>"001100101",
  8994=>"001011110",
  8995=>"111000000",
  8996=>"100000100",
  8997=>"111000011",
  8998=>"001000011",
  8999=>"001101101",
  9000=>"111011110",
  9001=>"011110101",
  9002=>"001101011",
  9003=>"010011010",
  9004=>"010111111",
  9005=>"000001010",
  9006=>"000011010",
  9007=>"111000010",
  9008=>"001000100",
  9009=>"110110010",
  9010=>"110110100",
  9011=>"011100100",
  9012=>"101011111",
  9013=>"010011011",
  9014=>"000011000",
  9015=>"000110010",
  9016=>"000001010",
  9017=>"001000000",
  9018=>"010000110",
  9019=>"110010000",
  9020=>"001110101",
  9021=>"001010111",
  9022=>"000000001",
  9023=>"011000110",
  9024=>"000101110",
  9025=>"100001110",
  9026=>"011101100",
  9027=>"001000111",
  9028=>"000100111",
  9029=>"001101101",
  9030=>"100100100",
  9031=>"100101111",
  9032=>"010111110",
  9033=>"000001011",
  9034=>"000100011",
  9035=>"010110001",
  9036=>"110101001",
  9037=>"111100101",
  9038=>"001110000",
  9039=>"001001001",
  9040=>"010011000",
  9041=>"000100111",
  9042=>"100000111",
  9043=>"110011100",
  9044=>"100111111",
  9045=>"001001100",
  9046=>"110101111",
  9047=>"000100010",
  9048=>"100110100",
  9049=>"111011111",
  9050=>"000110100",
  9051=>"000101101",
  9052=>"111001100",
  9053=>"000100001",
  9054=>"000101100",
  9055=>"100001110",
  9056=>"100101000",
  9057=>"111101100",
  9058=>"101110001",
  9059=>"110111011",
  9060=>"110001110",
  9061=>"110100000",
  9062=>"000100011",
  9063=>"001010110",
  9064=>"110100011",
  9065=>"001001110",
  9066=>"001010101",
  9067=>"011100000",
  9068=>"000110100",
  9069=>"000100101",
  9070=>"010001010",
  9071=>"001101101",
  9072=>"101001111",
  9073=>"100111011",
  9074=>"101001001",
  9075=>"010111011",
  9076=>"000100100",
  9077=>"010000010",
  9078=>"011000010",
  9079=>"100101000",
  9080=>"111100101",
  9081=>"010100001",
  9082=>"000101101",
  9083=>"001011000",
  9084=>"011111101",
  9085=>"101010100",
  9086=>"111011011",
  9087=>"100111010",
  9088=>"110010100",
  9089=>"110000110",
  9090=>"100001100",
  9091=>"001101100",
  9092=>"000010101",
  9093=>"101110001",
  9094=>"000011000",
  9095=>"100011100",
  9096=>"111010011",
  9097=>"110110100",
  9098=>"110111010",
  9099=>"110010010",
  9100=>"101011111",
  9101=>"011001110",
  9102=>"001101011",
  9103=>"011001011",
  9104=>"100001110",
  9105=>"000010101",
  9106=>"100110110",
  9107=>"100010111",
  9108=>"110111000",
  9109=>"111001101",
  9110=>"011101100",
  9111=>"001101000",
  9112=>"111010011",
  9113=>"011111011",
  9114=>"110000001",
  9115=>"101001110",
  9116=>"010111101",
  9117=>"001100000",
  9118=>"001000000",
  9119=>"110011111",
  9120=>"001000101",
  9121=>"000011001",
  9122=>"001101000",
  9123=>"111010000",
  9124=>"110001111",
  9125=>"001010100",
  9126=>"000101111",
  9127=>"101011101",
  9128=>"110011000",
  9129=>"011000000",
  9130=>"110010011",
  9131=>"101100010",
  9132=>"010100011",
  9133=>"101001011",
  9134=>"101110010",
  9135=>"110000100",
  9136=>"010000111",
  9137=>"111101001",
  9138=>"000100001",
  9139=>"000101100",
  9140=>"000101111",
  9141=>"000111000",
  9142=>"111011010",
  9143=>"011101101",
  9144=>"011011000",
  9145=>"011100000",
  9146=>"010111000",
  9147=>"110101010",
  9148=>"000000010",
  9149=>"110111010",
  9150=>"001001010",
  9151=>"001100110",
  9152=>"000111100",
  9153=>"010111101",
  9154=>"000101000",
  9155=>"000100110",
  9156=>"001001011",
  9157=>"101100011",
  9158=>"101110010",
  9159=>"110001011",
  9160=>"111111111",
  9161=>"101110110",
  9162=>"101110001",
  9163=>"100110111",
  9164=>"001011001",
  9165=>"011001101",
  9166=>"001001001",
  9167=>"000010100",
  9168=>"101101010",
  9169=>"010011111",
  9170=>"101101001",
  9171=>"101111000",
  9172=>"011010011",
  9173=>"011011010",
  9174=>"011001101",
  9175=>"000101001",
  9176=>"011001011",
  9177=>"000010101",
  9178=>"110010000",
  9179=>"111110000",
  9180=>"101000000",
  9181=>"100010100",
  9182=>"101000110",
  9183=>"110110111",
  9184=>"110100000",
  9185=>"110110111",
  9186=>"101010010",
  9187=>"110111101",
  9188=>"110000001",
  9189=>"100111011",
  9190=>"000100010",
  9191=>"100101100",
  9192=>"101101001",
  9193=>"111000010",
  9194=>"011000100",
  9195=>"110011001",
  9196=>"010111111",
  9197=>"011100011",
  9198=>"011100110",
  9199=>"110111110",
  9200=>"110010100",
  9201=>"110101110",
  9202=>"100101001",
  9203=>"111000000",
  9204=>"011110111",
  9205=>"110111100",
  9206=>"110011011",
  9207=>"111011100",
  9208=>"001111110",
  9209=>"010100111",
  9210=>"111010010",
  9211=>"111000001",
  9212=>"111100001",
  9213=>"010000101",
  9214=>"000101100",
  9215=>"001010001",
  9216=>"010101100",
  9217=>"011011110",
  9218=>"110101111",
  9219=>"010001010",
  9220=>"010010101",
  9221=>"110100001",
  9222=>"111110100",
  9223=>"110111011",
  9224=>"011001101",
  9225=>"101101010",
  9226=>"111011000",
  9227=>"010011010",
  9228=>"110010100",
  9229=>"000101000",
  9230=>"001111100",
  9231=>"100111110",
  9232=>"000111101",
  9233=>"111000010",
  9234=>"000100110",
  9235=>"101110100",
  9236=>"101000001",
  9237=>"100011101",
  9238=>"000000011",
  9239=>"111111011",
  9240=>"100010001",
  9241=>"010101001",
  9242=>"111111010",
  9243=>"111111111",
  9244=>"111110000",
  9245=>"101110101",
  9246=>"001100110",
  9247=>"001010101",
  9248=>"100110111",
  9249=>"100110010",
  9250=>"110110000",
  9251=>"100000111",
  9252=>"100110100",
  9253=>"011010000",
  9254=>"111110000",
  9255=>"011110110",
  9256=>"010011000",
  9257=>"101001001",
  9258=>"001010000",
  9259=>"001010011",
  9260=>"101000111",
  9261=>"011110001",
  9262=>"110010101",
  9263=>"100011010",
  9264=>"011110110",
  9265=>"111010010",
  9266=>"110101110",
  9267=>"110101001",
  9268=>"111110111",
  9269=>"001000011",
  9270=>"111011011",
  9271=>"110110001",
  9272=>"001010010",
  9273=>"110111110",
  9274=>"011010000",
  9275=>"011010100",
  9276=>"000110001",
  9277=>"000100010",
  9278=>"111010101",
  9279=>"110110100",
  9280=>"111000110",
  9281=>"010010110",
  9282=>"011010001",
  9283=>"011100001",
  9284=>"000100010",
  9285=>"011111111",
  9286=>"111110110",
  9287=>"001100000",
  9288=>"000011001",
  9289=>"111011101",
  9290=>"001101000",
  9291=>"100011001",
  9292=>"100001110",
  9293=>"101101000",
  9294=>"100101000",
  9295=>"100111101",
  9296=>"010111000",
  9297=>"111101001",
  9298=>"101101111",
  9299=>"001011110",
  9300=>"111000111",
  9301=>"111100100",
  9302=>"101000111",
  9303=>"011110111",
  9304=>"001100011",
  9305=>"101111010",
  9306=>"001111000",
  9307=>"000101011",
  9308=>"011101110",
  9309=>"111100010",
  9310=>"110010010",
  9311=>"110000101",
  9312=>"000000110",
  9313=>"101100010",
  9314=>"010111000",
  9315=>"000001000",
  9316=>"000100000",
  9317=>"100100100",
  9318=>"011101100",
  9319=>"111010100",
  9320=>"011101000",
  9321=>"111101000",
  9322=>"111110000",
  9323=>"001110000",
  9324=>"011100100",
  9325=>"100110011",
  9326=>"101100000",
  9327=>"011110000",
  9328=>"101000110",
  9329=>"100100001",
  9330=>"111010110",
  9331=>"000110001",
  9332=>"110110100",
  9333=>"010111000",
  9334=>"011000010",
  9335=>"111101101",
  9336=>"111001011",
  9337=>"111001011",
  9338=>"011110110",
  9339=>"100010100",
  9340=>"101101011",
  9341=>"010111000",
  9342=>"100110110",
  9343=>"010011001",
  9344=>"110111011",
  9345=>"010101110",
  9346=>"110010001",
  9347=>"101110110",
  9348=>"111010000",
  9349=>"000101001",
  9350=>"111110100",
  9351=>"100010111",
  9352=>"001111110",
  9353=>"010000110",
  9354=>"100111110",
  9355=>"110111101",
  9356=>"010000101",
  9357=>"100100011",
  9358=>"100000011",
  9359=>"100001001",
  9360=>"011100000",
  9361=>"011000111",
  9362=>"000001101",
  9363=>"010011011",
  9364=>"000011010",
  9365=>"100110000",
  9366=>"111110111",
  9367=>"011001100",
  9368=>"011011000",
  9369=>"100001111",
  9370=>"111101011",
  9371=>"000001110",
  9372=>"111100000",
  9373=>"010111000",
  9374=>"101001010",
  9375=>"010110010",
  9376=>"111101011",
  9377=>"000010101",
  9378=>"010111111",
  9379=>"100010010",
  9380=>"110110110",
  9381=>"110100111",
  9382=>"000100010",
  9383=>"111100010",
  9384=>"010111100",
  9385=>"111110111",
  9386=>"011001001",
  9387=>"001110001",
  9388=>"011011100",
  9389=>"101010001",
  9390=>"101010011",
  9391=>"110011111",
  9392=>"111110111",
  9393=>"010011000",
  9394=>"101101100",
  9395=>"100000001",
  9396=>"000000000",
  9397=>"000000000",
  9398=>"101011110",
  9399=>"101111101",
  9400=>"010011000",
  9401=>"001001010",
  9402=>"111101000",
  9403=>"110110001",
  9404=>"011100100",
  9405=>"000101010",
  9406=>"110011101",
  9407=>"100111011",
  9408=>"100010011",
  9409=>"110111000",
  9410=>"011111111",
  9411=>"110101110",
  9412=>"010100101",
  9413=>"110010011",
  9414=>"000110011",
  9415=>"100000111",
  9416=>"010100111",
  9417=>"111110110",
  9418=>"111110001",
  9419=>"011000111",
  9420=>"100000000",
  9421=>"010111111",
  9422=>"111010101",
  9423=>"011100111",
  9424=>"101011011",
  9425=>"000111101",
  9426=>"001101000",
  9427=>"100000010",
  9428=>"111000000",
  9429=>"010011111",
  9430=>"101010111",
  9431=>"100011000",
  9432=>"000110011",
  9433=>"111001011",
  9434=>"000110100",
  9435=>"111110011",
  9436=>"001001000",
  9437=>"111111101",
  9438=>"011001111",
  9439=>"000011111",
  9440=>"010111101",
  9441=>"001101111",
  9442=>"011111010",
  9443=>"110111000",
  9444=>"001100100",
  9445=>"000101111",
  9446=>"010010000",
  9447=>"001111111",
  9448=>"001101110",
  9449=>"101000011",
  9450=>"111010111",
  9451=>"000110000",
  9452=>"100110101",
  9453=>"001101101",
  9454=>"000000001",
  9455=>"110000000",
  9456=>"000101101",
  9457=>"010101001",
  9458=>"000011010",
  9459=>"010100001",
  9460=>"110101100",
  9461=>"111111111",
  9462=>"010100000",
  9463=>"111111101",
  9464=>"100011100",
  9465=>"000011000",
  9466=>"000101100",
  9467=>"001011010",
  9468=>"011011010",
  9469=>"011000100",
  9470=>"111011110",
  9471=>"110100010",
  9472=>"000001110",
  9473=>"110011111",
  9474=>"000111100",
  9475=>"011110000",
  9476=>"000000111",
  9477=>"000101010",
  9478=>"011101110",
  9479=>"000110000",
  9480=>"011001110",
  9481=>"001101011",
  9482=>"110101001",
  9483=>"001010001",
  9484=>"111111111",
  9485=>"110110001",
  9486=>"001110100",
  9487=>"011101101",
  9488=>"000010111",
  9489=>"110011011",
  9490=>"010101100",
  9491=>"110010010",
  9492=>"100100101",
  9493=>"000010001",
  9494=>"111111010",
  9495=>"100010100",
  9496=>"111100001",
  9497=>"110001000",
  9498=>"111101111",
  9499=>"001101111",
  9500=>"110111101",
  9501=>"100011111",
  9502=>"101110010",
  9503=>"101101101",
  9504=>"010001111",
  9505=>"010011100",
  9506=>"110011001",
  9507=>"101001010",
  9508=>"000101000",
  9509=>"100010001",
  9510=>"001000010",
  9511=>"110011011",
  9512=>"000000100",
  9513=>"100101001",
  9514=>"110001010",
  9515=>"100101101",
  9516=>"000000111",
  9517=>"010001101",
  9518=>"011111101",
  9519=>"101001110",
  9520=>"001100110",
  9521=>"001010101",
  9522=>"110100110",
  9523=>"101100110",
  9524=>"010100000",
  9525=>"100111100",
  9526=>"001011000",
  9527=>"010101101",
  9528=>"000000110",
  9529=>"010100011",
  9530=>"010000000",
  9531=>"011000010",
  9532=>"000000100",
  9533=>"101111010",
  9534=>"000001011",
  9535=>"010001110",
  9536=>"111000101",
  9537=>"001111111",
  9538=>"001011100",
  9539=>"111110011",
  9540=>"011000111",
  9541=>"101011000",
  9542=>"001011000",
  9543=>"110000000",
  9544=>"000100010",
  9545=>"000100011",
  9546=>"100010000",
  9547=>"111111111",
  9548=>"011011111",
  9549=>"111010100",
  9550=>"001000010",
  9551=>"010010000",
  9552=>"011101011",
  9553=>"011101110",
  9554=>"000111101",
  9555=>"001111011",
  9556=>"111000101",
  9557=>"110101011",
  9558=>"011101110",
  9559=>"111000001",
  9560=>"101000101",
  9561=>"001000101",
  9562=>"000111000",
  9563=>"111000110",
  9564=>"110101001",
  9565=>"000011010",
  9566=>"101000000",
  9567=>"011101111",
  9568=>"111100111",
  9569=>"111001010",
  9570=>"101110111",
  9571=>"010111110",
  9572=>"100010110",
  9573=>"010001101",
  9574=>"000100001",
  9575=>"011110001",
  9576=>"011011100",
  9577=>"011110111",
  9578=>"001101110",
  9579=>"010110101",
  9580=>"011011111",
  9581=>"011111111",
  9582=>"011110100",
  9583=>"010110100",
  9584=>"010011111",
  9585=>"000001110",
  9586=>"011111011",
  9587=>"001001100",
  9588=>"110010101",
  9589=>"101000000",
  9590=>"101000011",
  9591=>"100000110",
  9592=>"100000101",
  9593=>"001010011",
  9594=>"110011001",
  9595=>"010101011",
  9596=>"111000010",
  9597=>"010100110",
  9598=>"000000010",
  9599=>"010111111",
  9600=>"101101000",
  9601=>"001000100",
  9602=>"001101101",
  9603=>"011011111",
  9604=>"001000010",
  9605=>"010110000",
  9606=>"100100100",
  9607=>"011000110",
  9608=>"110001101",
  9609=>"100000000",
  9610=>"111101100",
  9611=>"000110100",
  9612=>"101111110",
  9613=>"011100000",
  9614=>"011011110",
  9615=>"001101001",
  9616=>"011010100",
  9617=>"110010000",
  9618=>"110100110",
  9619=>"101010100",
  9620=>"001000100",
  9621=>"100100001",
  9622=>"011001010",
  9623=>"111011011",
  9624=>"011110011",
  9625=>"101011110",
  9626=>"101100000",
  9627=>"101011110",
  9628=>"001101111",
  9629=>"101110110",
  9630=>"011010011",
  9631=>"111010110",
  9632=>"110011011",
  9633=>"001001000",
  9634=>"001010101",
  9635=>"100100001",
  9636=>"101000000",
  9637=>"000001010",
  9638=>"001010100",
  9639=>"110111110",
  9640=>"001001011",
  9641=>"010001000",
  9642=>"000010111",
  9643=>"101011000",
  9644=>"000011101",
  9645=>"000100000",
  9646=>"010100111",
  9647=>"000001000",
  9648=>"001011000",
  9649=>"000110011",
  9650=>"100011010",
  9651=>"101101000",
  9652=>"101000001",
  9653=>"111001101",
  9654=>"011001010",
  9655=>"100001100",
  9656=>"110111001",
  9657=>"011101111",
  9658=>"011011111",
  9659=>"111110000",
  9660=>"000110101",
  9661=>"110000111",
  9662=>"001101010",
  9663=>"101100101",
  9664=>"100010010",
  9665=>"101100100",
  9666=>"010100010",
  9667=>"011011000",
  9668=>"011110111",
  9669=>"111011111",
  9670=>"111111110",
  9671=>"000000001",
  9672=>"010110110",
  9673=>"001010110",
  9674=>"100000101",
  9675=>"110010111",
  9676=>"011010111",
  9677=>"011000110",
  9678=>"010001011",
  9679=>"011010111",
  9680=>"011111100",
  9681=>"111010110",
  9682=>"100001111",
  9683=>"100101101",
  9684=>"001001110",
  9685=>"000110100",
  9686=>"011110100",
  9687=>"011111011",
  9688=>"111011001",
  9689=>"011111100",
  9690=>"110000101",
  9691=>"111111000",
  9692=>"010110100",
  9693=>"000010111",
  9694=>"000111110",
  9695=>"011011110",
  9696=>"001011101",
  9697=>"000001001",
  9698=>"000101001",
  9699=>"011010000",
  9700=>"000011010",
  9701=>"000110101",
  9702=>"100110101",
  9703=>"111101000",
  9704=>"010111110",
  9705=>"000101000",
  9706=>"011101100",
  9707=>"110000010",
  9708=>"001100000",
  9709=>"111111011",
  9710=>"010001101",
  9711=>"010011000",
  9712=>"010010101",
  9713=>"001110111",
  9714=>"110101111",
  9715=>"010001000",
  9716=>"010001001",
  9717=>"000011000",
  9718=>"000011011",
  9719=>"101101011",
  9720=>"110000111",
  9721=>"000110110",
  9722=>"111100101",
  9723=>"011010011",
  9724=>"010011110",
  9725=>"101110101",
  9726=>"010101000",
  9727=>"110001000",
  9728=>"001010110",
  9729=>"011110111",
  9730=>"110100000",
  9731=>"011000001",
  9732=>"011010010",
  9733=>"010000000",
  9734=>"010100101",
  9735=>"101111101",
  9736=>"100110001",
  9737=>"100111101",
  9738=>"010110000",
  9739=>"110011101",
  9740=>"011101111",
  9741=>"111011011",
  9742=>"100101011",
  9743=>"011111001",
  9744=>"000100110",
  9745=>"111110110",
  9746=>"101000010",
  9747=>"101110001",
  9748=>"000000010",
  9749=>"010000010",
  9750=>"111011110",
  9751=>"111100011",
  9752=>"111100111",
  9753=>"000100001",
  9754=>"110010011",
  9755=>"111000101",
  9756=>"001101001",
  9757=>"000000110",
  9758=>"011000111",
  9759=>"010111010",
  9760=>"010010000",
  9761=>"110100001",
  9762=>"100101000",
  9763=>"110111011",
  9764=>"100000011",
  9765=>"001000010",
  9766=>"101000011",
  9767=>"001000010",
  9768=>"000000100",
  9769=>"010000000",
  9770=>"010110100",
  9771=>"111100100",
  9772=>"001100111",
  9773=>"011110010",
  9774=>"101100100",
  9775=>"100001100",
  9776=>"101011001",
  9777=>"100111011",
  9778=>"100010110",
  9779=>"011110111",
  9780=>"001110011",
  9781=>"000111110",
  9782=>"110001100",
  9783=>"010100000",
  9784=>"001100001",
  9785=>"001110011",
  9786=>"011001101",
  9787=>"110100101",
  9788=>"101111000",
  9789=>"111110001",
  9790=>"000110111",
  9791=>"001001111",
  9792=>"000001011",
  9793=>"001100010",
  9794=>"011000000",
  9795=>"010100110",
  9796=>"010010100",
  9797=>"010001010",
  9798=>"110011111",
  9799=>"100000000",
  9800=>"111110001",
  9801=>"010011011",
  9802=>"110000111",
  9803=>"000001000",
  9804=>"000101000",
  9805=>"101001110",
  9806=>"110000100",
  9807=>"101001001",
  9808=>"001001011",
  9809=>"101100011",
  9810=>"101001100",
  9811=>"010011001",
  9812=>"100101001",
  9813=>"111111100",
  9814=>"011100110",
  9815=>"110010001",
  9816=>"101110010",
  9817=>"001010100",
  9818=>"000010001",
  9819=>"000000000",
  9820=>"001101010",
  9821=>"111000000",
  9822=>"100010111",
  9823=>"110101100",
  9824=>"011010100",
  9825=>"010001100",
  9826=>"010011010",
  9827=>"100111111",
  9828=>"011010000",
  9829=>"100000000",
  9830=>"000001101",
  9831=>"010011011",
  9832=>"101011011",
  9833=>"100101001",
  9834=>"001011110",
  9835=>"111101000",
  9836=>"010100110",
  9837=>"101111010",
  9838=>"000010101",
  9839=>"100001000",
  9840=>"000110000",
  9841=>"110110100",
  9842=>"011111100",
  9843=>"111101101",
  9844=>"000000010",
  9845=>"110001100",
  9846=>"000111000",
  9847=>"100011001",
  9848=>"111111010",
  9849=>"100110001",
  9850=>"010100001",
  9851=>"000001001",
  9852=>"100101000",
  9853=>"001100100",
  9854=>"100111101",
  9855=>"100000100",
  9856=>"001000000",
  9857=>"111111000",
  9858=>"100100110",
  9859=>"010010011",
  9860=>"011011110",
  9861=>"010110011",
  9862=>"011000111",
  9863=>"010110010",
  9864=>"010001111",
  9865=>"010010110",
  9866=>"100101101",
  9867=>"110000010",
  9868=>"010000111",
  9869=>"100011111",
  9870=>"011111010",
  9871=>"001100010",
  9872=>"101010100",
  9873=>"010000010",
  9874=>"100100101",
  9875=>"100010010",
  9876=>"101110010",
  9877=>"010110111",
  9878=>"000111100",
  9879=>"001110001",
  9880=>"111000101",
  9881=>"010011111",
  9882=>"101010001",
  9883=>"001010101",
  9884=>"101111000",
  9885=>"010100011",
  9886=>"001000000",
  9887=>"010011010",
  9888=>"100001010",
  9889=>"101010001",
  9890=>"001010000",
  9891=>"101011001",
  9892=>"011010101",
  9893=>"000111111",
  9894=>"001000100",
  9895=>"100001011",
  9896=>"010001100",
  9897=>"101010010",
  9898=>"111100001",
  9899=>"100000110",
  9900=>"000100111",
  9901=>"111010101",
  9902=>"100001011",
  9903=>"010111000",
  9904=>"001111101",
  9905=>"010101011",
  9906=>"111001010",
  9907=>"101011001",
  9908=>"011111110",
  9909=>"010010110",
  9910=>"100000111",
  9911=>"010011011",
  9912=>"111111100",
  9913=>"111000110",
  9914=>"001111101",
  9915=>"110111001",
  9916=>"101101100",
  9917=>"001101011",
  9918=>"111011001",
  9919=>"000001111",
  9920=>"011011001",
  9921=>"011111100",
  9922=>"110010100",
  9923=>"010100011",
  9924=>"100100000",
  9925=>"110101111",
  9926=>"001100100",
  9927=>"101100010",
  9928=>"101101111",
  9929=>"010001111",
  9930=>"011010010",
  9931=>"000110001",
  9932=>"101110011",
  9933=>"100010011",
  9934=>"101011000",
  9935=>"111011100",
  9936=>"000111100",
  9937=>"100110001",
  9938=>"100101110",
  9939=>"010110101",
  9940=>"010111111",
  9941=>"111001000",
  9942=>"011000011",
  9943=>"011001000",
  9944=>"000111000",
  9945=>"111101001",
  9946=>"111100010",
  9947=>"001100010",
  9948=>"110010101",
  9949=>"011000000",
  9950=>"100000000",
  9951=>"000001110",
  9952=>"000111010",
  9953=>"001001101",
  9954=>"000000111",
  9955=>"100011001",
  9956=>"101000001",
  9957=>"111110001",
  9958=>"001000101",
  9959=>"110001001",
  9960=>"000101001",
  9961=>"100010000",
  9962=>"011001110",
  9963=>"011010010",
  9964=>"000000010",
  9965=>"111101011",
  9966=>"000110001",
  9967=>"111111111",
  9968=>"001100001",
  9969=>"110101000",
  9970=>"011100100",
  9971=>"011001111",
  9972=>"101001100",
  9973=>"101000101",
  9974=>"011000000",
  9975=>"110010001",
  9976=>"011110111",
  9977=>"001101110",
  9978=>"000111100",
  9979=>"000000011",
  9980=>"010011011",
  9981=>"101111001",
  9982=>"110001001",
  9983=>"111110010",
  9984=>"111110111",
  9985=>"111000111",
  9986=>"011100000",
  9987=>"100110010",
  9988=>"111010000",
  9989=>"111001111",
  9990=>"001000101",
  9991=>"011001011",
  9992=>"110100101",
  9993=>"001010001",
  9994=>"001001111",
  9995=>"000101010",
  9996=>"111101111",
  9997=>"011001101",
  9998=>"100011101",
  9999=>"111101011",
  10000=>"100010110",
  10001=>"000000000",
  10002=>"000010100",
  10003=>"001000001",
  10004=>"010000100",
  10005=>"101101011",
  10006=>"000110111",
  10007=>"001011100",
  10008=>"001110101",
  10009=>"010101110",
  10010=>"100011000",
  10011=>"010001000",
  10012=>"011100000",
  10013=>"110000110",
  10014=>"010110011",
  10015=>"111011101",
  10016=>"011001110",
  10017=>"100000001",
  10018=>"111000000",
  10019=>"101100011",
  10020=>"110111010",
  10021=>"101110001",
  10022=>"101100110",
  10023=>"001101010",
  10024=>"100001111",
  10025=>"011110111",
  10026=>"101111001",
  10027=>"001000100",
  10028=>"000100110",
  10029=>"001001000",
  10030=>"111010110",
  10031=>"011111111",
  10032=>"011010111",
  10033=>"111010101",
  10034=>"000101011",
  10035=>"000000110",
  10036=>"011111000",
  10037=>"101001000",
  10038=>"100011010",
  10039=>"111101000",
  10040=>"111100010",
  10041=>"001010001",
  10042=>"011010000",
  10043=>"111110111",
  10044=>"101101110",
  10045=>"010001000",
  10046=>"000111110",
  10047=>"100000101",
  10048=>"000010100",
  10049=>"000110000",
  10050=>"001111010",
  10051=>"101011001",
  10052=>"011010101",
  10053=>"011101011",
  10054=>"000110111",
  10055=>"011101111",
  10056=>"101100001",
  10057=>"111011111",
  10058=>"101111101",
  10059=>"000110110",
  10060=>"011010110",
  10061=>"101110000",
  10062=>"101011001",
  10063=>"101101110",
  10064=>"111011001",
  10065=>"001111000",
  10066=>"111101000",
  10067=>"111010001",
  10068=>"101111111",
  10069=>"111101111",
  10070=>"001111101",
  10071=>"101010010",
  10072=>"011100101",
  10073=>"010100100",
  10074=>"100001011",
  10075=>"111100110",
  10076=>"110010010",
  10077=>"111000010",
  10078=>"110000100",
  10079=>"110001101",
  10080=>"111010110",
  10081=>"100010000",
  10082=>"001000000",
  10083=>"011110011",
  10084=>"001111111",
  10085=>"100000010",
  10086=>"111001010",
  10087=>"101100000",
  10088=>"000110000",
  10089=>"110101101",
  10090=>"111001010",
  10091=>"001001001",
  10092=>"000111111",
  10093=>"110111110",
  10094=>"000110101",
  10095=>"010001110",
  10096=>"010011010",
  10097=>"101110010",
  10098=>"001010000",
  10099=>"110010000",
  10100=>"001001001",
  10101=>"101001011",
  10102=>"000111001",
  10103=>"011011101",
  10104=>"101100011",
  10105=>"011100110",
  10106=>"010000110",
  10107=>"111101100",
  10108=>"100011100",
  10109=>"000011100",
  10110=>"001110111",
  10111=>"101110100",
  10112=>"111110101",
  10113=>"000110001",
  10114=>"000010010",
  10115=>"000100111",
  10116=>"010011001",
  10117=>"000010101",
  10118=>"000001011",
  10119=>"001011110",
  10120=>"000011111",
  10121=>"111010110",
  10122=>"000010001",
  10123=>"101110101",
  10124=>"111000111",
  10125=>"111101011",
  10126=>"010000101",
  10127=>"101110001",
  10128=>"000000010",
  10129=>"011001000",
  10130=>"011010001",
  10131=>"000011000",
  10132=>"111100101",
  10133=>"001010000",
  10134=>"001001111",
  10135=>"110110000",
  10136=>"100100010",
  10137=>"000011001",
  10138=>"100010101",
  10139=>"000000111",
  10140=>"001001000",
  10141=>"011011111",
  10142=>"111111100",
  10143=>"100100100",
  10144=>"001010100",
  10145=>"011111010",
  10146=>"001001011",
  10147=>"111000010",
  10148=>"000110111",
  10149=>"001101000",
  10150=>"100001000",
  10151=>"001110110",
  10152=>"000110011",
  10153=>"001111001",
  10154=>"010110010",
  10155=>"101000001",
  10156=>"111001101",
  10157=>"101110100",
  10158=>"011010111",
  10159=>"001011101",
  10160=>"111010100",
  10161=>"011110100",
  10162=>"101101001",
  10163=>"101011110",
  10164=>"011011111",
  10165=>"001011010",
  10166=>"011101110",
  10167=>"000101011",
  10168=>"111101010",
  10169=>"011011110",
  10170=>"101000100",
  10171=>"010000011",
  10172=>"100011011",
  10173=>"111011111",
  10174=>"111010101",
  10175=>"001001000",
  10176=>"000001000",
  10177=>"001100010",
  10178=>"010011111",
  10179=>"000100001",
  10180=>"100101011",
  10181=>"001011010",
  10182=>"111000101",
  10183=>"001101100",
  10184=>"011011001",
  10185=>"000000010",
  10186=>"101001001",
  10187=>"000001101",
  10188=>"111100000",
  10189=>"001111000",
  10190=>"100000101",
  10191=>"100000010",
  10192=>"011000010",
  10193=>"010000111",
  10194=>"101011101",
  10195=>"001110000",
  10196=>"110111010",
  10197=>"111101101",
  10198=>"000011001",
  10199=>"101011011",
  10200=>"011011101",
  10201=>"101110101",
  10202=>"101000000",
  10203=>"111001000",
  10204=>"001000010",
  10205=>"111001010",
  10206=>"001110100",
  10207=>"001101101",
  10208=>"111111010",
  10209=>"000000100",
  10210=>"111101111",
  10211=>"000001000",
  10212=>"101001000",
  10213=>"110001001",
  10214=>"111000110",
  10215=>"101001100",
  10216=>"000111101",
  10217=>"000111110",
  10218=>"100010100",
  10219=>"110100111",
  10220=>"101111111",
  10221=>"101001111",
  10222=>"101101000",
  10223=>"001110111",
  10224=>"000001101",
  10225=>"010011101",
  10226=>"110110111",
  10227=>"100100000",
  10228=>"001001111",
  10229=>"110111111",
  10230=>"111110010",
  10231=>"001101111",
  10232=>"010001010",
  10233=>"010001100",
  10234=>"111011100",
  10235=>"111000111",
  10236=>"011001001",
  10237=>"110111100",
  10238=>"011011011",
  10239=>"101100110",
  10240=>"110100111",
  10241=>"000101011",
  10242=>"010011101",
  10243=>"110001100",
  10244=>"101101100",
  10245=>"111011100",
  10246=>"010011110",
  10247=>"001001010",
  10248=>"010010110",
  10249=>"110101000",
  10250=>"100011111",
  10251=>"011110011",
  10252=>"000110000",
  10253=>"111010010",
  10254=>"010100010",
  10255=>"101010000",
  10256=>"111111110",
  10257=>"101101101",
  10258=>"111001001",
  10259=>"100001010",
  10260=>"110101111",
  10261=>"101110011",
  10262=>"010110100",
  10263=>"101101000",
  10264=>"100010100",
  10265=>"111011010",
  10266=>"101001100",
  10267=>"000110110",
  10268=>"111010101",
  10269=>"110001100",
  10270=>"101111000",
  10271=>"101101000",
  10272=>"000010000",
  10273=>"111011101",
  10274=>"000010011",
  10275=>"111010111",
  10276=>"101101110",
  10277=>"110111100",
  10278=>"001101001",
  10279=>"000011010",
  10280=>"100001010",
  10281=>"001111101",
  10282=>"010100001",
  10283=>"011110111",
  10284=>"110001010",
  10285=>"100000010",
  10286=>"001000011",
  10287=>"010110100",
  10288=>"111101010",
  10289=>"000011111",
  10290=>"111010110",
  10291=>"000010001",
  10292=>"011010100",
  10293=>"110010000",
  10294=>"001100100",
  10295=>"011011101",
  10296=>"011011101",
  10297=>"000010110",
  10298=>"001110001",
  10299=>"010111101",
  10300=>"001101101",
  10301=>"011110011",
  10302=>"010001000",
  10303=>"011100110",
  10304=>"110001001",
  10305=>"001111010",
  10306=>"100001001",
  10307=>"011101110",
  10308=>"101001101",
  10309=>"100101010",
  10310=>"000010111",
  10311=>"110001101",
  10312=>"100000111",
  10313=>"100101101",
  10314=>"100001000",
  10315=>"110111001",
  10316=>"011101011",
  10317=>"101100100",
  10318=>"110100000",
  10319=>"000011000",
  10320=>"011100101",
  10321=>"001100010",
  10322=>"111100101",
  10323=>"110101110",
  10324=>"001101100",
  10325=>"111001010",
  10326=>"001101011",
  10327=>"010011010",
  10328=>"000001110",
  10329=>"111110000",
  10330=>"110011101",
  10331=>"001101011",
  10332=>"100100110",
  10333=>"101000110",
  10334=>"111000101",
  10335=>"101101101",
  10336=>"010011101",
  10337=>"110000111",
  10338=>"101011001",
  10339=>"101011110",
  10340=>"110000110",
  10341=>"101001111",
  10342=>"110011000",
  10343=>"111010111",
  10344=>"101111001",
  10345=>"000010000",
  10346=>"010111010",
  10347=>"110100000",
  10348=>"111101001",
  10349=>"110110111",
  10350=>"010100100",
  10351=>"001111001",
  10352=>"010111011",
  10353=>"001110001",
  10354=>"001001100",
  10355=>"101100100",
  10356=>"101111000",
  10357=>"101010000",
  10358=>"001011001",
  10359=>"000000001",
  10360=>"110001010",
  10361=>"011111000",
  10362=>"011000011",
  10363=>"011010010",
  10364=>"110101111",
  10365=>"101001101",
  10366=>"000011000",
  10367=>"010010010",
  10368=>"110010011",
  10369=>"110111111",
  10370=>"101100000",
  10371=>"010001110",
  10372=>"111110111",
  10373=>"001101000",
  10374=>"101100111",
  10375=>"111001100",
  10376=>"111010000",
  10377=>"111111010",
  10378=>"111100000",
  10379=>"011010100",
  10380=>"100010110",
  10381=>"101110010",
  10382=>"111011100",
  10383=>"010010101",
  10384=>"010111000",
  10385=>"011001001",
  10386=>"110111001",
  10387=>"011100010",
  10388=>"100000010",
  10389=>"110000000",
  10390=>"100000110",
  10391=>"100111001",
  10392=>"001101110",
  10393=>"000010011",
  10394=>"111001111",
  10395=>"111100110",
  10396=>"011011100",
  10397=>"110101101",
  10398=>"011111011",
  10399=>"001010000",
  10400=>"001110001",
  10401=>"111111000",
  10402=>"011000001",
  10403=>"010110111",
  10404=>"110011111",
  10405=>"111111111",
  10406=>"010111001",
  10407=>"110111111",
  10408=>"110001100",
  10409=>"011011010",
  10410=>"111100110",
  10411=>"101010111",
  10412=>"011011011",
  10413=>"011011101",
  10414=>"001000010",
  10415=>"100010000",
  10416=>"001101010",
  10417=>"000111111",
  10418=>"111110011",
  10419=>"001100010",
  10420=>"011000011",
  10421=>"111111110",
  10422=>"110010110",
  10423=>"000000010",
  10424=>"010010111",
  10425=>"000001111",
  10426=>"111010101",
  10427=>"001011000",
  10428=>"001101010",
  10429=>"000001101",
  10430=>"111100001",
  10431=>"000010111",
  10432=>"010101111",
  10433=>"000001110",
  10434=>"111111111",
  10435=>"100000111",
  10436=>"111101100",
  10437=>"100010110",
  10438=>"001011100",
  10439=>"010111001",
  10440=>"101101101",
  10441=>"011010011",
  10442=>"011011001",
  10443=>"011100100",
  10444=>"101111000",
  10445=>"011010100",
  10446=>"000001111",
  10447=>"010110001",
  10448=>"101111111",
  10449=>"001101100",
  10450=>"110011000",
  10451=>"110001000",
  10452=>"100011011",
  10453=>"001001010",
  10454=>"001010101",
  10455=>"111010001",
  10456=>"000001111",
  10457=>"010110100",
  10458=>"101010011",
  10459=>"011000000",
  10460=>"000001001",
  10461=>"111001100",
  10462=>"100111100",
  10463=>"111001100",
  10464=>"010011111",
  10465=>"110001101",
  10466=>"011010100",
  10467=>"111100100",
  10468=>"100011111",
  10469=>"001101010",
  10470=>"111000011",
  10471=>"011001010",
  10472=>"000001100",
  10473=>"111010101",
  10474=>"011110001",
  10475=>"011111110",
  10476=>"010100001",
  10477=>"101001110",
  10478=>"111011111",
  10479=>"110101011",
  10480=>"011101110",
  10481=>"010111101",
  10482=>"111110000",
  10483=>"000001001",
  10484=>"110011011",
  10485=>"001011110",
  10486=>"110011000",
  10487=>"000101100",
  10488=>"110101111",
  10489=>"000100001",
  10490=>"111100111",
  10491=>"111011101",
  10492=>"010101011",
  10493=>"010010010",
  10494=>"011100100",
  10495=>"010001011",
  10496=>"101000110",
  10497=>"101110001",
  10498=>"001000010",
  10499=>"001001110",
  10500=>"011010001",
  10501=>"101101110",
  10502=>"011110010",
  10503=>"011010110",
  10504=>"111101000",
  10505=>"111001011",
  10506=>"001000001",
  10507=>"001101001",
  10508=>"011001001",
  10509=>"111010110",
  10510=>"000011100",
  10511=>"000011010",
  10512=>"011000111",
  10513=>"011011010",
  10514=>"011001000",
  10515=>"011011010",
  10516=>"111110001",
  10517=>"011110010",
  10518=>"001010000",
  10519=>"111101010",
  10520=>"110100000",
  10521=>"111100111",
  10522=>"111010010",
  10523=>"100011100",
  10524=>"000010001",
  10525=>"111001011",
  10526=>"110010011",
  10527=>"000010010",
  10528=>"111100111",
  10529=>"111010001",
  10530=>"111111110",
  10531=>"101001000",
  10532=>"111001111",
  10533=>"000101000",
  10534=>"010000011",
  10535=>"011000110",
  10536=>"111011110",
  10537=>"100000000",
  10538=>"100000001",
  10539=>"110100011",
  10540=>"001101100",
  10541=>"001001000",
  10542=>"111100010",
  10543=>"001000110",
  10544=>"110111111",
  10545=>"110011111",
  10546=>"111010110",
  10547=>"111110110",
  10548=>"011001011",
  10549=>"000000000",
  10550=>"010011100",
  10551=>"100110101",
  10552=>"111111001",
  10553=>"001101110",
  10554=>"101101000",
  10555=>"110101001",
  10556=>"101110100",
  10557=>"001100000",
  10558=>"100010100",
  10559=>"101101111",
  10560=>"111111111",
  10561=>"111110011",
  10562=>"000001111",
  10563=>"011110100",
  10564=>"011101101",
  10565=>"111100010",
  10566=>"100010001",
  10567=>"101100101",
  10568=>"111011101",
  10569=>"000000111",
  10570=>"100010000",
  10571=>"101000000",
  10572=>"001100010",
  10573=>"101110111",
  10574=>"010111101",
  10575=>"111111010",
  10576=>"001110100",
  10577=>"101001000",
  10578=>"100001101",
  10579=>"100010000",
  10580=>"011111001",
  10581=>"100100000",
  10582=>"010111010",
  10583=>"110110001",
  10584=>"101001101",
  10585=>"101001000",
  10586=>"010111001",
  10587=>"011100101",
  10588=>"001111011",
  10589=>"110011011",
  10590=>"111100101",
  10591=>"000111001",
  10592=>"010111010",
  10593=>"010110110",
  10594=>"000101011",
  10595=>"110011110",
  10596=>"000110101",
  10597=>"100001111",
  10598=>"111010010",
  10599=>"000010010",
  10600=>"111011111",
  10601=>"100010100",
  10602=>"011100100",
  10603=>"111000101",
  10604=>"111000111",
  10605=>"100111111",
  10606=>"111111110",
  10607=>"110101101",
  10608=>"000011110",
  10609=>"010001001",
  10610=>"110011010",
  10611=>"000010001",
  10612=>"000001000",
  10613=>"111001000",
  10614=>"011000101",
  10615=>"110000001",
  10616=>"010001101",
  10617=>"010100110",
  10618=>"110101010",
  10619=>"100001110",
  10620=>"001010001",
  10621=>"100101111",
  10622=>"101001011",
  10623=>"000010110",
  10624=>"101110111",
  10625=>"010001101",
  10626=>"111010111",
  10627=>"001001011",
  10628=>"110110011",
  10629=>"010011010",
  10630=>"010111000",
  10631=>"010101001",
  10632=>"111010001",
  10633=>"011110100",
  10634=>"010110001",
  10635=>"110001111",
  10636=>"011100111",
  10637=>"010011100",
  10638=>"011100000",
  10639=>"101001101",
  10640=>"010111100",
  10641=>"101101001",
  10642=>"100110011",
  10643=>"111111011",
  10644=>"111011010",
  10645=>"110001011",
  10646=>"000000010",
  10647=>"101010001",
  10648=>"100010100",
  10649=>"001101111",
  10650=>"111011011",
  10651=>"010010010",
  10652=>"001001001",
  10653=>"110110111",
  10654=>"100011111",
  10655=>"000110001",
  10656=>"001101011",
  10657=>"001000110",
  10658=>"111001110",
  10659=>"100000001",
  10660=>"011110010",
  10661=>"100101111",
  10662=>"101000111",
  10663=>"010111011",
  10664=>"000000011",
  10665=>"010000000",
  10666=>"010101111",
  10667=>"100001010",
  10668=>"111101000",
  10669=>"100000101",
  10670=>"100111111",
  10671=>"101110100",
  10672=>"111110001",
  10673=>"110000110",
  10674=>"011110110",
  10675=>"001010001",
  10676=>"111101110",
  10677=>"000010011",
  10678=>"000000010",
  10679=>"101010011",
  10680=>"100001111",
  10681=>"100010111",
  10682=>"110000110",
  10683=>"011110011",
  10684=>"000111100",
  10685=>"111011111",
  10686=>"110101111",
  10687=>"100011100",
  10688=>"010010001",
  10689=>"111100100",
  10690=>"110000101",
  10691=>"110001101",
  10692=>"101110011",
  10693=>"000100110",
  10694=>"011110101",
  10695=>"001111111",
  10696=>"100011101",
  10697=>"111100000",
  10698=>"111111111",
  10699=>"010100000",
  10700=>"101111010",
  10701=>"101011011",
  10702=>"000111111",
  10703=>"011110110",
  10704=>"110010011",
  10705=>"101011010",
  10706=>"001010000",
  10707=>"111001010",
  10708=>"011000100",
  10709=>"111010111",
  10710=>"001010101",
  10711=>"001111101",
  10712=>"110011011",
  10713=>"000100100",
  10714=>"110101000",
  10715=>"011100000",
  10716=>"101110100",
  10717=>"000100100",
  10718=>"111010111",
  10719=>"001000011",
  10720=>"111111111",
  10721=>"000001100",
  10722=>"000101110",
  10723=>"010101111",
  10724=>"000011011",
  10725=>"000100100",
  10726=>"100100100",
  10727=>"101110101",
  10728=>"111011110",
  10729=>"011100010",
  10730=>"000001110",
  10731=>"111010110",
  10732=>"111111111",
  10733=>"011110100",
  10734=>"111001111",
  10735=>"101100110",
  10736=>"001111011",
  10737=>"111111110",
  10738=>"111111101",
  10739=>"011010011",
  10740=>"101000000",
  10741=>"000011011",
  10742=>"101111011",
  10743=>"000000010",
  10744=>"001001111",
  10745=>"010001000",
  10746=>"111000110",
  10747=>"010100010",
  10748=>"101010110",
  10749=>"111111000",
  10750=>"100011000",
  10751=>"001000111",
  10752=>"011111100",
  10753=>"011101111",
  10754=>"111111110",
  10755=>"101001110",
  10756=>"000011000",
  10757=>"011101000",
  10758=>"011001010",
  10759=>"011011100",
  10760=>"100100011",
  10761=>"000001100",
  10762=>"111100011",
  10763=>"101110100",
  10764=>"010000000",
  10765=>"100010100",
  10766=>"010001010",
  10767=>"011101101",
  10768=>"100010001",
  10769=>"101110010",
  10770=>"100110000",
  10771=>"110100100",
  10772=>"110101001",
  10773=>"000111010",
  10774=>"001001010",
  10775=>"111001101",
  10776=>"001100011",
  10777=>"001100010",
  10778=>"100001010",
  10779=>"101010010",
  10780=>"111011001",
  10781=>"010100111",
  10782=>"110001110",
  10783=>"111000100",
  10784=>"110111110",
  10785=>"001001111",
  10786=>"001000111",
  10787=>"010111101",
  10788=>"110011011",
  10789=>"100010111",
  10790=>"011111101",
  10791=>"000001000",
  10792=>"000011000",
  10793=>"101101100",
  10794=>"011101010",
  10795=>"100001100",
  10796=>"011101100",
  10797=>"010011010",
  10798=>"001000001",
  10799=>"001011011",
  10800=>"101100111",
  10801=>"110000001",
  10802=>"010110100",
  10803=>"000101110",
  10804=>"011111111",
  10805=>"100001010",
  10806=>"000010110",
  10807=>"101111100",
  10808=>"100010010",
  10809=>"100011000",
  10810=>"111001100",
  10811=>"110010001",
  10812=>"111101100",
  10813=>"011001010",
  10814=>"100011111",
  10815=>"100100001",
  10816=>"100110001",
  10817=>"100010010",
  10818=>"101100101",
  10819=>"001000011",
  10820=>"100111110",
  10821=>"000001011",
  10822=>"001010000",
  10823=>"011010001",
  10824=>"111010000",
  10825=>"000011000",
  10826=>"011000010",
  10827=>"111111110",
  10828=>"100101100",
  10829=>"001111000",
  10830=>"010101111",
  10831=>"111101101",
  10832=>"000001000",
  10833=>"111110000",
  10834=>"111001110",
  10835=>"111101111",
  10836=>"000100010",
  10837=>"100111111",
  10838=>"111101011",
  10839=>"001011111",
  10840=>"001010111",
  10841=>"001001011",
  10842=>"111110100",
  10843=>"111111001",
  10844=>"000010010",
  10845=>"110110111",
  10846=>"101111101",
  10847=>"101010101",
  10848=>"101000001",
  10849=>"111011010",
  10850=>"111000111",
  10851=>"000100101",
  10852=>"110100010",
  10853=>"011100001",
  10854=>"001000000",
  10855=>"110101001",
  10856=>"010010001",
  10857=>"001010100",
  10858=>"110100001",
  10859=>"101010100",
  10860=>"001010000",
  10861=>"010011010",
  10862=>"111010010",
  10863=>"110001100",
  10864=>"000000110",
  10865=>"101001110",
  10866=>"010010010",
  10867=>"100000011",
  10868=>"000100000",
  10869=>"101001010",
  10870=>"111110111",
  10871=>"101011100",
  10872=>"110011111",
  10873=>"000100010",
  10874=>"010000100",
  10875=>"111111110",
  10876=>"110000110",
  10877=>"000010010",
  10878=>"101000000",
  10879=>"001110110",
  10880=>"110010111",
  10881=>"001001000",
  10882=>"111111000",
  10883=>"111111001",
  10884=>"111011100",
  10885=>"000110001",
  10886=>"111101100",
  10887=>"100100110",
  10888=>"010101011",
  10889=>"101011001",
  10890=>"111011010",
  10891=>"100111110",
  10892=>"010100111",
  10893=>"000101101",
  10894=>"010111110",
  10895=>"111100010",
  10896=>"010001000",
  10897=>"010010011",
  10898=>"100000110",
  10899=>"101001000",
  10900=>"111101001",
  10901=>"010101010",
  10902=>"001001001",
  10903=>"110100010",
  10904=>"111100101",
  10905=>"000101001",
  10906=>"111111001",
  10907=>"111011101",
  10908=>"111001000",
  10909=>"101100011",
  10910=>"000110101",
  10911=>"011011111",
  10912=>"101000110",
  10913=>"000001101",
  10914=>"001010101",
  10915=>"011011001",
  10916=>"111101011",
  10917=>"101011010",
  10918=>"111001101",
  10919=>"111101101",
  10920=>"010010001",
  10921=>"101010100",
  10922=>"101000111",
  10923=>"000001110",
  10924=>"111000010",
  10925=>"110101001",
  10926=>"010101000",
  10927=>"110100101",
  10928=>"101110011",
  10929=>"101001110",
  10930=>"101010011",
  10931=>"111010111",
  10932=>"111001001",
  10933=>"011001111",
  10934=>"010000101",
  10935=>"101111111",
  10936=>"011101010",
  10937=>"011111110",
  10938=>"110110000",
  10939=>"101001010",
  10940=>"001101111",
  10941=>"110110111",
  10942=>"010101111",
  10943=>"101100100",
  10944=>"010001101",
  10945=>"100110010",
  10946=>"100000011",
  10947=>"011111101",
  10948=>"100001111",
  10949=>"111010100",
  10950=>"101110101",
  10951=>"010010000",
  10952=>"010010111",
  10953=>"000101000",
  10954=>"010000000",
  10955=>"111111100",
  10956=>"101100101",
  10957=>"001111101",
  10958=>"011110110",
  10959=>"000010000",
  10960=>"101011101",
  10961=>"001100111",
  10962=>"101110110",
  10963=>"001111111",
  10964=>"101001000",
  10965=>"111110110",
  10966=>"000000111",
  10967=>"110110001",
  10968=>"000000011",
  10969=>"100101110",
  10970=>"110111101",
  10971=>"011111011",
  10972=>"101011011",
  10973=>"100100010",
  10974=>"010101100",
  10975=>"011111011",
  10976=>"101110011",
  10977=>"111000111",
  10978=>"011010011",
  10979=>"011011001",
  10980=>"001011011",
  10981=>"001010111",
  10982=>"111111111",
  10983=>"010010011",
  10984=>"101010100",
  10985=>"010111000",
  10986=>"111101010",
  10987=>"100001101",
  10988=>"001101100",
  10989=>"011101000",
  10990=>"011111110",
  10991=>"110100110",
  10992=>"000000011",
  10993=>"101100110",
  10994=>"001101101",
  10995=>"010000000",
  10996=>"111100101",
  10997=>"000011100",
  10998=>"000001110",
  10999=>"101001111",
  11000=>"010010111",
  11001=>"111100001",
  11002=>"000001001",
  11003=>"101100110",
  11004=>"101100100",
  11005=>"101101111",
  11006=>"101001010",
  11007=>"100110100",
  11008=>"111010100",
  11009=>"110000011",
  11010=>"000101011",
  11011=>"011011010",
  11012=>"010100011",
  11013=>"101011001",
  11014=>"001110011",
  11015=>"100001011",
  11016=>"111001000",
  11017=>"010101110",
  11018=>"000000001",
  11019=>"010000101",
  11020=>"010010110",
  11021=>"000011110",
  11022=>"000100010",
  11023=>"001010110",
  11024=>"111011101",
  11025=>"110100011",
  11026=>"010101010",
  11027=>"000000010",
  11028=>"110000010",
  11029=>"011001010",
  11030=>"011110100",
  11031=>"110001101",
  11032=>"101111101",
  11033=>"010011001",
  11034=>"011110111",
  11035=>"100110010",
  11036=>"101000010",
  11037=>"011101110",
  11038=>"011111101",
  11039=>"110110101",
  11040=>"111011111",
  11041=>"001000000",
  11042=>"001100100",
  11043=>"010011100",
  11044=>"111001010",
  11045=>"110110011",
  11046=>"111011000",
  11047=>"110000010",
  11048=>"111011101",
  11049=>"110111011",
  11050=>"011111000",
  11051=>"011101011",
  11052=>"111111110",
  11053=>"110110001",
  11054=>"000100111",
  11055=>"100100110",
  11056=>"001000110",
  11057=>"100010001",
  11058=>"001011111",
  11059=>"101110100",
  11060=>"010001101",
  11061=>"010001100",
  11062=>"110101000",
  11063=>"010000101",
  11064=>"011110110",
  11065=>"011100001",
  11066=>"110111001",
  11067=>"010011101",
  11068=>"001111011",
  11069=>"111010010",
  11070=>"110001111",
  11071=>"000001000",
  11072=>"100000011",
  11073=>"100100111",
  11074=>"100110101",
  11075=>"001110100",
  11076=>"111101000",
  11077=>"001100011",
  11078=>"000010100",
  11079=>"100001100",
  11080=>"000101001",
  11081=>"100011111",
  11082=>"101100101",
  11083=>"110001110",
  11084=>"000100011",
  11085=>"101010110",
  11086=>"011101111",
  11087=>"001011001",
  11088=>"101101111",
  11089=>"111110010",
  11090=>"101100011",
  11091=>"100111010",
  11092=>"001010000",
  11093=>"011101000",
  11094=>"101011001",
  11095=>"010011000",
  11096=>"001010001",
  11097=>"101000101",
  11098=>"111010110",
  11099=>"001101011",
  11100=>"010010010",
  11101=>"011010111",
  11102=>"101011110",
  11103=>"000110101",
  11104=>"101011111",
  11105=>"111010010",
  11106=>"101011010",
  11107=>"001000101",
  11108=>"101010001",
  11109=>"000001001",
  11110=>"000111111",
  11111=>"111101011",
  11112=>"011000110",
  11113=>"101010111",
  11114=>"101011100",
  11115=>"000100000",
  11116=>"000110101",
  11117=>"000011000",
  11118=>"011101110",
  11119=>"101010001",
  11120=>"110000111",
  11121=>"111111001",
  11122=>"111010101",
  11123=>"111100111",
  11124=>"010001110",
  11125=>"101010100",
  11126=>"110111011",
  11127=>"101011111",
  11128=>"011101111",
  11129=>"001000010",
  11130=>"011000011",
  11131=>"101010101",
  11132=>"000101011",
  11133=>"001000011",
  11134=>"011001100",
  11135=>"010100011",
  11136=>"010110011",
  11137=>"111110000",
  11138=>"111101001",
  11139=>"000100000",
  11140=>"111110000",
  11141=>"000100010",
  11142=>"010001100",
  11143=>"110000100",
  11144=>"111010010",
  11145=>"000001110",
  11146=>"000110010",
  11147=>"111011111",
  11148=>"111001010",
  11149=>"000100011",
  11150=>"001110001",
  11151=>"100110110",
  11152=>"111010111",
  11153=>"100010000",
  11154=>"001010011",
  11155=>"110100001",
  11156=>"000111101",
  11157=>"001011111",
  11158=>"001110000",
  11159=>"000010100",
  11160=>"000101000",
  11161=>"001001000",
  11162=>"101111111",
  11163=>"000010111",
  11164=>"000111110",
  11165=>"111001110",
  11166=>"110111101",
  11167=>"010100100",
  11168=>"010000111",
  11169=>"111000010",
  11170=>"000101100",
  11171=>"100100111",
  11172=>"110001101",
  11173=>"001000001",
  11174=>"001011110",
  11175=>"110000101",
  11176=>"001010111",
  11177=>"110110110",
  11178=>"001101101",
  11179=>"010110101",
  11180=>"101100111",
  11181=>"101001111",
  11182=>"000011011",
  11183=>"101101010",
  11184=>"111001101",
  11185=>"111110100",
  11186=>"111010000",
  11187=>"011000101",
  11188=>"000010001",
  11189=>"111100111",
  11190=>"010011010",
  11191=>"111001010",
  11192=>"110100011",
  11193=>"000011001",
  11194=>"011000100",
  11195=>"011100010",
  11196=>"101001011",
  11197=>"011110000",
  11198=>"010001010",
  11199=>"000001111",
  11200=>"011110010",
  11201=>"000110100",
  11202=>"100010111",
  11203=>"100010000",
  11204=>"111100011",
  11205=>"001000101",
  11206=>"111110101",
  11207=>"010101110",
  11208=>"011100100",
  11209=>"101101000",
  11210=>"111010100",
  11211=>"100100000",
  11212=>"011111011",
  11213=>"110000111",
  11214=>"110000011",
  11215=>"000110001",
  11216=>"011011101",
  11217=>"101110101",
  11218=>"001111001",
  11219=>"000011111",
  11220=>"001100111",
  11221=>"010000011",
  11222=>"111101111",
  11223=>"101010010",
  11224=>"000010110",
  11225=>"100111110",
  11226=>"101110101",
  11227=>"110011001",
  11228=>"111111111",
  11229=>"111111101",
  11230=>"110010110",
  11231=>"000000011",
  11232=>"001010010",
  11233=>"001111000",
  11234=>"001011111",
  11235=>"101100100",
  11236=>"111110010",
  11237=>"000111101",
  11238=>"110010010",
  11239=>"111111101",
  11240=>"100011111",
  11241=>"111011110",
  11242=>"001110000",
  11243=>"100001001",
  11244=>"000100111",
  11245=>"001100011",
  11246=>"000001111",
  11247=>"100111110",
  11248=>"001110100",
  11249=>"100111000",
  11250=>"101100011",
  11251=>"110011110",
  11252=>"011110001",
  11253=>"111000101",
  11254=>"111010010",
  11255=>"110111101",
  11256=>"101101111",
  11257=>"011101110",
  11258=>"000101101",
  11259=>"111000000",
  11260=>"011010010",
  11261=>"010111111",
  11262=>"001100111",
  11263=>"000101111",
  11264=>"001000100",
  11265=>"011101110",
  11266=>"001011010",
  11267=>"011110101",
  11268=>"101100000",
  11269=>"010011010",
  11270=>"000001011",
  11271=>"001100110",
  11272=>"101000010",
  11273=>"010100100",
  11274=>"010001000",
  11275=>"010100011",
  11276=>"100100010",
  11277=>"011101011",
  11278=>"011010000",
  11279=>"111001010",
  11280=>"101100101",
  11281=>"010111001",
  11282=>"001110100",
  11283=>"111101111",
  11284=>"000111001",
  11285=>"111010010",
  11286=>"100111011",
  11287=>"101000101",
  11288=>"100010100",
  11289=>"001000011",
  11290=>"000011101",
  11291=>"001011001",
  11292=>"100001111",
  11293=>"111111011",
  11294=>"010100100",
  11295=>"111111111",
  11296=>"011010100",
  11297=>"100111111",
  11298=>"000001110",
  11299=>"111000101",
  11300=>"001011000",
  11301=>"101100000",
  11302=>"100011101",
  11303=>"010100101",
  11304=>"100100100",
  11305=>"101000101",
  11306=>"001111101",
  11307=>"100111011",
  11308=>"101000100",
  11309=>"101110111",
  11310=>"000010011",
  11311=>"110011010",
  11312=>"011110000",
  11313=>"110001101",
  11314=>"100100011",
  11315=>"110011001",
  11316=>"011000110",
  11317=>"011100001",
  11318=>"110111011",
  11319=>"011001011",
  11320=>"011110111",
  11321=>"100101010",
  11322=>"010110100",
  11323=>"000011011",
  11324=>"000111011",
  11325=>"111011011",
  11326=>"000110110",
  11327=>"011101001",
  11328=>"001000100",
  11329=>"001010011",
  11330=>"101000100",
  11331=>"110111000",
  11332=>"111010110",
  11333=>"001111010",
  11334=>"111010100",
  11335=>"110000000",
  11336=>"001101001",
  11337=>"000100110",
  11338=>"001100001",
  11339=>"100111110",
  11340=>"011101001",
  11341=>"110011111",
  11342=>"011100001",
  11343=>"100110011",
  11344=>"101101101",
  11345=>"000101100",
  11346=>"100101111",
  11347=>"001101110",
  11348=>"000111011",
  11349=>"100010000",
  11350=>"000000110",
  11351=>"101010111",
  11352=>"011111111",
  11353=>"000110111",
  11354=>"011110010",
  11355=>"101101000",
  11356=>"010111100",
  11357=>"100110111",
  11358=>"101100010",
  11359=>"001000111",
  11360=>"010100101",
  11361=>"111101111",
  11362=>"101011111",
  11363=>"011001011",
  11364=>"111010001",
  11365=>"100011110",
  11366=>"010011100",
  11367=>"001001011",
  11368=>"110010101",
  11369=>"001111111",
  11370=>"011000011",
  11371=>"001111010",
  11372=>"110011100",
  11373=>"101111110",
  11374=>"100010011",
  11375=>"111110010",
  11376=>"111111000",
  11377=>"010111100",
  11378=>"100110011",
  11379=>"010100001",
  11380=>"010000011",
  11381=>"111000010",
  11382=>"101011100",
  11383=>"110110000",
  11384=>"110010010",
  11385=>"000010011",
  11386=>"001101101",
  11387=>"011100101",
  11388=>"101010000",
  11389=>"101011010",
  11390=>"010110000",
  11391=>"111110101",
  11392=>"100000010",
  11393=>"011011010",
  11394=>"010010110",
  11395=>"100101101",
  11396=>"011100110",
  11397=>"011011100",
  11398=>"111110111",
  11399=>"110011111",
  11400=>"000001111",
  11401=>"100010000",
  11402=>"100011101",
  11403=>"000110011",
  11404=>"101001100",
  11405=>"110100100",
  11406=>"001000001",
  11407=>"100000100",
  11408=>"101010011",
  11409=>"100010010",
  11410=>"010110010",
  11411=>"111010011",
  11412=>"010110010",
  11413=>"010000001",
  11414=>"001111100",
  11415=>"001011100",
  11416=>"010111010",
  11417=>"000011100",
  11418=>"001011000",
  11419=>"101011110",
  11420=>"001110101",
  11421=>"011100000",
  11422=>"011011010",
  11423=>"101110100",
  11424=>"010000010",
  11425=>"111110001",
  11426=>"111000101",
  11427=>"000001111",
  11428=>"111101001",
  11429=>"101110111",
  11430=>"110010000",
  11431=>"011001100",
  11432=>"010101100",
  11433=>"011010001",
  11434=>"010111100",
  11435=>"001001001",
  11436=>"000011111",
  11437=>"011100010",
  11438=>"101001000",
  11439=>"111101100",
  11440=>"010101111",
  11441=>"110010101",
  11442=>"000000110",
  11443=>"100010010",
  11444=>"001101000",
  11445=>"001110011",
  11446=>"110001101",
  11447=>"010111001",
  11448=>"110010011",
  11449=>"000110000",
  11450=>"111100001",
  11451=>"100111111",
  11452=>"111001110",
  11453=>"111010100",
  11454=>"100101110",
  11455=>"001011101",
  11456=>"111001110",
  11457=>"101000110",
  11458=>"000010101",
  11459=>"011011110",
  11460=>"101101100",
  11461=>"001111111",
  11462=>"101101110",
  11463=>"001100000",
  11464=>"011001010",
  11465=>"010111101",
  11466=>"001110100",
  11467=>"110000111",
  11468=>"000000001",
  11469=>"110111000",
  11470=>"001101000",
  11471=>"010100000",
  11472=>"011101010",
  11473=>"111001101",
  11474=>"001010000",
  11475=>"111111001",
  11476=>"110000111",
  11477=>"001100101",
  11478=>"110111000",
  11479=>"101100111",
  11480=>"001001100",
  11481=>"011010000",
  11482=>"000001000",
  11483=>"001001000",
  11484=>"110010011",
  11485=>"111101010",
  11486=>"110001110",
  11487=>"111010101",
  11488=>"100110111",
  11489=>"010011010",
  11490=>"011011110",
  11491=>"100101111",
  11492=>"001100010",
  11493=>"100001011",
  11494=>"100011110",
  11495=>"110011111",
  11496=>"011011000",
  11497=>"001111000",
  11498=>"011000000",
  11499=>"101101011",
  11500=>"001001101",
  11501=>"001000000",
  11502=>"001101100",
  11503=>"010110111",
  11504=>"111011011",
  11505=>"100111100",
  11506=>"010001001",
  11507=>"110000111",
  11508=>"110101100",
  11509=>"011101010",
  11510=>"110000111",
  11511=>"010000011",
  11512=>"101001110",
  11513=>"110110000",
  11514=>"110011110",
  11515=>"111110010",
  11516=>"010000000",
  11517=>"000111011",
  11518=>"000000110",
  11519=>"001111111",
  11520=>"101101000",
  11521=>"010110010",
  11522=>"110111110",
  11523=>"000100111",
  11524=>"100010001",
  11525=>"110110000",
  11526=>"001101011",
  11527=>"101010111",
  11528=>"000001000",
  11529=>"001010111",
  11530=>"110100000",
  11531=>"101011000",
  11532=>"000101100",
  11533=>"100011011",
  11534=>"000010000",
  11535=>"000110000",
  11536=>"111101101",
  11537=>"110101010",
  11538=>"000001110",
  11539=>"001100010",
  11540=>"001001111",
  11541=>"011001110",
  11542=>"010110010",
  11543=>"011100100",
  11544=>"010010100",
  11545=>"110101101",
  11546=>"110100100",
  11547=>"110011001",
  11548=>"011100101",
  11549=>"110001100",
  11550=>"110111010",
  11551=>"001111000",
  11552=>"000010001",
  11553=>"000011011",
  11554=>"101101010",
  11555=>"011001101",
  11556=>"000110010",
  11557=>"011111000",
  11558=>"101011101",
  11559=>"110101100",
  11560=>"101100100",
  11561=>"100101100",
  11562=>"100000010",
  11563=>"100001111",
  11564=>"011010010",
  11565=>"001010100",
  11566=>"101001111",
  11567=>"001011000",
  11568=>"011010000",
  11569=>"011010011",
  11570=>"100111111",
  11571=>"111000010",
  11572=>"110100001",
  11573=>"111011101",
  11574=>"000000000",
  11575=>"011100001",
  11576=>"000001100",
  11577=>"110011100",
  11578=>"111101001",
  11579=>"101000110",
  11580=>"111010110",
  11581=>"111011001",
  11582=>"111111100",
  11583=>"000101000",
  11584=>"000111010",
  11585=>"111100000",
  11586=>"011110000",
  11587=>"101001000",
  11588=>"000101010",
  11589=>"100011010",
  11590=>"010011010",
  11591=>"100011100",
  11592=>"000000110",
  11593=>"110000110",
  11594=>"010110001",
  11595=>"110011000",
  11596=>"101111011",
  11597=>"001011101",
  11598=>"101100100",
  11599=>"100110111",
  11600=>"011001000",
  11601=>"111011101",
  11602=>"000000000",
  11603=>"010001110",
  11604=>"011100010",
  11605=>"100100110",
  11606=>"000100101",
  11607=>"101101001",
  11608=>"110111011",
  11609=>"000110001",
  11610=>"100000111",
  11611=>"000001111",
  11612=>"110011001",
  11613=>"000010010",
  11614=>"110100111",
  11615=>"100000101",
  11616=>"001101100",
  11617=>"010000101",
  11618=>"010010101",
  11619=>"000111111",
  11620=>"000101011",
  11621=>"100011100",
  11622=>"010000011",
  11623=>"000010010",
  11624=>"001100000",
  11625=>"111001101",
  11626=>"111010100",
  11627=>"101010110",
  11628=>"101100001",
  11629=>"101111100",
  11630=>"111110111",
  11631=>"101001111",
  11632=>"001101101",
  11633=>"011101010",
  11634=>"011000101",
  11635=>"011101110",
  11636=>"110011001",
  11637=>"111000011",
  11638=>"001101001",
  11639=>"001110100",
  11640=>"001001011",
  11641=>"011110111",
  11642=>"001111101",
  11643=>"111101010",
  11644=>"111011011",
  11645=>"000101100",
  11646=>"010011100",
  11647=>"110101011",
  11648=>"110101011",
  11649=>"110100101",
  11650=>"100110000",
  11651=>"000001011",
  11652=>"011010001",
  11653=>"000100000",
  11654=>"011110010",
  11655=>"000010101",
  11656=>"000010010",
  11657=>"001100101",
  11658=>"100101100",
  11659=>"000111111",
  11660=>"011101011",
  11661=>"000010110",
  11662=>"000011100",
  11663=>"101000001",
  11664=>"111111111",
  11665=>"000001110",
  11666=>"110100011",
  11667=>"111010101",
  11668=>"011101010",
  11669=>"010110100",
  11670=>"000100101",
  11671=>"101101100",
  11672=>"111011000",
  11673=>"001100010",
  11674=>"001011100",
  11675=>"101110111",
  11676=>"100100100",
  11677=>"100011110",
  11678=>"111101000",
  11679=>"111000001",
  11680=>"101001000",
  11681=>"100010111",
  11682=>"100110100",
  11683=>"101000100",
  11684=>"110001011",
  11685=>"100101100",
  11686=>"110011000",
  11687=>"001100000",
  11688=>"100001101",
  11689=>"001111101",
  11690=>"110100010",
  11691=>"010100010",
  11692=>"011101110",
  11693=>"111110100",
  11694=>"010101001",
  11695=>"010110000",
  11696=>"000100101",
  11697=>"000100000",
  11698=>"100001101",
  11699=>"110000011",
  11700=>"110010111",
  11701=>"111010111",
  11702=>"110001010",
  11703=>"001110100",
  11704=>"011101100",
  11705=>"000011010",
  11706=>"011001000",
  11707=>"111000011",
  11708=>"100100111",
  11709=>"000010001",
  11710=>"101001001",
  11711=>"101000111",
  11712=>"110000001",
  11713=>"101000101",
  11714=>"100011101",
  11715=>"111000000",
  11716=>"111100001",
  11717=>"101001111",
  11718=>"010001111",
  11719=>"000000001",
  11720=>"001110101",
  11721=>"100100101",
  11722=>"000001001",
  11723=>"111101110",
  11724=>"111001100",
  11725=>"110111101",
  11726=>"100101111",
  11727=>"101100100",
  11728=>"100001111",
  11729=>"001100010",
  11730=>"110101001",
  11731=>"110110111",
  11732=>"101011111",
  11733=>"000000110",
  11734=>"010110001",
  11735=>"100101010",
  11736=>"011000011",
  11737=>"100110011",
  11738=>"010110011",
  11739=>"011110011",
  11740=>"100001111",
  11741=>"110100010",
  11742=>"111111101",
  11743=>"100101101",
  11744=>"111011011",
  11745=>"111100011",
  11746=>"110011101",
  11747=>"101101100",
  11748=>"000010111",
  11749=>"010011000",
  11750=>"101011001",
  11751=>"100000111",
  11752=>"111010010",
  11753=>"010110010",
  11754=>"001100000",
  11755=>"000011101",
  11756=>"011011100",
  11757=>"000100100",
  11758=>"101010110",
  11759=>"110010000",
  11760=>"101011010",
  11761=>"110011110",
  11762=>"010001011",
  11763=>"100001101",
  11764=>"111000000",
  11765=>"100000010",
  11766=>"010011111",
  11767=>"011010101",
  11768=>"011010011",
  11769=>"000110011",
  11770=>"100010111",
  11771=>"100111101",
  11772=>"101111111",
  11773=>"000111011",
  11774=>"000110100",
  11775=>"110101001",
  11776=>"001101110",
  11777=>"100101000",
  11778=>"000010101",
  11779=>"011111001",
  11780=>"100001111",
  11781=>"010100010",
  11782=>"000110000",
  11783=>"110111111",
  11784=>"000000001",
  11785=>"000101000",
  11786=>"001100100",
  11787=>"001010100",
  11788=>"111101110",
  11789=>"000101000",
  11790=>"110100001",
  11791=>"101000111",
  11792=>"001111110",
  11793=>"110110010",
  11794=>"000000000",
  11795=>"100011001",
  11796=>"100000011",
  11797=>"110001000",
  11798=>"011101001",
  11799=>"110000001",
  11800=>"010000101",
  11801=>"110101111",
  11802=>"000001011",
  11803=>"100011110",
  11804=>"011110100",
  11805=>"001111111",
  11806=>"101001111",
  11807=>"111111010",
  11808=>"001011000",
  11809=>"000111000",
  11810=>"001000111",
  11811=>"000001110",
  11812=>"110111010",
  11813=>"100111100",
  11814=>"100100010",
  11815=>"111101010",
  11816=>"100111110",
  11817=>"101101111",
  11818=>"101010011",
  11819=>"111011000",
  11820=>"000010010",
  11821=>"100100010",
  11822=>"110110110",
  11823=>"101101010",
  11824=>"010111100",
  11825=>"011011100",
  11826=>"100010111",
  11827=>"110010001",
  11828=>"000000011",
  11829=>"111001000",
  11830=>"100111001",
  11831=>"000010111",
  11832=>"101010100",
  11833=>"111011000",
  11834=>"100011010",
  11835=>"101101001",
  11836=>"101110001",
  11837=>"101111000",
  11838=>"010111001",
  11839=>"010100000",
  11840=>"000000100",
  11841=>"111011010",
  11842=>"010110111",
  11843=>"011000101",
  11844=>"000011110",
  11845=>"001001101",
  11846=>"100000011",
  11847=>"101110110",
  11848=>"010100111",
  11849=>"100101010",
  11850=>"010111100",
  11851=>"000010000",
  11852=>"110010100",
  11853=>"001011011",
  11854=>"010110101",
  11855=>"011111100",
  11856=>"110001011",
  11857=>"110000011",
  11858=>"111010000",
  11859=>"110010100",
  11860=>"101011000",
  11861=>"100100011",
  11862=>"010010010",
  11863=>"110000010",
  11864=>"111100111",
  11865=>"110100101",
  11866=>"001000001",
  11867=>"100101000",
  11868=>"110100100",
  11869=>"000101001",
  11870=>"110111111",
  11871=>"101110001",
  11872=>"011011000",
  11873=>"010110001",
  11874=>"100010110",
  11875=>"011100100",
  11876=>"011010110",
  11877=>"010000100",
  11878=>"001001011",
  11879=>"101010100",
  11880=>"011000001",
  11881=>"011111000",
  11882=>"111110010",
  11883=>"100100000",
  11884=>"110000011",
  11885=>"110010101",
  11886=>"010011111",
  11887=>"100100110",
  11888=>"011011011",
  11889=>"000010001",
  11890=>"111101011",
  11891=>"010110111",
  11892=>"100011010",
  11893=>"001000111",
  11894=>"000010110",
  11895=>"100010010",
  11896=>"001111001",
  11897=>"111000110",
  11898=>"101011000",
  11899=>"110111101",
  11900=>"101100100",
  11901=>"011010110",
  11902=>"110111011",
  11903=>"101000000",
  11904=>"111110100",
  11905=>"111101000",
  11906=>"000111001",
  11907=>"101011111",
  11908=>"101001100",
  11909=>"111010001",
  11910=>"111111111",
  11911=>"000101111",
  11912=>"100101101",
  11913=>"000000001",
  11914=>"011100111",
  11915=>"011001010",
  11916=>"000011000",
  11917=>"001000110",
  11918=>"010010110",
  11919=>"100110010",
  11920=>"100001101",
  11921=>"001010110",
  11922=>"110111011",
  11923=>"111111111",
  11924=>"010010000",
  11925=>"110010101",
  11926=>"010000111",
  11927=>"011100010",
  11928=>"100110001",
  11929=>"010101101",
  11930=>"011110110",
  11931=>"011011101",
  11932=>"010111011",
  11933=>"001111000",
  11934=>"100101111",
  11935=>"110110101",
  11936=>"011010010",
  11937=>"001110100",
  11938=>"101111111",
  11939=>"100100111",
  11940=>"110001000",
  11941=>"010010000",
  11942=>"100100011",
  11943=>"000100000",
  11944=>"100100010",
  11945=>"100001011",
  11946=>"101100000",
  11947=>"010101010",
  11948=>"000110001",
  11949=>"100101011",
  11950=>"010001111",
  11951=>"111101111",
  11952=>"011110001",
  11953=>"100110100",
  11954=>"100111010",
  11955=>"000100101",
  11956=>"110001111",
  11957=>"011110101",
  11958=>"110111000",
  11959=>"000111001",
  11960=>"001101110",
  11961=>"110101100",
  11962=>"101110110",
  11963=>"010011111",
  11964=>"011100001",
  11965=>"110001010",
  11966=>"001010111",
  11967=>"000000011",
  11968=>"110010001",
  11969=>"001110010",
  11970=>"011100011",
  11971=>"010100010",
  11972=>"100111000",
  11973=>"110101110",
  11974=>"100110110",
  11975=>"001100111",
  11976=>"000100110",
  11977=>"101100011",
  11978=>"010101011",
  11979=>"110101011",
  11980=>"011000010",
  11981=>"000010101",
  11982=>"011110000",
  11983=>"000101110",
  11984=>"110000110",
  11985=>"100100001",
  11986=>"001110001",
  11987=>"000010001",
  11988=>"011110001",
  11989=>"001110111",
  11990=>"000100000",
  11991=>"011000000",
  11992=>"010111011",
  11993=>"010010011",
  11994=>"110000100",
  11995=>"111110000",
  11996=>"000111011",
  11997=>"100010111",
  11998=>"101000101",
  11999=>"010011010",
  12000=>"101011001",
  12001=>"000111100",
  12002=>"011001011",
  12003=>"000110110",
  12004=>"101011000",
  12005=>"001101111",
  12006=>"110111100",
  12007=>"001110011",
  12008=>"000110001",
  12009=>"101101010",
  12010=>"110111000",
  12011=>"110011010",
  12012=>"111010010",
  12013=>"100100011",
  12014=>"110100010",
  12015=>"111001011",
  12016=>"000011111",
  12017=>"101010110",
  12018=>"011011010",
  12019=>"111011111",
  12020=>"011001010",
  12021=>"110100111",
  12022=>"101001111",
  12023=>"000000110",
  12024=>"010100100",
  12025=>"000100101",
  12026=>"001111010",
  12027=>"101011000",
  12028=>"101001101",
  12029=>"100100000",
  12030=>"001000000",
  12031=>"110110001",
  12032=>"010110000",
  12033=>"010000000",
  12034=>"110101001",
  12035=>"001100011",
  12036=>"011100011",
  12037=>"001110101",
  12038=>"101010101",
  12039=>"011010110",
  12040=>"001111100",
  12041=>"001100111",
  12042=>"100111011",
  12043=>"110110111",
  12044=>"100000100",
  12045=>"110011110",
  12046=>"000111100",
  12047=>"000111111",
  12048=>"001101111",
  12049=>"000111110",
  12050=>"001111100",
  12051=>"001110111",
  12052=>"100011100",
  12053=>"101100001",
  12054=>"100101100",
  12055=>"011101010",
  12056=>"111000010",
  12057=>"010011110",
  12058=>"001001010",
  12059=>"101111101",
  12060=>"010010001",
  12061=>"001011100",
  12062=>"100100100",
  12063=>"010111011",
  12064=>"001100101",
  12065=>"101110111",
  12066=>"100011111",
  12067=>"011001011",
  12068=>"010000001",
  12069=>"110110111",
  12070=>"000010000",
  12071=>"000111011",
  12072=>"001001111",
  12073=>"001100010",
  12074=>"100000101",
  12075=>"001011011",
  12076=>"010111011",
  12077=>"100000101",
  12078=>"101001100",
  12079=>"111011100",
  12080=>"011000000",
  12081=>"111001010",
  12082=>"011000010",
  12083=>"111000011",
  12084=>"000111100",
  12085=>"010010111",
  12086=>"101101001",
  12087=>"011101010",
  12088=>"100101001",
  12089=>"010111011",
  12090=>"100110000",
  12091=>"101011111",
  12092=>"100011100",
  12093=>"011010000",
  12094=>"010100010",
  12095=>"000000011",
  12096=>"101011010",
  12097=>"001010101",
  12098=>"011111100",
  12099=>"001100111",
  12100=>"011101110",
  12101=>"011110000",
  12102=>"000011110",
  12103=>"101001101",
  12104=>"001100010",
  12105=>"101100011",
  12106=>"101111110",
  12107=>"000010111",
  12108=>"001111000",
  12109=>"111100000",
  12110=>"110011101",
  12111=>"001001110",
  12112=>"001000011",
  12113=>"011010100",
  12114=>"010000001",
  12115=>"111000010",
  12116=>"000010101",
  12117=>"010011100",
  12118=>"000100101",
  12119=>"111111100",
  12120=>"110110100",
  12121=>"100000100",
  12122=>"111010010",
  12123=>"110011111",
  12124=>"010000010",
  12125=>"101001110",
  12126=>"100011011",
  12127=>"000000010",
  12128=>"101011010",
  12129=>"011101010",
  12130=>"011100101",
  12131=>"110101000",
  12132=>"010111010",
  12133=>"111010100",
  12134=>"001110011",
  12135=>"100011001",
  12136=>"100101000",
  12137=>"101000000",
  12138=>"100000101",
  12139=>"111100101",
  12140=>"101000011",
  12141=>"011001000",
  12142=>"101110101",
  12143=>"101110101",
  12144=>"100110001",
  12145=>"011011101",
  12146=>"010010000",
  12147=>"100011010",
  12148=>"101010010",
  12149=>"010010000",
  12150=>"110110011",
  12151=>"100011100",
  12152=>"101011111",
  12153=>"000111110",
  12154=>"111111011",
  12155=>"101101101",
  12156=>"010011010",
  12157=>"001001010",
  12158=>"011100000",
  12159=>"010101101",
  12160=>"000111111",
  12161=>"001100111",
  12162=>"101111000",
  12163=>"010011000",
  12164=>"000110101",
  12165=>"110001000",
  12166=>"000000000",
  12167=>"001101100",
  12168=>"110001110",
  12169=>"101001010",
  12170=>"001111010",
  12171=>"110011111",
  12172=>"010101000",
  12173=>"101000110",
  12174=>"110110010",
  12175=>"001110101",
  12176=>"001001000",
  12177=>"111101001",
  12178=>"001100011",
  12179=>"010011101",
  12180=>"010110011",
  12181=>"011001100",
  12182=>"001011111",
  12183=>"011001011",
  12184=>"100110011",
  12185=>"011001011",
  12186=>"101110010",
  12187=>"100001011",
  12188=>"010101000",
  12189=>"011010100",
  12190=>"101000010",
  12191=>"111101101",
  12192=>"000100101",
  12193=>"111110101",
  12194=>"000010011",
  12195=>"011101011",
  12196=>"001001001",
  12197=>"101010111",
  12198=>"100100100",
  12199=>"000111111",
  12200=>"010100111",
  12201=>"000001011",
  12202=>"001110110",
  12203=>"001001110",
  12204=>"001001100",
  12205=>"000011010",
  12206=>"110100111",
  12207=>"000111010",
  12208=>"010001010",
  12209=>"100111111",
  12210=>"101010101",
  12211=>"101101110",
  12212=>"001100101",
  12213=>"110010001",
  12214=>"010010001",
  12215=>"010001011",
  12216=>"010011001",
  12217=>"101110101",
  12218=>"001101011",
  12219=>"110111111",
  12220=>"100001110",
  12221=>"010011100",
  12222=>"111010100",
  12223=>"100101101",
  12224=>"001100001",
  12225=>"001000100",
  12226=>"001100110",
  12227=>"011101011",
  12228=>"000000110",
  12229=>"011110101",
  12230=>"110101010",
  12231=>"111000010",
  12232=>"001110110",
  12233=>"101111111",
  12234=>"110100111",
  12235=>"110101101",
  12236=>"110011000",
  12237=>"010111100",
  12238=>"011110001",
  12239=>"101101101",
  12240=>"111010000",
  12241=>"100000001",
  12242=>"101101111",
  12243=>"001001100",
  12244=>"011110111",
  12245=>"001100010",
  12246=>"101010010",
  12247=>"001010001",
  12248=>"011111111",
  12249=>"100111101",
  12250=>"101011001",
  12251=>"101111001",
  12252=>"101111011",
  12253=>"111100010",
  12254=>"000110110",
  12255=>"100001011",
  12256=>"110111110",
  12257=>"111011101",
  12258=>"001011101",
  12259=>"000110010",
  12260=>"000001010",
  12261=>"101101111",
  12262=>"001111010",
  12263=>"000101100",
  12264=>"000100001",
  12265=>"010110010",
  12266=>"001101000",
  12267=>"000011010",
  12268=>"101100000",
  12269=>"010001000",
  12270=>"000000111",
  12271=>"100001110",
  12272=>"000110010",
  12273=>"100011110",
  12274=>"010111001",
  12275=>"111100001",
  12276=>"101101000",
  12277=>"001011100",
  12278=>"000000011",
  12279=>"001010111",
  12280=>"010100001",
  12281=>"011000100",
  12282=>"000000100",
  12283=>"001111101",
  12284=>"011101111",
  12285=>"010110011",
  12286=>"010101100",
  12287=>"010100111",
  12288=>"110100110",
  12289=>"110100110",
  12290=>"010000100",
  12291=>"010100010",
  12292=>"001111101",
  12293=>"001110011",
  12294=>"011000101",
  12295=>"000010001",
  12296=>"110101100",
  12297=>"100011010",
  12298=>"000110110",
  12299=>"101100011",
  12300=>"110110110",
  12301=>"100101001",
  12302=>"100100000",
  12303=>"100101100",
  12304=>"000010111",
  12305=>"110010000",
  12306=>"010000000",
  12307=>"010010000",
  12308=>"000010011",
  12309=>"000111010",
  12310=>"001110010",
  12311=>"110001001",
  12312=>"111101110",
  12313=>"100011100",
  12314=>"100000101",
  12315=>"111011101",
  12316=>"110101000",
  12317=>"111010001",
  12318=>"001111100",
  12319=>"010001000",
  12320=>"110000011",
  12321=>"000010001",
  12322=>"111101010",
  12323=>"101010001",
  12324=>"010001010",
  12325=>"101110111",
  12326=>"101111101",
  12327=>"100011100",
  12328=>"011101111",
  12329=>"000011111",
  12330=>"101000011",
  12331=>"101010111",
  12332=>"101011010",
  12333=>"111100000",
  12334=>"000000000",
  12335=>"100101110",
  12336=>"001000111",
  12337=>"111100000",
  12338=>"101100110",
  12339=>"000110100",
  12340=>"101001010",
  12341=>"000001000",
  12342=>"000100000",
  12343=>"001101111",
  12344=>"000001010",
  12345=>"000001000",
  12346=>"101010010",
  12347=>"001001110",
  12348=>"111010101",
  12349=>"111000101",
  12350=>"010011001",
  12351=>"011011011",
  12352=>"001110100",
  12353=>"100100000",
  12354=>"000100001",
  12355=>"010111111",
  12356=>"111111000",
  12357=>"001011010",
  12358=>"001000100",
  12359=>"010001000",
  12360=>"000110011",
  12361=>"000000010",
  12362=>"011001110",
  12363=>"001101010",
  12364=>"000100100",
  12365=>"001100111",
  12366=>"100110001",
  12367=>"101011000",
  12368=>"100100001",
  12369=>"000100011",
  12370=>"100100001",
  12371=>"000000111",
  12372=>"000111001",
  12373=>"110010000",
  12374=>"011100110",
  12375=>"010010011",
  12376=>"100010001",
  12377=>"010000010",
  12378=>"011101100",
  12379=>"000100011",
  12380=>"110001111",
  12381=>"100000011",
  12382=>"000001000",
  12383=>"001001110",
  12384=>"010111011",
  12385=>"001011010",
  12386=>"000010101",
  12387=>"111000010",
  12388=>"000010111",
  12389=>"101101100",
  12390=>"101000001",
  12391=>"000101100",
  12392=>"001101100",
  12393=>"011101011",
  12394=>"100111001",
  12395=>"001001100",
  12396=>"000111000",
  12397=>"110110101",
  12398=>"010000101",
  12399=>"111110100",
  12400=>"101101010",
  12401=>"001010001",
  12402=>"011110100",
  12403=>"000111101",
  12404=>"011110010",
  12405=>"100011101",
  12406=>"001011111",
  12407=>"001000100",
  12408=>"000000001",
  12409=>"000110110",
  12410=>"011100101",
  12411=>"101001101",
  12412=>"110110011",
  12413=>"111100100",
  12414=>"011010000",
  12415=>"111001101",
  12416=>"110100110",
  12417=>"001111110",
  12418=>"010000111",
  12419=>"100101101",
  12420=>"100001100",
  12421=>"000100001",
  12422=>"010101110",
  12423=>"100000110",
  12424=>"000011011",
  12425=>"100000100",
  12426=>"110001000",
  12427=>"100010010",
  12428=>"000111000",
  12429=>"000000101",
  12430=>"111001001",
  12431=>"010001110",
  12432=>"010100000",
  12433=>"111011111",
  12434=>"111101111",
  12435=>"110110001",
  12436=>"100111000",
  12437=>"100011110",
  12438=>"111011000",
  12439=>"011110100",
  12440=>"010100110",
  12441=>"010000000",
  12442=>"111001111",
  12443=>"100101010",
  12444=>"001010110",
  12445=>"001000100",
  12446=>"110010011",
  12447=>"111001100",
  12448=>"111011111",
  12449=>"110010001",
  12450=>"101001001",
  12451=>"010111010",
  12452=>"101100100",
  12453=>"110111100",
  12454=>"000100011",
  12455=>"110010010",
  12456=>"001000111",
  12457=>"101001101",
  12458=>"111111011",
  12459=>"010001001",
  12460=>"001000101",
  12461=>"000011000",
  12462=>"110001110",
  12463=>"011101001",
  12464=>"001010001",
  12465=>"111010000",
  12466=>"011011111",
  12467=>"000011111",
  12468=>"101110000",
  12469=>"110011001",
  12470=>"100110010",
  12471=>"010110110",
  12472=>"000001001",
  12473=>"100100110",
  12474=>"100111011",
  12475=>"000001101",
  12476=>"101001111",
  12477=>"110001000",
  12478=>"001111001",
  12479=>"011100110",
  12480=>"100010110",
  12481=>"111100010",
  12482=>"000111111",
  12483=>"010010100",
  12484=>"010110110",
  12485=>"000010001",
  12486=>"101101011",
  12487=>"010110000",
  12488=>"011010010",
  12489=>"100111100",
  12490=>"110001001",
  12491=>"101100110",
  12492=>"100000100",
  12493=>"101000011",
  12494=>"001010110",
  12495=>"110000000",
  12496=>"001110111",
  12497=>"001100110",
  12498=>"100000101",
  12499=>"110001101",
  12500=>"010111011",
  12501=>"011111101",
  12502=>"110101001",
  12503=>"100001101",
  12504=>"101011110",
  12505=>"010001010",
  12506=>"000111111",
  12507=>"110111110",
  12508=>"011000101",
  12509=>"010000101",
  12510=>"000000011",
  12511=>"111011001",
  12512=>"110010011",
  12513=>"100101011",
  12514=>"111000000",
  12515=>"010000111",
  12516=>"100001111",
  12517=>"010010101",
  12518=>"011010011",
  12519=>"100111001",
  12520=>"110100001",
  12521=>"000101100",
  12522=>"010001101",
  12523=>"001001101",
  12524=>"100000000",
  12525=>"001000110",
  12526=>"010001010",
  12527=>"010001000",
  12528=>"011010010",
  12529=>"100011101",
  12530=>"010100100",
  12531=>"001111101",
  12532=>"111110011",
  12533=>"001011111",
  12534=>"101010100",
  12535=>"000111110",
  12536=>"011100111",
  12537=>"001000001",
  12538=>"100111111",
  12539=>"000100100",
  12540=>"101111111",
  12541=>"110000011",
  12542=>"100000011",
  12543=>"110110011",
  12544=>"001001000",
  12545=>"100011001",
  12546=>"101101110",
  12547=>"011000000",
  12548=>"111001001",
  12549=>"101100000",
  12550=>"011011011",
  12551=>"010011010",
  12552=>"111010001",
  12553=>"000000001",
  12554=>"011010000",
  12555=>"011101011",
  12556=>"110100110",
  12557=>"001100110",
  12558=>"101000001",
  12559=>"101101111",
  12560=>"001101000",
  12561=>"100000001",
  12562=>"000101011",
  12563=>"110111111",
  12564=>"111111111",
  12565=>"010000011",
  12566=>"000011111",
  12567=>"100010101",
  12568=>"100100101",
  12569=>"011001101",
  12570=>"110001110",
  12571=>"101001110",
  12572=>"001011101",
  12573=>"101010101",
  12574=>"010111011",
  12575=>"001000001",
  12576=>"100100000",
  12577=>"100100001",
  12578=>"100100000",
  12579=>"001110110",
  12580=>"111111011",
  12581=>"011111000",
  12582=>"100011001",
  12583=>"001101010",
  12584=>"001111000",
  12585=>"011111111",
  12586=>"101111001",
  12587=>"111100111",
  12588=>"110010001",
  12589=>"111011100",
  12590=>"100101100",
  12591=>"101111101",
  12592=>"100100000",
  12593=>"101110000",
  12594=>"001001100",
  12595=>"011010000",
  12596=>"100100000",
  12597=>"000000100",
  12598=>"000111101",
  12599=>"101110111",
  12600=>"100011001",
  12601=>"100100000",
  12602=>"100101111",
  12603=>"101001100",
  12604=>"000011101",
  12605=>"101100010",
  12606=>"100011100",
  12607=>"001010001",
  12608=>"101011011",
  12609=>"011111111",
  12610=>"000110001",
  12611=>"000100001",
  12612=>"000111100",
  12613=>"010001010",
  12614=>"101001101",
  12615=>"100001100",
  12616=>"010110110",
  12617=>"000110001",
  12618=>"110100110",
  12619=>"001111100",
  12620=>"011000111",
  12621=>"110010110",
  12622=>"111000011",
  12623=>"110110100",
  12624=>"101111101",
  12625=>"011010000",
  12626=>"000001101",
  12627=>"110100100",
  12628=>"100100000",
  12629=>"100001011",
  12630=>"001101000",
  12631=>"000000010",
  12632=>"000000111",
  12633=>"100101001",
  12634=>"100010110",
  12635=>"000111000",
  12636=>"101000010",
  12637=>"011110001",
  12638=>"010101111",
  12639=>"100110111",
  12640=>"000000000",
  12641=>"010111001",
  12642=>"000111111",
  12643=>"000000001",
  12644=>"110011010",
  12645=>"010010001",
  12646=>"001111100",
  12647=>"111010011",
  12648=>"001001011",
  12649=>"000000000",
  12650=>"101010101",
  12651=>"001010111",
  12652=>"010101000",
  12653=>"110011110",
  12654=>"100111110",
  12655=>"101111101",
  12656=>"000100101",
  12657=>"010010001",
  12658=>"101111001",
  12659=>"101110010",
  12660=>"011100011",
  12661=>"010110000",
  12662=>"001101110",
  12663=>"010001011",
  12664=>"011001100",
  12665=>"111111100",
  12666=>"110111011",
  12667=>"011100110",
  12668=>"010000001",
  12669=>"010000000",
  12670=>"011110101",
  12671=>"000110011",
  12672=>"111100111",
  12673=>"111110001",
  12674=>"101010110",
  12675=>"111111011",
  12676=>"110001101",
  12677=>"101101110",
  12678=>"101101010",
  12679=>"010101000",
  12680=>"100111111",
  12681=>"100010111",
  12682=>"110111010",
  12683=>"011010011",
  12684=>"101111010",
  12685=>"111001001",
  12686=>"000000000",
  12687=>"011110001",
  12688=>"001111111",
  12689=>"010010101",
  12690=>"000101000",
  12691=>"111111111",
  12692=>"000010000",
  12693=>"111000001",
  12694=>"111111011",
  12695=>"101000110",
  12696=>"110111011",
  12697=>"001010001",
  12698=>"011111100",
  12699=>"010010111",
  12700=>"011000001",
  12701=>"101110011",
  12702=>"001111100",
  12703=>"111100010",
  12704=>"001001111",
  12705=>"100001100",
  12706=>"000110010",
  12707=>"011110010",
  12708=>"001110101",
  12709=>"001101111",
  12710=>"000010011",
  12711=>"001110000",
  12712=>"100111001",
  12713=>"001100001",
  12714=>"011001010",
  12715=>"001111001",
  12716=>"000011011",
  12717=>"110001111",
  12718=>"111001001",
  12719=>"000000010",
  12720=>"011001010",
  12721=>"011111100",
  12722=>"010011001",
  12723=>"100010001",
  12724=>"000101100",
  12725=>"010001100",
  12726=>"011111001",
  12727=>"001110001",
  12728=>"100010101",
  12729=>"100000001",
  12730=>"000110110",
  12731=>"000101111",
  12732=>"010110110",
  12733=>"111100110",
  12734=>"111000111",
  12735=>"111010101",
  12736=>"110010000",
  12737=>"110110000",
  12738=>"111001101",
  12739=>"111001100",
  12740=>"100000000",
  12741=>"110110110",
  12742=>"010111010",
  12743=>"010101010",
  12744=>"000111100",
  12745=>"111000101",
  12746=>"011000101",
  12747=>"101111001",
  12748=>"011011110",
  12749=>"010011110",
  12750=>"000000100",
  12751=>"100000000",
  12752=>"001001010",
  12753=>"011011011",
  12754=>"111010000",
  12755=>"010111000",
  12756=>"001111100",
  12757=>"001000000",
  12758=>"111101111",
  12759=>"001110111",
  12760=>"011000101",
  12761=>"110100010",
  12762=>"000111000",
  12763=>"100000001",
  12764=>"100011111",
  12765=>"111010011",
  12766=>"001001110",
  12767=>"101101100",
  12768=>"110011110",
  12769=>"101101010",
  12770=>"010010101",
  12771=>"001010000",
  12772=>"000000111",
  12773=>"001111100",
  12774=>"001011101",
  12775=>"001101111",
  12776=>"011000011",
  12777=>"110010110",
  12778=>"110000000",
  12779=>"000011110",
  12780=>"000001001",
  12781=>"101101110",
  12782=>"000100001",
  12783=>"001000000",
  12784=>"011001001",
  12785=>"110100001",
  12786=>"001000010",
  12787=>"000101110",
  12788=>"110010101",
  12789=>"001110101",
  12790=>"101110010",
  12791=>"100101100",
  12792=>"110011011",
  12793=>"111110001",
  12794=>"111001110",
  12795=>"110100110",
  12796=>"101011101",
  12797=>"011100011",
  12798=>"000011111",
  12799=>"001111101",
  12800=>"000101010",
  12801=>"000111100",
  12802=>"110010100",
  12803=>"000010000",
  12804=>"010111011",
  12805=>"101011000",
  12806=>"101111000",
  12807=>"101011111",
  12808=>"010001000",
  12809=>"011111001",
  12810=>"111100110",
  12811=>"001111100",
  12812=>"001110101",
  12813=>"010001000",
  12814=>"000111011",
  12815=>"011000100",
  12816=>"010000001",
  12817=>"001001111",
  12818=>"111110010",
  12819=>"110101000",
  12820=>"001010000",
  12821=>"100111000",
  12822=>"111010110",
  12823=>"010001101",
  12824=>"010011000",
  12825=>"010100011",
  12826=>"001001010",
  12827=>"011100000",
  12828=>"010110110",
  12829=>"100110101",
  12830=>"000011011",
  12831=>"101100011",
  12832=>"010101101",
  12833=>"011010000",
  12834=>"000011001",
  12835=>"001010010",
  12836=>"111110000",
  12837=>"010100010",
  12838=>"111100000",
  12839=>"001101000",
  12840=>"101111101",
  12841=>"001000011",
  12842=>"000101101",
  12843=>"000110010",
  12844=>"101110111",
  12845=>"000110011",
  12846=>"100001101",
  12847=>"110011100",
  12848=>"110010011",
  12849=>"111010101",
  12850=>"001000111",
  12851=>"110110111",
  12852=>"001011111",
  12853=>"001110000",
  12854=>"110100001",
  12855=>"000000000",
  12856=>"111010101",
  12857=>"100101110",
  12858=>"000100011",
  12859=>"110111100",
  12860=>"101101111",
  12861=>"111011000",
  12862=>"111111111",
  12863=>"000001001",
  12864=>"101000101",
  12865=>"001000110",
  12866=>"010001110",
  12867=>"011000110",
  12868=>"111100010",
  12869=>"101100001",
  12870=>"000001011",
  12871=>"011010100",
  12872=>"110000111",
  12873=>"001111011",
  12874=>"101111010",
  12875=>"110101001",
  12876=>"011011111",
  12877=>"101011110",
  12878=>"001110100",
  12879=>"111000010",
  12880=>"010110001",
  12881=>"101001010",
  12882=>"111110001",
  12883=>"100111001",
  12884=>"011011110",
  12885=>"000101101",
  12886=>"111110001",
  12887=>"100011100",
  12888=>"001010111",
  12889=>"000111110",
  12890=>"111110011",
  12891=>"010111100",
  12892=>"100001001",
  12893=>"101000101",
  12894=>"101100100",
  12895=>"010010001",
  12896=>"001110111",
  12897=>"110111001",
  12898=>"101011011",
  12899=>"100000000",
  12900=>"110011000",
  12901=>"010010010",
  12902=>"101110001",
  12903=>"000110111",
  12904=>"101110110",
  12905=>"000001010",
  12906=>"010111001",
  12907=>"001110111",
  12908=>"101001011",
  12909=>"101110011",
  12910=>"011001111",
  12911=>"111001011",
  12912=>"110111011",
  12913=>"001011111",
  12914=>"111000111",
  12915=>"000001110",
  12916=>"111100010",
  12917=>"000001110",
  12918=>"000000011",
  12919=>"010111100",
  12920=>"001100111",
  12921=>"000110000",
  12922=>"100010011",
  12923=>"011000010",
  12924=>"111000100",
  12925=>"100101001",
  12926=>"011011011",
  12927=>"100110000",
  12928=>"110111111",
  12929=>"000011001",
  12930=>"101101010",
  12931=>"000010000",
  12932=>"100010110",
  12933=>"100111101",
  12934=>"111110000",
  12935=>"011000111",
  12936=>"001011101",
  12937=>"000011011",
  12938=>"000010000",
  12939=>"010001011",
  12940=>"110100010",
  12941=>"011111111",
  12942=>"101000111",
  12943=>"001110001",
  12944=>"000101111",
  12945=>"011000111",
  12946=>"010010111",
  12947=>"010000000",
  12948=>"100000001",
  12949=>"101000000",
  12950=>"000010110",
  12951=>"001000100",
  12952=>"011100011",
  12953=>"011110110",
  12954=>"100010110",
  12955=>"011111111",
  12956=>"011001011",
  12957=>"110100110",
  12958=>"101001001",
  12959=>"100111010",
  12960=>"010101100",
  12961=>"011010011",
  12962=>"111001001",
  12963=>"001111000",
  12964=>"010101000",
  12965=>"111110000",
  12966=>"010011110",
  12967=>"110101101",
  12968=>"100010101",
  12969=>"000000111",
  12970=>"100101100",
  12971=>"100111111",
  12972=>"101110100",
  12973=>"111111001",
  12974=>"101011011",
  12975=>"010101100",
  12976=>"111111110",
  12977=>"001001111",
  12978=>"100011100",
  12979=>"010100000",
  12980=>"101100001",
  12981=>"101111110",
  12982=>"110111010",
  12983=>"101111001",
  12984=>"110000001",
  12985=>"111000011",
  12986=>"011001111",
  12987=>"101110101",
  12988=>"000011001",
  12989=>"001011101",
  12990=>"000110000",
  12991=>"011011001",
  12992=>"111110111",
  12993=>"011000100",
  12994=>"110011100",
  12995=>"000101011",
  12996=>"000010100",
  12997=>"111110110",
  12998=>"001111000",
  12999=>"111100000",
  13000=>"111010101",
  13001=>"001101000",
  13002=>"001001011",
  13003=>"100011011",
  13004=>"110101101",
  13005=>"000111101",
  13006=>"000000000",
  13007=>"010110000",
  13008=>"110001111",
  13009=>"011110001",
  13010=>"111110001",
  13011=>"000001001",
  13012=>"111000010",
  13013=>"010101000",
  13014=>"111001010",
  13015=>"000110010",
  13016=>"110011010",
  13017=>"001111011",
  13018=>"001001111",
  13019=>"111010011",
  13020=>"000110100",
  13021=>"111110100",
  13022=>"010001110",
  13023=>"100000100",
  13024=>"011001011",
  13025=>"001100110",
  13026=>"100100010",
  13027=>"101011011",
  13028=>"101110101",
  13029=>"100010001",
  13030=>"010101000",
  13031=>"010010101",
  13032=>"001001000",
  13033=>"010101000",
  13034=>"100101101",
  13035=>"000111010",
  13036=>"000011000",
  13037=>"100011010",
  13038=>"010011010",
  13039=>"100011010",
  13040=>"011011001",
  13041=>"011010100",
  13042=>"100100010",
  13043=>"100001111",
  13044=>"100111101",
  13045=>"001110110",
  13046=>"000000011",
  13047=>"111010011",
  13048=>"000110101",
  13049=>"101100111",
  13050=>"101011011",
  13051=>"000100000",
  13052=>"000010111",
  13053=>"111001111",
  13054=>"010011010",
  13055=>"010101010",
  13056=>"101111000",
  13057=>"000111111",
  13058=>"101111111",
  13059=>"010000000",
  13060=>"001001010",
  13061=>"010000110",
  13062=>"011101110",
  13063=>"100111000",
  13064=>"101011110",
  13065=>"101101101",
  13066=>"001100111",
  13067=>"000100011",
  13068=>"000100011",
  13069=>"100111000",
  13070=>"110000110",
  13071=>"100110000",
  13072=>"010011011",
  13073=>"010001011",
  13074=>"101100100",
  13075=>"111011011",
  13076=>"001001000",
  13077=>"001010011",
  13078=>"011110111",
  13079=>"001101100",
  13080=>"111001111",
  13081=>"010000101",
  13082=>"010001101",
  13083=>"100100101",
  13084=>"000101011",
  13085=>"000100000",
  13086=>"001000000",
  13087=>"111001111",
  13088=>"010001000",
  13089=>"101010010",
  13090=>"010110000",
  13091=>"100000100",
  13092=>"000011010",
  13093=>"001111010",
  13094=>"111100000",
  13095=>"011101010",
  13096=>"111001011",
  13097=>"000101000",
  13098=>"111111111",
  13099=>"001001001",
  13100=>"111010001",
  13101=>"000101101",
  13102=>"011010101",
  13103=>"100100111",
  13104=>"101011010",
  13105=>"110011011",
  13106=>"010000110",
  13107=>"101111000",
  13108=>"100111010",
  13109=>"011101000",
  13110=>"110100110",
  13111=>"010111111",
  13112=>"010010010",
  13113=>"111011011",
  13114=>"000000110",
  13115=>"101001111",
  13116=>"110010111",
  13117=>"011000011",
  13118=>"110010001",
  13119=>"110011000",
  13120=>"010001110",
  13121=>"001001000",
  13122=>"110000010",
  13123=>"010000000",
  13124=>"010001111",
  13125=>"010101100",
  13126=>"011011111",
  13127=>"001111101",
  13128=>"110010000",
  13129=>"111011100",
  13130=>"000001011",
  13131=>"111010011",
  13132=>"000000100",
  13133=>"100010101",
  13134=>"000100111",
  13135=>"111111100",
  13136=>"010001111",
  13137=>"100010110",
  13138=>"001111100",
  13139=>"110100000",
  13140=>"101000011",
  13141=>"001001010",
  13142=>"101110000",
  13143=>"101001101",
  13144=>"100110111",
  13145=>"010111000",
  13146=>"011000110",
  13147=>"010110001",
  13148=>"011111010",
  13149=>"111111101",
  13150=>"101111111",
  13151=>"111000100",
  13152=>"011101010",
  13153=>"100011110",
  13154=>"101000000",
  13155=>"001110100",
  13156=>"010101110",
  13157=>"110011011",
  13158=>"110100100",
  13159=>"010101111",
  13160=>"000000101",
  13161=>"001111110",
  13162=>"010010101",
  13163=>"010101010",
  13164=>"101101011",
  13165=>"111010100",
  13166=>"010100110",
  13167=>"111001100",
  13168=>"111111110",
  13169=>"100000000",
  13170=>"100100100",
  13171=>"101010010",
  13172=>"101000101",
  13173=>"011101011",
  13174=>"010110000",
  13175=>"100110111",
  13176=>"111000010",
  13177=>"011101001",
  13178=>"110111100",
  13179=>"001010100",
  13180=>"000000000",
  13181=>"011000000",
  13182=>"001001000",
  13183=>"101110011",
  13184=>"000010100",
  13185=>"011011000",
  13186=>"101010010",
  13187=>"110111100",
  13188=>"111000010",
  13189=>"111011100",
  13190=>"001011000",
  13191=>"010110011",
  13192=>"001000000",
  13193=>"100100100",
  13194=>"010110000",
  13195=>"000110000",
  13196=>"101011010",
  13197=>"101011010",
  13198=>"111110001",
  13199=>"000000011",
  13200=>"001001001",
  13201=>"000001110",
  13202=>"100100111",
  13203=>"001010100",
  13204=>"100010110",
  13205=>"110110010",
  13206=>"000001000",
  13207=>"000111001",
  13208=>"010101101",
  13209=>"100001010",
  13210=>"010101111",
  13211=>"001100101",
  13212=>"110011000",
  13213=>"101111100",
  13214=>"111000011",
  13215=>"001001101",
  13216=>"111110111",
  13217=>"111011001",
  13218=>"100011000",
  13219=>"001100101",
  13220=>"111101001",
  13221=>"010011101",
  13222=>"111110010",
  13223=>"000000111",
  13224=>"101101100",
  13225=>"011100100",
  13226=>"111010000",
  13227=>"101000011",
  13228=>"010100110",
  13229=>"111100100",
  13230=>"000001011",
  13231=>"000100010",
  13232=>"000101000",
  13233=>"111111100",
  13234=>"001101000",
  13235=>"101100011",
  13236=>"000010010",
  13237=>"000001001",
  13238=>"011001000",
  13239=>"110110100",
  13240=>"110010101",
  13241=>"110010101",
  13242=>"101110111",
  13243=>"001000000",
  13244=>"100001111",
  13245=>"011111001",
  13246=>"111110011",
  13247=>"101110101",
  13248=>"100000101",
  13249=>"111100111",
  13250=>"100111110",
  13251=>"011111011",
  13252=>"010111100",
  13253=>"000110011",
  13254=>"100011100",
  13255=>"100000101",
  13256=>"000100110",
  13257=>"000111010",
  13258=>"110011010",
  13259=>"111110010",
  13260=>"010110010",
  13261=>"010110000",
  13262=>"011111000",
  13263=>"101110000",
  13264=>"110110010",
  13265=>"010110111",
  13266=>"010100101",
  13267=>"000111111",
  13268=>"011010110",
  13269=>"001100001",
  13270=>"010000010",
  13271=>"010101001",
  13272=>"100100000",
  13273=>"100111111",
  13274=>"101100101",
  13275=>"001000110",
  13276=>"001001111",
  13277=>"000110011",
  13278=>"101010100",
  13279=>"100000110",
  13280=>"110010010",
  13281=>"100011101",
  13282=>"011010000",
  13283=>"001110100",
  13284=>"010010010",
  13285=>"011110100",
  13286=>"010101111",
  13287=>"011000100",
  13288=>"100100011",
  13289=>"100011111",
  13290=>"001111011",
  13291=>"110001101",
  13292=>"101001100",
  13293=>"010010111",
  13294=>"011010101",
  13295=>"011001010",
  13296=>"010001001",
  13297=>"000010110",
  13298=>"010100100",
  13299=>"000010000",
  13300=>"111011111",
  13301=>"011010111",
  13302=>"100110000",
  13303=>"111110101",
  13304=>"100000101",
  13305=>"011011011",
  13306=>"011111000",
  13307=>"011001111",
  13308=>"100010011",
  13309=>"010100011",
  13310=>"011101000",
  13311=>"111100111",
  13312=>"001101011",
  13313=>"101010001",
  13314=>"010011101",
  13315=>"100000010",
  13316=>"100111000",
  13317=>"001100011",
  13318=>"000010100",
  13319=>"011101000",
  13320=>"110001110",
  13321=>"001001011",
  13322=>"100111011",
  13323=>"110110000",
  13324=>"100100010",
  13325=>"001110000",
  13326=>"011101000",
  13327=>"011011100",
  13328=>"000100101",
  13329=>"000001100",
  13330=>"000101000",
  13331=>"001001100",
  13332=>"110111101",
  13333=>"010000101",
  13334=>"101110101",
  13335=>"111111001",
  13336=>"101100111",
  13337=>"111000001",
  13338=>"110000101",
  13339=>"000000111",
  13340=>"001000100",
  13341=>"111100101",
  13342=>"001010010",
  13343=>"101010011",
  13344=>"101000101",
  13345=>"000010010",
  13346=>"011010000",
  13347=>"110111000",
  13348=>"101001000",
  13349=>"101101100",
  13350=>"010100111",
  13351=>"101111000",
  13352=>"111110111",
  13353=>"110101111",
  13354=>"111010011",
  13355=>"000011111",
  13356=>"000101101",
  13357=>"111010000",
  13358=>"001001010",
  13359=>"110011010",
  13360=>"111101010",
  13361=>"111010111",
  13362=>"101010110",
  13363=>"100011110",
  13364=>"010110111",
  13365=>"111001111",
  13366=>"100110110",
  13367=>"001100110",
  13368=>"000110001",
  13369=>"100011101",
  13370=>"000010010",
  13371=>"011010000",
  13372=>"100100010",
  13373=>"111001100",
  13374=>"010011001",
  13375=>"011000100",
  13376=>"011001011",
  13377=>"010011101",
  13378=>"001100011",
  13379=>"010111011",
  13380=>"001110100",
  13381=>"110010010",
  13382=>"110101000",
  13383=>"110011001",
  13384=>"101010110",
  13385=>"101100110",
  13386=>"000101001",
  13387=>"101001101",
  13388=>"100010101",
  13389=>"100110010",
  13390=>"000011001",
  13391=>"010100001",
  13392=>"100000110",
  13393=>"000000111",
  13394=>"010001010",
  13395=>"101010100",
  13396=>"010001011",
  13397=>"000010010",
  13398=>"000011001",
  13399=>"101111011",
  13400=>"101011111",
  13401=>"100000010",
  13402=>"101010110",
  13403=>"110010000",
  13404=>"110010111",
  13405=>"001111100",
  13406=>"001011001",
  13407=>"101010110",
  13408=>"111111011",
  13409=>"111100101",
  13410=>"000011001",
  13411=>"100101111",
  13412=>"110000001",
  13413=>"000011001",
  13414=>"110000100",
  13415=>"101011000",
  13416=>"000110101",
  13417=>"111010001",
  13418=>"100110110",
  13419=>"000001100",
  13420=>"110111111",
  13421=>"000000011",
  13422=>"111001111",
  13423=>"000010011",
  13424=>"101110110",
  13425=>"100101100",
  13426=>"111010110",
  13427=>"011100101",
  13428=>"011111111",
  13429=>"110110111",
  13430=>"001000000",
  13431=>"100110001",
  13432=>"111111100",
  13433=>"101000001",
  13434=>"110100011",
  13435=>"011000010",
  13436=>"000111001",
  13437=>"110011010",
  13438=>"111101101",
  13439=>"111011100",
  13440=>"000010001",
  13441=>"001000010",
  13442=>"101100110",
  13443=>"010101000",
  13444=>"110111010",
  13445=>"111110010",
  13446=>"001111011",
  13447=>"100001011",
  13448=>"000111111",
  13449=>"111001110",
  13450=>"010000011",
  13451=>"100111110",
  13452=>"001000001",
  13453=>"100110111",
  13454=>"010011110",
  13455=>"001110110",
  13456=>"011100011",
  13457=>"010010000",
  13458=>"000111010",
  13459=>"010100010",
  13460=>"001000111",
  13461=>"000101110",
  13462=>"000000100",
  13463=>"110100001",
  13464=>"000001100",
  13465=>"111010100",
  13466=>"111010100",
  13467=>"001011110",
  13468=>"100001001",
  13469=>"000000111",
  13470=>"010011101",
  13471=>"100110110",
  13472=>"110101110",
  13473=>"100101111",
  13474=>"111001011",
  13475=>"111101001",
  13476=>"111111111",
  13477=>"000001000",
  13478=>"000001010",
  13479=>"100100011",
  13480=>"010111111",
  13481=>"111001000",
  13482=>"100000011",
  13483=>"101100111",
  13484=>"111011011",
  13485=>"110010011",
  13486=>"111101011",
  13487=>"111011010",
  13488=>"111111011",
  13489=>"011010000",
  13490=>"000010111",
  13491=>"000100011",
  13492=>"010100001",
  13493=>"010000100",
  13494=>"000111100",
  13495=>"010110011",
  13496=>"001011100",
  13497=>"000000110",
  13498=>"110001001",
  13499=>"000010111",
  13500=>"111100110",
  13501=>"001001001",
  13502=>"101010001",
  13503=>"111101001",
  13504=>"111111100",
  13505=>"011001001",
  13506=>"110011001",
  13507=>"111001111",
  13508=>"100001010",
  13509=>"010100111",
  13510=>"110000011",
  13511=>"010010011",
  13512=>"010010000",
  13513=>"111001111",
  13514=>"001000001",
  13515=>"011111101",
  13516=>"000011000",
  13517=>"101101001",
  13518=>"110111111",
  13519=>"010111001",
  13520=>"001010000",
  13521=>"001100000",
  13522=>"101110110",
  13523=>"110011001",
  13524=>"011010110",
  13525=>"010010010",
  13526=>"101100101",
  13527=>"001110100",
  13528=>"111001100",
  13529=>"011000110",
  13530=>"010111111",
  13531=>"011000011",
  13532=>"110011111",
  13533=>"101010110",
  13534=>"000011100",
  13535=>"110011010",
  13536=>"010011111",
  13537=>"000001111",
  13538=>"111110100",
  13539=>"111011010",
  13540=>"001011110",
  13541=>"101011111",
  13542=>"011000011",
  13543=>"000100001",
  13544=>"011000110",
  13545=>"111100111",
  13546=>"100000100",
  13547=>"001000011",
  13548=>"011011011",
  13549=>"011010000",
  13550=>"000111010",
  13551=>"111011000",
  13552=>"001111110",
  13553=>"101011110",
  13554=>"000010000",
  13555=>"101000100",
  13556=>"111110101",
  13557=>"111101000",
  13558=>"111010010",
  13559=>"111111111",
  13560=>"111111011",
  13561=>"100000011",
  13562=>"010001110",
  13563=>"100011111",
  13564=>"000000001",
  13565=>"010011110",
  13566=>"011100001",
  13567=>"000011110",
  13568=>"000100101",
  13569=>"110101111",
  13570=>"100110110",
  13571=>"000011011",
  13572=>"111101011",
  13573=>"001011000",
  13574=>"000101100",
  13575=>"000001001",
  13576=>"110000100",
  13577=>"100110110",
  13578=>"101011010",
  13579=>"101000111",
  13580=>"011011000",
  13581=>"011001011",
  13582=>"011000001",
  13583=>"001101000",
  13584=>"000100011",
  13585=>"101000111",
  13586=>"011000101",
  13587=>"111101010",
  13588=>"100110111",
  13589=>"000100100",
  13590=>"101110011",
  13591=>"011001010",
  13592=>"110010001",
  13593=>"000101001",
  13594=>"100010001",
  13595=>"100000001",
  13596=>"011011110",
  13597=>"010011100",
  13598=>"101000110",
  13599=>"101111001",
  13600=>"010000011",
  13601=>"010111000",
  13602=>"011110111",
  13603=>"000110100",
  13604=>"110101010",
  13605=>"101101100",
  13606=>"110111110",
  13607=>"100100010",
  13608=>"111011010",
  13609=>"111001011",
  13610=>"110001101",
  13611=>"100000111",
  13612=>"110001010",
  13613=>"110011100",
  13614=>"001101100",
  13615=>"101100011",
  13616=>"010011100",
  13617=>"011101010",
  13618=>"010000000",
  13619=>"001010111",
  13620=>"000110000",
  13621=>"001000111",
  13622=>"101110111",
  13623=>"000011010",
  13624=>"001011011",
  13625=>"000101010",
  13626=>"000000111",
  13627=>"111100111",
  13628=>"010110001",
  13629=>"011101100",
  13630=>"011001001",
  13631=>"001101101",
  13632=>"111111001",
  13633=>"010000100",
  13634=>"001001101",
  13635=>"100011010",
  13636=>"010100010",
  13637=>"001100011",
  13638=>"011101111",
  13639=>"001101101",
  13640=>"100000000",
  13641=>"000010100",
  13642=>"101111100",
  13643=>"110011100",
  13644=>"100010111",
  13645=>"011000010",
  13646=>"010000111",
  13647=>"110101010",
  13648=>"001111110",
  13649=>"010010001",
  13650=>"011000110",
  13651=>"001001000",
  13652=>"110010010",
  13653=>"101110000",
  13654=>"011011001",
  13655=>"001001101",
  13656=>"100101011",
  13657=>"000101101",
  13658=>"011010000",
  13659=>"110001000",
  13660=>"100110101",
  13661=>"101011011",
  13662=>"010011100",
  13663=>"100101011",
  13664=>"110110100",
  13665=>"001011000",
  13666=>"100110010",
  13667=>"010000001",
  13668=>"111101001",
  13669=>"100000110",
  13670=>"101011110",
  13671=>"100010100",
  13672=>"111011111",
  13673=>"001000000",
  13674=>"110010110",
  13675=>"100001000",
  13676=>"000101111",
  13677=>"010010111",
  13678=>"011010110",
  13679=>"001101100",
  13680=>"011001110",
  13681=>"100101110",
  13682=>"110100000",
  13683=>"011101001",
  13684=>"111001001",
  13685=>"011100100",
  13686=>"011101010",
  13687=>"100100110",
  13688=>"000111110",
  13689=>"010001010",
  13690=>"101100011",
  13691=>"110100011",
  13692=>"000010000",
  13693=>"010000110",
  13694=>"010101100",
  13695=>"101000101",
  13696=>"100001010",
  13697=>"010111001",
  13698=>"101011100",
  13699=>"110110111",
  13700=>"100111111",
  13701=>"010010110",
  13702=>"100000101",
  13703=>"011000001",
  13704=>"000010001",
  13705=>"111111010",
  13706=>"000000001",
  13707=>"010000000",
  13708=>"010010010",
  13709=>"010101011",
  13710=>"010110011",
  13711=>"000100010",
  13712=>"111111111",
  13713=>"000010001",
  13714=>"011000001",
  13715=>"100011011",
  13716=>"101101000",
  13717=>"001010010",
  13718=>"010000010",
  13719=>"000111110",
  13720=>"010010101",
  13721=>"000110100",
  13722=>"000110110",
  13723=>"100110111",
  13724=>"011000010",
  13725=>"000111100",
  13726=>"001000101",
  13727=>"101100101",
  13728=>"010000011",
  13729=>"010010000",
  13730=>"011111000",
  13731=>"101001011",
  13732=>"101100010",
  13733=>"101111000",
  13734=>"101110000",
  13735=>"111010111",
  13736=>"010000010",
  13737=>"001001001",
  13738=>"010100111",
  13739=>"011110001",
  13740=>"111101111",
  13741=>"101001000",
  13742=>"100100000",
  13743=>"101000100",
  13744=>"001010101",
  13745=>"000110001",
  13746=>"110110110",
  13747=>"101011111",
  13748=>"010100100",
  13749=>"011001100",
  13750=>"111010110",
  13751=>"110111000",
  13752=>"011111010",
  13753=>"110010110",
  13754=>"010011001",
  13755=>"111111101",
  13756=>"110110001",
  13757=>"111011000",
  13758=>"001100011",
  13759=>"010101100",
  13760=>"010000110",
  13761=>"011010001",
  13762=>"011010011",
  13763=>"011111110",
  13764=>"010010100",
  13765=>"001101100",
  13766=>"011100110",
  13767=>"001010111",
  13768=>"000000000",
  13769=>"111111111",
  13770=>"000011100",
  13771=>"001100110",
  13772=>"111001001",
  13773=>"110001100",
  13774=>"010100011",
  13775=>"000100010",
  13776=>"101001111",
  13777=>"011001111",
  13778=>"110001110",
  13779=>"001110001",
  13780=>"110111101",
  13781=>"100101001",
  13782=>"101001111",
  13783=>"100011000",
  13784=>"001010101",
  13785=>"010000011",
  13786=>"000011001",
  13787=>"001110000",
  13788=>"000011100",
  13789=>"101001101",
  13790=>"011111100",
  13791=>"101010001",
  13792=>"010000111",
  13793=>"001011100",
  13794=>"000100110",
  13795=>"000001000",
  13796=>"010101100",
  13797=>"110111001",
  13798=>"101011111",
  13799=>"011001100",
  13800=>"010000100",
  13801=>"000111111",
  13802=>"100000010",
  13803=>"100110001",
  13804=>"011001011",
  13805=>"111101010",
  13806=>"001100010",
  13807=>"000010111",
  13808=>"100101011",
  13809=>"001110001",
  13810=>"100110110",
  13811=>"000010000",
  13812=>"000111101",
  13813=>"000001010",
  13814=>"110011110",
  13815=>"100001101",
  13816=>"001000001",
  13817=>"111001000",
  13818=>"001001110",
  13819=>"101001000",
  13820=>"111110001",
  13821=>"111011100",
  13822=>"110011000",
  13823=>"111000100",
  13824=>"111000101",
  13825=>"000101110",
  13826=>"011110011",
  13827=>"010101011",
  13828=>"100000001",
  13829=>"011100010",
  13830=>"101101111",
  13831=>"000010001",
  13832=>"101110111",
  13833=>"011010001",
  13834=>"111101101",
  13835=>"010000110",
  13836=>"000001011",
  13837=>"110010101",
  13838=>"101011110",
  13839=>"000110001",
  13840=>"110100111",
  13841=>"101011000",
  13842=>"100101100",
  13843=>"011011101",
  13844=>"100101000",
  13845=>"111001000",
  13846=>"101000011",
  13847=>"101110010",
  13848=>"110001110",
  13849=>"010100010",
  13850=>"101000001",
  13851=>"001000111",
  13852=>"100101110",
  13853=>"000110001",
  13854=>"001110000",
  13855=>"111010010",
  13856=>"010111001",
  13857=>"111001111",
  13858=>"100000010",
  13859=>"110101011",
  13860=>"111000100",
  13861=>"110000111",
  13862=>"011100100",
  13863=>"100000111",
  13864=>"001000000",
  13865=>"110101011",
  13866=>"110010001",
  13867=>"101000010",
  13868=>"001100111",
  13869=>"100110111",
  13870=>"001000000",
  13871=>"110010011",
  13872=>"111001001",
  13873=>"101010000",
  13874=>"011100000",
  13875=>"010001111",
  13876=>"111110111",
  13877=>"100111111",
  13878=>"000111110",
  13879=>"110110001",
  13880=>"010000011",
  13881=>"000111100",
  13882=>"100100101",
  13883=>"100010111",
  13884=>"000000100",
  13885=>"011101001",
  13886=>"010011000",
  13887=>"000101010",
  13888=>"100110000",
  13889=>"010010100",
  13890=>"000110011",
  13891=>"001111111",
  13892=>"101001101",
  13893=>"111001111",
  13894=>"001001111",
  13895=>"101001001",
  13896=>"111011101",
  13897=>"111101000",
  13898=>"000111001",
  13899=>"110100111",
  13900=>"001001111",
  13901=>"110010010",
  13902=>"000000010",
  13903=>"000011011",
  13904=>"111110000",
  13905=>"011010000",
  13906=>"001010011",
  13907=>"011101001",
  13908=>"001100111",
  13909=>"110111000",
  13910=>"011001000",
  13911=>"001111110",
  13912=>"001000010",
  13913=>"100010000",
  13914=>"110011011",
  13915=>"011010100",
  13916=>"000010010",
  13917=>"101010100",
  13918=>"110111001",
  13919=>"101111101",
  13920=>"001011101",
  13921=>"011110001",
  13922=>"010111101",
  13923=>"110010101",
  13924=>"101011000",
  13925=>"101111000",
  13926=>"000110011",
  13927=>"010010001",
  13928=>"010100000",
  13929=>"000000110",
  13930=>"110100011",
  13931=>"010000111",
  13932=>"000111101",
  13933=>"101100001",
  13934=>"000110010",
  13935=>"110100110",
  13936=>"000101111",
  13937=>"011101110",
  13938=>"000011000",
  13939=>"111100000",
  13940=>"010000110",
  13941=>"110111000",
  13942=>"001011110",
  13943=>"011011111",
  13944=>"110000100",
  13945=>"000101011",
  13946=>"100010111",
  13947=>"000100011",
  13948=>"001101101",
  13949=>"001011000",
  13950=>"011110010",
  13951=>"001110111",
  13952=>"000110010",
  13953=>"100110100",
  13954=>"111011010",
  13955=>"000001001",
  13956=>"010110000",
  13957=>"010001011",
  13958=>"010000000",
  13959=>"101010101",
  13960=>"011001111",
  13961=>"000010110",
  13962=>"111000001",
  13963=>"101001011",
  13964=>"010111110",
  13965=>"110000011",
  13966=>"000001010",
  13967=>"110111000",
  13968=>"100111000",
  13969=>"110000010",
  13970=>"100100111",
  13971=>"101001001",
  13972=>"001000101",
  13973=>"111011110",
  13974=>"111000100",
  13975=>"110111101",
  13976=>"010100011",
  13977=>"000001000",
  13978=>"001111000",
  13979=>"100000110",
  13980=>"111000110",
  13981=>"100011101",
  13982=>"000000110",
  13983=>"111001000",
  13984=>"111111110",
  13985=>"011000111",
  13986=>"000101010",
  13987=>"011000110",
  13988=>"011101101",
  13989=>"000111011",
  13990=>"000011111",
  13991=>"001010011",
  13992=>"010111000",
  13993=>"100001110",
  13994=>"011100110",
  13995=>"000000100",
  13996=>"101000001",
  13997=>"101010000",
  13998=>"010110111",
  13999=>"011100000",
  14000=>"101000101",
  14001=>"000100100",
  14002=>"010101100",
  14003=>"011011011",
  14004=>"010010001",
  14005=>"101011010",
  14006=>"000001110",
  14007=>"100101001",
  14008=>"011111100",
  14009=>"010011111",
  14010=>"011101000",
  14011=>"001111011",
  14012=>"001110100",
  14013=>"011000000",
  14014=>"001000000",
  14015=>"111010011",
  14016=>"110110000",
  14017=>"101101110",
  14018=>"110101001",
  14019=>"111011101",
  14020=>"111010100",
  14021=>"001110011",
  14022=>"001100001",
  14023=>"000000000",
  14024=>"000000000",
  14025=>"110111011",
  14026=>"110101001",
  14027=>"000000111",
  14028=>"100111011",
  14029=>"111101110",
  14030=>"101110101",
  14031=>"000010010",
  14032=>"011111111",
  14033=>"011000001",
  14034=>"010100000",
  14035=>"001011101",
  14036=>"010111001",
  14037=>"000010111",
  14038=>"101100110",
  14039=>"000001101",
  14040=>"010000110",
  14041=>"111100000",
  14042=>"010001101",
  14043=>"111011111",
  14044=>"101100111",
  14045=>"111000010",
  14046=>"000000011",
  14047=>"111110001",
  14048=>"101011110",
  14049=>"101001111",
  14050=>"101101010",
  14051=>"101101001",
  14052=>"110111111",
  14053=>"010111101",
  14054=>"111100100",
  14055=>"101100000",
  14056=>"101001100",
  14057=>"010000001",
  14058=>"010111110",
  14059=>"011011000",
  14060=>"100110000",
  14061=>"110100100",
  14062=>"111100100",
  14063=>"000101100",
  14064=>"010010101",
  14065=>"111110000",
  14066=>"101101001",
  14067=>"001101000",
  14068=>"000111011",
  14069=>"100100011",
  14070=>"101101011",
  14071=>"010000010",
  14072=>"000101111",
  14073=>"001111100",
  14074=>"111011110",
  14075=>"000111101",
  14076=>"011001111",
  14077=>"110101111",
  14078=>"110101111",
  14079=>"000010100",
  14080=>"100101110",
  14081=>"101011101",
  14082=>"101101100",
  14083=>"110100100",
  14084=>"010111101",
  14085=>"101011011",
  14086=>"101010010",
  14087=>"111000100",
  14088=>"001111111",
  14089=>"000100000",
  14090=>"110010101",
  14091=>"111011100",
  14092=>"111000000",
  14093=>"011101100",
  14094=>"110111001",
  14095=>"010100010",
  14096=>"111110001",
  14097=>"111111101",
  14098=>"111011000",
  14099=>"100010101",
  14100=>"110000010",
  14101=>"110110100",
  14102=>"011111110",
  14103=>"001001110",
  14104=>"000001100",
  14105=>"101000100",
  14106=>"110111011",
  14107=>"000000000",
  14108=>"000111111",
  14109=>"001010101",
  14110=>"011011101",
  14111=>"010111110",
  14112=>"001101100",
  14113=>"111100010",
  14114=>"111110000",
  14115=>"111111000",
  14116=>"110000101",
  14117=>"000000111",
  14118=>"000001101",
  14119=>"111001100",
  14120=>"110101101",
  14121=>"001100000",
  14122=>"000100101",
  14123=>"100110000",
  14124=>"111111000",
  14125=>"001010111",
  14126=>"010000100",
  14127=>"101110001",
  14128=>"000011101",
  14129=>"101111110",
  14130=>"000000000",
  14131=>"000011111",
  14132=>"010110001",
  14133=>"001000101",
  14134=>"011000001",
  14135=>"011001000",
  14136=>"100110111",
  14137=>"001101001",
  14138=>"101100111",
  14139=>"110000001",
  14140=>"111011000",
  14141=>"101011110",
  14142=>"101001000",
  14143=>"000101100",
  14144=>"101101101",
  14145=>"100001100",
  14146=>"100100110",
  14147=>"011111011",
  14148=>"010111010",
  14149=>"010101111",
  14150=>"001011101",
  14151=>"111100000",
  14152=>"001010101",
  14153=>"110111010",
  14154=>"011011011",
  14155=>"101110110",
  14156=>"001010100",
  14157=>"110000101",
  14158=>"101101110",
  14159=>"010111001",
  14160=>"010100000",
  14161=>"111000110",
  14162=>"110111000",
  14163=>"100111111",
  14164=>"010001101",
  14165=>"101011010",
  14166=>"100001111",
  14167=>"111011011",
  14168=>"110110010",
  14169=>"010010010",
  14170=>"110001000",
  14171=>"100001101",
  14172=>"010010101",
  14173=>"011110101",
  14174=>"111101110",
  14175=>"111111111",
  14176=>"001110101",
  14177=>"000011010",
  14178=>"010010001",
  14179=>"110011110",
  14180=>"101100101",
  14181=>"010110001",
  14182=>"011001111",
  14183=>"100011101",
  14184=>"111111000",
  14185=>"111100000",
  14186=>"001101001",
  14187=>"111000000",
  14188=>"011101011",
  14189=>"100101001",
  14190=>"001111100",
  14191=>"111110100",
  14192=>"010000001",
  14193=>"111000001",
  14194=>"110001100",
  14195=>"011100111",
  14196=>"011111110",
  14197=>"100101100",
  14198=>"000100010",
  14199=>"110011101",
  14200=>"101111100",
  14201=>"101110111",
  14202=>"000110010",
  14203=>"110111110",
  14204=>"010101000",
  14205=>"100011011",
  14206=>"111011100",
  14207=>"010100011",
  14208=>"111001001",
  14209=>"000010111",
  14210=>"100011001",
  14211=>"011010110",
  14212=>"111001101",
  14213=>"000101100",
  14214=>"100100111",
  14215=>"000100011",
  14216=>"101111011",
  14217=>"100101100",
  14218=>"001010100",
  14219=>"001000001",
  14220=>"000101111",
  14221=>"011111111",
  14222=>"101100111",
  14223=>"001000011",
  14224=>"110010101",
  14225=>"100010011",
  14226=>"001011011",
  14227=>"000101111",
  14228=>"110100100",
  14229=>"011110000",
  14230=>"011100110",
  14231=>"001011001",
  14232=>"000100000",
  14233=>"110111111",
  14234=>"101110110",
  14235=>"010011100",
  14236=>"110011000",
  14237=>"001000111",
  14238=>"111010101",
  14239=>"011000111",
  14240=>"001101100",
  14241=>"101000110",
  14242=>"100010000",
  14243=>"100000101",
  14244=>"111111000",
  14245=>"101100100",
  14246=>"111001110",
  14247=>"010110101",
  14248=>"110110000",
  14249=>"111011100",
  14250=>"011011111",
  14251=>"100100101",
  14252=>"011001000",
  14253=>"100110010",
  14254=>"011001010",
  14255=>"110010001",
  14256=>"101100001",
  14257=>"001010111",
  14258=>"100110000",
  14259=>"000101111",
  14260=>"100101110",
  14261=>"110001001",
  14262=>"111111010",
  14263=>"111110101",
  14264=>"010001010",
  14265=>"000111001",
  14266=>"101011011",
  14267=>"000111100",
  14268=>"010110001",
  14269=>"101100001",
  14270=>"100101000",
  14271=>"000010110",
  14272=>"000111111",
  14273=>"101100001",
  14274=>"001101011",
  14275=>"000001101",
  14276=>"000110111",
  14277=>"100001011",
  14278=>"111101110",
  14279=>"100000110",
  14280=>"100000110",
  14281=>"000001011",
  14282=>"010000001",
  14283=>"100010010",
  14284=>"111110111",
  14285=>"101100001",
  14286=>"110011110",
  14287=>"100011000",
  14288=>"010110010",
  14289=>"001010000",
  14290=>"100100011",
  14291=>"111001011",
  14292=>"001100010",
  14293=>"110001001",
  14294=>"000101101",
  14295=>"100011111",
  14296=>"011010111",
  14297=>"011000010",
  14298=>"110001000",
  14299=>"001001011",
  14300=>"000010001",
  14301=>"011000101",
  14302=>"000111100",
  14303=>"100001111",
  14304=>"001011101",
  14305=>"000110010",
  14306=>"000100111",
  14307=>"111100100",
  14308=>"000001101",
  14309=>"000111101",
  14310=>"000010110",
  14311=>"000000100",
  14312=>"000001000",
  14313=>"010001100",
  14314=>"100100001",
  14315=>"101110010",
  14316=>"001101001",
  14317=>"100010010",
  14318=>"010000011",
  14319=>"000110011",
  14320=>"110000110",
  14321=>"111100111",
  14322=>"100000001",
  14323=>"111010100",
  14324=>"111011100",
  14325=>"011000001",
  14326=>"001001110",
  14327=>"000000001",
  14328=>"001000110",
  14329=>"100111011",
  14330=>"100010101",
  14331=>"011110100",
  14332=>"010000101",
  14333=>"011101111",
  14334=>"000101101",
  14335=>"101010001",
  14336=>"010000111",
  14337=>"000011010",
  14338=>"000100000",
  14339=>"100010110",
  14340=>"000001101",
  14341=>"010010101",
  14342=>"011000010",
  14343=>"110011110",
  14344=>"111010101",
  14345=>"010111111",
  14346=>"100001110",
  14347=>"110111001",
  14348=>"011010010",
  14349=>"000001010",
  14350=>"110111110",
  14351=>"111000110",
  14352=>"010001110",
  14353=>"001110100",
  14354=>"100010100",
  14355=>"111101101",
  14356=>"001011001",
  14357=>"000000100",
  14358=>"010100000",
  14359=>"001011101",
  14360=>"010011001",
  14361=>"110010001",
  14362=>"011100001",
  14363=>"000011011",
  14364=>"000010010",
  14365=>"101011000",
  14366=>"010110110",
  14367=>"001000000",
  14368=>"111110111",
  14369=>"000111110",
  14370=>"000010000",
  14371=>"011000000",
  14372=>"111100100",
  14373=>"101111101",
  14374=>"100011000",
  14375=>"110100111",
  14376=>"001010111",
  14377=>"101100111",
  14378=>"100101001",
  14379=>"111000000",
  14380=>"011010100",
  14381=>"100111110",
  14382=>"101010011",
  14383=>"101111100",
  14384=>"100100101",
  14385=>"010101000",
  14386=>"000101110",
  14387=>"011010100",
  14388=>"111000000",
  14389=>"010011101",
  14390=>"010100001",
  14391=>"000111010",
  14392=>"100100111",
  14393=>"110000100",
  14394=>"011010011",
  14395=>"000011110",
  14396=>"111111000",
  14397=>"000000110",
  14398=>"111111000",
  14399=>"111110110",
  14400=>"010101101",
  14401=>"100000101",
  14402=>"000100101",
  14403=>"000110101",
  14404=>"000110001",
  14405=>"000000001",
  14406=>"001011111",
  14407=>"101110100",
  14408=>"010010000",
  14409=>"011000101",
  14410=>"100010000",
  14411=>"011010100",
  14412=>"000000110",
  14413=>"101101001",
  14414=>"101111011",
  14415=>"011111110",
  14416=>"011000010",
  14417=>"100011101",
  14418=>"101010101",
  14419=>"011100000",
  14420=>"110100001",
  14421=>"111110101",
  14422=>"011001111",
  14423=>"100011101",
  14424=>"111111101",
  14425=>"101111001",
  14426=>"110000100",
  14427=>"001000101",
  14428=>"000111110",
  14429=>"001110100",
  14430=>"010000011",
  14431=>"001000011",
  14432=>"101001110",
  14433=>"111011100",
  14434=>"101010110",
  14435=>"001101110",
  14436=>"011001011",
  14437=>"011001111",
  14438=>"111010100",
  14439=>"110001100",
  14440=>"010001101",
  14441=>"111110010",
  14442=>"000000000",
  14443=>"001011011",
  14444=>"110101101",
  14445=>"101101110",
  14446=>"101001011",
  14447=>"011011010",
  14448=>"001101001",
  14449=>"011011110",
  14450=>"111101101",
  14451=>"011111100",
  14452=>"011010111",
  14453=>"011111000",
  14454=>"001100001",
  14455=>"000111000",
  14456=>"010100011",
  14457=>"100001101",
  14458=>"110110101",
  14459=>"000010100",
  14460=>"100101000",
  14461=>"001100001",
  14462=>"111001111",
  14463=>"001000000",
  14464=>"011110000",
  14465=>"111101101",
  14466=>"010000011",
  14467=>"000011000",
  14468=>"010001101",
  14469=>"010100111",
  14470=>"010101000",
  14471=>"111111110",
  14472=>"110011100",
  14473=>"101001001",
  14474=>"100001111",
  14475=>"000011100",
  14476=>"111111100",
  14477=>"000011101",
  14478=>"110101001",
  14479=>"110010110",
  14480=>"111111110",
  14481=>"101010111",
  14482=>"001100100",
  14483=>"001010111",
  14484=>"011001001",
  14485=>"011101111",
  14486=>"111010000",
  14487=>"001011111",
  14488=>"100010100",
  14489=>"010111101",
  14490=>"000010011",
  14491=>"010101000",
  14492=>"001111101",
  14493=>"001000011",
  14494=>"101000100",
  14495=>"101011010",
  14496=>"001001010",
  14497=>"001010101",
  14498=>"001100111",
  14499=>"010110001",
  14500=>"011011000",
  14501=>"111001111",
  14502=>"110000010",
  14503=>"101100010",
  14504=>"100010011",
  14505=>"011110000",
  14506=>"100001000",
  14507=>"000100011",
  14508=>"111111010",
  14509=>"000101011",
  14510=>"001010111",
  14511=>"110100110",
  14512=>"101010011",
  14513=>"011010100",
  14514=>"000101001",
  14515=>"001100111",
  14516=>"110011101",
  14517=>"000000010",
  14518=>"100111101",
  14519=>"010100001",
  14520=>"100011111",
  14521=>"101001000",
  14522=>"000101100",
  14523=>"101110001",
  14524=>"100101001",
  14525=>"010100111",
  14526=>"111111111",
  14527=>"101010000",
  14528=>"000000000",
  14529=>"000010111",
  14530=>"001101100",
  14531=>"000000101",
  14532=>"111001001",
  14533=>"011000011",
  14534=>"110010000",
  14535=>"101011101",
  14536=>"111101110",
  14537=>"010110000",
  14538=>"011101101",
  14539=>"001100010",
  14540=>"110011111",
  14541=>"011110011",
  14542=>"100101011",
  14543=>"101010000",
  14544=>"011110001",
  14545=>"100000111",
  14546=>"000101100",
  14547=>"001000100",
  14548=>"101100000",
  14549=>"111010111",
  14550=>"110010111",
  14551=>"001000000",
  14552=>"000000010",
  14553=>"110101100",
  14554=>"000101100",
  14555=>"011010101",
  14556=>"001101110",
  14557=>"100101101",
  14558=>"000101001",
  14559=>"111000010",
  14560=>"011010101",
  14561=>"001011001",
  14562=>"111000110",
  14563=>"000111100",
  14564=>"010101110",
  14565=>"011000100",
  14566=>"101001010",
  14567=>"111010101",
  14568=>"011001010",
  14569=>"001001000",
  14570=>"111011110",
  14571=>"011010001",
  14572=>"110101000",
  14573=>"011000011",
  14574=>"001000010",
  14575=>"111110000",
  14576=>"001001011",
  14577=>"111011100",
  14578=>"000001111",
  14579=>"001000011",
  14580=>"110100000",
  14581=>"001100000",
  14582=>"100000010",
  14583=>"100000100",
  14584=>"000011000",
  14585=>"001100000",
  14586=>"110001101",
  14587=>"100100000",
  14588=>"000110001",
  14589=>"110101000",
  14590=>"101111111",
  14591=>"011000100",
  14592=>"011000000",
  14593=>"001001100",
  14594=>"001101010",
  14595=>"110110110",
  14596=>"011100001",
  14597=>"100000110",
  14598=>"000001000",
  14599=>"011101001",
  14600=>"000000000",
  14601=>"000011111",
  14602=>"111011001",
  14603=>"101110001",
  14604=>"011110011",
  14605=>"100001000",
  14606=>"001001001",
  14607=>"101011010",
  14608=>"010000101",
  14609=>"000101001",
  14610=>"110101101",
  14611=>"110011000",
  14612=>"100001110",
  14613=>"000010000",
  14614=>"111110010",
  14615=>"100011010",
  14616=>"101100110",
  14617=>"001110000",
  14618=>"010000110",
  14619=>"100011000",
  14620=>"101101000",
  14621=>"110001110",
  14622=>"101111000",
  14623=>"111010101",
  14624=>"001001011",
  14625=>"110111100",
  14626=>"001001010",
  14627=>"000111100",
  14628=>"001001100",
  14629=>"000111100",
  14630=>"101100010",
  14631=>"110011100",
  14632=>"011000101",
  14633=>"101010011",
  14634=>"010001001",
  14635=>"101011000",
  14636=>"000011000",
  14637=>"101100001",
  14638=>"110111100",
  14639=>"000100101",
  14640=>"111101010",
  14641=>"001001110",
  14642=>"001110101",
  14643=>"000110111",
  14644=>"011001001",
  14645=>"001001010",
  14646=>"110111110",
  14647=>"001100001",
  14648=>"100000111",
  14649=>"001100010",
  14650=>"010110001",
  14651=>"101000101",
  14652=>"011110111",
  14653=>"101000011",
  14654=>"001010001",
  14655=>"100101101",
  14656=>"100000011",
  14657=>"001101111",
  14658=>"000010000",
  14659=>"010110000",
  14660=>"100111001",
  14661=>"100010110",
  14662=>"101001101",
  14663=>"101001000",
  14664=>"011010101",
  14665=>"001011000",
  14666=>"110111011",
  14667=>"001110001",
  14668=>"110000010",
  14669=>"110110001",
  14670=>"100001111",
  14671=>"001001011",
  14672=>"111110011",
  14673=>"010001010",
  14674=>"011100101",
  14675=>"100100000",
  14676=>"111111110",
  14677=>"000011011",
  14678=>"010101011",
  14679=>"100001100",
  14680=>"010101101",
  14681=>"110011011",
  14682=>"001101001",
  14683=>"101000101",
  14684=>"111000010",
  14685=>"100100001",
  14686=>"000110101",
  14687=>"111001010",
  14688=>"111011000",
  14689=>"000100000",
  14690=>"011010001",
  14691=>"100010110",
  14692=>"101001100",
  14693=>"100000101",
  14694=>"001000100",
  14695=>"000000001",
  14696=>"001000101",
  14697=>"100110111",
  14698=>"100111101",
  14699=>"001111110",
  14700=>"100010010",
  14701=>"101110111",
  14702=>"010111010",
  14703=>"001001111",
  14704=>"000101010",
  14705=>"111100110",
  14706=>"001010001",
  14707=>"100110001",
  14708=>"111100001",
  14709=>"000011000",
  14710=>"100000110",
  14711=>"000100110",
  14712=>"011101001",
  14713=>"111001010",
  14714=>"110110010",
  14715=>"100001110",
  14716=>"100111110",
  14717=>"000110110",
  14718=>"100001000",
  14719=>"010100001",
  14720=>"010011101",
  14721=>"110010000",
  14722=>"001001101",
  14723=>"100000111",
  14724=>"111011101",
  14725=>"011101110",
  14726=>"001011001",
  14727=>"000011101",
  14728=>"001011001",
  14729=>"010101100",
  14730=>"000010010",
  14731=>"010000101",
  14732=>"100100110",
  14733=>"110001101",
  14734=>"010100101",
  14735=>"011101010",
  14736=>"011100000",
  14737=>"001001111",
  14738=>"111101010",
  14739=>"111001100",
  14740=>"101011000",
  14741=>"100000110",
  14742=>"110011010",
  14743=>"110101000",
  14744=>"011101101",
  14745=>"100110101",
  14746=>"111001100",
  14747=>"010100010",
  14748=>"111101001",
  14749=>"001000001",
  14750=>"100111000",
  14751=>"010101011",
  14752=>"010100101",
  14753=>"101101000",
  14754=>"000111100",
  14755=>"011011010",
  14756=>"101100100",
  14757=>"101111011",
  14758=>"000011001",
  14759=>"000001101",
  14760=>"110000010",
  14761=>"101010011",
  14762=>"100001001",
  14763=>"000101001",
  14764=>"111100011",
  14765=>"011111100",
  14766=>"010011111",
  14767=>"000010010",
  14768=>"000001111",
  14769=>"100010000",
  14770=>"100100101",
  14771=>"100010111",
  14772=>"011100001",
  14773=>"110100111",
  14774=>"100101100",
  14775=>"000111101",
  14776=>"110101110",
  14777=>"010111001",
  14778=>"110011010",
  14779=>"001000010",
  14780=>"000011010",
  14781=>"110110110",
  14782=>"001100000",
  14783=>"010111011",
  14784=>"101000000",
  14785=>"111111110",
  14786=>"000111010",
  14787=>"111011011",
  14788=>"101100100",
  14789=>"011001110",
  14790=>"100001100",
  14791=>"010011001",
  14792=>"001111000",
  14793=>"010000010",
  14794=>"011010100",
  14795=>"000011000",
  14796=>"011010001",
  14797=>"110111101",
  14798=>"100101010",
  14799=>"001001110",
  14800=>"110001001",
  14801=>"010110011",
  14802=>"101101010",
  14803=>"101110001",
  14804=>"010111011",
  14805=>"010011011",
  14806=>"000000110",
  14807=>"000000010",
  14808=>"001011000",
  14809=>"000111010",
  14810=>"110000010",
  14811=>"000011110",
  14812=>"100101000",
  14813=>"001001110",
  14814=>"101000001",
  14815=>"101111111",
  14816=>"110000011",
  14817=>"000000001",
  14818=>"111000100",
  14819=>"101100111",
  14820=>"000111001",
  14821=>"001010101",
  14822=>"001011100",
  14823=>"000100000",
  14824=>"101111111",
  14825=>"111011011",
  14826=>"110010010",
  14827=>"001000101",
  14828=>"010000111",
  14829=>"101001000",
  14830=>"110010100",
  14831=>"000100010",
  14832=>"011011011",
  14833=>"100011101",
  14834=>"000101110",
  14835=>"001101000",
  14836=>"100000100",
  14837=>"100111101",
  14838=>"001001000",
  14839=>"100001010",
  14840=>"101101010",
  14841=>"001110011",
  14842=>"011000100",
  14843=>"010001001",
  14844=>"011110111",
  14845=>"010001100",
  14846=>"101010001",
  14847=>"011010100",
  14848=>"111011110",
  14849=>"001001001",
  14850=>"001110110",
  14851=>"101100111",
  14852=>"110111101",
  14853=>"000111110",
  14854=>"000111011",
  14855=>"110010101",
  14856=>"110001100",
  14857=>"111010000",
  14858=>"100011100",
  14859=>"101111100",
  14860=>"001011000",
  14861=>"100000010",
  14862=>"011101101",
  14863=>"001111101",
  14864=>"010001111",
  14865=>"000000000",
  14866=>"011111010",
  14867=>"111101011",
  14868=>"101101111",
  14869=>"010111111",
  14870=>"000100010",
  14871=>"011011101",
  14872=>"011000000",
  14873=>"010110010",
  14874=>"011001110",
  14875=>"100110000",
  14876=>"000111101",
  14877=>"100010000",
  14878=>"101110100",
  14879=>"011000110",
  14880=>"010010110",
  14881=>"110000010",
  14882=>"110110100",
  14883=>"101001110",
  14884=>"001001111",
  14885=>"011001101",
  14886=>"011010110",
  14887=>"011010000",
  14888=>"100101100",
  14889=>"010100101",
  14890=>"011011000",
  14891=>"111011001",
  14892=>"110001100",
  14893=>"100101001",
  14894=>"010101000",
  14895=>"011011010",
  14896=>"000101110",
  14897=>"100101000",
  14898=>"010110101",
  14899=>"110000110",
  14900=>"110000101",
  14901=>"111011010",
  14902=>"010010110",
  14903=>"101000010",
  14904=>"101010000",
  14905=>"101110000",
  14906=>"011011000",
  14907=>"101010100",
  14908=>"010001011",
  14909=>"011101000",
  14910=>"010011000",
  14911=>"111100110",
  14912=>"110100010",
  14913=>"101001010",
  14914=>"000110000",
  14915=>"000010001",
  14916=>"011111010",
  14917=>"100011101",
  14918=>"111010011",
  14919=>"001000111",
  14920=>"110111111",
  14921=>"000100111",
  14922=>"100000001",
  14923=>"101111100",
  14924=>"101110111",
  14925=>"100100000",
  14926=>"100010001",
  14927=>"100110101",
  14928=>"000111000",
  14929=>"101101011",
  14930=>"100011010",
  14931=>"101011000",
  14932=>"000001011",
  14933=>"001110110",
  14934=>"111100101",
  14935=>"110001011",
  14936=>"111011000",
  14937=>"100111010",
  14938=>"101101001",
  14939=>"100000001",
  14940=>"110101100",
  14941=>"110010111",
  14942=>"101110001",
  14943=>"001111010",
  14944=>"110000000",
  14945=>"000110001",
  14946=>"110111011",
  14947=>"110110000",
  14948=>"111111011",
  14949=>"000001000",
  14950=>"100000000",
  14951=>"111000000",
  14952=>"100001101",
  14953=>"111100001",
  14954=>"011101111",
  14955=>"110001111",
  14956=>"100101000",
  14957=>"110011111",
  14958=>"110101111",
  14959=>"001001110",
  14960=>"001001000",
  14961=>"000011110",
  14962=>"110101000",
  14963=>"100010110",
  14964=>"100010000",
  14965=>"101010000",
  14966=>"001000101",
  14967=>"101000000",
  14968=>"010001000",
  14969=>"110001011",
  14970=>"010001111",
  14971=>"000000110",
  14972=>"011010101",
  14973=>"110011111",
  14974=>"110111100",
  14975=>"100000110",
  14976=>"111000001",
  14977=>"001110000",
  14978=>"111111010",
  14979=>"000001001",
  14980=>"010011100",
  14981=>"010100101",
  14982=>"001111101",
  14983=>"110010111",
  14984=>"010000101",
  14985=>"011000101",
  14986=>"000011101",
  14987=>"111111000",
  14988=>"000101101",
  14989=>"101101111",
  14990=>"001000010",
  14991=>"001000001",
  14992=>"110010100",
  14993=>"110000100",
  14994=>"000010011",
  14995=>"101111100",
  14996=>"110110110",
  14997=>"110000011",
  14998=>"111100001",
  14999=>"010111000",
  15000=>"001000101",
  15001=>"100111110",
  15002=>"000010001",
  15003=>"100001111",
  15004=>"010110100",
  15005=>"011110111",
  15006=>"111111111",
  15007=>"000010001",
  15008=>"011100101",
  15009=>"100110110",
  15010=>"111111101",
  15011=>"100111111",
  15012=>"010110100",
  15013=>"100111101",
  15014=>"011011011",
  15015=>"101100000",
  15016=>"010010100",
  15017=>"000100101",
  15018=>"111011000",
  15019=>"101101101",
  15020=>"110000011",
  15021=>"111010001",
  15022=>"010000000",
  15023=>"011111111",
  15024=>"010001111",
  15025=>"100101110",
  15026=>"110010111",
  15027=>"000110011",
  15028=>"011001001",
  15029=>"000100110",
  15030=>"001100100",
  15031=>"000111100",
  15032=>"101011101",
  15033=>"100100101",
  15034=>"111010110",
  15035=>"000001011",
  15036=>"101100110",
  15037=>"110000010",
  15038=>"000100111",
  15039=>"111110110",
  15040=>"110001100",
  15041=>"110100110",
  15042=>"000011110",
  15043=>"110000111",
  15044=>"000111111",
  15045=>"111010011",
  15046=>"011000011",
  15047=>"100100111",
  15048=>"101100011",
  15049=>"101001010",
  15050=>"001011010",
  15051=>"110001101",
  15052=>"100111111",
  15053=>"010000000",
  15054=>"100010001",
  15055=>"110010110",
  15056=>"001101011",
  15057=>"110011001",
  15058=>"101111100",
  15059=>"001010110",
  15060=>"110000101",
  15061=>"010100010",
  15062=>"111011010",
  15063=>"111101110",
  15064=>"111110010",
  15065=>"100000101",
  15066=>"101000011",
  15067=>"101110001",
  15068=>"001001100",
  15069=>"000000000",
  15070=>"101001111",
  15071=>"101100010",
  15072=>"001001011",
  15073=>"001010010",
  15074=>"111010111",
  15075=>"110101110",
  15076=>"111000111",
  15077=>"101100100",
  15078=>"001101010",
  15079=>"111100101",
  15080=>"110011000",
  15081=>"110011111",
  15082=>"111110110",
  15083=>"000100011",
  15084=>"001000101",
  15085=>"001010110",
  15086=>"001001100",
  15087=>"110110011",
  15088=>"011000101",
  15089=>"011011110",
  15090=>"111111011",
  15091=>"001100010",
  15092=>"111111000",
  15093=>"000001101",
  15094=>"101000100",
  15095=>"110000110",
  15096=>"011111101",
  15097=>"000010011",
  15098=>"011100101",
  15099=>"000100010",
  15100=>"000010000",
  15101=>"000011000",
  15102=>"001000000",
  15103=>"100010110",
  15104=>"110000010",
  15105=>"011101101",
  15106=>"101000001",
  15107=>"110100110",
  15108=>"001000111",
  15109=>"100000001",
  15110=>"011111000",
  15111=>"000010011",
  15112=>"101011100",
  15113=>"001111100",
  15114=>"000101010",
  15115=>"000010101",
  15116=>"111110111",
  15117=>"011011110",
  15118=>"110000100",
  15119=>"100100110",
  15120=>"111010110",
  15121=>"110011010",
  15122=>"001001111",
  15123=>"101100101",
  15124=>"101011010",
  15125=>"011000010",
  15126=>"011100100",
  15127=>"110111100",
  15128=>"110010000",
  15129=>"110011110",
  15130=>"000000101",
  15131=>"010101111",
  15132=>"101001000",
  15133=>"110110111",
  15134=>"010010010",
  15135=>"111011011",
  15136=>"110010001",
  15137=>"100001001",
  15138=>"101100101",
  15139=>"101100011",
  15140=>"000111011",
  15141=>"101100011",
  15142=>"011000101",
  15143=>"101110111",
  15144=>"011010000",
  15145=>"110001001",
  15146=>"001000010",
  15147=>"011001100",
  15148=>"000010010",
  15149=>"110100110",
  15150=>"100010110",
  15151=>"111111111",
  15152=>"101111000",
  15153=>"100001100",
  15154=>"111100111",
  15155=>"011000101",
  15156=>"110100011",
  15157=>"111101000",
  15158=>"000011010",
  15159=>"110100001",
  15160=>"101100111",
  15161=>"110100101",
  15162=>"011011000",
  15163=>"010011101",
  15164=>"011101000",
  15165=>"110011101",
  15166=>"001001010",
  15167=>"111111000",
  15168=>"000001011",
  15169=>"111000011",
  15170=>"011010011",
  15171=>"100101011",
  15172=>"100000010",
  15173=>"011101000",
  15174=>"001000111",
  15175=>"110010101",
  15176=>"110011010",
  15177=>"101010100",
  15178=>"011111001",
  15179=>"001100101",
  15180=>"101101000",
  15181=>"001111110",
  15182=>"010111110",
  15183=>"011011101",
  15184=>"110101010",
  15185=>"001111001",
  15186=>"000010110",
  15187=>"110101110",
  15188=>"111111111",
  15189=>"001010101",
  15190=>"110000110",
  15191=>"010100011",
  15192=>"000000010",
  15193=>"111010001",
  15194=>"010110100",
  15195=>"001100101",
  15196=>"010100010",
  15197=>"011100010",
  15198=>"010110110",
  15199=>"100001010",
  15200=>"001101001",
  15201=>"110100010",
  15202=>"101001111",
  15203=>"111111100",
  15204=>"011011111",
  15205=>"111110000",
  15206=>"001011100",
  15207=>"000101000",
  15208=>"111000000",
  15209=>"001111000",
  15210=>"001011100",
  15211=>"010110100",
  15212=>"011111100",
  15213=>"001001000",
  15214=>"001110111",
  15215=>"001010101",
  15216=>"111100001",
  15217=>"011111101",
  15218=>"100111000",
  15219=>"100110110",
  15220=>"000010110",
  15221=>"111010101",
  15222=>"110011010",
  15223=>"001000101",
  15224=>"100111001",
  15225=>"010000001",
  15226=>"010011000",
  15227=>"001111110",
  15228=>"111111110",
  15229=>"101100010",
  15230=>"110110010",
  15231=>"110011001",
  15232=>"101100100",
  15233=>"101100000",
  15234=>"000111010",
  15235=>"011110100",
  15236=>"100000101",
  15237=>"001000001",
  15238=>"111100110",
  15239=>"100101001",
  15240=>"101010101",
  15241=>"111101101",
  15242=>"001010111",
  15243=>"111110100",
  15244=>"110000001",
  15245=>"111011111",
  15246=>"111011100",
  15247=>"110101010",
  15248=>"110011011",
  15249=>"110110001",
  15250=>"100101001",
  15251=>"100010010",
  15252=>"010011110",
  15253=>"111101100",
  15254=>"110001100",
  15255=>"111100100",
  15256=>"000000111",
  15257=>"000111000",
  15258=>"111100000",
  15259=>"101110010",
  15260=>"101111101",
  15261=>"111111010",
  15262=>"000111000",
  15263=>"001001110",
  15264=>"101000010",
  15265=>"010000110",
  15266=>"110101011",
  15267=>"011010000",
  15268=>"000110101",
  15269=>"000010101",
  15270=>"011000100",
  15271=>"101010001",
  15272=>"100000110",
  15273=>"110000000",
  15274=>"101101011",
  15275=>"001011110",
  15276=>"000000110",
  15277=>"100000011",
  15278=>"100000011",
  15279=>"001010110",
  15280=>"111000001",
  15281=>"101001010",
  15282=>"100101110",
  15283=>"100000101",
  15284=>"011110010",
  15285=>"000100110",
  15286=>"110101011",
  15287=>"000011001",
  15288=>"111101110",
  15289=>"100001100",
  15290=>"100011100",
  15291=>"001101001",
  15292=>"001011001",
  15293=>"111110001",
  15294=>"010100011",
  15295=>"100100100",
  15296=>"101101001",
  15297=>"100101111",
  15298=>"001001110",
  15299=>"110101001",
  15300=>"111000011",
  15301=>"011011111",
  15302=>"101100001",
  15303=>"100101111",
  15304=>"001111101",
  15305=>"101101011",
  15306=>"101100111",
  15307=>"011001001",
  15308=>"110000110",
  15309=>"110100101",
  15310=>"010110100",
  15311=>"100000110",
  15312=>"110000101",
  15313=>"011110000",
  15314=>"001101010",
  15315=>"001101110",
  15316=>"000110001",
  15317=>"100011100",
  15318=>"001010011",
  15319=>"011010001",
  15320=>"001000101",
  15321=>"111101110",
  15322=>"001000100",
  15323=>"010111110",
  15324=>"110000100",
  15325=>"000100101",
  15326=>"100100011",
  15327=>"111110001",
  15328=>"000000110",
  15329=>"001101111",
  15330=>"010001101",
  15331=>"011011010",
  15332=>"010110000",
  15333=>"100100111",
  15334=>"010011011",
  15335=>"000000000",
  15336=>"101001001",
  15337=>"111010110",
  15338=>"100000011",
  15339=>"101100011",
  15340=>"100101000",
  15341=>"101111111",
  15342=>"010010000",
  15343=>"111000111",
  15344=>"000100010",
  15345=>"100011100",
  15346=>"001000001",
  15347=>"001001000",
  15348=>"110011001",
  15349=>"111010010",
  15350=>"000001000",
  15351=>"011000100",
  15352=>"000100010",
  15353=>"111100000",
  15354=>"000011100",
  15355=>"010011000",
  15356=>"111100011",
  15357=>"010101000",
  15358=>"101111000",
  15359=>"011011101",
  15360=>"010100110",
  15361=>"101110111",
  15362=>"000101111",
  15363=>"101011000",
  15364=>"000010010",
  15365=>"000110101",
  15366=>"111000011",
  15367=>"010011000",
  15368=>"100101100",
  15369=>"001100001",
  15370=>"010011011",
  15371=>"100011100",
  15372=>"100001111",
  15373=>"001111010",
  15374=>"000100010",
  15375=>"001011010",
  15376=>"110010110",
  15377=>"011110110",
  15378=>"011010010",
  15379=>"001011001",
  15380=>"101100100",
  15381=>"111011001",
  15382=>"001011111",
  15383=>"001100011",
  15384=>"111111111",
  15385=>"010000101",
  15386=>"111110110",
  15387=>"100111010",
  15388=>"111101101",
  15389=>"000010110",
  15390=>"001000010",
  15391=>"111011001",
  15392=>"101101001",
  15393=>"000101111",
  15394=>"111110110",
  15395=>"001111110",
  15396=>"011001110",
  15397=>"111111001",
  15398=>"101111110",
  15399=>"110111100",
  15400=>"100110001",
  15401=>"111000010",
  15402=>"011100110",
  15403=>"100111010",
  15404=>"000110011",
  15405=>"011110000",
  15406=>"001010110",
  15407=>"011110110",
  15408=>"110001110",
  15409=>"111111101",
  15410=>"010010000",
  15411=>"001110100",
  15412=>"010101000",
  15413=>"011100000",
  15414=>"001110110",
  15415=>"000011110",
  15416=>"101111111",
  15417=>"101100000",
  15418=>"110111111",
  15419=>"100000101",
  15420=>"011101100",
  15421=>"100000000",
  15422=>"101111111",
  15423=>"010111010",
  15424=>"000001010",
  15425=>"000010000",
  15426=>"000010111",
  15427=>"101110000",
  15428=>"100010100",
  15429=>"101011100",
  15430=>"100111010",
  15431=>"000000001",
  15432=>"101110100",
  15433=>"011001001",
  15434=>"100100011",
  15435=>"000000000",
  15436=>"010000101",
  15437=>"111110110",
  15438=>"010100000",
  15439=>"111111111",
  15440=>"110111000",
  15441=>"001100000",
  15442=>"001111010",
  15443=>"111101110",
  15444=>"100100101",
  15445=>"100011000",
  15446=>"011011000",
  15447=>"101010010",
  15448=>"101011000",
  15449=>"010100010",
  15450=>"010001001",
  15451=>"010100100",
  15452=>"011000010",
  15453=>"100101000",
  15454=>"000111000",
  15455=>"000001100",
  15456=>"000001001",
  15457=>"110011111",
  15458=>"010100111",
  15459=>"100111010",
  15460=>"001000100",
  15461=>"010000001",
  15462=>"100101111",
  15463=>"111001011",
  15464=>"010000011",
  15465=>"101011101",
  15466=>"001110001",
  15467=>"001110011",
  15468=>"001111001",
  15469=>"010110000",
  15470=>"110111010",
  15471=>"010000101",
  15472=>"100000000",
  15473=>"010110000",
  15474=>"111001010",
  15475=>"000101110",
  15476=>"010000100",
  15477=>"101000000",
  15478=>"111011011",
  15479=>"000001100",
  15480=>"010011101",
  15481=>"001000000",
  15482=>"001001101",
  15483=>"100000101",
  15484=>"011010000",
  15485=>"010111000",
  15486=>"000000001",
  15487=>"010001011",
  15488=>"111100111",
  15489=>"000000111",
  15490=>"010100010",
  15491=>"001100000",
  15492=>"100110110",
  15493=>"101001010",
  15494=>"001110000",
  15495=>"101001110",
  15496=>"011011010",
  15497=>"101100110",
  15498=>"101011101",
  15499=>"011010000",
  15500=>"000000010",
  15501=>"100100001",
  15502=>"000011001",
  15503=>"010101111",
  15504=>"010001001",
  15505=>"111111101",
  15506=>"001000101",
  15507=>"000100000",
  15508=>"101111000",
  15509=>"011000011",
  15510=>"111111100",
  15511=>"001111111",
  15512=>"001101111",
  15513=>"101010010",
  15514=>"011111011",
  15515=>"001111101",
  15516=>"000110100",
  15517=>"011011111",
  15518=>"001010111",
  15519=>"000100000",
  15520=>"010101101",
  15521=>"001111111",
  15522=>"110010011",
  15523=>"010100101",
  15524=>"111011011",
  15525=>"100011110",
  15526=>"100110011",
  15527=>"001100110",
  15528=>"101001000",
  15529=>"111011111",
  15530=>"101110001",
  15531=>"100000101",
  15532=>"101001101",
  15533=>"111111100",
  15534=>"011111011",
  15535=>"111000011",
  15536=>"101101010",
  15537=>"000110000",
  15538=>"101110111",
  15539=>"010011000",
  15540=>"001100011",
  15541=>"111010101",
  15542=>"000000110",
  15543=>"100111001",
  15544=>"010110110",
  15545=>"111001010",
  15546=>"000100001",
  15547=>"110110011",
  15548=>"011100001",
  15549=>"100100111",
  15550=>"100011101",
  15551=>"101110111",
  15552=>"001101110",
  15553=>"001000111",
  15554=>"111010010",
  15555=>"001001111",
  15556=>"111100101",
  15557=>"010110111",
  15558=>"010000100",
  15559=>"000010110",
  15560=>"101011110",
  15561=>"101011111",
  15562=>"000110111",
  15563=>"000101011",
  15564=>"001010110",
  15565=>"011010001",
  15566=>"000000000",
  15567=>"010010011",
  15568=>"011000000",
  15569=>"101011110",
  15570=>"010101110",
  15571=>"011101111",
  15572=>"001000111",
  15573=>"010100010",
  15574=>"010010010",
  15575=>"100101011",
  15576=>"100100000",
  15577=>"001111000",
  15578=>"011100110",
  15579=>"100000111",
  15580=>"110001000",
  15581=>"101011000",
  15582=>"010101111",
  15583=>"000000001",
  15584=>"011100101",
  15585=>"101011000",
  15586=>"001110111",
  15587=>"000000001",
  15588=>"000010000",
  15589=>"110111101",
  15590=>"111111101",
  15591=>"001111101",
  15592=>"101100000",
  15593=>"111111100",
  15594=>"110111011",
  15595=>"011100010",
  15596=>"010010101",
  15597=>"000101111",
  15598=>"101000011",
  15599=>"000010100",
  15600=>"111100111",
  15601=>"110111011",
  15602=>"101010000",
  15603=>"110100110",
  15604=>"010110001",
  15605=>"111001111",
  15606=>"001000101",
  15607=>"111010001",
  15608=>"100001100",
  15609=>"100010101",
  15610=>"001101000",
  15611=>"000011000",
  15612=>"000011101",
  15613=>"000100001",
  15614=>"001001111",
  15615=>"100111110",
  15616=>"111011000",
  15617=>"110100110",
  15618=>"000000001",
  15619=>"001011110",
  15620=>"101111001",
  15621=>"010101110",
  15622=>"000001010",
  15623=>"110010110",
  15624=>"111001111",
  15625=>"111100010",
  15626=>"110011011",
  15627=>"000001101",
  15628=>"001011101",
  15629=>"110010111",
  15630=>"111000010",
  15631=>"000101001",
  15632=>"101101010",
  15633=>"101011111",
  15634=>"100011011",
  15635=>"110011001",
  15636=>"111001101",
  15637=>"000000000",
  15638=>"001000110",
  15639=>"011110000",
  15640=>"100011111",
  15641=>"101100011",
  15642=>"110110010",
  15643=>"110110111",
  15644=>"101001010",
  15645=>"100101000",
  15646=>"111101001",
  15647=>"110101001",
  15648=>"111000001",
  15649=>"101010011",
  15650=>"001100011",
  15651=>"111111011",
  15652=>"000111001",
  15653=>"100001011",
  15654=>"111000000",
  15655=>"100110010",
  15656=>"010000111",
  15657=>"000010100",
  15658=>"011110010",
  15659=>"000001100",
  15660=>"000110010",
  15661=>"010100111",
  15662=>"010001010",
  15663=>"001011100",
  15664=>"100110010",
  15665=>"000001110",
  15666=>"101110001",
  15667=>"010100000",
  15668=>"011011000",
  15669=>"011000101",
  15670=>"001100100",
  15671=>"000001010",
  15672=>"101000101",
  15673=>"001100101",
  15674=>"000011110",
  15675=>"111111010",
  15676=>"110100110",
  15677=>"010100101",
  15678=>"101110100",
  15679=>"000000100",
  15680=>"100100110",
  15681=>"011111001",
  15682=>"111000111",
  15683=>"111011101",
  15684=>"110010111",
  15685=>"100101111",
  15686=>"000100101",
  15687=>"001101001",
  15688=>"101101111",
  15689=>"010011111",
  15690=>"000001001",
  15691=>"110001000",
  15692=>"110101000",
  15693=>"110111110",
  15694=>"110100000",
  15695=>"101011011",
  15696=>"111000001",
  15697=>"001010110",
  15698=>"110100000",
  15699=>"111000011",
  15700=>"000000010",
  15701=>"101100111",
  15702=>"110011111",
  15703=>"000011010",
  15704=>"011010100",
  15705=>"011111010",
  15706=>"000010111",
  15707=>"101000110",
  15708=>"010011001",
  15709=>"010101100",
  15710=>"001101001",
  15711=>"000001001",
  15712=>"110011100",
  15713=>"001001101",
  15714=>"111010011",
  15715=>"011011000",
  15716=>"001000100",
  15717=>"001010111",
  15718=>"001001100",
  15719=>"011111110",
  15720=>"011011111",
  15721=>"010110000",
  15722=>"001011010",
  15723=>"010010101",
  15724=>"100000000",
  15725=>"111111100",
  15726=>"001111110",
  15727=>"010100000",
  15728=>"010100001",
  15729=>"111000000",
  15730=>"111101110",
  15731=>"101010100",
  15732=>"110010011",
  15733=>"101111101",
  15734=>"111110010",
  15735=>"001100010",
  15736=>"000000011",
  15737=>"111001111",
  15738=>"010000010",
  15739=>"100110011",
  15740=>"111010011",
  15741=>"101110101",
  15742=>"101011010",
  15743=>"101001010",
  15744=>"011110000",
  15745=>"000001101",
  15746=>"110111101",
  15747=>"001010010",
  15748=>"000110001",
  15749=>"000000100",
  15750=>"010101111",
  15751=>"111101001",
  15752=>"111001101",
  15753=>"111111011",
  15754=>"101101011",
  15755=>"111001011",
  15756=>"000111101",
  15757=>"010011001",
  15758=>"000101010",
  15759=>"001010001",
  15760=>"010101001",
  15761=>"110000000",
  15762=>"001111010",
  15763=>"011001111",
  15764=>"101001111",
  15765=>"100100110",
  15766=>"010100110",
  15767=>"000110100",
  15768=>"110010001",
  15769=>"000111010",
  15770=>"001001001",
  15771=>"101001001",
  15772=>"111101101",
  15773=>"100100000",
  15774=>"000110101",
  15775=>"111011111",
  15776=>"101101100",
  15777=>"111111111",
  15778=>"011101001",
  15779=>"001000110",
  15780=>"101110000",
  15781=>"000001011",
  15782=>"110010010",
  15783=>"011101001",
  15784=>"010001101",
  15785=>"111000111",
  15786=>"101110111",
  15787=>"101001111",
  15788=>"101010110",
  15789=>"101110010",
  15790=>"110101111",
  15791=>"000111110",
  15792=>"111110011",
  15793=>"011110100",
  15794=>"011110011",
  15795=>"010110010",
  15796=>"010000001",
  15797=>"100000100",
  15798=>"110011011",
  15799=>"001100101",
  15800=>"100100000",
  15801=>"000110111",
  15802=>"000011001",
  15803=>"000001001",
  15804=>"001111001",
  15805=>"010101001",
  15806=>"000010000",
  15807=>"010101111",
  15808=>"110101111",
  15809=>"100001011",
  15810=>"100101001",
  15811=>"011111101",
  15812=>"011010101",
  15813=>"000000010",
  15814=>"000000001",
  15815=>"101110000",
  15816=>"001011110",
  15817=>"100110011",
  15818=>"010000000",
  15819=>"100000100",
  15820=>"111110111",
  15821=>"100010101",
  15822=>"000001111",
  15823=>"000010011",
  15824=>"010110010",
  15825=>"010010010",
  15826=>"001000010",
  15827=>"111100110",
  15828=>"000001011",
  15829=>"101000001",
  15830=>"010000010",
  15831=>"000100110",
  15832=>"100010101",
  15833=>"101001111",
  15834=>"101010100",
  15835=>"100010110",
  15836=>"010100101",
  15837=>"101111001",
  15838=>"010100110",
  15839=>"010011101",
  15840=>"100110100",
  15841=>"100111100",
  15842=>"000001110",
  15843=>"001001001",
  15844=>"001010101",
  15845=>"000110001",
  15846=>"110001100",
  15847=>"101011000",
  15848=>"110001011",
  15849=>"111011111",
  15850=>"011010101",
  15851=>"111011001",
  15852=>"101110101",
  15853=>"001011101",
  15854=>"011100011",
  15855=>"110111000",
  15856=>"010010010",
  15857=>"010110111",
  15858=>"110111101",
  15859=>"000000001",
  15860=>"111101000",
  15861=>"011010011",
  15862=>"000011111",
  15863=>"000100100",
  15864=>"111111010",
  15865=>"110101110",
  15866=>"000011101",
  15867=>"101010011",
  15868=>"101011001",
  15869=>"010101011",
  15870=>"100100010",
  15871=>"111111111",
  15872=>"001111000",
  15873=>"010101110",
  15874=>"001010010",
  15875=>"000000000",
  15876=>"001010010",
  15877=>"110110110",
  15878=>"010000010",
  15879=>"101001111",
  15880=>"010111111",
  15881=>"010110100",
  15882=>"000101001",
  15883=>"000100011",
  15884=>"100110011",
  15885=>"110100001",
  15886=>"100010001",
  15887=>"101100101",
  15888=>"101110110",
  15889=>"110001110",
  15890=>"011111110",
  15891=>"101001110",
  15892=>"110101010",
  15893=>"100101000",
  15894=>"111101001",
  15895=>"101001010",
  15896=>"011000000",
  15897=>"001110011",
  15898=>"000101011",
  15899=>"011000011",
  15900=>"000000000",
  15901=>"000010100",
  15902=>"010110110",
  15903=>"101100101",
  15904=>"101000001",
  15905=>"100101100",
  15906=>"111010111",
  15907=>"011110000",
  15908=>"111011001",
  15909=>"110111111",
  15910=>"010111001",
  15911=>"111101011",
  15912=>"111111100",
  15913=>"110110100",
  15914=>"111000011",
  15915=>"000100111",
  15916=>"011110001",
  15917=>"000001010",
  15918=>"111100110",
  15919=>"001000100",
  15920=>"011100110",
  15921=>"111111101",
  15922=>"101011010",
  15923=>"111011101",
  15924=>"101110110",
  15925=>"000001100",
  15926=>"101000001",
  15927=>"100010110",
  15928=>"000011111",
  15929=>"100101101",
  15930=>"100110111",
  15931=>"001100111",
  15932=>"110000010",
  15933=>"000001001",
  15934=>"000010110",
  15935=>"101111000",
  15936=>"001000100",
  15937=>"111010111",
  15938=>"010011001",
  15939=>"000000111",
  15940=>"010010001",
  15941=>"011001110",
  15942=>"010110010",
  15943=>"010111010",
  15944=>"001111111",
  15945=>"110101111",
  15946=>"100001011",
  15947=>"001101000",
  15948=>"110101111",
  15949=>"101011100",
  15950=>"110000101",
  15951=>"110110100",
  15952=>"111011000",
  15953=>"001101001",
  15954=>"001110011",
  15955=>"011101000",
  15956=>"010101110",
  15957=>"010101011",
  15958=>"000001100",
  15959=>"111110011",
  15960=>"000000110",
  15961=>"100011111",
  15962=>"100111110",
  15963=>"100010001",
  15964=>"111011011",
  15965=>"010101001",
  15966=>"111010110",
  15967=>"000110101",
  15968=>"000000000",
  15969=>"010101010",
  15970=>"100100100",
  15971=>"100011111",
  15972=>"100001110",
  15973=>"011100101",
  15974=>"010000111",
  15975=>"111011111",
  15976=>"001011000",
  15977=>"000101100",
  15978=>"011100111",
  15979=>"000100000",
  15980=>"011010001",
  15981=>"111011110",
  15982=>"000010111",
  15983=>"000111010",
  15984=>"111100001",
  15985=>"100100010",
  15986=>"000011010",
  15987=>"000110101",
  15988=>"000100001",
  15989=>"001111010",
  15990=>"001001011",
  15991=>"101100101",
  15992=>"010011000",
  15993=>"011111000",
  15994=>"011110101",
  15995=>"010011011",
  15996=>"000101001",
  15997=>"110100001",
  15998=>"110011100",
  15999=>"000000010",
  16000=>"011001011",
  16001=>"001001111",
  16002=>"001101111",
  16003=>"111101111",
  16004=>"010001011",
  16005=>"000110011",
  16006=>"110100010",
  16007=>"101001000",
  16008=>"011010000",
  16009=>"111000101",
  16010=>"110011011",
  16011=>"100000001",
  16012=>"010100000",
  16013=>"111011100",
  16014=>"001000001",
  16015=>"111111001",
  16016=>"010000011",
  16017=>"100110111",
  16018=>"000101111",
  16019=>"011101001",
  16020=>"001011011",
  16021=>"111010010",
  16022=>"100011010",
  16023=>"110111110",
  16024=>"111011111",
  16025=>"101001011",
  16026=>"110000000",
  16027=>"001111010",
  16028=>"101100100",
  16029=>"100000001",
  16030=>"010010011",
  16031=>"111011000",
  16032=>"010011110",
  16033=>"100100110",
  16034=>"000000101",
  16035=>"110111011",
  16036=>"101101000",
  16037=>"100110010",
  16038=>"001110011",
  16039=>"011110010",
  16040=>"010010001",
  16041=>"000000000",
  16042=>"101110101",
  16043=>"111101011",
  16044=>"000000100",
  16045=>"000100011",
  16046=>"000011010",
  16047=>"001011001",
  16048=>"001100100",
  16049=>"001001001",
  16050=>"011001000",
  16051=>"001001100",
  16052=>"110000101",
  16053=>"110110100",
  16054=>"100000101",
  16055=>"101001101",
  16056=>"000101101",
  16057=>"011001010",
  16058=>"111011111",
  16059=>"100100101",
  16060=>"001001000",
  16061=>"010001101",
  16062=>"000010001",
  16063=>"101101001",
  16064=>"100001010",
  16065=>"010101101",
  16066=>"000000111",
  16067=>"110110101",
  16068=>"000011001",
  16069=>"100100110",
  16070=>"010111101",
  16071=>"010111000",
  16072=>"101100011",
  16073=>"001010001",
  16074=>"001101000",
  16075=>"000100110",
  16076=>"110101111",
  16077=>"111111110",
  16078=>"110101001",
  16079=>"110110111",
  16080=>"100001011",
  16081=>"010001100",
  16082=>"010100010",
  16083=>"111010110",
  16084=>"011010000",
  16085=>"001000101",
  16086=>"011110000",
  16087=>"010100100",
  16088=>"100110100",
  16089=>"101001010",
  16090=>"000110110",
  16091=>"100001011",
  16092=>"101011100",
  16093=>"000010110",
  16094=>"110010010",
  16095=>"000000100",
  16096=>"110010010",
  16097=>"100001001",
  16098=>"010100001",
  16099=>"001011100",
  16100=>"000000000",
  16101=>"001101011",
  16102=>"010000000",
  16103=>"010001011",
  16104=>"101010010",
  16105=>"010100100",
  16106=>"000000001",
  16107=>"111110011",
  16108=>"010110011",
  16109=>"010110100",
  16110=>"111100011",
  16111=>"001010000",
  16112=>"100110110",
  16113=>"110001010",
  16114=>"011001101",
  16115=>"011111111",
  16116=>"000000110",
  16117=>"011001001",
  16118=>"001101110",
  16119=>"011110010",
  16120=>"001111001",
  16121=>"000100110",
  16122=>"000111110",
  16123=>"010011001",
  16124=>"110111100",
  16125=>"100001001",
  16126=>"110011111",
  16127=>"010111001",
  16128=>"110010001",
  16129=>"101001000",
  16130=>"111110111",
  16131=>"100010011",
  16132=>"000011001",
  16133=>"100000000",
  16134=>"110100100",
  16135=>"101110011",
  16136=>"000010001",
  16137=>"001101100",
  16138=>"111110110",
  16139=>"010100000",
  16140=>"010001000",
  16141=>"110010110",
  16142=>"111011011",
  16143=>"110101100",
  16144=>"000100001",
  16145=>"111111011",
  16146=>"100010000",
  16147=>"011100100",
  16148=>"100110101",
  16149=>"001100001",
  16150=>"010100010",
  16151=>"000001100",
  16152=>"111100101",
  16153=>"101101101",
  16154=>"101000100",
  16155=>"111011110",
  16156=>"000000001",
  16157=>"111110011",
  16158=>"011000100",
  16159=>"100101010",
  16160=>"110011101",
  16161=>"010110100",
  16162=>"111111011",
  16163=>"101110101",
  16164=>"110011110",
  16165=>"100010110",
  16166=>"110011111",
  16167=>"111101111",
  16168=>"100001110",
  16169=>"001000101",
  16170=>"111011001",
  16171=>"110111111",
  16172=>"110101110",
  16173=>"010001011",
  16174=>"011010011",
  16175=>"001111010",
  16176=>"001110111",
  16177=>"100100100",
  16178=>"110111111",
  16179=>"110101110",
  16180=>"010100010",
  16181=>"111101000",
  16182=>"101111110",
  16183=>"100001010",
  16184=>"110001110",
  16185=>"111110100",
  16186=>"110111000",
  16187=>"011001001",
  16188=>"101101001",
  16189=>"101010000",
  16190=>"010011101",
  16191=>"100110011",
  16192=>"010110000",
  16193=>"101001111",
  16194=>"101000100",
  16195=>"111011000",
  16196=>"100101110",
  16197=>"110001011",
  16198=>"110100001",
  16199=>"010111100",
  16200=>"101010000",
  16201=>"110101001",
  16202=>"000010001",
  16203=>"000001000",
  16204=>"001100011",
  16205=>"001010110",
  16206=>"101100110",
  16207=>"010101101",
  16208=>"001010011",
  16209=>"101011110",
  16210=>"000011100",
  16211=>"110001011",
  16212=>"100010110",
  16213=>"111010011",
  16214=>"110000011",
  16215=>"000000110",
  16216=>"011001010",
  16217=>"010010110",
  16218=>"100010101",
  16219=>"111111110",
  16220=>"011000110",
  16221=>"101010000",
  16222=>"000001100",
  16223=>"010010000",
  16224=>"001000001",
  16225=>"110111000",
  16226=>"010001011",
  16227=>"110010101",
  16228=>"111110010",
  16229=>"111100100",
  16230=>"101111111",
  16231=>"111111100",
  16232=>"011100011",
  16233=>"011111101",
  16234=>"000111001",
  16235=>"110111000",
  16236=>"110111010",
  16237=>"111110011",
  16238=>"001111101",
  16239=>"110111111",
  16240=>"000001000",
  16241=>"011101010",
  16242=>"011111100",
  16243=>"101010111",
  16244=>"001001000",
  16245=>"010001000",
  16246=>"000101110",
  16247=>"100110000",
  16248=>"011010011",
  16249=>"010100001",
  16250=>"100001110",
  16251=>"010001000",
  16252=>"000000001",
  16253=>"100101111",
  16254=>"101101011",
  16255=>"001111010",
  16256=>"100101100",
  16257=>"111001111",
  16258=>"111011101",
  16259=>"100111111",
  16260=>"100111011",
  16261=>"110101000",
  16262=>"000111101",
  16263=>"000100111",
  16264=>"001111011",
  16265=>"110111000",
  16266=>"111010000",
  16267=>"101111011",
  16268=>"111111100",
  16269=>"000011000",
  16270=>"111101011",
  16271=>"001001110",
  16272=>"111111011",
  16273=>"101100110",
  16274=>"011010011",
  16275=>"111000100",
  16276=>"001011110",
  16277=>"000000010",
  16278=>"111001111",
  16279=>"010000100",
  16280=>"111000010",
  16281=>"110101110",
  16282=>"111110110",
  16283=>"110010010",
  16284=>"011101100",
  16285=>"110011010",
  16286=>"011011010",
  16287=>"111101110",
  16288=>"111110001",
  16289=>"101100111",
  16290=>"100110110",
  16291=>"001101000",
  16292=>"101111010",
  16293=>"111010111",
  16294=>"110001101",
  16295=>"111001111",
  16296=>"101011111",
  16297=>"011100111",
  16298=>"111101011",
  16299=>"001111011",
  16300=>"110110011",
  16301=>"000001010",
  16302=>"100101000",
  16303=>"010100101",
  16304=>"101100110",
  16305=>"111101010",
  16306=>"101000101",
  16307=>"111111000",
  16308=>"000101110",
  16309=>"100100110",
  16310=>"101100011",
  16311=>"100010011",
  16312=>"010010001",
  16313=>"100111101",
  16314=>"100101100",
  16315=>"111011000",
  16316=>"111001100",
  16317=>"010101001",
  16318=>"000001001",
  16319=>"111110101",
  16320=>"010101010",
  16321=>"001100010",
  16322=>"111110000",
  16323=>"111010000",
  16324=>"100010101",
  16325=>"011111110",
  16326=>"011011000",
  16327=>"000001100",
  16328=>"000001110",
  16329=>"001000010",
  16330=>"010001101",
  16331=>"110000010",
  16332=>"001011000",
  16333=>"000000010",
  16334=>"111010011",
  16335=>"100000111",
  16336=>"111000000",
  16337=>"000111001",
  16338=>"000001000",
  16339=>"000010011",
  16340=>"000100000",
  16341=>"100011110",
  16342=>"110000110",
  16343=>"111000101",
  16344=>"001001101",
  16345=>"001111000",
  16346=>"111101111",
  16347=>"110000100",
  16348=>"110001011",
  16349=>"101110101",
  16350=>"010011011",
  16351=>"010011100",
  16352=>"110110001",
  16353=>"110010111",
  16354=>"011000001",
  16355=>"000001111",
  16356=>"101100100",
  16357=>"100111000",
  16358=>"111110110",
  16359=>"011010000",
  16360=>"111011101",
  16361=>"010101000",
  16362=>"110101100",
  16363=>"000000111",
  16364=>"011010100",
  16365=>"011111101",
  16366=>"001000111",
  16367=>"101110100",
  16368=>"010000110",
  16369=>"001110101",
  16370=>"010100010",
  16371=>"110110000",
  16372=>"101110000",
  16373=>"000101110",
  16374=>"000010110",
  16375=>"111010011",
  16376=>"010101111",
  16377=>"111011101",
  16378=>"100100100",
  16379=>"111000011",
  16380=>"111010101",
  16381=>"110000000",
  16382=>"111010100",
  16383=>"001111000",
  16384=>"010000001",
  16385=>"100011101",
  16386=>"010100000",
  16387=>"110010101",
  16388=>"110101101",
  16389=>"101001011",
  16390=>"101110010",
  16391=>"010001011",
  16392=>"100010000",
  16393=>"100010011",
  16394=>"111011011",
  16395=>"101100010",
  16396=>"000111000",
  16397=>"010011011",
  16398=>"100101010",
  16399=>"101110111",
  16400=>"010110100",
  16401=>"100100110",
  16402=>"110100111",
  16403=>"110101111",
  16404=>"010011001",
  16405=>"000010101",
  16406=>"101110000",
  16407=>"000000011",
  16408=>"100111001",
  16409=>"000010110",
  16410=>"011101100",
  16411=>"100100111",
  16412=>"100010010",
  16413=>"110101010",
  16414=>"010010101",
  16415=>"100111010",
  16416=>"000110100",
  16417=>"100101011",
  16418=>"110011000",
  16419=>"111001000",
  16420=>"101011010",
  16421=>"010101111",
  16422=>"110111100",
  16423=>"110011010",
  16424=>"010010100",
  16425=>"111010010",
  16426=>"001000101",
  16427=>"010110001",
  16428=>"010101011",
  16429=>"000000110",
  16430=>"001010111",
  16431=>"111111011",
  16432=>"100001111",
  16433=>"011100000",
  16434=>"011011000",
  16435=>"010111000",
  16436=>"111101111",
  16437=>"110100111",
  16438=>"100001000",
  16439=>"011011011",
  16440=>"000110010",
  16441=>"010111011",
  16442=>"000110011",
  16443=>"110100010",
  16444=>"010001100",
  16445=>"001000111",
  16446=>"110000100",
  16447=>"100010101",
  16448=>"011001010",
  16449=>"101001100",
  16450=>"001100000",
  16451=>"011101001",
  16452=>"010001001",
  16453=>"000010001",
  16454=>"001001101",
  16455=>"010011100",
  16456=>"001001110",
  16457=>"100111011",
  16458=>"100110111",
  16459=>"111110001",
  16460=>"010010101",
  16461=>"001011001",
  16462=>"000010010",
  16463=>"100000011",
  16464=>"000011110",
  16465=>"000011101",
  16466=>"011001111",
  16467=>"101100101",
  16468=>"111000110",
  16469=>"001000111",
  16470=>"000011011",
  16471=>"000000010",
  16472=>"000011010",
  16473=>"011011101",
  16474=>"000010010",
  16475=>"011100001",
  16476=>"111100010",
  16477=>"011011010",
  16478=>"100111101",
  16479=>"100000011",
  16480=>"101100001",
  16481=>"111001000",
  16482=>"011111001",
  16483=>"011111110",
  16484=>"011000001",
  16485=>"111111110",
  16486=>"001010110",
  16487=>"011110111",
  16488=>"000110111",
  16489=>"000111000",
  16490=>"101010101",
  16491=>"000101000",
  16492=>"011000100",
  16493=>"010101101",
  16494=>"100100011",
  16495=>"110100100",
  16496=>"110000000",
  16497=>"000000010",
  16498=>"000010101",
  16499=>"101101100",
  16500=>"011001010",
  16501=>"010110011",
  16502=>"110000100",
  16503=>"111110011",
  16504=>"000111001",
  16505=>"000110010",
  16506=>"010101011",
  16507=>"101001100",
  16508=>"010000100",
  16509=>"100100000",
  16510=>"100100010",
  16511=>"101110000",
  16512=>"001101000",
  16513=>"011111100",
  16514=>"101001101",
  16515=>"111011110",
  16516=>"100000100",
  16517=>"110100110",
  16518=>"000001001",
  16519=>"101111000",
  16520=>"000100101",
  16521=>"110101001",
  16522=>"000000010",
  16523=>"000001101",
  16524=>"111101011",
  16525=>"000011001",
  16526=>"001001110",
  16527=>"100011000",
  16528=>"101100110",
  16529=>"100111000",
  16530=>"001110101",
  16531=>"111100111",
  16532=>"110101111",
  16533=>"100110000",
  16534=>"000001000",
  16535=>"110101111",
  16536=>"000001010",
  16537=>"001010110",
  16538=>"101111101",
  16539=>"110011001",
  16540=>"001101111",
  16541=>"100010010",
  16542=>"010100110",
  16543=>"011010110",
  16544=>"101000011",
  16545=>"101100010",
  16546=>"100011111",
  16547=>"001110010",
  16548=>"001001111",
  16549=>"001000011",
  16550=>"100100011",
  16551=>"001110010",
  16552=>"010001110",
  16553=>"101111010",
  16554=>"000000000",
  16555=>"110111100",
  16556=>"001001001",
  16557=>"001111100",
  16558=>"010001011",
  16559=>"001010100",
  16560=>"110101010",
  16561=>"111110011",
  16562=>"100101010",
  16563=>"000101011",
  16564=>"101000111",
  16565=>"001110111",
  16566=>"011000001",
  16567=>"101111111",
  16568=>"011011111",
  16569=>"100000010",
  16570=>"110000110",
  16571=>"111111011",
  16572=>"010010001",
  16573=>"010100010",
  16574=>"010001011",
  16575=>"000110110",
  16576=>"001010001",
  16577=>"000011010",
  16578=>"100001100",
  16579=>"000110111",
  16580=>"010001100",
  16581=>"110010011",
  16582=>"111111100",
  16583=>"001101110",
  16584=>"111000001",
  16585=>"111100000",
  16586=>"010011010",
  16587=>"110001110",
  16588=>"000111100",
  16589=>"000000010",
  16590=>"011011000",
  16591=>"111001010",
  16592=>"111010001",
  16593=>"101110110",
  16594=>"001000001",
  16595=>"000101101",
  16596=>"100010111",
  16597=>"001110000",
  16598=>"110111001",
  16599=>"001010000",
  16600=>"001010011",
  16601=>"110001000",
  16602=>"011101101",
  16603=>"000011001",
  16604=>"010011110",
  16605=>"101000100",
  16606=>"010011000",
  16607=>"011111100",
  16608=>"110111011",
  16609=>"110101011",
  16610=>"100001001",
  16611=>"110101001",
  16612=>"010101101",
  16613=>"101101110",
  16614=>"110110101",
  16615=>"111111111",
  16616=>"111110011",
  16617=>"111111000",
  16618=>"000110100",
  16619=>"101000010",
  16620=>"101110110",
  16621=>"000111000",
  16622=>"011000001",
  16623=>"110000110",
  16624=>"010001110",
  16625=>"010100110",
  16626=>"011100001",
  16627=>"110000000",
  16628=>"001001010",
  16629=>"110110010",
  16630=>"011111011",
  16631=>"010000010",
  16632=>"110101111",
  16633=>"010100011",
  16634=>"001100001",
  16635=>"010000000",
  16636=>"000101001",
  16637=>"011011110",
  16638=>"010101010",
  16639=>"000000101",
  16640=>"000001100",
  16641=>"000000000",
  16642=>"001110111",
  16643=>"011011011",
  16644=>"110010001",
  16645=>"010110101",
  16646=>"111000101",
  16647=>"001000110",
  16648=>"000111111",
  16649=>"001001101",
  16650=>"100101111",
  16651=>"101001001",
  16652=>"001101001",
  16653=>"000100111",
  16654=>"000001110",
  16655=>"000100101",
  16656=>"110111101",
  16657=>"001110001",
  16658=>"010011000",
  16659=>"101110001",
  16660=>"110101110",
  16661=>"001001110",
  16662=>"111111110",
  16663=>"110111111",
  16664=>"000111011",
  16665=>"000000100",
  16666=>"111101011",
  16667=>"100011110",
  16668=>"001000010",
  16669=>"110110100",
  16670=>"010001011",
  16671=>"110001000",
  16672=>"010101000",
  16673=>"000000000",
  16674=>"010010100",
  16675=>"000000101",
  16676=>"000000111",
  16677=>"100000111",
  16678=>"110110011",
  16679=>"011001011",
  16680=>"011001010",
  16681=>"000001111",
  16682=>"101001001",
  16683=>"010111110",
  16684=>"001110100",
  16685=>"011001010",
  16686=>"111010110",
  16687=>"111110001",
  16688=>"100110010",
  16689=>"111001111",
  16690=>"001010000",
  16691=>"001011011",
  16692=>"010111110",
  16693=>"010111110",
  16694=>"110000100",
  16695=>"111000000",
  16696=>"110101000",
  16697=>"100000001",
  16698=>"110100010",
  16699=>"100110110",
  16700=>"110011100",
  16701=>"110101111",
  16702=>"100111001",
  16703=>"111101000",
  16704=>"001111111",
  16705=>"001011110",
  16706=>"000010110",
  16707=>"111100011",
  16708=>"111111011",
  16709=>"000010110",
  16710=>"011100010",
  16711=>"110011101",
  16712=>"111010101",
  16713=>"011010100",
  16714=>"000010101",
  16715=>"000001101",
  16716=>"101000000",
  16717=>"000010010",
  16718=>"101111110",
  16719=>"101001010",
  16720=>"111000000",
  16721=>"110100011",
  16722=>"000001010",
  16723=>"001110001",
  16724=>"111010011",
  16725=>"000010101",
  16726=>"101111001",
  16727=>"011011110",
  16728=>"010110011",
  16729=>"111000111",
  16730=>"001010010",
  16731=>"111010011",
  16732=>"101011101",
  16733=>"011111111",
  16734=>"110101010",
  16735=>"110110111",
  16736=>"110111000",
  16737=>"111011011",
  16738=>"101011001",
  16739=>"111110100",
  16740=>"101111111",
  16741=>"010011100",
  16742=>"010001110",
  16743=>"001111110",
  16744=>"011011111",
  16745=>"011101101",
  16746=>"101010101",
  16747=>"111001000",
  16748=>"100101110",
  16749=>"011111011",
  16750=>"111001011",
  16751=>"010110000",
  16752=>"010001100",
  16753=>"001001010",
  16754=>"101000011",
  16755=>"110100000",
  16756=>"110001001",
  16757=>"100101011",
  16758=>"100111111",
  16759=>"111111111",
  16760=>"010000101",
  16761=>"010001110",
  16762=>"000000001",
  16763=>"111100111",
  16764=>"011011101",
  16765=>"111111110",
  16766=>"110010101",
  16767=>"000010011",
  16768=>"100001110",
  16769=>"100111100",
  16770=>"101000101",
  16771=>"011001011",
  16772=>"000010011",
  16773=>"010110101",
  16774=>"001000100",
  16775=>"001100110",
  16776=>"011011010",
  16777=>"010000101",
  16778=>"111110011",
  16779=>"111100100",
  16780=>"000011100",
  16781=>"010101101",
  16782=>"011101000",
  16783=>"111010001",
  16784=>"010011001",
  16785=>"000001000",
  16786=>"111010110",
  16787=>"000001001",
  16788=>"110100111",
  16789=>"111101011",
  16790=>"111111110",
  16791=>"111111100",
  16792=>"001111111",
  16793=>"010000101",
  16794=>"101100010",
  16795=>"001011101",
  16796=>"100010101",
  16797=>"000110110",
  16798=>"000000110",
  16799=>"111101111",
  16800=>"000010010",
  16801=>"101111111",
  16802=>"001101011",
  16803=>"000011010",
  16804=>"001111100",
  16805=>"101110100",
  16806=>"011011100",
  16807=>"100010100",
  16808=>"111010111",
  16809=>"110000010",
  16810=>"100000000",
  16811=>"100100100",
  16812=>"110011100",
  16813=>"111101101",
  16814=>"001000100",
  16815=>"000000010",
  16816=>"000001101",
  16817=>"110101111",
  16818=>"100101110",
  16819=>"101010000",
  16820=>"000010000",
  16821=>"010010010",
  16822=>"010010111",
  16823=>"110010000",
  16824=>"010100101",
  16825=>"110010000",
  16826=>"101100100",
  16827=>"011010000",
  16828=>"101010101",
  16829=>"110110110",
  16830=>"001111011",
  16831=>"100010000",
  16832=>"000110001",
  16833=>"000011110",
  16834=>"010110010",
  16835=>"011001101",
  16836=>"001110011",
  16837=>"011100101",
  16838=>"101001011",
  16839=>"001100000",
  16840=>"110011101",
  16841=>"101111010",
  16842=>"101100110",
  16843=>"101010000",
  16844=>"111111101",
  16845=>"001101011",
  16846=>"111100001",
  16847=>"111000001",
  16848=>"100000000",
  16849=>"010101111",
  16850=>"100111101",
  16851=>"001001010",
  16852=>"001100101",
  16853=>"110010101",
  16854=>"100000000",
  16855=>"000110100",
  16856=>"001100110",
  16857=>"000011011",
  16858=>"001100101",
  16859=>"000001111",
  16860=>"010011100",
  16861=>"000110111",
  16862=>"110110000",
  16863=>"110110100",
  16864=>"110110100",
  16865=>"001111011",
  16866=>"111011111",
  16867=>"111110101",
  16868=>"100000000",
  16869=>"101010011",
  16870=>"101110001",
  16871=>"111011110",
  16872=>"000000010",
  16873=>"101001111",
  16874=>"011100100",
  16875=>"110110000",
  16876=>"000010100",
  16877=>"110000100",
  16878=>"011010000",
  16879=>"101011111",
  16880=>"101001001",
  16881=>"000101000",
  16882=>"111001100",
  16883=>"111000001",
  16884=>"100110100",
  16885=>"101001101",
  16886=>"101011110",
  16887=>"000011000",
  16888=>"010101100",
  16889=>"110011110",
  16890=>"010000000",
  16891=>"011010100",
  16892=>"100010111",
  16893=>"011101111",
  16894=>"011000100",
  16895=>"001001001",
  16896=>"100000010",
  16897=>"111011011",
  16898=>"110111100",
  16899=>"010101111",
  16900=>"011100010",
  16901=>"010101001",
  16902=>"010000111",
  16903=>"001010111",
  16904=>"010100101",
  16905=>"100101110",
  16906=>"001000101",
  16907=>"100110000",
  16908=>"101000010",
  16909=>"010110001",
  16910=>"110010111",
  16911=>"010100010",
  16912=>"111000010",
  16913=>"110001011",
  16914=>"000001000",
  16915=>"010111011",
  16916=>"010100100",
  16917=>"110000101",
  16918=>"100100101",
  16919=>"100011101",
  16920=>"100001010",
  16921=>"000111001",
  16922=>"001110100",
  16923=>"111110110",
  16924=>"110101100",
  16925=>"001010011",
  16926=>"101111000",
  16927=>"000101000",
  16928=>"000011110",
  16929=>"101110101",
  16930=>"110101101",
  16931=>"101110010",
  16932=>"010011000",
  16933=>"010010101",
  16934=>"010111110",
  16935=>"011110101",
  16936=>"000000100",
  16937=>"011011110",
  16938=>"001111000",
  16939=>"001001010",
  16940=>"011110000",
  16941=>"100001000",
  16942=>"111011110",
  16943=>"101001010",
  16944=>"100000001",
  16945=>"000101101",
  16946=>"101101110",
  16947=>"011000101",
  16948=>"010001001",
  16949=>"000001100",
  16950=>"111100100",
  16951=>"001111111",
  16952=>"100111110",
  16953=>"110110100",
  16954=>"110011001",
  16955=>"101100111",
  16956=>"111111010",
  16957=>"000110100",
  16958=>"101000010",
  16959=>"010000001",
  16960=>"110110100",
  16961=>"001001011",
  16962=>"101010100",
  16963=>"000101011",
  16964=>"110110101",
  16965=>"011001101",
  16966=>"100000100",
  16967=>"000011011",
  16968=>"001010110",
  16969=>"101001001",
  16970=>"111000100",
  16971=>"000101100",
  16972=>"111100011",
  16973=>"101101101",
  16974=>"110011111",
  16975=>"101011010",
  16976=>"110001001",
  16977=>"111011010",
  16978=>"100010000",
  16979=>"100001010",
  16980=>"110000010",
  16981=>"110100110",
  16982=>"010110011",
  16983=>"111010111",
  16984=>"100101110",
  16985=>"011101101",
  16986=>"000001100",
  16987=>"101101110",
  16988=>"101111001",
  16989=>"001011001",
  16990=>"110111101",
  16991=>"000011000",
  16992=>"100000110",
  16993=>"000011111",
  16994=>"101001101",
  16995=>"000010000",
  16996=>"100111101",
  16997=>"100010011",
  16998=>"011100001",
  16999=>"010100010",
  17000=>"110001010",
  17001=>"100101101",
  17002=>"100111110",
  17003=>"111001110",
  17004=>"110100001",
  17005=>"101000110",
  17006=>"111000001",
  17007=>"010011010",
  17008=>"000001110",
  17009=>"001110000",
  17010=>"111000000",
  17011=>"110100100",
  17012=>"100100010",
  17013=>"001011111",
  17014=>"111000010",
  17015=>"010011101",
  17016=>"111001110",
  17017=>"000011001",
  17018=>"001110011",
  17019=>"000100111",
  17020=>"110101001",
  17021=>"000010101",
  17022=>"001000001",
  17023=>"010101001",
  17024=>"100010110",
  17025=>"111110110",
  17026=>"000100000",
  17027=>"001101000",
  17028=>"110111111",
  17029=>"101001011",
  17030=>"010100001",
  17031=>"110111111",
  17032=>"100011110",
  17033=>"001010101",
  17034=>"000101100",
  17035=>"101011101",
  17036=>"011101011",
  17037=>"101001111",
  17038=>"100111101",
  17039=>"010000111",
  17040=>"101011001",
  17041=>"011000100",
  17042=>"010100011",
  17043=>"101101011",
  17044=>"111110010",
  17045=>"001111100",
  17046=>"111111101",
  17047=>"101000100",
  17048=>"011100111",
  17049=>"110011110",
  17050=>"110101000",
  17051=>"100101110",
  17052=>"101110001",
  17053=>"001111110",
  17054=>"111111000",
  17055=>"000000000",
  17056=>"111111101",
  17057=>"001111011",
  17058=>"010001000",
  17059=>"111010100",
  17060=>"100000101",
  17061=>"111111101",
  17062=>"010111110",
  17063=>"111111000",
  17064=>"101001111",
  17065=>"001110010",
  17066=>"111011010",
  17067=>"010100011",
  17068=>"001110001",
  17069=>"010010101",
  17070=>"101111000",
  17071=>"101000001",
  17072=>"010010011",
  17073=>"011011001",
  17074=>"111101010",
  17075=>"000001111",
  17076=>"010001100",
  17077=>"101000101",
  17078=>"100111011",
  17079=>"100010010",
  17080=>"011100010",
  17081=>"110001100",
  17082=>"100000100",
  17083=>"110011010",
  17084=>"000110001",
  17085=>"000110001",
  17086=>"011110100",
  17087=>"100100001",
  17088=>"000010011",
  17089=>"110011111",
  17090=>"111111100",
  17091=>"010100001",
  17092=>"111001010",
  17093=>"011101111",
  17094=>"010111011",
  17095=>"010000111",
  17096=>"000110010",
  17097=>"000111001",
  17098=>"111111011",
  17099=>"010000001",
  17100=>"111110101",
  17101=>"110101101",
  17102=>"001010111",
  17103=>"101110111",
  17104=>"110111101",
  17105=>"111100011",
  17106=>"110001000",
  17107=>"010101111",
  17108=>"010000010",
  17109=>"000110001",
  17110=>"100011000",
  17111=>"100101001",
  17112=>"011111000",
  17113=>"011101000",
  17114=>"010010001",
  17115=>"000111111",
  17116=>"011111011",
  17117=>"011110101",
  17118=>"011110011",
  17119=>"001000001",
  17120=>"100110100",
  17121=>"010010011",
  17122=>"110011110",
  17123=>"010111000",
  17124=>"111000110",
  17125=>"101101011",
  17126=>"100100000",
  17127=>"010111010",
  17128=>"000101101",
  17129=>"100101001",
  17130=>"000110011",
  17131=>"010011110",
  17132=>"010000001",
  17133=>"010001010",
  17134=>"111011100",
  17135=>"111000011",
  17136=>"100111111",
  17137=>"001101001",
  17138=>"011001010",
  17139=>"010011000",
  17140=>"000001101",
  17141=>"011010011",
  17142=>"011101100",
  17143=>"001101100",
  17144=>"000011111",
  17145=>"100000011",
  17146=>"010010000",
  17147=>"001110111",
  17148=>"111111100",
  17149=>"111010110",
  17150=>"110001010",
  17151=>"110010001",
  17152=>"100011111",
  17153=>"001010101",
  17154=>"000110000",
  17155=>"000001001",
  17156=>"001100111",
  17157=>"011100000",
  17158=>"101010100",
  17159=>"101100001",
  17160=>"111010011",
  17161=>"110111110",
  17162=>"111011000",
  17163=>"000000111",
  17164=>"000110110",
  17165=>"000001011",
  17166=>"111100011",
  17167=>"000011110",
  17168=>"011111110",
  17169=>"001100111",
  17170=>"001100001",
  17171=>"000101011",
  17172=>"010000101",
  17173=>"011001111",
  17174=>"100010101",
  17175=>"110010101",
  17176=>"011001100",
  17177=>"010110111",
  17178=>"010001101",
  17179=>"111101000",
  17180=>"111111010",
  17181=>"010101000",
  17182=>"010110100",
  17183=>"100101011",
  17184=>"001000001",
  17185=>"000101011",
  17186=>"001100011",
  17187=>"100001011",
  17188=>"000110100",
  17189=>"110111111",
  17190=>"111110001",
  17191=>"011111111",
  17192=>"010111111",
  17193=>"000010011",
  17194=>"011111010",
  17195=>"010011000",
  17196=>"100100110",
  17197=>"110100000",
  17198=>"101011000",
  17199=>"001000111",
  17200=>"100100010",
  17201=>"110111001",
  17202=>"101011000",
  17203=>"011100000",
  17204=>"000010111",
  17205=>"011010101",
  17206=>"100111100",
  17207=>"110010000",
  17208=>"101011010",
  17209=>"110011111",
  17210=>"011001011",
  17211=>"101010101",
  17212=>"001111100",
  17213=>"101000011",
  17214=>"000010110",
  17215=>"010111110",
  17216=>"011101110",
  17217=>"111001100",
  17218=>"000000001",
  17219=>"100011111",
  17220=>"110001001",
  17221=>"100000101",
  17222=>"111100010",
  17223=>"100111001",
  17224=>"110101111",
  17225=>"000101010",
  17226=>"101010110",
  17227=>"111010100",
  17228=>"000011110",
  17229=>"000100111",
  17230=>"001000110",
  17231=>"101010000",
  17232=>"011010000",
  17233=>"000000111",
  17234=>"000111010",
  17235=>"001000011",
  17236=>"000110111",
  17237=>"110001110",
  17238=>"000111001",
  17239=>"111111110",
  17240=>"110000111",
  17241=>"001101111",
  17242=>"001000010",
  17243=>"111000101",
  17244=>"101101011",
  17245=>"001110100",
  17246=>"000101110",
  17247=>"111111101",
  17248=>"001010010",
  17249=>"010100111",
  17250=>"111101011",
  17251=>"000011101",
  17252=>"101111011",
  17253=>"110001110",
  17254=>"011010010",
  17255=>"000101101",
  17256=>"010001110",
  17257=>"001100000",
  17258=>"110111010",
  17259=>"001000111",
  17260=>"000100001",
  17261=>"010110000",
  17262=>"110001110",
  17263=>"000110000",
  17264=>"110110101",
  17265=>"100100000",
  17266=>"000100001",
  17267=>"100111000",
  17268=>"001000101",
  17269=>"100010110",
  17270=>"110010110",
  17271=>"101101110",
  17272=>"010011110",
  17273=>"101111101",
  17274=>"110001100",
  17275=>"100111110",
  17276=>"000110110",
  17277=>"000100000",
  17278=>"001011010",
  17279=>"000001011",
  17280=>"100010010",
  17281=>"101000110",
  17282=>"011001011",
  17283=>"011111111",
  17284=>"001111110",
  17285=>"111001101",
  17286=>"010110011",
  17287=>"001111011",
  17288=>"010001000",
  17289=>"101000100",
  17290=>"111110011",
  17291=>"000100010",
  17292=>"101100011",
  17293=>"100001111",
  17294=>"100100000",
  17295=>"101010010",
  17296=>"010000010",
  17297=>"110111110",
  17298=>"001010111",
  17299=>"110100101",
  17300=>"101000111",
  17301=>"111101110",
  17302=>"000111010",
  17303=>"000101101",
  17304=>"101111000",
  17305=>"001100100",
  17306=>"111100000",
  17307=>"110111010",
  17308=>"010000001",
  17309=>"001101000",
  17310=>"110100010",
  17311=>"101101011",
  17312=>"101011001",
  17313=>"110000011",
  17314=>"001111010",
  17315=>"110000001",
  17316=>"100101111",
  17317=>"011001100",
  17318=>"101101011",
  17319=>"000011010",
  17320=>"001001100",
  17321=>"000010011",
  17322=>"110000110",
  17323=>"111110010",
  17324=>"011000000",
  17325=>"001011000",
  17326=>"111101100",
  17327=>"010111110",
  17328=>"010001001",
  17329=>"011011110",
  17330=>"000111010",
  17331=>"010001100",
  17332=>"011011010",
  17333=>"111001000",
  17334=>"000110110",
  17335=>"001100000",
  17336=>"100001000",
  17337=>"111101111",
  17338=>"010101101",
  17339=>"011100110",
  17340=>"111110001",
  17341=>"001000101",
  17342=>"000010001",
  17343=>"010000110",
  17344=>"000100011",
  17345=>"010100101",
  17346=>"111110100",
  17347=>"010011001",
  17348=>"101111111",
  17349=>"100101010",
  17350=>"110110110",
  17351=>"000001011",
  17352=>"110000001",
  17353=>"010110001",
  17354=>"010000110",
  17355=>"100011000",
  17356=>"100010101",
  17357=>"000111100",
  17358=>"111000011",
  17359=>"001111000",
  17360=>"011110101",
  17361=>"011001010",
  17362=>"110010001",
  17363=>"100001100",
  17364=>"011111100",
  17365=>"111000001",
  17366=>"010000101",
  17367=>"101101100",
  17368=>"001011110",
  17369=>"101100101",
  17370=>"000110111",
  17371=>"001001001",
  17372=>"101001001",
  17373=>"010010011",
  17374=>"100011101",
  17375=>"100011001",
  17376=>"100111111",
  17377=>"000011110",
  17378=>"010011001",
  17379=>"001001010",
  17380=>"110100000",
  17381=>"110011011",
  17382=>"011100000",
  17383=>"000100010",
  17384=>"010011011",
  17385=>"011101000",
  17386=>"100010011",
  17387=>"101001111",
  17388=>"010101010",
  17389=>"111101101",
  17390=>"010001101",
  17391=>"101010000",
  17392=>"010101001",
  17393=>"000101010",
  17394=>"110100001",
  17395=>"011101010",
  17396=>"100001111",
  17397=>"000100010",
  17398=>"111001001",
  17399=>"001011100",
  17400=>"110000000",
  17401=>"010100000",
  17402=>"011011101",
  17403=>"100000011",
  17404=>"010000011",
  17405=>"000001100",
  17406=>"101110110",
  17407=>"100110100",
  17408=>"010101000",
  17409=>"100011001",
  17410=>"110111110",
  17411=>"011000001",
  17412=>"000110101",
  17413=>"010000001",
  17414=>"010100000",
  17415=>"110110110",
  17416=>"101100011",
  17417=>"001100011",
  17418=>"010110100",
  17419=>"111011110",
  17420=>"011110110",
  17421=>"101001110",
  17422=>"000000101",
  17423=>"001100100",
  17424=>"110000111",
  17425=>"111011000",
  17426=>"111101000",
  17427=>"110011111",
  17428=>"000100001",
  17429=>"010111010",
  17430=>"010111110",
  17431=>"110011111",
  17432=>"110000110",
  17433=>"000100110",
  17434=>"110111010",
  17435=>"101101111",
  17436=>"001010101",
  17437=>"001010111",
  17438=>"011100010",
  17439=>"111110010",
  17440=>"111101100",
  17441=>"100101111",
  17442=>"111110101",
  17443=>"011010000",
  17444=>"110110111",
  17445=>"000011111",
  17446=>"101111010",
  17447=>"110110101",
  17448=>"100000010",
  17449=>"001111111",
  17450=>"011011000",
  17451=>"001010000",
  17452=>"101101111",
  17453=>"000101101",
  17454=>"010100100",
  17455=>"110000110",
  17456=>"110010011",
  17457=>"000011010",
  17458=>"000001101",
  17459=>"101001110",
  17460=>"111100101",
  17461=>"101110000",
  17462=>"111110110",
  17463=>"001001001",
  17464=>"011010011",
  17465=>"011000001",
  17466=>"111011000",
  17467=>"110110111",
  17468=>"011100000",
  17469=>"101111011",
  17470=>"001010000",
  17471=>"111100101",
  17472=>"111110001",
  17473=>"111001001",
  17474=>"010001011",
  17475=>"111011000",
  17476=>"001001001",
  17477=>"000110101",
  17478=>"111100101",
  17479=>"101110110",
  17480=>"010001011",
  17481=>"011111011",
  17482=>"001010001",
  17483=>"001011111",
  17484=>"101011011",
  17485=>"111000111",
  17486=>"010010100",
  17487=>"100111000",
  17488=>"001111100",
  17489=>"101100100",
  17490=>"000001010",
  17491=>"100001001",
  17492=>"011011000",
  17493=>"011000100",
  17494=>"010110011",
  17495=>"101101001",
  17496=>"011010010",
  17497=>"011101110",
  17498=>"110011000",
  17499=>"100001110",
  17500=>"000101010",
  17501=>"001101010",
  17502=>"100111000",
  17503=>"110110101",
  17504=>"110100011",
  17505=>"011111011",
  17506=>"011100100",
  17507=>"001011011",
  17508=>"110010011",
  17509=>"010001010",
  17510=>"100011111",
  17511=>"010111000",
  17512=>"010101001",
  17513=>"010001110",
  17514=>"001101000",
  17515=>"111110110",
  17516=>"001100111",
  17517=>"000110011",
  17518=>"010110011",
  17519=>"101000110",
  17520=>"110001011",
  17521=>"100100101",
  17522=>"011100101",
  17523=>"101100100",
  17524=>"010100001",
  17525=>"001100001",
  17526=>"111010100",
  17527=>"001111110",
  17528=>"000100100",
  17529=>"010100110",
  17530=>"111001010",
  17531=>"000001000",
  17532=>"000100011",
  17533=>"111100110",
  17534=>"000000100",
  17535=>"111111010",
  17536=>"001110011",
  17537=>"101111111",
  17538=>"111101011",
  17539=>"110000011",
  17540=>"101110111",
  17541=>"000111001",
  17542=>"001001001",
  17543=>"111101001",
  17544=>"110001111",
  17545=>"101000011",
  17546=>"100001011",
  17547=>"000111000",
  17548=>"111010000",
  17549=>"101000010",
  17550=>"010100010",
  17551=>"000010001",
  17552=>"011110010",
  17553=>"001101111",
  17554=>"111011001",
  17555=>"000001110",
  17556=>"011001010",
  17557=>"101111010",
  17558=>"111101101",
  17559=>"100000010",
  17560=>"010001111",
  17561=>"101100111",
  17562=>"010100001",
  17563=>"000001010",
  17564=>"010000101",
  17565=>"110011101",
  17566=>"110111100",
  17567=>"110011010",
  17568=>"111100011",
  17569=>"101100110",
  17570=>"010111111",
  17571=>"001110010",
  17572=>"010011101",
  17573=>"001001000",
  17574=>"010000110",
  17575=>"100011111",
  17576=>"011011010",
  17577=>"101010010",
  17578=>"110000010",
  17579=>"000111111",
  17580=>"111111011",
  17581=>"100101100",
  17582=>"110110100",
  17583=>"111011100",
  17584=>"111101110",
  17585=>"110000011",
  17586=>"110111001",
  17587=>"001101010",
  17588=>"001001001",
  17589=>"011000010",
  17590=>"000001101",
  17591=>"011010001",
  17592=>"110111111",
  17593=>"011011100",
  17594=>"100101111",
  17595=>"110111110",
  17596=>"010011101",
  17597=>"000010101",
  17598=>"101011101",
  17599=>"011010001",
  17600=>"011001111",
  17601=>"010000110",
  17602=>"100000111",
  17603=>"000111111",
  17604=>"111110100",
  17605=>"100111000",
  17606=>"000000001",
  17607=>"011110101",
  17608=>"010010011",
  17609=>"100100110",
  17610=>"011010110",
  17611=>"000010011",
  17612=>"001101100",
  17613=>"001100100",
  17614=>"000100101",
  17615=>"001001100",
  17616=>"001001010",
  17617=>"011101110",
  17618=>"100110011",
  17619=>"010101111",
  17620=>"111101001",
  17621=>"011011100",
  17622=>"010000101",
  17623=>"000010010",
  17624=>"100110001",
  17625=>"110010100",
  17626=>"111001001",
  17627=>"100111100",
  17628=>"010101111",
  17629=>"100011010",
  17630=>"110101110",
  17631=>"011110101",
  17632=>"110110110",
  17633=>"111111011",
  17634=>"111000110",
  17635=>"001110100",
  17636=>"000001000",
  17637=>"100100100",
  17638=>"010011110",
  17639=>"110011001",
  17640=>"000101001",
  17641=>"011011001",
  17642=>"000010100",
  17643=>"100101101",
  17644=>"100010000",
  17645=>"110010100",
  17646=>"000001010",
  17647=>"111101000",
  17648=>"011010000",
  17649=>"111111011",
  17650=>"101000101",
  17651=>"101000110",
  17652=>"100110011",
  17653=>"011110111",
  17654=>"110001010",
  17655=>"110100100",
  17656=>"110101110",
  17657=>"100001100",
  17658=>"110001000",
  17659=>"100100110",
  17660=>"110011000",
  17661=>"001010101",
  17662=>"011010110",
  17663=>"110101101",
  17664=>"111111111",
  17665=>"111000000",
  17666=>"011010100",
  17667=>"011010110",
  17668=>"011001011",
  17669=>"010001111",
  17670=>"001111010",
  17671=>"100000001",
  17672=>"000010010",
  17673=>"000110100",
  17674=>"010011011",
  17675=>"100000111",
  17676=>"110000011",
  17677=>"101010001",
  17678=>"101010110",
  17679=>"010000100",
  17680=>"110011010",
  17681=>"100110110",
  17682=>"100111111",
  17683=>"010100011",
  17684=>"101001011",
  17685=>"010011010",
  17686=>"111111110",
  17687=>"110100001",
  17688=>"111011000",
  17689=>"100101111",
  17690=>"011000010",
  17691=>"101011101",
  17692=>"001110011",
  17693=>"000110110",
  17694=>"100011000",
  17695=>"000101101",
  17696=>"000101000",
  17697=>"011100001",
  17698=>"111011111",
  17699=>"011111000",
  17700=>"110110110",
  17701=>"011111101",
  17702=>"010000001",
  17703=>"000001101",
  17704=>"011111110",
  17705=>"111000100",
  17706=>"110111111",
  17707=>"101111011",
  17708=>"110000110",
  17709=>"111000101",
  17710=>"001111011",
  17711=>"000101110",
  17712=>"101000101",
  17713=>"011111011",
  17714=>"100000010",
  17715=>"011011011",
  17716=>"010010001",
  17717=>"111011110",
  17718=>"000111010",
  17719=>"100001000",
  17720=>"110111000",
  17721=>"000111110",
  17722=>"000100111",
  17723=>"111101110",
  17724=>"111011001",
  17725=>"110000011",
  17726=>"111110010",
  17727=>"110001101",
  17728=>"000000000",
  17729=>"100101010",
  17730=>"110011111",
  17731=>"100011000",
  17732=>"010001110",
  17733=>"001100111",
  17734=>"101111110",
  17735=>"011000110",
  17736=>"110110101",
  17737=>"110100001",
  17738=>"000100010",
  17739=>"010001100",
  17740=>"010011010",
  17741=>"000001110",
  17742=>"001100111",
  17743=>"001011010",
  17744=>"111101010",
  17745=>"010010100",
  17746=>"001101010",
  17747=>"000110000",
  17748=>"000000000",
  17749=>"111110101",
  17750=>"110010000",
  17751=>"000111100",
  17752=>"010101101",
  17753=>"110011011",
  17754=>"111110011",
  17755=>"001001001",
  17756=>"110100001",
  17757=>"110010011",
  17758=>"010011100",
  17759=>"110010111",
  17760=>"110000100",
  17761=>"001000111",
  17762=>"000000101",
  17763=>"000000101",
  17764=>"011010001",
  17765=>"100010100",
  17766=>"100100011",
  17767=>"010010001",
  17768=>"000100110",
  17769=>"001000010",
  17770=>"000011011",
  17771=>"000001001",
  17772=>"000111111",
  17773=>"111111011",
  17774=>"000100011",
  17775=>"101001101",
  17776=>"110001001",
  17777=>"100000001",
  17778=>"011101110",
  17779=>"110001010",
  17780=>"010110011",
  17781=>"011010110",
  17782=>"001100110",
  17783=>"101100000",
  17784=>"001010100",
  17785=>"100111100",
  17786=>"100001010",
  17787=>"101110000",
  17788=>"100100011",
  17789=>"010111101",
  17790=>"101111111",
  17791=>"110000001",
  17792=>"011111000",
  17793=>"010100000",
  17794=>"111101010",
  17795=>"101111111",
  17796=>"110001000",
  17797=>"100101010",
  17798=>"001000010",
  17799=>"001100000",
  17800=>"111000011",
  17801=>"001011101",
  17802=>"011001001",
  17803=>"101000011",
  17804=>"011011000",
  17805=>"011001111",
  17806=>"111001000",
  17807=>"111110010",
  17808=>"010100111",
  17809=>"000100001",
  17810=>"000011011",
  17811=>"101111111",
  17812=>"100010000",
  17813=>"111000010",
  17814=>"100000101",
  17815=>"010100110",
  17816=>"001111101",
  17817=>"111001000",
  17818=>"100000101",
  17819=>"110110000",
  17820=>"101000000",
  17821=>"000011100",
  17822=>"001111000",
  17823=>"110101111",
  17824=>"111110000",
  17825=>"000001111",
  17826=>"010000001",
  17827=>"110100001",
  17828=>"100000100",
  17829=>"110000001",
  17830=>"110000100",
  17831=>"110100100",
  17832=>"001111101",
  17833=>"010101010",
  17834=>"000101110",
  17835=>"111010100",
  17836=>"011111110",
  17837=>"110110000",
  17838=>"100001000",
  17839=>"011000110",
  17840=>"111101000",
  17841=>"001000010",
  17842=>"010110000",
  17843=>"101100011",
  17844=>"110000001",
  17845=>"010101011",
  17846=>"010101011",
  17847=>"011011000",
  17848=>"110010110",
  17849=>"001001111",
  17850=>"000110011",
  17851=>"001010100",
  17852=>"110001011",
  17853=>"111100111",
  17854=>"111001011",
  17855=>"101001000",
  17856=>"010001101",
  17857=>"111110001",
  17858=>"011110100",
  17859=>"011110111",
  17860=>"111101000",
  17861=>"110110001",
  17862=>"110101000",
  17863=>"111110100",
  17864=>"001100011",
  17865=>"100110110",
  17866=>"000000101",
  17867=>"010101011",
  17868=>"001010000",
  17869=>"011110000",
  17870=>"100100110",
  17871=>"000110100",
  17872=>"111011111",
  17873=>"111011100",
  17874=>"111110010",
  17875=>"110111111",
  17876=>"010110111",
  17877=>"001101001",
  17878=>"100111100",
  17879=>"000101010",
  17880=>"111000011",
  17881=>"111011100",
  17882=>"111001001",
  17883=>"001011101",
  17884=>"100000111",
  17885=>"011111001",
  17886=>"010011000",
  17887=>"111000011",
  17888=>"001011110",
  17889=>"010011001",
  17890=>"101010010",
  17891=>"000111010",
  17892=>"101011001",
  17893=>"011101110",
  17894=>"100100100",
  17895=>"011110111",
  17896=>"011110011",
  17897=>"101001010",
  17898=>"100110011",
  17899=>"101000110",
  17900=>"100110100",
  17901=>"100000010",
  17902=>"101101001",
  17903=>"111010001",
  17904=>"000110111",
  17905=>"000001001",
  17906=>"100100100",
  17907=>"101111101",
  17908=>"101110111",
  17909=>"110101001",
  17910=>"010101000",
  17911=>"011010100",
  17912=>"111000011",
  17913=>"100110001",
  17914=>"111011111",
  17915=>"010110001",
  17916=>"101001001",
  17917=>"001000100",
  17918=>"100001111",
  17919=>"011100011",
  17920=>"111010110",
  17921=>"010110100",
  17922=>"110010000",
  17923=>"011001111",
  17924=>"011011111",
  17925=>"101111001",
  17926=>"111111110",
  17927=>"011110010",
  17928=>"100010010",
  17929=>"000101000",
  17930=>"101011000",
  17931=>"011010011",
  17932=>"111111010",
  17933=>"011111010",
  17934=>"111000010",
  17935=>"110111001",
  17936=>"000010011",
  17937=>"101011110",
  17938=>"101111000",
  17939=>"100011101",
  17940=>"000101000",
  17941=>"000010000",
  17942=>"100101010",
  17943=>"010110000",
  17944=>"110001000",
  17945=>"101100101",
  17946=>"000111110",
  17947=>"010010110",
  17948=>"011110101",
  17949=>"110001010",
  17950=>"001001110",
  17951=>"011101101",
  17952=>"111001000",
  17953=>"001100100",
  17954=>"010101110",
  17955=>"010111111",
  17956=>"011001000",
  17957=>"110100110",
  17958=>"101011111",
  17959=>"101110100",
  17960=>"100100000",
  17961=>"100011000",
  17962=>"011100001",
  17963=>"101100000",
  17964=>"000000100",
  17965=>"011000000",
  17966=>"111101010",
  17967=>"110001010",
  17968=>"101010101",
  17969=>"111100000",
  17970=>"011000101",
  17971=>"110111010",
  17972=>"010100111",
  17973=>"011000111",
  17974=>"001110111",
  17975=>"011000010",
  17976=>"010110100",
  17977=>"101000000",
  17978=>"011000101",
  17979=>"111110011",
  17980=>"110011010",
  17981=>"011001111",
  17982=>"011110010",
  17983=>"100111110",
  17984=>"110100110",
  17985=>"001110000",
  17986=>"010100000",
  17987=>"001111110",
  17988=>"101100111",
  17989=>"000110111",
  17990=>"100000101",
  17991=>"111101000",
  17992=>"111001111",
  17993=>"100101101",
  17994=>"101101001",
  17995=>"011101011",
  17996=>"000101111",
  17997=>"100111111",
  17998=>"001000010",
  17999=>"010100010",
  18000=>"111110000",
  18001=>"111001010",
  18002=>"100100100",
  18003=>"001101100",
  18004=>"110100111",
  18005=>"010101111",
  18006=>"011000011",
  18007=>"111101100",
  18008=>"010001101",
  18009=>"001101111",
  18010=>"000101110",
  18011=>"011010001",
  18012=>"111110010",
  18013=>"011110000",
  18014=>"000011111",
  18015=>"111000000",
  18016=>"010111111",
  18017=>"010100101",
  18018=>"100010001",
  18019=>"110110110",
  18020=>"101011001",
  18021=>"110110010",
  18022=>"110001111",
  18023=>"110101111",
  18024=>"001110010",
  18025=>"011000110",
  18026=>"100000101",
  18027=>"110011010",
  18028=>"011000101",
  18029=>"100011001",
  18030=>"011011010",
  18031=>"111000100",
  18032=>"000010110",
  18033=>"000010001",
  18034=>"101001101",
  18035=>"001100111",
  18036=>"001000000",
  18037=>"110101011",
  18038=>"110111100",
  18039=>"101101000",
  18040=>"110100001",
  18041=>"111100001",
  18042=>"010101011",
  18043=>"000010011",
  18044=>"101100001",
  18045=>"001010101",
  18046=>"011010010",
  18047=>"101000011",
  18048=>"011000101",
  18049=>"000011011",
  18050=>"010101011",
  18051=>"111101110",
  18052=>"101111101",
  18053=>"101101110",
  18054=>"111111000",
  18055=>"010011001",
  18056=>"001100010",
  18057=>"000001010",
  18058=>"001100111",
  18059=>"010100110",
  18060=>"111100100",
  18061=>"011111000",
  18062=>"001001001",
  18063=>"000110101",
  18064=>"111010100",
  18065=>"111010001",
  18066=>"111100001",
  18067=>"111011110",
  18068=>"011100000",
  18069=>"111010110",
  18070=>"010100111",
  18071=>"000100101",
  18072=>"010101000",
  18073=>"001000111",
  18074=>"110101100",
  18075=>"010101110",
  18076=>"110100011",
  18077=>"100100110",
  18078=>"011100111",
  18079=>"101110001",
  18080=>"110111100",
  18081=>"100010000",
  18082=>"101010101",
  18083=>"000111010",
  18084=>"001101001",
  18085=>"001101101",
  18086=>"100101000",
  18087=>"110111011",
  18088=>"011100110",
  18089=>"001000001",
  18090=>"100001111",
  18091=>"011110110",
  18092=>"101010011",
  18093=>"001001100",
  18094=>"111011011",
  18095=>"000010000",
  18096=>"101000110",
  18097=>"101010100",
  18098=>"100000011",
  18099=>"100111101",
  18100=>"100001100",
  18101=>"001111110",
  18102=>"110100000",
  18103=>"101111001",
  18104=>"010100011",
  18105=>"011010111",
  18106=>"111011111",
  18107=>"001001001",
  18108=>"111010000",
  18109=>"011011110",
  18110=>"100100101",
  18111=>"000111111",
  18112=>"111000101",
  18113=>"001100011",
  18114=>"101110101",
  18115=>"100010101",
  18116=>"010000101",
  18117=>"100011000",
  18118=>"011001001",
  18119=>"101111111",
  18120=>"001100011",
  18121=>"001011010",
  18122=>"101100111",
  18123=>"000100101",
  18124=>"100110110",
  18125=>"001100111",
  18126=>"100001101",
  18127=>"101100111",
  18128=>"011101111",
  18129=>"101011100",
  18130=>"111001111",
  18131=>"011011101",
  18132=>"111101111",
  18133=>"000100001",
  18134=>"001000010",
  18135=>"001001100",
  18136=>"101010010",
  18137=>"001010111",
  18138=>"000011000",
  18139=>"111111101",
  18140=>"001101100",
  18141=>"010101010",
  18142=>"010110010",
  18143=>"011011110",
  18144=>"110110010",
  18145=>"010010001",
  18146=>"111100100",
  18147=>"111101101",
  18148=>"000110101",
  18149=>"100110010",
  18150=>"100110110",
  18151=>"001110011",
  18152=>"001001001",
  18153=>"010101001",
  18154=>"010100100",
  18155=>"101000001",
  18156=>"011101001",
  18157=>"100011110",
  18158=>"001111001",
  18159=>"000001010",
  18160=>"100101110",
  18161=>"001110000",
  18162=>"010000000",
  18163=>"010100111",
  18164=>"001110011",
  18165=>"110111011",
  18166=>"000000110",
  18167=>"100111000",
  18168=>"011101111",
  18169=>"111111100",
  18170=>"111010111",
  18171=>"010010011",
  18172=>"010100110",
  18173=>"001001011",
  18174=>"100101110",
  18175=>"000011110",
  18176=>"101100011",
  18177=>"001111110",
  18178=>"111111010",
  18179=>"001001010",
  18180=>"111110001",
  18181=>"110001000",
  18182=>"000001011",
  18183=>"011010001",
  18184=>"000101000",
  18185=>"010100010",
  18186=>"100001100",
  18187=>"001101101",
  18188=>"111101110",
  18189=>"010100110",
  18190=>"111010111",
  18191=>"000001011",
  18192=>"010010011",
  18193=>"001100111",
  18194=>"100101101",
  18195=>"011011101",
  18196=>"000011111",
  18197=>"010001111",
  18198=>"000011000",
  18199=>"000001011",
  18200=>"111010101",
  18201=>"111100110",
  18202=>"110000101",
  18203=>"100000110",
  18204=>"000100010",
  18205=>"011000111",
  18206=>"001110000",
  18207=>"001100111",
  18208=>"100010101",
  18209=>"111001001",
  18210=>"001111100",
  18211=>"110000110",
  18212=>"010000000",
  18213=>"010111011",
  18214=>"100101101",
  18215=>"000011110",
  18216=>"100101001",
  18217=>"000100110",
  18218=>"110010100",
  18219=>"111001100",
  18220=>"101110111",
  18221=>"001110110",
  18222=>"000011000",
  18223=>"010011000",
  18224=>"101100100",
  18225=>"111100000",
  18226=>"000010101",
  18227=>"000110111",
  18228=>"101100011",
  18229=>"110111100",
  18230=>"111100110",
  18231=>"110101100",
  18232=>"000100000",
  18233=>"111000010",
  18234=>"010001110",
  18235=>"010101101",
  18236=>"000011110",
  18237=>"011101111",
  18238=>"111110000",
  18239=>"010110000",
  18240=>"100101110",
  18241=>"010001100",
  18242=>"010001100",
  18243=>"011001000",
  18244=>"001010011",
  18245=>"011110101",
  18246=>"010101101",
  18247=>"110101010",
  18248=>"111001010",
  18249=>"111101101",
  18250=>"010101011",
  18251=>"010010000",
  18252=>"000011001",
  18253=>"110011011",
  18254=>"010000010",
  18255=>"100001011",
  18256=>"010001001",
  18257=>"101101111",
  18258=>"001011000",
  18259=>"011101001",
  18260=>"100100101",
  18261=>"000000110",
  18262=>"101010010",
  18263=>"111010001",
  18264=>"111101110",
  18265=>"101100101",
  18266=>"000000011",
  18267=>"010000100",
  18268=>"111001000",
  18269=>"110111101",
  18270=>"011110011",
  18271=>"011111010",
  18272=>"001010110",
  18273=>"111100100",
  18274=>"000100100",
  18275=>"010110001",
  18276=>"101011101",
  18277=>"011100111",
  18278=>"000011001",
  18279=>"010000101",
  18280=>"000010000",
  18281=>"100001001",
  18282=>"000101000",
  18283=>"100011000",
  18284=>"001011001",
  18285=>"111111011",
  18286=>"011000110",
  18287=>"110101111",
  18288=>"011101110",
  18289=>"100000000",
  18290=>"111111100",
  18291=>"100001001",
  18292=>"111000110",
  18293=>"110001010",
  18294=>"000001100",
  18295=>"110100101",
  18296=>"111110110",
  18297=>"111010110",
  18298=>"011000110",
  18299=>"110101000",
  18300=>"011110011",
  18301=>"111000111",
  18302=>"011110101",
  18303=>"001010000",
  18304=>"010011100",
  18305=>"000111011",
  18306=>"001100111",
  18307=>"010100101",
  18308=>"010010001",
  18309=>"111111100",
  18310=>"111011001",
  18311=>"110011101",
  18312=>"110111100",
  18313=>"101111111",
  18314=>"111100100",
  18315=>"110011000",
  18316=>"001110110",
  18317=>"111001110",
  18318=>"100011100",
  18319=>"011101000",
  18320=>"110001001",
  18321=>"000010000",
  18322=>"111100001",
  18323=>"001110101",
  18324=>"001001001",
  18325=>"110001110",
  18326=>"001001000",
  18327=>"011001000",
  18328=>"111110110",
  18329=>"110110100",
  18330=>"101011100",
  18331=>"100000111",
  18332=>"111000001",
  18333=>"110000100",
  18334=>"000010110",
  18335=>"000001111",
  18336=>"110101110",
  18337=>"000000010",
  18338=>"111000011",
  18339=>"000001111",
  18340=>"101111010",
  18341=>"100110110",
  18342=>"001111101",
  18343=>"011000111",
  18344=>"010001101",
  18345=>"101011100",
  18346=>"101110011",
  18347=>"000010110",
  18348=>"101000101",
  18349=>"010111000",
  18350=>"001111001",
  18351=>"010011011",
  18352=>"110100111",
  18353=>"010000000",
  18354=>"100100011",
  18355=>"001111001",
  18356=>"000000011",
  18357=>"111110000",
  18358=>"010010010",
  18359=>"110101011",
  18360=>"111001000",
  18361=>"101100000",
  18362=>"010010100",
  18363=>"010001010",
  18364=>"111100100",
  18365=>"001101110",
  18366=>"111010100",
  18367=>"010101001",
  18368=>"111001110",
  18369=>"001000000",
  18370=>"011100100",
  18371=>"111001011",
  18372=>"011000110",
  18373=>"011001111",
  18374=>"100001110",
  18375=>"110011001",
  18376=>"000000010",
  18377=>"101110100",
  18378=>"101111101",
  18379=>"001001101",
  18380=>"110011101",
  18381=>"001111110",
  18382=>"000100100",
  18383=>"011011010",
  18384=>"111011111",
  18385=>"100111001",
  18386=>"000100110",
  18387=>"011111011",
  18388=>"010101100",
  18389=>"100110111",
  18390=>"010010001",
  18391=>"111111010",
  18392=>"100001001",
  18393=>"111001000",
  18394=>"111110000",
  18395=>"001000100",
  18396=>"101110101",
  18397=>"010111000",
  18398=>"000011011",
  18399=>"011000100",
  18400=>"001111100",
  18401=>"000111000",
  18402=>"000110110",
  18403=>"000110010",
  18404=>"011001001",
  18405=>"001010111",
  18406=>"111010110",
  18407=>"001000101",
  18408=>"011010100",
  18409=>"001100111",
  18410=>"010010111",
  18411=>"001111111",
  18412=>"011110110",
  18413=>"100101000",
  18414=>"100010111",
  18415=>"111110101",
  18416=>"100000111",
  18417=>"100011110",
  18418=>"111101010",
  18419=>"000000000",
  18420=>"000000010",
  18421=>"101001001",
  18422=>"001110010",
  18423=>"011000111",
  18424=>"011011001",
  18425=>"100110110",
  18426=>"011000001",
  18427=>"000100000",
  18428=>"010101100",
  18429=>"011011100",
  18430=>"011111010",
  18431=>"000101100",
  18432=>"000110111",
  18433=>"000101000",
  18434=>"001011100",
  18435=>"100111011",
  18436=>"000111010",
  18437=>"000100011",
  18438=>"000010011",
  18439=>"011010011",
  18440=>"110001011",
  18441=>"000011000",
  18442=>"100001001",
  18443=>"011100001",
  18444=>"100100011",
  18445=>"101010110",
  18446=>"101001100",
  18447=>"000100100",
  18448=>"100000011",
  18449=>"101000101",
  18450=>"100001100",
  18451=>"011010000",
  18452=>"000001000",
  18453=>"101001100",
  18454=>"001101010",
  18455=>"000111001",
  18456=>"010001111",
  18457=>"110110101",
  18458=>"001010111",
  18459=>"011011100",
  18460=>"001110101",
  18461=>"000001010",
  18462=>"000011001",
  18463=>"110100011",
  18464=>"110010001",
  18465=>"010100100",
  18466=>"100100110",
  18467=>"100011111",
  18468=>"001111011",
  18469=>"010000111",
  18470=>"011001011",
  18471=>"000101100",
  18472=>"011010000",
  18473=>"000101001",
  18474=>"111011111",
  18475=>"011110010",
  18476=>"011101000",
  18477=>"111111001",
  18478=>"000101001",
  18479=>"100100011",
  18480=>"110111110",
  18481=>"011101000",
  18482=>"011100000",
  18483=>"010000001",
  18484=>"010101001",
  18485=>"100001101",
  18486=>"010111110",
  18487=>"001001111",
  18488=>"011101010",
  18489=>"111110100",
  18490=>"101001101",
  18491=>"010111010",
  18492=>"010001101",
  18493=>"010010101",
  18494=>"101101011",
  18495=>"001100101",
  18496=>"000001011",
  18497=>"000000100",
  18498=>"010010101",
  18499=>"110100101",
  18500=>"110101101",
  18501=>"100011011",
  18502=>"001101101",
  18503=>"001011101",
  18504=>"011010011",
  18505=>"011110101",
  18506=>"001110100",
  18507=>"011000101",
  18508=>"001110110",
  18509=>"010111111",
  18510=>"110001000",
  18511=>"100101001",
  18512=>"111100010",
  18513=>"010011011",
  18514=>"110110001",
  18515=>"011001101",
  18516=>"110110010",
  18517=>"001001000",
  18518=>"001111110",
  18519=>"001000100",
  18520=>"110010000",
  18521=>"110101110",
  18522=>"011101001",
  18523=>"111100011",
  18524=>"010101011",
  18525=>"101111001",
  18526=>"100100011",
  18527=>"000000000",
  18528=>"100101000",
  18529=>"101000100",
  18530=>"100100001",
  18531=>"001100011",
  18532=>"101000100",
  18533=>"111010000",
  18534=>"010000011",
  18535=>"001100000",
  18536=>"100001111",
  18537=>"010000110",
  18538=>"010000011",
  18539=>"001000001",
  18540=>"000100011",
  18541=>"000111101",
  18542=>"001100100",
  18543=>"001111010",
  18544=>"011100111",
  18545=>"001110100",
  18546=>"110111111",
  18547=>"010000010",
  18548=>"001100101",
  18549=>"001101000",
  18550=>"011101011",
  18551=>"000011011",
  18552=>"001110101",
  18553=>"001110100",
  18554=>"001110011",
  18555=>"011011010",
  18556=>"010000111",
  18557=>"100000111",
  18558=>"010100111",
  18559=>"000011010",
  18560=>"001010110",
  18561=>"001100101",
  18562=>"111000001",
  18563=>"101110001",
  18564=>"110110011",
  18565=>"100001001",
  18566=>"001010101",
  18567=>"101000000",
  18568=>"001100010",
  18569=>"101011010",
  18570=>"001011100",
  18571=>"010111011",
  18572=>"011101000",
  18573=>"100010000",
  18574=>"000101110",
  18575=>"000000100",
  18576=>"111000001",
  18577=>"100110101",
  18578=>"011011100",
  18579=>"111011101",
  18580=>"100101100",
  18581=>"000101001",
  18582=>"011111011",
  18583=>"001101110",
  18584=>"110111011",
  18585=>"110100111",
  18586=>"101101101",
  18587=>"011011111",
  18588=>"010010000",
  18589=>"000100011",
  18590=>"110111100",
  18591=>"110101000",
  18592=>"001110111",
  18593=>"110011101",
  18594=>"011001001",
  18595=>"100001101",
  18596=>"000110000",
  18597=>"110100100",
  18598=>"101101100",
  18599=>"010001100",
  18600=>"010010100",
  18601=>"011111111",
  18602=>"111101001",
  18603=>"101000101",
  18604=>"100010111",
  18605=>"100011000",
  18606=>"010011111",
  18607=>"011001110",
  18608=>"101011101",
  18609=>"110110001",
  18610=>"111100001",
  18611=>"011011011",
  18612=>"111010111",
  18613=>"011111100",
  18614=>"000000111",
  18615=>"010110010",
  18616=>"011010010",
  18617=>"011011000",
  18618=>"001010100",
  18619=>"010011111",
  18620=>"011010010",
  18621=>"000011001",
  18622=>"011110001",
  18623=>"010100000",
  18624=>"010000000",
  18625=>"001111111",
  18626=>"111110000",
  18627=>"110101111",
  18628=>"010101001",
  18629=>"110010000",
  18630=>"111001001",
  18631=>"000000000",
  18632=>"011110100",
  18633=>"101010001",
  18634=>"110110011",
  18635=>"001111110",
  18636=>"100100000",
  18637=>"111110100",
  18638=>"001110111",
  18639=>"000101001",
  18640=>"000000100",
  18641=>"000011011",
  18642=>"000011110",
  18643=>"110000111",
  18644=>"101010011",
  18645=>"010101011",
  18646=>"000011100",
  18647=>"001100101",
  18648=>"111100111",
  18649=>"000101011",
  18650=>"001000001",
  18651=>"110010110",
  18652=>"000110010",
  18653=>"111010001",
  18654=>"011010100",
  18655=>"001111111",
  18656=>"110010110",
  18657=>"011110110",
  18658=>"010110001",
  18659=>"010101000",
  18660=>"001101000",
  18661=>"010001110",
  18662=>"100111100",
  18663=>"011001010",
  18664=>"111101011",
  18665=>"111111100",
  18666=>"011100000",
  18667=>"101001001",
  18668=>"110101001",
  18669=>"101011100",
  18670=>"100000010",
  18671=>"100001000",
  18672=>"010010000",
  18673=>"100100001",
  18674=>"000101111",
  18675=>"111100001",
  18676=>"101101001",
  18677=>"101110010",
  18678=>"011001101",
  18679=>"000011011",
  18680=>"000111111",
  18681=>"111000101",
  18682=>"001000010",
  18683=>"011001001",
  18684=>"111111111",
  18685=>"110010000",
  18686=>"010110011",
  18687=>"010110011",
  18688=>"111000010",
  18689=>"110001010",
  18690=>"011011111",
  18691=>"111010001",
  18692=>"011011111",
  18693=>"000111011",
  18694=>"010000101",
  18695=>"100011100",
  18696=>"011101110",
  18697=>"000111011",
  18698=>"011111111",
  18699=>"011111111",
  18700=>"010101101",
  18701=>"000000101",
  18702=>"111010000",
  18703=>"110101001",
  18704=>"111010110",
  18705=>"100110001",
  18706=>"100000111",
  18707=>"011101110",
  18708=>"100001111",
  18709=>"001011001",
  18710=>"101001001",
  18711=>"000101100",
  18712=>"000000001",
  18713=>"100101110",
  18714=>"000101011",
  18715=>"000000011",
  18716=>"011110000",
  18717=>"010000100",
  18718=>"101010110",
  18719=>"001010111",
  18720=>"010010100",
  18721=>"100011000",
  18722=>"000111010",
  18723=>"110011011",
  18724=>"010110111",
  18725=>"100010100",
  18726=>"001010101",
  18727=>"001010011",
  18728=>"001000001",
  18729=>"011010011",
  18730=>"110111111",
  18731=>"001010010",
  18732=>"000110101",
  18733=>"100111100",
  18734=>"000011010",
  18735=>"000011110",
  18736=>"000011000",
  18737=>"101001111",
  18738=>"011101001",
  18739=>"010000110",
  18740=>"011110111",
  18741=>"100011101",
  18742=>"001111000",
  18743=>"101101111",
  18744=>"000010001",
  18745=>"010110110",
  18746=>"101111110",
  18747=>"001000101",
  18748=>"100111101",
  18749=>"001111110",
  18750=>"101110101",
  18751=>"111111010",
  18752=>"011101011",
  18753=>"000110100",
  18754=>"010100100",
  18755=>"100101001",
  18756=>"111001111",
  18757=>"000011100",
  18758=>"001010000",
  18759=>"001111001",
  18760=>"111000111",
  18761=>"000100011",
  18762=>"001101111",
  18763=>"011111000",
  18764=>"111000111",
  18765=>"100100000",
  18766=>"010100110",
  18767=>"110110010",
  18768=>"100100001",
  18769=>"101111000",
  18770=>"110100100",
  18771=>"110101011",
  18772=>"001010001",
  18773=>"010000001",
  18774=>"011010000",
  18775=>"110110001",
  18776=>"100100110",
  18777=>"100010010",
  18778=>"000101111",
  18779=>"000100011",
  18780=>"011111111",
  18781=>"011101111",
  18782=>"111110100",
  18783=>"100101000",
  18784=>"010000100",
  18785=>"001010111",
  18786=>"010011110",
  18787=>"110000000",
  18788=>"011100001",
  18789=>"110110010",
  18790=>"111000001",
  18791=>"111000011",
  18792=>"000001010",
  18793=>"110111010",
  18794=>"000100111",
  18795=>"000111001",
  18796=>"111001010",
  18797=>"111100000",
  18798=>"101000101",
  18799=>"000000101",
  18800=>"001000011",
  18801=>"000110101",
  18802=>"111001110",
  18803=>"100101111",
  18804=>"010001111",
  18805=>"001001111",
  18806=>"100100111",
  18807=>"000010110",
  18808=>"000110110",
  18809=>"011100010",
  18810=>"001010011",
  18811=>"111111110",
  18812=>"000110110",
  18813=>"110101100",
  18814=>"111100110",
  18815=>"011111011",
  18816=>"000110110",
  18817=>"000000110",
  18818=>"001000000",
  18819=>"010100110",
  18820=>"110001101",
  18821=>"111100111",
  18822=>"010111001",
  18823=>"111110001",
  18824=>"110111110",
  18825=>"100001000",
  18826=>"100110010",
  18827=>"110000010",
  18828=>"001110100",
  18829=>"001101001",
  18830=>"101110000",
  18831=>"010110101",
  18832=>"101010101",
  18833=>"001000110",
  18834=>"010001111",
  18835=>"101101100",
  18836=>"111110100",
  18837=>"110101000",
  18838=>"110011001",
  18839=>"011111110",
  18840=>"100010111",
  18841=>"011111010",
  18842=>"101001001",
  18843=>"010010000",
  18844=>"111000111",
  18845=>"111111000",
  18846=>"010110111",
  18847=>"011001010",
  18848=>"100010011",
  18849=>"101000111",
  18850=>"101100111",
  18851=>"111101011",
  18852=>"011101111",
  18853=>"011100101",
  18854=>"010111010",
  18855=>"011010000",
  18856=>"000001101",
  18857=>"110000101",
  18858=>"111101000",
  18859=>"010110110",
  18860=>"010010110",
  18861=>"110110000",
  18862=>"000010100",
  18863=>"111111010",
  18864=>"100111000",
  18865=>"000000010",
  18866=>"011010100",
  18867=>"001001011",
  18868=>"011010111",
  18869=>"001010000",
  18870=>"111101011",
  18871=>"101010000",
  18872=>"111010010",
  18873=>"111101111",
  18874=>"000010100",
  18875=>"010011001",
  18876=>"100111110",
  18877=>"101111111",
  18878=>"110101111",
  18879=>"011001001",
  18880=>"010011000",
  18881=>"000100010",
  18882=>"101010010",
  18883=>"101100000",
  18884=>"111011110",
  18885=>"011000011",
  18886=>"011011100",
  18887=>"110011100",
  18888=>"000001000",
  18889=>"111101101",
  18890=>"011001110",
  18891=>"110101111",
  18892=>"010010010",
  18893=>"100000001",
  18894=>"101010100",
  18895=>"010110001",
  18896=>"001110101",
  18897=>"001101001",
  18898=>"100001101",
  18899=>"011010000",
  18900=>"000101101",
  18901=>"100100100",
  18902=>"111000000",
  18903=>"001011110",
  18904=>"000111101",
  18905=>"111001111",
  18906=>"011010111",
  18907=>"010000000",
  18908=>"101111001",
  18909=>"100000000",
  18910=>"010010001",
  18911=>"111101001",
  18912=>"100100010",
  18913=>"100100110",
  18914=>"110101100",
  18915=>"010011001",
  18916=>"011101100",
  18917=>"001001000",
  18918=>"111100001",
  18919=>"100111011",
  18920=>"010101000",
  18921=>"010110010",
  18922=>"011001010",
  18923=>"000011101",
  18924=>"011010101",
  18925=>"001110010",
  18926=>"010001101",
  18927=>"011101000",
  18928=>"111010010",
  18929=>"011011101",
  18930=>"000000010",
  18931=>"011100110",
  18932=>"011001011",
  18933=>"101100100",
  18934=>"110001100",
  18935=>"010100000",
  18936=>"101000001",
  18937=>"010111111",
  18938=>"111101011",
  18939=>"000101110",
  18940=>"100100111",
  18941=>"101100111",
  18942=>"010000111",
  18943=>"101011001",
  18944=>"000011001",
  18945=>"101101111",
  18946=>"011101111",
  18947=>"011100010",
  18948=>"101101110",
  18949=>"000010111",
  18950=>"000111000",
  18951=>"110110100",
  18952=>"011100010",
  18953=>"000100100",
  18954=>"110000001",
  18955=>"010001000",
  18956=>"101101001",
  18957=>"001001100",
  18958=>"100110100",
  18959=>"011101000",
  18960=>"101111101",
  18961=>"001100111",
  18962=>"000111000",
  18963=>"010111010",
  18964=>"001101101",
  18965=>"010100010",
  18966=>"110110001",
  18967=>"111010111",
  18968=>"001011011",
  18969=>"111111000",
  18970=>"011110111",
  18971=>"100011110",
  18972=>"001011101",
  18973=>"000111010",
  18974=>"001010000",
  18975=>"001011011",
  18976=>"101110100",
  18977=>"111011101",
  18978=>"001001100",
  18979=>"110001011",
  18980=>"111101010",
  18981=>"001000011",
  18982=>"011010000",
  18983=>"010101100",
  18984=>"111111001",
  18985=>"111001000",
  18986=>"011100110",
  18987=>"101111000",
  18988=>"111101110",
  18989=>"011101111",
  18990=>"000010010",
  18991=>"101001011",
  18992=>"011010100",
  18993=>"000101110",
  18994=>"000000101",
  18995=>"010010111",
  18996=>"011010000",
  18997=>"111010000",
  18998=>"101110010",
  18999=>"011010110",
  19000=>"001000000",
  19001=>"011111010",
  19002=>"110100101",
  19003=>"001100100",
  19004=>"010100010",
  19005=>"001101011",
  19006=>"001100110",
  19007=>"001111011",
  19008=>"100011001",
  19009=>"110110111",
  19010=>"100011011",
  19011=>"001011000",
  19012=>"101000110",
  19013=>"001000111",
  19014=>"111101101",
  19015=>"101000011",
  19016=>"000011000",
  19017=>"111000101",
  19018=>"101000000",
  19019=>"001110100",
  19020=>"110000100",
  19021=>"000001001",
  19022=>"010111001",
  19023=>"001110000",
  19024=>"001010111",
  19025=>"011010001",
  19026=>"000110000",
  19027=>"100000001",
  19028=>"001110100",
  19029=>"101111101",
  19030=>"011110100",
  19031=>"000110011",
  19032=>"011110110",
  19033=>"001111101",
  19034=>"001110100",
  19035=>"101110110",
  19036=>"000101111",
  19037=>"101001010",
  19038=>"000101110",
  19039=>"011001000",
  19040=>"011110000",
  19041=>"010000101",
  19042=>"010111111",
  19043=>"101001101",
  19044=>"001101110",
  19045=>"110000111",
  19046=>"010001100",
  19047=>"110000011",
  19048=>"111010000",
  19049=>"110001100",
  19050=>"001011010",
  19051=>"100011000",
  19052=>"001000101",
  19053=>"100001110",
  19054=>"110000010",
  19055=>"010101010",
  19056=>"111001001",
  19057=>"100000101",
  19058=>"101110001",
  19059=>"100001110",
  19060=>"001011111",
  19061=>"100111010",
  19062=>"110011011",
  19063=>"000010010",
  19064=>"001001010",
  19065=>"110101011",
  19066=>"110100111",
  19067=>"111100000",
  19068=>"010101101",
  19069=>"110001001",
  19070=>"100100110",
  19071=>"110110111",
  19072=>"111100111",
  19073=>"101100000",
  19074=>"110101001",
  19075=>"000010010",
  19076=>"000001011",
  19077=>"000010011",
  19078=>"011000010",
  19079=>"001101010",
  19080=>"010010010",
  19081=>"101111010",
  19082=>"110101001",
  19083=>"010011011",
  19084=>"101111000",
  19085=>"011000101",
  19086=>"100111111",
  19087=>"100111010",
  19088=>"111100000",
  19089=>"110101111",
  19090=>"110110000",
  19091=>"001111101",
  19092=>"010000000",
  19093=>"011010111",
  19094=>"111100001",
  19095=>"010000000",
  19096=>"011110000",
  19097=>"111111110",
  19098=>"101110110",
  19099=>"111000000",
  19100=>"010100111",
  19101=>"001111111",
  19102=>"000110011",
  19103=>"101100101",
  19104=>"010101011",
  19105=>"110001010",
  19106=>"100010111",
  19107=>"000101000",
  19108=>"111111011",
  19109=>"101011010",
  19110=>"111110100",
  19111=>"001000000",
  19112=>"100010101",
  19113=>"001101100",
  19114=>"101010000",
  19115=>"101011011",
  19116=>"011001100",
  19117=>"000010000",
  19118=>"001101001",
  19119=>"011101101",
  19120=>"000010100",
  19121=>"010011101",
  19122=>"110000000",
  19123=>"111000110",
  19124=>"111111010",
  19125=>"111101011",
  19126=>"001111100",
  19127=>"010010111",
  19128=>"111000000",
  19129=>"100110111",
  19130=>"000110100",
  19131=>"001010111",
  19132=>"101011000",
  19133=>"011010010",
  19134=>"000111010",
  19135=>"100000001",
  19136=>"000110011",
  19137=>"101110001",
  19138=>"010101111",
  19139=>"111100001",
  19140=>"111011111",
  19141=>"110101100",
  19142=>"001001111",
  19143=>"000110000",
  19144=>"001101111",
  19145=>"110100000",
  19146=>"000001111",
  19147=>"001000100",
  19148=>"010001101",
  19149=>"110000010",
  19150=>"011110110",
  19151=>"010000111",
  19152=>"101001110",
  19153=>"100111100",
  19154=>"100001010",
  19155=>"001010001",
  19156=>"100011011",
  19157=>"101000001",
  19158=>"011010011",
  19159=>"010010000",
  19160=>"011000000",
  19161=>"110111001",
  19162=>"010010100",
  19163=>"110011100",
  19164=>"001100111",
  19165=>"111000001",
  19166=>"110101000",
  19167=>"100101000",
  19168=>"111011001",
  19169=>"011100101",
  19170=>"000111110",
  19171=>"100100001",
  19172=>"010100111",
  19173=>"001111001",
  19174=>"001010100",
  19175=>"000101000",
  19176=>"011010110",
  19177=>"100100110",
  19178=>"111111000",
  19179=>"010100001",
  19180=>"101100010",
  19181=>"010001000",
  19182=>"111111001",
  19183=>"011000110",
  19184=>"010101110",
  19185=>"011011010",
  19186=>"110001100",
  19187=>"101001010",
  19188=>"001101111",
  19189=>"001101011",
  19190=>"000010011",
  19191=>"000010001",
  19192=>"011100110",
  19193=>"011111100",
  19194=>"000100111",
  19195=>"110010000",
  19196=>"000101001",
  19197=>"101000011",
  19198=>"100001010",
  19199=>"101101101",
  19200=>"100000000",
  19201=>"000000010",
  19202=>"000110110",
  19203=>"110100110",
  19204=>"001001101",
  19205=>"100011000",
  19206=>"110101111",
  19207=>"111010100",
  19208=>"010011111",
  19209=>"000101111",
  19210=>"011000101",
  19211=>"100011000",
  19212=>"010001011",
  19213=>"111111010",
  19214=>"110110111",
  19215=>"100010110",
  19216=>"010011000",
  19217=>"110100101",
  19218=>"111101110",
  19219=>"111100101",
  19220=>"100000000",
  19221=>"111100011",
  19222=>"000000010",
  19223=>"110101000",
  19224=>"010111000",
  19225=>"010011001",
  19226=>"011110111",
  19227=>"110100001",
  19228=>"001110110",
  19229=>"001001010",
  19230=>"011110001",
  19231=>"001100011",
  19232=>"100000001",
  19233=>"001110000",
  19234=>"000001110",
  19235=>"000100010",
  19236=>"110100110",
  19237=>"100001001",
  19238=>"011110100",
  19239=>"001001011",
  19240=>"000101011",
  19241=>"110101111",
  19242=>"100111101",
  19243=>"011010010",
  19244=>"011111011",
  19245=>"000011110",
  19246=>"001110110",
  19247=>"101001000",
  19248=>"100011110",
  19249=>"100011000",
  19250=>"000011001",
  19251=>"001110000",
  19252=>"101100001",
  19253=>"100010000",
  19254=>"110110010",
  19255=>"110001101",
  19256=>"100010000",
  19257=>"101010000",
  19258=>"011010010",
  19259=>"011100101",
  19260=>"001110010",
  19261=>"001101010",
  19262=>"000001000",
  19263=>"010001110",
  19264=>"111100000",
  19265=>"010110001",
  19266=>"110011010",
  19267=>"101011010",
  19268=>"000000011",
  19269=>"100101110",
  19270=>"111110011",
  19271=>"010100010",
  19272=>"000111011",
  19273=>"000000010",
  19274=>"001011010",
  19275=>"011011011",
  19276=>"111101100",
  19277=>"111100000",
  19278=>"001001001",
  19279=>"000100000",
  19280=>"000010010",
  19281=>"101110110",
  19282=>"100000101",
  19283=>"011000010",
  19284=>"001011110",
  19285=>"100101101",
  19286=>"011011111",
  19287=>"111101100",
  19288=>"001110110",
  19289=>"010110100",
  19290=>"111010010",
  19291=>"101100100",
  19292=>"011001101",
  19293=>"000010001",
  19294=>"111101100",
  19295=>"001001101",
  19296=>"001101001",
  19297=>"000000001",
  19298=>"101001110",
  19299=>"101011011",
  19300=>"011101110",
  19301=>"010111110",
  19302=>"100101010",
  19303=>"010111010",
  19304=>"001000110",
  19305=>"000000101",
  19306=>"110010010",
  19307=>"001000101",
  19308=>"000101100",
  19309=>"000110000",
  19310=>"101101111",
  19311=>"110100111",
  19312=>"001111001",
  19313=>"011010111",
  19314=>"101101111",
  19315=>"001110111",
  19316=>"110010011",
  19317=>"011010011",
  19318=>"111000000",
  19319=>"001111000",
  19320=>"000001000",
  19321=>"000111100",
  19322=>"101010011",
  19323=>"110001001",
  19324=>"000000000",
  19325=>"001100010",
  19326=>"001000100",
  19327=>"110010111",
  19328=>"011100011",
  19329=>"100111101",
  19330=>"000010000",
  19331=>"110010000",
  19332=>"011010111",
  19333=>"000000011",
  19334=>"001110000",
  19335=>"000011111",
  19336=>"110110011",
  19337=>"000001000",
  19338=>"101101101",
  19339=>"101000101",
  19340=>"000100011",
  19341=>"011101001",
  19342=>"000111111",
  19343=>"011011110",
  19344=>"000101110",
  19345=>"000111111",
  19346=>"001101001",
  19347=>"001111100",
  19348=>"010100011",
  19349=>"010110100",
  19350=>"111011100",
  19351=>"000111110",
  19352=>"001110000",
  19353=>"100110111",
  19354=>"111100011",
  19355=>"111011011",
  19356=>"011101000",
  19357=>"000100000",
  19358=>"000001000",
  19359=>"000010000",
  19360=>"111111110",
  19361=>"000110101",
  19362=>"111010000",
  19363=>"011100101",
  19364=>"000010000",
  19365=>"110001001",
  19366=>"001011111",
  19367=>"101111001",
  19368=>"110111011",
  19369=>"110001101",
  19370=>"100101111",
  19371=>"001011010",
  19372=>"111101111",
  19373=>"110010100",
  19374=>"110011110",
  19375=>"001000010",
  19376=>"011011011",
  19377=>"111101001",
  19378=>"010101111",
  19379=>"011001000",
  19380=>"110001000",
  19381=>"100010100",
  19382=>"100100000",
  19383=>"000000110",
  19384=>"101111011",
  19385=>"101011000",
  19386=>"011110001",
  19387=>"100010010",
  19388=>"010111011",
  19389=>"101010100",
  19390=>"110101101",
  19391=>"110000101",
  19392=>"011111010",
  19393=>"101100111",
  19394=>"000100000",
  19395=>"011000110",
  19396=>"000010100",
  19397=>"000101100",
  19398=>"000010110",
  19399=>"000010101",
  19400=>"000001101",
  19401=>"001000001",
  19402=>"101100101",
  19403=>"001111000",
  19404=>"010101111",
  19405=>"000100001",
  19406=>"100011100",
  19407=>"110010111",
  19408=>"011010111",
  19409=>"100100010",
  19410=>"111010010",
  19411=>"101010110",
  19412=>"001001100",
  19413=>"001001110",
  19414=>"101010101",
  19415=>"000000010",
  19416=>"100101111",
  19417=>"000000010",
  19418=>"010010101",
  19419=>"100010111",
  19420=>"001011000",
  19421=>"101110110",
  19422=>"010111110",
  19423=>"000010110",
  19424=>"110011010",
  19425=>"110110011",
  19426=>"111011001",
  19427=>"111110011",
  19428=>"111010101",
  19429=>"000011110",
  19430=>"111011000",
  19431=>"010001110",
  19432=>"101111100",
  19433=>"111011011",
  19434=>"101001010",
  19435=>"000000110",
  19436=>"010110101",
  19437=>"001101000",
  19438=>"001000010",
  19439=>"100010000",
  19440=>"110001011",
  19441=>"100011001",
  19442=>"011110111",
  19443=>"101011001",
  19444=>"100101100",
  19445=>"001000101",
  19446=>"100110110",
  19447=>"000001011",
  19448=>"011001100",
  19449=>"000000111",
  19450=>"001110110",
  19451=>"100011111",
  19452=>"110000001",
  19453=>"010001010",
  19454=>"010000000",
  19455=>"010010110",
  19456=>"010000000",
  19457=>"111101110",
  19458=>"000101110",
  19459=>"100001100",
  19460=>"001100000",
  19461=>"001000000",
  19462=>"010111101",
  19463=>"111111111",
  19464=>"100000011",
  19465=>"011110010",
  19466=>"100101001",
  19467=>"101101111",
  19468=>"110001111",
  19469=>"000111110",
  19470=>"110101010",
  19471=>"001001010",
  19472=>"001010101",
  19473=>"010000100",
  19474=>"000011010",
  19475=>"001000001",
  19476=>"001111000",
  19477=>"010101100",
  19478=>"000110010",
  19479=>"111011010",
  19480=>"101100000",
  19481=>"111010001",
  19482=>"000101001",
  19483=>"010111110",
  19484=>"100100101",
  19485=>"101000110",
  19486=>"001010111",
  19487=>"010010001",
  19488=>"100011001",
  19489=>"000111110",
  19490=>"000111101",
  19491=>"010000010",
  19492=>"110100000",
  19493=>"000101101",
  19494=>"100001010",
  19495=>"111111010",
  19496=>"010010111",
  19497=>"101011000",
  19498=>"011101001",
  19499=>"000000110",
  19500=>"000110000",
  19501=>"000011000",
  19502=>"010111000",
  19503=>"110011100",
  19504=>"011010000",
  19505=>"010010011",
  19506=>"000110110",
  19507=>"010110100",
  19508=>"100101011",
  19509=>"000000000",
  19510=>"000100000",
  19511=>"100111010",
  19512=>"001111111",
  19513=>"000000111",
  19514=>"110010000",
  19515=>"000010000",
  19516=>"001010000",
  19517=>"100100100",
  19518=>"000101110",
  19519=>"101100100",
  19520=>"111001000",
  19521=>"001000010",
  19522=>"111001001",
  19523=>"110111010",
  19524=>"001111011",
  19525=>"001001110",
  19526=>"100110110",
  19527=>"111100111",
  19528=>"110111101",
  19529=>"100111001",
  19530=>"111100101",
  19531=>"000000000",
  19532=>"100100000",
  19533=>"101100010",
  19534=>"000101000",
  19535=>"111110010",
  19536=>"110101100",
  19537=>"001001101",
  19538=>"110001100",
  19539=>"101010111",
  19540=>"111100110",
  19541=>"011111111",
  19542=>"111100100",
  19543=>"001010001",
  19544=>"000101100",
  19545=>"000011011",
  19546=>"011011010",
  19547=>"000101100",
  19548=>"001011010",
  19549=>"110000111",
  19550=>"010101110",
  19551=>"110000001",
  19552=>"100000000",
  19553=>"000110010",
  19554=>"111101011",
  19555=>"110011010",
  19556=>"000011001",
  19557=>"000011010",
  19558=>"010100011",
  19559=>"111000101",
  19560=>"001110000",
  19561=>"111101011",
  19562=>"101011101",
  19563=>"110001011",
  19564=>"110010110",
  19565=>"000010010",
  19566=>"000100010",
  19567=>"100000111",
  19568=>"100010000",
  19569=>"000001100",
  19570=>"100000011",
  19571=>"010111110",
  19572=>"011101110",
  19573=>"011000011",
  19574=>"111110011",
  19575=>"000110000",
  19576=>"010101110",
  19577=>"010011111",
  19578=>"011000001",
  19579=>"100011100",
  19580=>"011101101",
  19581=>"111000000",
  19582=>"011111100",
  19583=>"101011111",
  19584=>"001001111",
  19585=>"101011110",
  19586=>"011000101",
  19587=>"000011111",
  19588=>"000111100",
  19589=>"110001100",
  19590=>"101101000",
  19591=>"000001001",
  19592=>"001111001",
  19593=>"111001100",
  19594=>"101001110",
  19595=>"101010100",
  19596=>"010110111",
  19597=>"101110101",
  19598=>"110100101",
  19599=>"010111101",
  19600=>"111001101",
  19601=>"111100100",
  19602=>"110000001",
  19603=>"001010111",
  19604=>"100000000",
  19605=>"110000110",
  19606=>"001100111",
  19607=>"010010101",
  19608=>"111101101",
  19609=>"001101110",
  19610=>"100010101",
  19611=>"000101010",
  19612=>"111111101",
  19613=>"011001101",
  19614=>"111010101",
  19615=>"010011010",
  19616=>"010011100",
  19617=>"011100101",
  19618=>"110000110",
  19619=>"001101100",
  19620=>"111101001",
  19621=>"100000100",
  19622=>"100100111",
  19623=>"011001100",
  19624=>"010001011",
  19625=>"110010001",
  19626=>"000110110",
  19627=>"111100111",
  19628=>"111000101",
  19629=>"110000101",
  19630=>"111010000",
  19631=>"011011000",
  19632=>"001001011",
  19633=>"110010011",
  19634=>"000010010",
  19635=>"111001000",
  19636=>"111100101",
  19637=>"101011100",
  19638=>"000000000",
  19639=>"110011101",
  19640=>"010000000",
  19641=>"111001111",
  19642=>"100001001",
  19643=>"011111100",
  19644=>"100110000",
  19645=>"111100011",
  19646=>"100101100",
  19647=>"001111001",
  19648=>"001101101",
  19649=>"001000111",
  19650=>"001001110",
  19651=>"001000001",
  19652=>"111111110",
  19653=>"111001101",
  19654=>"100011000",
  19655=>"011010111",
  19656=>"101110100",
  19657=>"001101001",
  19658=>"111000100",
  19659=>"001000010",
  19660=>"000010110",
  19661=>"001001001",
  19662=>"100000100",
  19663=>"000011011",
  19664=>"110001001",
  19665=>"110000001",
  19666=>"100010000",
  19667=>"010010110",
  19668=>"011000011",
  19669=>"100000001",
  19670=>"111000000",
  19671=>"111101110",
  19672=>"011100110",
  19673=>"011011111",
  19674=>"000010011",
  19675=>"000110100",
  19676=>"100010001",
  19677=>"111100010",
  19678=>"000001011",
  19679=>"111110010",
  19680=>"000000110",
  19681=>"000111100",
  19682=>"100001100",
  19683=>"000011011",
  19684=>"000101001",
  19685=>"101110010",
  19686=>"110001000",
  19687=>"111000111",
  19688=>"011111011",
  19689=>"110110010",
  19690=>"011000011",
  19691=>"010000010",
  19692=>"011100000",
  19693=>"011011000",
  19694=>"001001101",
  19695=>"010000000",
  19696=>"101100111",
  19697=>"010000011",
  19698=>"101001110",
  19699=>"110010111",
  19700=>"001111100",
  19701=>"001010001",
  19702=>"111111100",
  19703=>"011010011",
  19704=>"011100101",
  19705=>"000010101",
  19706=>"000001101",
  19707=>"001111111",
  19708=>"011010001",
  19709=>"011011010",
  19710=>"000011111",
  19711=>"100000010",
  19712=>"010101111",
  19713=>"110101100",
  19714=>"001110001",
  19715=>"100100100",
  19716=>"111011000",
  19717=>"011001001",
  19718=>"111101010",
  19719=>"010010011",
  19720=>"110010100",
  19721=>"111010111",
  19722=>"110010101",
  19723=>"110100000",
  19724=>"011101000",
  19725=>"101100110",
  19726=>"000100110",
  19727=>"011001100",
  19728=>"010111100",
  19729=>"101101000",
  19730=>"001101101",
  19731=>"101111000",
  19732=>"110010111",
  19733=>"111101111",
  19734=>"010000000",
  19735=>"001101100",
  19736=>"001110010",
  19737=>"010000001",
  19738=>"000011101",
  19739=>"000110000",
  19740=>"000101001",
  19741=>"100011110",
  19742=>"111100111",
  19743=>"000000011",
  19744=>"011000000",
  19745=>"100011000",
  19746=>"011010101",
  19747=>"111101001",
  19748=>"110011010",
  19749=>"010000000",
  19750=>"011010010",
  19751=>"001100001",
  19752=>"111111111",
  19753=>"010010110",
  19754=>"001100000",
  19755=>"111100011",
  19756=>"011011100",
  19757=>"100000010",
  19758=>"000101110",
  19759=>"000000101",
  19760=>"001011000",
  19761=>"100110000",
  19762=>"000000111",
  19763=>"000100100",
  19764=>"110011010",
  19765=>"110111101",
  19766=>"110011011",
  19767=>"111100111",
  19768=>"011111111",
  19769=>"011011111",
  19770=>"010000101",
  19771=>"000000001",
  19772=>"100001111",
  19773=>"111100000",
  19774=>"011101100",
  19775=>"111100001",
  19776=>"001100100",
  19777=>"101001011",
  19778=>"010111000",
  19779=>"010011010",
  19780=>"000100101",
  19781=>"111100101",
  19782=>"100000110",
  19783=>"001000000",
  19784=>"000010101",
  19785=>"001000101",
  19786=>"110101100",
  19787=>"000111010",
  19788=>"010110000",
  19789=>"111111001",
  19790=>"101100101",
  19791=>"001011001",
  19792=>"001000011",
  19793=>"111000001",
  19794=>"010001000",
  19795=>"010110010",
  19796=>"001010001",
  19797=>"000000100",
  19798=>"011111110",
  19799=>"010000010",
  19800=>"000011111",
  19801=>"110000000",
  19802=>"101001000",
  19803=>"100110100",
  19804=>"100001111",
  19805=>"111011100",
  19806=>"000001111",
  19807=>"111101111",
  19808=>"110111111",
  19809=>"001010100",
  19810=>"010011100",
  19811=>"001110101",
  19812=>"110110101",
  19813=>"111100111",
  19814=>"000110110",
  19815=>"000100100",
  19816=>"100011010",
  19817=>"000001101",
  19818=>"100011100",
  19819=>"000011011",
  19820=>"011010000",
  19821=>"000010101",
  19822=>"111101111",
  19823=>"101001010",
  19824=>"101000101",
  19825=>"011111001",
  19826=>"010111100",
  19827=>"000110000",
  19828=>"001001000",
  19829=>"000010011",
  19830=>"000111000",
  19831=>"101001111",
  19832=>"011111011",
  19833=>"000000111",
  19834=>"001010100",
  19835=>"010110001",
  19836=>"101011110",
  19837=>"101101111",
  19838=>"101001100",
  19839=>"001100111",
  19840=>"101100111",
  19841=>"100000011",
  19842=>"011010110",
  19843=>"101101000",
  19844=>"011100111",
  19845=>"000100101",
  19846=>"110111101",
  19847=>"101101101",
  19848=>"101000100",
  19849=>"100010110",
  19850=>"011001010",
  19851=>"101101010",
  19852=>"100011101",
  19853=>"001100010",
  19854=>"000001111",
  19855=>"000101011",
  19856=>"011101010",
  19857=>"111000111",
  19858=>"001000011",
  19859=>"101000010",
  19860=>"001011011",
  19861=>"100101011",
  19862=>"010010001",
  19863=>"001101001",
  19864=>"111101111",
  19865=>"100000111",
  19866=>"111010101",
  19867=>"111000010",
  19868=>"000001100",
  19869=>"101111100",
  19870=>"101101010",
  19871=>"110011101",
  19872=>"100101011",
  19873=>"101010000",
  19874=>"110011010",
  19875=>"101110110",
  19876=>"111011111",
  19877=>"000100101",
  19878=>"110011001",
  19879=>"001010000",
  19880=>"010100010",
  19881=>"011010001",
  19882=>"100000110",
  19883=>"011010010",
  19884=>"100010110",
  19885=>"010000011",
  19886=>"100010000",
  19887=>"011111010",
  19888=>"110011000",
  19889=>"101101101",
  19890=>"111111101",
  19891=>"101011100",
  19892=>"100101001",
  19893=>"000101100",
  19894=>"111011111",
  19895=>"011100010",
  19896=>"001001000",
  19897=>"110011111",
  19898=>"110000010",
  19899=>"010010011",
  19900=>"001001000",
  19901=>"000111010",
  19902=>"000110101",
  19903=>"111011011",
  19904=>"100000000",
  19905=>"000000001",
  19906=>"100111110",
  19907=>"010010001",
  19908=>"100111110",
  19909=>"010010010",
  19910=>"001011100",
  19911=>"100000000",
  19912=>"001111111",
  19913=>"001001011",
  19914=>"101000010",
  19915=>"000010001",
  19916=>"111101100",
  19917=>"111111101",
  19918=>"000111100",
  19919=>"100100010",
  19920=>"011011000",
  19921=>"110001110",
  19922=>"000001101",
  19923=>"100110101",
  19924=>"001001111",
  19925=>"000001110",
  19926=>"000010000",
  19927=>"100000011",
  19928=>"000000111",
  19929=>"000000010",
  19930=>"101000011",
  19931=>"100101111",
  19932=>"000111100",
  19933=>"111111111",
  19934=>"110011001",
  19935=>"100101110",
  19936=>"111111001",
  19937=>"001111011",
  19938=>"101111001",
  19939=>"101010110",
  19940=>"010111011",
  19941=>"111101101",
  19942=>"101100000",
  19943=>"101101001",
  19944=>"110001101",
  19945=>"111000100",
  19946=>"000001010",
  19947=>"111011101",
  19948=>"001001011",
  19949=>"010110111",
  19950=>"100000100",
  19951=>"101001110",
  19952=>"000011111",
  19953=>"101010011",
  19954=>"010101000",
  19955=>"000110111",
  19956=>"000110100",
  19957=>"000110010",
  19958=>"101101110",
  19959=>"000100010",
  19960=>"101111111",
  19961=>"111000100",
  19962=>"010110010",
  19963=>"000001110",
  19964=>"100101100",
  19965=>"110010000",
  19966=>"001010110",
  19967=>"110111011",
  19968=>"101101100",
  19969=>"001001011",
  19970=>"001110010",
  19971=>"111110110",
  19972=>"010011111",
  19973=>"100010110",
  19974=>"010100001",
  19975=>"110111100",
  19976=>"011010110",
  19977=>"110000011",
  19978=>"000010100",
  19979=>"000100111",
  19980=>"001001001",
  19981=>"111011100",
  19982=>"110010001",
  19983=>"100000011",
  19984=>"011000100",
  19985=>"110011111",
  19986=>"001010100",
  19987=>"011101100",
  19988=>"000010111",
  19989=>"111111001",
  19990=>"011011011",
  19991=>"001010100",
  19992=>"111111111",
  19993=>"001011110",
  19994=>"101000010",
  19995=>"010010011",
  19996=>"100010000",
  19997=>"001100101",
  19998=>"001010001",
  19999=>"001001110",
  20000=>"111100100",
  20001=>"111100001",
  20002=>"111100011",
  20003=>"110011110",
  20004=>"000000000",
  20005=>"001001011",
  20006=>"010011011",
  20007=>"110011000",
  20008=>"000111001",
  20009=>"011101100",
  20010=>"111101100",
  20011=>"000011111",
  20012=>"101101011",
  20013=>"111110100",
  20014=>"011000110",
  20015=>"011100010",
  20016=>"001110110",
  20017=>"100011110",
  20018=>"101011100",
  20019=>"000010111",
  20020=>"001010111",
  20021=>"010000001",
  20022=>"100011011",
  20023=>"010010111",
  20024=>"110000101",
  20025=>"110011010",
  20026=>"011101100",
  20027=>"101101010",
  20028=>"010000001",
  20029=>"111001101",
  20030=>"010110001",
  20031=>"110100000",
  20032=>"000010011",
  20033=>"111001010",
  20034=>"111101111",
  20035=>"010011110",
  20036=>"011011101",
  20037=>"011110100",
  20038=>"010101000",
  20039=>"100010011",
  20040=>"101011100",
  20041=>"010010010",
  20042=>"010110111",
  20043=>"100010001",
  20044=>"100001011",
  20045=>"111100010",
  20046=>"000000110",
  20047=>"111111110",
  20048=>"101111000",
  20049=>"101011001",
  20050=>"000100001",
  20051=>"001110000",
  20052=>"011110111",
  20053=>"010000111",
  20054=>"000000111",
  20055=>"101110001",
  20056=>"110110111",
  20057=>"011011011",
  20058=>"001001010",
  20059=>"101010000",
  20060=>"000100100",
  20061=>"000111010",
  20062=>"000010011",
  20063=>"111010011",
  20064=>"110111001",
  20065=>"010001011",
  20066=>"111000110",
  20067=>"011111100",
  20068=>"101010110",
  20069=>"000111100",
  20070=>"000101001",
  20071=>"101011100",
  20072=>"010100100",
  20073=>"110000010",
  20074=>"011110100",
  20075=>"000000000",
  20076=>"001100100",
  20077=>"011101011",
  20078=>"001111000",
  20079=>"001110010",
  20080=>"111010100",
  20081=>"110111011",
  20082=>"011101101",
  20083=>"110001101",
  20084=>"010001111",
  20085=>"000000100",
  20086=>"100010111",
  20087=>"111110100",
  20088=>"010111010",
  20089=>"011001110",
  20090=>"111110010",
  20091=>"000000001",
  20092=>"100100111",
  20093=>"011111101",
  20094=>"100010011",
  20095=>"001110111",
  20096=>"000000001",
  20097=>"101111101",
  20098=>"001110101",
  20099=>"011000000",
  20100=>"001101011",
  20101=>"011010011",
  20102=>"011011101",
  20103=>"001010000",
  20104=>"010000010",
  20105=>"111101010",
  20106=>"101101111",
  20107=>"100010101",
  20108=>"010000100",
  20109=>"001001100",
  20110=>"110010000",
  20111=>"110000100",
  20112=>"001000011",
  20113=>"001000111",
  20114=>"100111101",
  20115=>"000110101",
  20116=>"000101101",
  20117=>"010000000",
  20118=>"011100000",
  20119=>"000101101",
  20120=>"110011110",
  20121=>"110010111",
  20122=>"111001111",
  20123=>"110101011",
  20124=>"010011111",
  20125=>"110010000",
  20126=>"100110110",
  20127=>"110000011",
  20128=>"001101000",
  20129=>"011101001",
  20130=>"100010101",
  20131=>"100110011",
  20132=>"010101100",
  20133=>"110000000",
  20134=>"101011011",
  20135=>"000000000",
  20136=>"001011101",
  20137=>"110001101",
  20138=>"110101110",
  20139=>"000100000",
  20140=>"001000101",
  20141=>"100011101",
  20142=>"101001111",
  20143=>"101011111",
  20144=>"011111101",
  20145=>"001001001",
  20146=>"111110111",
  20147=>"000101001",
  20148=>"010101111",
  20149=>"010010001",
  20150=>"001001100",
  20151=>"100110110",
  20152=>"101101010",
  20153=>"011000111",
  20154=>"000001011",
  20155=>"111001000",
  20156=>"001101010",
  20157=>"101110100",
  20158=>"100001101",
  20159=>"011111110",
  20160=>"001001011",
  20161=>"011110101",
  20162=>"100011101",
  20163=>"011000111",
  20164=>"101111100",
  20165=>"001111100",
  20166=>"111001011",
  20167=>"101000000",
  20168=>"111011101",
  20169=>"011101111",
  20170=>"010001010",
  20171=>"110101110",
  20172=>"010100101",
  20173=>"010010000",
  20174=>"010110111",
  20175=>"101111001",
  20176=>"011100000",
  20177=>"011110100",
  20178=>"101111010",
  20179=>"111110011",
  20180=>"101100000",
  20181=>"111110110",
  20182=>"011010000",
  20183=>"110110101",
  20184=>"100000001",
  20185=>"010100011",
  20186=>"110101010",
  20187=>"000001011",
  20188=>"001000101",
  20189=>"111100001",
  20190=>"111000111",
  20191=>"110100010",
  20192=>"000000111",
  20193=>"010011100",
  20194=>"011101001",
  20195=>"111111011",
  20196=>"011001111",
  20197=>"000000100",
  20198=>"000011110",
  20199=>"110001000",
  20200=>"100010110",
  20201=>"010001110",
  20202=>"001111101",
  20203=>"000111011",
  20204=>"000010111",
  20205=>"001110100",
  20206=>"010110001",
  20207=>"001100010",
  20208=>"010000111",
  20209=>"001011000",
  20210=>"000010000",
  20211=>"110001000",
  20212=>"111110111",
  20213=>"101110001",
  20214=>"100110101",
  20215=>"110111000",
  20216=>"100111001",
  20217=>"100110000",
  20218=>"100110001",
  20219=>"000110010",
  20220=>"001111110",
  20221=>"011111011",
  20222=>"011010001",
  20223=>"100011010",
  20224=>"100001011",
  20225=>"010101101",
  20226=>"111110000",
  20227=>"101001111",
  20228=>"010010001",
  20229=>"000010000",
  20230=>"110100111",
  20231=>"001011111",
  20232=>"000100011",
  20233=>"000011000",
  20234=>"100000000",
  20235=>"100000001",
  20236=>"111011010",
  20237=>"000110111",
  20238=>"000011100",
  20239=>"011100111",
  20240=>"001011101",
  20241=>"111001101",
  20242=>"101100000",
  20243=>"110110001",
  20244=>"010000110",
  20245=>"110001001",
  20246=>"111000000",
  20247=>"110011101",
  20248=>"111100101",
  20249=>"000101100",
  20250=>"011100000",
  20251=>"010010011",
  20252=>"010001011",
  20253=>"000111100",
  20254=>"100000001",
  20255=>"000000000",
  20256=>"010101101",
  20257=>"110111011",
  20258=>"000111001",
  20259=>"011111111",
  20260=>"111001001",
  20261=>"000110001",
  20262=>"000111001",
  20263=>"101111011",
  20264=>"000001110",
  20265=>"101100101",
  20266=>"001101011",
  20267=>"100100010",
  20268=>"000101011",
  20269=>"011100000",
  20270=>"100001111",
  20271=>"010101001",
  20272=>"111000001",
  20273=>"111001011",
  20274=>"101101010",
  20275=>"100110100",
  20276=>"000010000",
  20277=>"001100111",
  20278=>"000000100",
  20279=>"110011101",
  20280=>"111110010",
  20281=>"000011101",
  20282=>"011011101",
  20283=>"000011001",
  20284=>"010110000",
  20285=>"001001000",
  20286=>"001111101",
  20287=>"111101000",
  20288=>"000100111",
  20289=>"100000010",
  20290=>"110111100",
  20291=>"000101101",
  20292=>"011000110",
  20293=>"111110001",
  20294=>"010001100",
  20295=>"111000011",
  20296=>"001001101",
  20297=>"011111010",
  20298=>"000010000",
  20299=>"001100100",
  20300=>"010100110",
  20301=>"111100101",
  20302=>"001000000",
  20303=>"011101001",
  20304=>"100110010",
  20305=>"001001110",
  20306=>"111000111",
  20307=>"000110101",
  20308=>"010100001",
  20309=>"000000110",
  20310=>"000010011",
  20311=>"010011101",
  20312=>"010111011",
  20313=>"011110010",
  20314=>"001011001",
  20315=>"000100010",
  20316=>"111001000",
  20317=>"010110100",
  20318=>"000100100",
  20319=>"111000101",
  20320=>"100001111",
  20321=>"001100101",
  20322=>"000111100",
  20323=>"011100101",
  20324=>"011111000",
  20325=>"010001011",
  20326=>"011111010",
  20327=>"011000000",
  20328=>"010010111",
  20329=>"110001011",
  20330=>"111001110",
  20331=>"011001000",
  20332=>"101011001",
  20333=>"001011101",
  20334=>"110110001",
  20335=>"111110110",
  20336=>"000010100",
  20337=>"001011110",
  20338=>"010110111",
  20339=>"111011001",
  20340=>"111101001",
  20341=>"110110001",
  20342=>"001100100",
  20343=>"000010110",
  20344=>"110010111",
  20345=>"110101001",
  20346=>"110110110",
  20347=>"111111001",
  20348=>"011001101",
  20349=>"011000010",
  20350=>"110101101",
  20351=>"111000001",
  20352=>"100100110",
  20353=>"100110011",
  20354=>"011111111",
  20355=>"111011110",
  20356=>"100101000",
  20357=>"000101100",
  20358=>"111011001",
  20359=>"111000100",
  20360=>"011100101",
  20361=>"000101000",
  20362=>"111111100",
  20363=>"111001010",
  20364=>"010011000",
  20365=>"001100110",
  20366=>"110000100",
  20367=>"000010101",
  20368=>"001001001",
  20369=>"101110101",
  20370=>"010101110",
  20371=>"000011100",
  20372=>"001011000",
  20373=>"101001011",
  20374=>"111010100",
  20375=>"110000100",
  20376=>"001101111",
  20377=>"111100110",
  20378=>"010101110",
  20379=>"110111110",
  20380=>"000000101",
  20381=>"100110011",
  20382=>"100011111",
  20383=>"000000101",
  20384=>"111010100",
  20385=>"100001101",
  20386=>"110100001",
  20387=>"110110101",
  20388=>"110001000",
  20389=>"101010010",
  20390=>"111011101",
  20391=>"111010111",
  20392=>"000100000",
  20393=>"101000000",
  20394=>"101110101",
  20395=>"001010000",
  20396=>"110011011",
  20397=>"000101100",
  20398=>"111111101",
  20399=>"100111000",
  20400=>"010110010",
  20401=>"001100101",
  20402=>"010000000",
  20403=>"111111110",
  20404=>"100001111",
  20405=>"000011011",
  20406=>"100101101",
  20407=>"100010111",
  20408=>"010011000",
  20409=>"100110011",
  20410=>"100000000",
  20411=>"010111001",
  20412=>"101010111",
  20413=>"010100010",
  20414=>"000010000",
  20415=>"000110110",
  20416=>"110110101",
  20417=>"110111110",
  20418=>"100001001",
  20419=>"001100111",
  20420=>"101010111",
  20421=>"101101010",
  20422=>"010011101",
  20423=>"100100010",
  20424=>"000010011",
  20425=>"110000111",
  20426=>"011010000",
  20427=>"001100011",
  20428=>"101000111",
  20429=>"000001010",
  20430=>"010001001",
  20431=>"101100111",
  20432=>"000001010",
  20433=>"111111001",
  20434=>"000010111",
  20435=>"110011001",
  20436=>"000010111",
  20437=>"001000010",
  20438=>"101000101",
  20439=>"101000001",
  20440=>"011111100",
  20441=>"101000110",
  20442=>"111101111",
  20443=>"111101010",
  20444=>"111010110",
  20445=>"100010111",
  20446=>"101011011",
  20447=>"110010111",
  20448=>"010011110",
  20449=>"101001001",
  20450=>"000110000",
  20451=>"001101000",
  20452=>"000101111",
  20453=>"111101001",
  20454=>"001110110",
  20455=>"011100111",
  20456=>"111101110",
  20457=>"010101111",
  20458=>"000100100",
  20459=>"100011011",
  20460=>"000100110",
  20461=>"111010110",
  20462=>"101001010",
  20463=>"100110011",
  20464=>"100001001",
  20465=>"101010011",
  20466=>"000001110",
  20467=>"101000111",
  20468=>"111100111",
  20469=>"111011001",
  20470=>"111110101",
  20471=>"101101111",
  20472=>"100100000",
  20473=>"000110110",
  20474=>"110100100",
  20475=>"010111001",
  20476=>"010110010",
  20477=>"100000000",
  20478=>"100000001",
  20479=>"000010001",
  20480=>"111010011",
  20481=>"011110110",
  20482=>"101100101",
  20483=>"010000101",
  20484=>"010110101",
  20485=>"111000101",
  20486=>"100101101",
  20487=>"000100000",
  20488=>"000010101",
  20489=>"101110110",
  20490=>"000010000",
  20491=>"101011011",
  20492=>"001001011",
  20493=>"010010101",
  20494=>"000111100",
  20495=>"000101101",
  20496=>"111101111",
  20497=>"111111111",
  20498=>"001110110",
  20499=>"001011001",
  20500=>"100000011",
  20501=>"111110101",
  20502=>"110000110",
  20503=>"011011010",
  20504=>"110111010",
  20505=>"000110011",
  20506=>"010100001",
  20507=>"011101000",
  20508=>"011000101",
  20509=>"101111101",
  20510=>"001110000",
  20511=>"011111101",
  20512=>"011011001",
  20513=>"101000100",
  20514=>"011011000",
  20515=>"110100001",
  20516=>"010100111",
  20517=>"100001110",
  20518=>"110011100",
  20519=>"110100110",
  20520=>"011001000",
  20521=>"101001000",
  20522=>"011010100",
  20523=>"110001100",
  20524=>"101001001",
  20525=>"110100001",
  20526=>"000110110",
  20527=>"111100100",
  20528=>"111011101",
  20529=>"100100100",
  20530=>"110011100",
  20531=>"101011000",
  20532=>"110111101",
  20533=>"001011000",
  20534=>"011111011",
  20535=>"010010100",
  20536=>"100100000",
  20537=>"011110011",
  20538=>"101001110",
  20539=>"011001100",
  20540=>"111100101",
  20541=>"010101110",
  20542=>"101010011",
  20543=>"000010100",
  20544=>"101000110",
  20545=>"001000010",
  20546=>"111110110",
  20547=>"110000110",
  20548=>"110001110",
  20549=>"001110000",
  20550=>"100101100",
  20551=>"010111011",
  20552=>"110010111",
  20553=>"101110010",
  20554=>"010011101",
  20555=>"000000110",
  20556=>"001010010",
  20557=>"011011100",
  20558=>"111000101",
  20559=>"110101010",
  20560=>"100011001",
  20561=>"110111111",
  20562=>"010000100",
  20563=>"001100111",
  20564=>"110100101",
  20565=>"101110111",
  20566=>"101100111",
  20567=>"110110111",
  20568=>"110110001",
  20569=>"110010011",
  20570=>"101000100",
  20571=>"010010001",
  20572=>"100011101",
  20573=>"000101010",
  20574=>"010010011",
  20575=>"100100000",
  20576=>"011111011",
  20577=>"100100001",
  20578=>"001001011",
  20579=>"101000110",
  20580=>"110011110",
  20581=>"111101110",
  20582=>"101000010",
  20583=>"101110000",
  20584=>"101001110",
  20585=>"111100111",
  20586=>"111100101",
  20587=>"010000010",
  20588=>"110111110",
  20589=>"000000101",
  20590=>"100101101",
  20591=>"000001001",
  20592=>"000111111",
  20593=>"100100111",
  20594=>"111010000",
  20595=>"010100111",
  20596=>"000001101",
  20597=>"111111000",
  20598=>"010100010",
  20599=>"111100011",
  20600=>"101101110",
  20601=>"010001101",
  20602=>"101000111",
  20603=>"010010010",
  20604=>"000100111",
  20605=>"001000110",
  20606=>"001011010",
  20607=>"111110111",
  20608=>"110001000",
  20609=>"001010011",
  20610=>"101110100",
  20611=>"001111000",
  20612=>"011010001",
  20613=>"101111011",
  20614=>"110010110",
  20615=>"111100110",
  20616=>"110101001",
  20617=>"101110100",
  20618=>"111011111",
  20619=>"001111111",
  20620=>"011000101",
  20621=>"110010101",
  20622=>"110110000",
  20623=>"101111010",
  20624=>"100100100",
  20625=>"110000100",
  20626=>"110001010",
  20627=>"100100010",
  20628=>"100000011",
  20629=>"001010111",
  20630=>"101110010",
  20631=>"000011011",
  20632=>"000001001",
  20633=>"111111001",
  20634=>"010100100",
  20635=>"110110101",
  20636=>"000001010",
  20637=>"001111110",
  20638=>"011001001",
  20639=>"100011001",
  20640=>"001110100",
  20641=>"101100000",
  20642=>"111000000",
  20643=>"111101111",
  20644=>"010000100",
  20645=>"111010010",
  20646=>"001000100",
  20647=>"110000000",
  20648=>"110011001",
  20649=>"000111111",
  20650=>"010010000",
  20651=>"010000101",
  20652=>"110010111",
  20653=>"001011000",
  20654=>"100101110",
  20655=>"111100100",
  20656=>"011010001",
  20657=>"110010001",
  20658=>"001000110",
  20659=>"111100100",
  20660=>"010101101",
  20661=>"010010101",
  20662=>"101011111",
  20663=>"110010011",
  20664=>"010001101",
  20665=>"010000111",
  20666=>"001100000",
  20667=>"011001011",
  20668=>"001010011",
  20669=>"001010001",
  20670=>"110100110",
  20671=>"100000011",
  20672=>"111101010",
  20673=>"011101001",
  20674=>"000110111",
  20675=>"100110011",
  20676=>"100000000",
  20677=>"100101010",
  20678=>"000000101",
  20679=>"101001110",
  20680=>"110011111",
  20681=>"011100001",
  20682=>"001000111",
  20683=>"110110010",
  20684=>"111101101",
  20685=>"101110111",
  20686=>"011110101",
  20687=>"101011100",
  20688=>"110011010",
  20689=>"010111000",
  20690=>"101101101",
  20691=>"000010110",
  20692=>"011001100",
  20693=>"101101111",
  20694=>"011011001",
  20695=>"000000000",
  20696=>"010001000",
  20697=>"111101000",
  20698=>"011011000",
  20699=>"110110000",
  20700=>"101001011",
  20701=>"100101110",
  20702=>"101100000",
  20703=>"001101100",
  20704=>"001011010",
  20705=>"100010110",
  20706=>"000010100",
  20707=>"111100101",
  20708=>"101101001",
  20709=>"011011101",
  20710=>"001011011",
  20711=>"001010110",
  20712=>"100110100",
  20713=>"100001110",
  20714=>"000010010",
  20715=>"010110110",
  20716=>"001011111",
  20717=>"110001010",
  20718=>"110000110",
  20719=>"111111000",
  20720=>"111110011",
  20721=>"100001000",
  20722=>"011111011",
  20723=>"001100011",
  20724=>"111011010",
  20725=>"000010010",
  20726=>"110010010",
  20727=>"000011111",
  20728=>"100101000",
  20729=>"100001011",
  20730=>"011101110",
  20731=>"110000000",
  20732=>"011011010",
  20733=>"011001110",
  20734=>"111101011",
  20735=>"100101111",
  20736=>"000010001",
  20737=>"011100001",
  20738=>"110100101",
  20739=>"110001111",
  20740=>"001111000",
  20741=>"111011001",
  20742=>"101000011",
  20743=>"111101001",
  20744=>"010101111",
  20745=>"000000111",
  20746=>"111011001",
  20747=>"000100101",
  20748=>"110001100",
  20749=>"000111101",
  20750=>"000100011",
  20751=>"110000110",
  20752=>"100000000",
  20753=>"100100101",
  20754=>"011000011",
  20755=>"111111110",
  20756=>"011011001",
  20757=>"100011100",
  20758=>"000111000",
  20759=>"100100001",
  20760=>"010011000",
  20761=>"101101001",
  20762=>"101001100",
  20763=>"110110110",
  20764=>"110010111",
  20765=>"111010000",
  20766=>"011010100",
  20767=>"110100001",
  20768=>"001010010",
  20769=>"010100001",
  20770=>"111011010",
  20771=>"010100101",
  20772=>"001011101",
  20773=>"110111011",
  20774=>"110110010",
  20775=>"010011011",
  20776=>"010100011",
  20777=>"101010110",
  20778=>"110001101",
  20779=>"101000000",
  20780=>"000000100",
  20781=>"011111011",
  20782=>"011101001",
  20783=>"010011010",
  20784=>"100111101",
  20785=>"011100100",
  20786=>"000101110",
  20787=>"100101111",
  20788=>"100011110",
  20789=>"100100011",
  20790=>"111000100",
  20791=>"011010000",
  20792=>"110111010",
  20793=>"100110001",
  20794=>"011101101",
  20795=>"010011101",
  20796=>"000110000",
  20797=>"011001001",
  20798=>"010101000",
  20799=>"110001011",
  20800=>"110111110",
  20801=>"011001011",
  20802=>"011111010",
  20803=>"111011010",
  20804=>"001101011",
  20805=>"111001010",
  20806=>"011011010",
  20807=>"000100101",
  20808=>"000010101",
  20809=>"010010011",
  20810=>"011110111",
  20811=>"001100001",
  20812=>"110011100",
  20813=>"100110111",
  20814=>"100100001",
  20815=>"011000001",
  20816=>"111011010",
  20817=>"111001110",
  20818=>"001000111",
  20819=>"111011111",
  20820=>"100011101",
  20821=>"111011110",
  20822=>"011101110",
  20823=>"100101000",
  20824=>"100101001",
  20825=>"101101100",
  20826=>"001100010",
  20827=>"111111001",
  20828=>"010110001",
  20829=>"100010100",
  20830=>"000010011",
  20831=>"011010000",
  20832=>"111011010",
  20833=>"010110000",
  20834=>"001100100",
  20835=>"001010101",
  20836=>"100110011",
  20837=>"111111110",
  20838=>"100011111",
  20839=>"011001101",
  20840=>"100110010",
  20841=>"111100111",
  20842=>"001011100",
  20843=>"100011111",
  20844=>"101110101",
  20845=>"101111111",
  20846=>"001101001",
  20847=>"101011111",
  20848=>"001001100",
  20849=>"000000101",
  20850=>"100110001",
  20851=>"001110011",
  20852=>"001111110",
  20853=>"111011001",
  20854=>"010010000",
  20855=>"011010111",
  20856=>"111000001",
  20857=>"110111000",
  20858=>"101100111",
  20859=>"100101111",
  20860=>"011010010",
  20861=>"010000001",
  20862=>"110011000",
  20863=>"011101101",
  20864=>"000000001",
  20865=>"100000101",
  20866=>"111111111",
  20867=>"000001000",
  20868=>"110001111",
  20869=>"010000111",
  20870=>"000011011",
  20871=>"000000100",
  20872=>"100110110",
  20873=>"100110000",
  20874=>"100111001",
  20875=>"000110000",
  20876=>"000111111",
  20877=>"011010110",
  20878=>"100111110",
  20879=>"011101110",
  20880=>"001011101",
  20881=>"000011100",
  20882=>"001110001",
  20883=>"100010111",
  20884=>"101010101",
  20885=>"000011100",
  20886=>"001101100",
  20887=>"101110111",
  20888=>"110010111",
  20889=>"001110000",
  20890=>"001110000",
  20891=>"110000100",
  20892=>"011100111",
  20893=>"010000110",
  20894=>"101111100",
  20895=>"000000010",
  20896=>"011110000",
  20897=>"111001001",
  20898=>"111010100",
  20899=>"000101100",
  20900=>"110110111",
  20901=>"111010000",
  20902=>"001001010",
  20903=>"111001000",
  20904=>"111011011",
  20905=>"111101001",
  20906=>"010110111",
  20907=>"001011000",
  20908=>"000110010",
  20909=>"000000000",
  20910=>"001010000",
  20911=>"110011101",
  20912=>"100010101",
  20913=>"001010000",
  20914=>"101111000",
  20915=>"110110010",
  20916=>"110101101",
  20917=>"011111011",
  20918=>"110010001",
  20919=>"101101001",
  20920=>"000001111",
  20921=>"100101100",
  20922=>"110111101",
  20923=>"110001001",
  20924=>"101011001",
  20925=>"000011000",
  20926=>"001101101",
  20927=>"010110010",
  20928=>"001000000",
  20929=>"111101110",
  20930=>"011111110",
  20931=>"010010111",
  20932=>"000110000",
  20933=>"011110010",
  20934=>"010111100",
  20935=>"110100111",
  20936=>"000011001",
  20937=>"111000110",
  20938=>"100100010",
  20939=>"010010001",
  20940=>"000100110",
  20941=>"101110000",
  20942=>"010110100",
  20943=>"010011011",
  20944=>"100111110",
  20945=>"101100000",
  20946=>"000001111",
  20947=>"001011111",
  20948=>"000110011",
  20949=>"011100000",
  20950=>"100101011",
  20951=>"100111000",
  20952=>"010010010",
  20953=>"011011100",
  20954=>"011010100",
  20955=>"000111101",
  20956=>"100010111",
  20957=>"001010010",
  20958=>"000010100",
  20959=>"100001101",
  20960=>"100110101",
  20961=>"001000110",
  20962=>"101000110",
  20963=>"011111001",
  20964=>"110010010",
  20965=>"101100000",
  20966=>"010101001",
  20967=>"011101011",
  20968=>"010001000",
  20969=>"010000110",
  20970=>"000101110",
  20971=>"111001111",
  20972=>"011000110",
  20973=>"010110111",
  20974=>"100110010",
  20975=>"110110010",
  20976=>"100010110",
  20977=>"111010001",
  20978=>"111010000",
  20979=>"001101100",
  20980=>"011010011",
  20981=>"000110111",
  20982=>"001110000",
  20983=>"101000110",
  20984=>"011110011",
  20985=>"011111000",
  20986=>"100000111",
  20987=>"101100101",
  20988=>"100010000",
  20989=>"111111011",
  20990=>"010001100",
  20991=>"011100010",
  20992=>"001111111",
  20993=>"111000111",
  20994=>"111010011",
  20995=>"011101111",
  20996=>"010000110",
  20997=>"110001011",
  20998=>"100100010",
  20999=>"010111010",
  21000=>"001101110",
  21001=>"000110010",
  21002=>"010101111",
  21003=>"110001010",
  21004=>"100110010",
  21005=>"011111111",
  21006=>"011111011",
  21007=>"100011010",
  21008=>"110101101",
  21009=>"000000101",
  21010=>"101001101",
  21011=>"110000001",
  21012=>"111111000",
  21013=>"001111100",
  21014=>"111001101",
  21015=>"011100100",
  21016=>"100001100",
  21017=>"101000110",
  21018=>"000001100",
  21019=>"000001100",
  21020=>"101001100",
  21021=>"100010101",
  21022=>"100100010",
  21023=>"011001000",
  21024=>"110010000",
  21025=>"111101100",
  21026=>"011110000",
  21027=>"001001101",
  21028=>"011001101",
  21029=>"110101011",
  21030=>"110101111",
  21031=>"100001010",
  21032=>"100000110",
  21033=>"000011000",
  21034=>"001011000",
  21035=>"001111001",
  21036=>"010100111",
  21037=>"111100000",
  21038=>"000110100",
  21039=>"010100101",
  21040=>"001111011",
  21041=>"001010111",
  21042=>"000001111",
  21043=>"011100111",
  21044=>"001000010",
  21045=>"111111100",
  21046=>"010000010",
  21047=>"111101010",
  21048=>"110111001",
  21049=>"001110100",
  21050=>"110111101",
  21051=>"100000010",
  21052=>"000100001",
  21053=>"101010110",
  21054=>"011000000",
  21055=>"111110011",
  21056=>"011011011",
  21057=>"001110001",
  21058=>"011000000",
  21059=>"011011100",
  21060=>"100101101",
  21061=>"101010011",
  21062=>"100001010",
  21063=>"111001000",
  21064=>"101001110",
  21065=>"010111101",
  21066=>"000101000",
  21067=>"000000101",
  21068=>"100100010",
  21069=>"010000010",
  21070=>"001001111",
  21071=>"010000000",
  21072=>"000001000",
  21073=>"001000111",
  21074=>"101000000",
  21075=>"101011001",
  21076=>"000000001",
  21077=>"000001111",
  21078=>"000000010",
  21079=>"011001101",
  21080=>"010111011",
  21081=>"110110001",
  21082=>"011111001",
  21083=>"101000000",
  21084=>"100011010",
  21085=>"111000000",
  21086=>"000010001",
  21087=>"101100101",
  21088=>"110000011",
  21089=>"101011001",
  21090=>"101010110",
  21091=>"011110011",
  21092=>"001111000",
  21093=>"000101101",
  21094=>"001001111",
  21095=>"001101011",
  21096=>"000101111",
  21097=>"101000000",
  21098=>"110010001",
  21099=>"010101110",
  21100=>"011000001",
  21101=>"000111110",
  21102=>"001101001",
  21103=>"100110111",
  21104=>"101011000",
  21105=>"000000111",
  21106=>"001011001",
  21107=>"111011100",
  21108=>"010111100",
  21109=>"011101000",
  21110=>"011101101",
  21111=>"011100010",
  21112=>"100000000",
  21113=>"111000011",
  21114=>"001111101",
  21115=>"011000001",
  21116=>"101001111",
  21117=>"001011001",
  21118=>"111110000",
  21119=>"111011010",
  21120=>"110010111",
  21121=>"110111011",
  21122=>"110110111",
  21123=>"000001101",
  21124=>"001100110",
  21125=>"101001100",
  21126=>"111101111",
  21127=>"101101000",
  21128=>"110110101",
  21129=>"111100110",
  21130=>"011010101",
  21131=>"100111010",
  21132=>"011000101",
  21133=>"110000101",
  21134=>"100010010",
  21135=>"110001111",
  21136=>"010111010",
  21137=>"111111111",
  21138=>"000010011",
  21139=>"110110111",
  21140=>"101110101",
  21141=>"101001110",
  21142=>"110001101",
  21143=>"001011011",
  21144=>"110000001",
  21145=>"110000011",
  21146=>"000000110",
  21147=>"100011000",
  21148=>"100101101",
  21149=>"100111101",
  21150=>"000110010",
  21151=>"001000011",
  21152=>"001001101",
  21153=>"101001000",
  21154=>"100000111",
  21155=>"010111110",
  21156=>"010100001",
  21157=>"011001100",
  21158=>"001111101",
  21159=>"111110110",
  21160=>"001100111",
  21161=>"001100101",
  21162=>"001001111",
  21163=>"110000111",
  21164=>"000110100",
  21165=>"101110010",
  21166=>"010110010",
  21167=>"010110010",
  21168=>"101110101",
  21169=>"011100111",
  21170=>"001010010",
  21171=>"111101001",
  21172=>"010000010",
  21173=>"000000011",
  21174=>"100111000",
  21175=>"110000110",
  21176=>"111000101",
  21177=>"011101001",
  21178=>"010000010",
  21179=>"001100000",
  21180=>"001100111",
  21181=>"001000001",
  21182=>"000111101",
  21183=>"010110110",
  21184=>"000110110",
  21185=>"011000101",
  21186=>"010111101",
  21187=>"001001101",
  21188=>"100010110",
  21189=>"000110000",
  21190=>"001101000",
  21191=>"111011110",
  21192=>"110111010",
  21193=>"010011001",
  21194=>"110000111",
  21195=>"001111110",
  21196=>"000001101",
  21197=>"001000101",
  21198=>"010101110",
  21199=>"000010001",
  21200=>"101010100",
  21201=>"000100000",
  21202=>"011000110",
  21203=>"000011010",
  21204=>"011001111",
  21205=>"010011001",
  21206=>"010101000",
  21207=>"101001111",
  21208=>"001000000",
  21209=>"010000110",
  21210=>"011011111",
  21211=>"011000111",
  21212=>"000110001",
  21213=>"101000111",
  21214=>"101110011",
  21215=>"001010100",
  21216=>"100001000",
  21217=>"101110001",
  21218=>"110101000",
  21219=>"001100000",
  21220=>"010010010",
  21221=>"101000010",
  21222=>"000111000",
  21223=>"001011000",
  21224=>"010010110",
  21225=>"000100011",
  21226=>"011010110",
  21227=>"110110111",
  21228=>"010001011",
  21229=>"110000001",
  21230=>"001010111",
  21231=>"010010100",
  21232=>"110100100",
  21233=>"101100010",
  21234=>"101111010",
  21235=>"111100010",
  21236=>"011111000",
  21237=>"110001000",
  21238=>"000110010",
  21239=>"000101000",
  21240=>"101000011",
  21241=>"000000100",
  21242=>"100110101",
  21243=>"101100000",
  21244=>"110010100",
  21245=>"011110011",
  21246=>"101010010",
  21247=>"101010001",
  21248=>"010011101",
  21249=>"100101110",
  21250=>"110010111",
  21251=>"110101101",
  21252=>"100100010",
  21253=>"111101010",
  21254=>"001001001",
  21255=>"000011110",
  21256=>"010101000",
  21257=>"101010011",
  21258=>"101101001",
  21259=>"111100001",
  21260=>"101100111",
  21261=>"111011010",
  21262=>"010000101",
  21263=>"110101000",
  21264=>"110111000",
  21265=>"000000110",
  21266=>"001000010",
  21267=>"100010001",
  21268=>"011110100",
  21269=>"000010010",
  21270=>"000100100",
  21271=>"110000010",
  21272=>"111101101",
  21273=>"010011001",
  21274=>"000110000",
  21275=>"011101111",
  21276=>"111011100",
  21277=>"001001111",
  21278=>"011010000",
  21279=>"100101000",
  21280=>"101110110",
  21281=>"001010100",
  21282=>"100001011",
  21283=>"100010011",
  21284=>"010001100",
  21285=>"111010010",
  21286=>"010010000",
  21287=>"111110011",
  21288=>"000000101",
  21289=>"100000010",
  21290=>"111110001",
  21291=>"110111100",
  21292=>"010010101",
  21293=>"010100001",
  21294=>"110011100",
  21295=>"011000100",
  21296=>"001011100",
  21297=>"110101100",
  21298=>"010100000",
  21299=>"101001111",
  21300=>"001111101",
  21301=>"100010110",
  21302=>"111111010",
  21303=>"001101111",
  21304=>"010100011",
  21305=>"010000001",
  21306=>"111000001",
  21307=>"010101100",
  21308=>"001101011",
  21309=>"010010111",
  21310=>"011111111",
  21311=>"110111110",
  21312=>"001000111",
  21313=>"011100010",
  21314=>"110001101",
  21315=>"100010000",
  21316=>"111111001",
  21317=>"010100111",
  21318=>"110000010",
  21319=>"110010101",
  21320=>"100000011",
  21321=>"010001011",
  21322=>"001001100",
  21323=>"000011101",
  21324=>"001111110",
  21325=>"101001000",
  21326=>"000010100",
  21327=>"100001110",
  21328=>"110101011",
  21329=>"010000011",
  21330=>"110110010",
  21331=>"110101000",
  21332=>"001010001",
  21333=>"111011100",
  21334=>"110100101",
  21335=>"101110000",
  21336=>"010101010",
  21337=>"011100110",
  21338=>"010001100",
  21339=>"001001100",
  21340=>"111000111",
  21341=>"011000100",
  21342=>"000000001",
  21343=>"110100000",
  21344=>"000100010",
  21345=>"000001111",
  21346=>"010010111",
  21347=>"000100001",
  21348=>"011111010",
  21349=>"100100110",
  21350=>"011100100",
  21351=>"001100001",
  21352=>"001000111",
  21353=>"010010011",
  21354=>"001101000",
  21355=>"000011011",
  21356=>"010010011",
  21357=>"011100011",
  21358=>"011100101",
  21359=>"001110011",
  21360=>"000011110",
  21361=>"100111001",
  21362=>"110100000",
  21363=>"100010001",
  21364=>"101000001",
  21365=>"010001000",
  21366=>"111000010",
  21367=>"110100111",
  21368=>"111101000",
  21369=>"011110011",
  21370=>"010100111",
  21371=>"010100000",
  21372=>"011000011",
  21373=>"000110001",
  21374=>"100000010",
  21375=>"101110100",
  21376=>"101111011",
  21377=>"110011111",
  21378=>"101010111",
  21379=>"000100000",
  21380=>"111001110",
  21381=>"011000100",
  21382=>"001000011",
  21383=>"100011110",
  21384=>"010011000",
  21385=>"000000011",
  21386=>"111111111",
  21387=>"111010101",
  21388=>"001111010",
  21389=>"111011000",
  21390=>"011100011",
  21391=>"010100101",
  21392=>"101101110",
  21393=>"011110001",
  21394=>"000100101",
  21395=>"011010100",
  21396=>"011111000",
  21397=>"111011110",
  21398=>"000110111",
  21399=>"010001011",
  21400=>"110001010",
  21401=>"001000001",
  21402=>"101010101",
  21403=>"011111111",
  21404=>"010101001",
  21405=>"000011000",
  21406=>"110110011",
  21407=>"010100010",
  21408=>"001001011",
  21409=>"101001010",
  21410=>"100101100",
  21411=>"011101000",
  21412=>"100000000",
  21413=>"110010100",
  21414=>"000000010",
  21415=>"001011011",
  21416=>"110001011",
  21417=>"001111000",
  21418=>"111011110",
  21419=>"111001000",
  21420=>"011100101",
  21421=>"010001000",
  21422=>"000111001",
  21423=>"010011010",
  21424=>"001010001",
  21425=>"010011100",
  21426=>"010011101",
  21427=>"000111010",
  21428=>"101000010",
  21429=>"101011010",
  21430=>"011000111",
  21431=>"101011111",
  21432=>"111011010",
  21433=>"100011101",
  21434=>"010000111",
  21435=>"101111100",
  21436=>"101111011",
  21437=>"111101000",
  21438=>"101110001",
  21439=>"001011111",
  21440=>"010110111",
  21441=>"011100001",
  21442=>"110100011",
  21443=>"001001100",
  21444=>"011101111",
  21445=>"000101001",
  21446=>"010101001",
  21447=>"110100100",
  21448=>"000001000",
  21449=>"001010101",
  21450=>"001000001",
  21451=>"001010100",
  21452=>"011010011",
  21453=>"001101100",
  21454=>"011100100",
  21455=>"010100011",
  21456=>"011101100",
  21457=>"011010011",
  21458=>"111111001",
  21459=>"001000101",
  21460=>"111111100",
  21461=>"010111100",
  21462=>"111101000",
  21463=>"110110110",
  21464=>"000010111",
  21465=>"000100010",
  21466=>"111111011",
  21467=>"100101010",
  21468=>"101010100",
  21469=>"110000100",
  21470=>"100110110",
  21471=>"010010001",
  21472=>"010001000",
  21473=>"110011001",
  21474=>"100010011",
  21475=>"010011000",
  21476=>"011010110",
  21477=>"001000110",
  21478=>"110100100",
  21479=>"101101010",
  21480=>"000010001",
  21481=>"111110000",
  21482=>"101111010",
  21483=>"010000111",
  21484=>"101011101",
  21485=>"110001101",
  21486=>"110111000",
  21487=>"110000010",
  21488=>"101100101",
  21489=>"001000001",
  21490=>"001000001",
  21491=>"111100111",
  21492=>"010100100",
  21493=>"101100110",
  21494=>"001010010",
  21495=>"010111111",
  21496=>"111000001",
  21497=>"100100110",
  21498=>"111101000",
  21499=>"110111101",
  21500=>"110000101",
  21501=>"010000011",
  21502=>"110010000",
  21503=>"111111111",
  21504=>"111010100",
  21505=>"010100000",
  21506=>"101001110",
  21507=>"000001111",
  21508=>"011110010",
  21509=>"011000000",
  21510=>"101100100",
  21511=>"000011111",
  21512=>"011000011",
  21513=>"010000010",
  21514=>"010000000",
  21515=>"101001111",
  21516=>"011101101",
  21517=>"011011110",
  21518=>"001011110",
  21519=>"011011111",
  21520=>"100010001",
  21521=>"101001000",
  21522=>"001010010",
  21523=>"111000110",
  21524=>"000110000",
  21525=>"111010101",
  21526=>"111111101",
  21527=>"000000010",
  21528=>"001101100",
  21529=>"000111000",
  21530=>"101101001",
  21531=>"100100110",
  21532=>"010110110",
  21533=>"101101110",
  21534=>"000000110",
  21535=>"100011101",
  21536=>"001011110",
  21537=>"111110110",
  21538=>"000001110",
  21539=>"011010100",
  21540=>"001110111",
  21541=>"010111111",
  21542=>"010100110",
  21543=>"100100110",
  21544=>"111000101",
  21545=>"010000110",
  21546=>"101110010",
  21547=>"001000000",
  21548=>"000111101",
  21549=>"111110101",
  21550=>"100101111",
  21551=>"010001101",
  21552=>"011001000",
  21553=>"101011110",
  21554=>"010000100",
  21555=>"101111000",
  21556=>"011011101",
  21557=>"100010000",
  21558=>"001110001",
  21559=>"000101111",
  21560=>"011011111",
  21561=>"110001000",
  21562=>"000100110",
  21563=>"101000001",
  21564=>"000100001",
  21565=>"101111101",
  21566=>"101010100",
  21567=>"011111101",
  21568=>"010010111",
  21569=>"000000000",
  21570=>"101000101",
  21571=>"010011010",
  21572=>"110101101",
  21573=>"000010011",
  21574=>"001011010",
  21575=>"100001010",
  21576=>"101101010",
  21577=>"110010010",
  21578=>"100000000",
  21579=>"110111001",
  21580=>"100011001",
  21581=>"101001110",
  21582=>"011000001",
  21583=>"101100101",
  21584=>"111010101",
  21585=>"001001100",
  21586=>"100101011",
  21587=>"000010101",
  21588=>"001011001",
  21589=>"001000100",
  21590=>"001010111",
  21591=>"010110000",
  21592=>"010101111",
  21593=>"001100011",
  21594=>"100100111",
  21595=>"101101100",
  21596=>"101000011",
  21597=>"100101110",
  21598=>"101100010",
  21599=>"011011000",
  21600=>"110110011",
  21601=>"110111101",
  21602=>"011001001",
  21603=>"000100111",
  21604=>"001100100",
  21605=>"111100000",
  21606=>"000110011",
  21607=>"000011100",
  21608=>"001111001",
  21609=>"100011110",
  21610=>"100111110",
  21611=>"011111101",
  21612=>"011110010",
  21613=>"110000011",
  21614=>"111010110",
  21615=>"101011010",
  21616=>"110011011",
  21617=>"101110000",
  21618=>"110111110",
  21619=>"001001011",
  21620=>"101101111",
  21621=>"101011000",
  21622=>"111010001",
  21623=>"100100010",
  21624=>"001111000",
  21625=>"101101111",
  21626=>"110011001",
  21627=>"000101101",
  21628=>"111101011",
  21629=>"010101010",
  21630=>"011001110",
  21631=>"110110100",
  21632=>"000101100",
  21633=>"100010010",
  21634=>"111110010",
  21635=>"010111110",
  21636=>"000101111",
  21637=>"011101000",
  21638=>"111111000",
  21639=>"100011100",
  21640=>"000011000",
  21641=>"011010100",
  21642=>"111011010",
  21643=>"111110101",
  21644=>"011111101",
  21645=>"101110110",
  21646=>"000101110",
  21647=>"000010011",
  21648=>"001010101",
  21649=>"011101110",
  21650=>"000011101",
  21651=>"000010010",
  21652=>"011101111",
  21653=>"001100110",
  21654=>"010111110",
  21655=>"110110010",
  21656=>"000101011",
  21657=>"101110100",
  21658=>"010011101",
  21659=>"111110000",
  21660=>"111101011",
  21661=>"000001110",
  21662=>"000100001",
  21663=>"010100000",
  21664=>"110101101",
  21665=>"101100010",
  21666=>"111110111",
  21667=>"100001110",
  21668=>"111110101",
  21669=>"100010000",
  21670=>"011101110",
  21671=>"100101110",
  21672=>"111011010",
  21673=>"110000110",
  21674=>"010101100",
  21675=>"100010001",
  21676=>"101101101",
  21677=>"101010111",
  21678=>"110111110",
  21679=>"100100000",
  21680=>"111001111",
  21681=>"000110101",
  21682=>"111111100",
  21683=>"000100110",
  21684=>"101000001",
  21685=>"110111011",
  21686=>"111010110",
  21687=>"110011011",
  21688=>"000011001",
  21689=>"010111111",
  21690=>"101001110",
  21691=>"010000100",
  21692=>"000110010",
  21693=>"001011000",
  21694=>"101101101",
  21695=>"011000101",
  21696=>"010010010",
  21697=>"110110101",
  21698=>"000001011",
  21699=>"001000101",
  21700=>"001101000",
  21701=>"110110000",
  21702=>"010010110",
  21703=>"101111111",
  21704=>"001011100",
  21705=>"101111010",
  21706=>"010011111",
  21707=>"001001111",
  21708=>"101110111",
  21709=>"011010111",
  21710=>"010010101",
  21711=>"110010000",
  21712=>"000000100",
  21713=>"000001100",
  21714=>"001101100",
  21715=>"011111001",
  21716=>"100101110",
  21717=>"101001111",
  21718=>"111110010",
  21719=>"010110011",
  21720=>"010000100",
  21721=>"100000101",
  21722=>"001001000",
  21723=>"001010011",
  21724=>"001011100",
  21725=>"100101100",
  21726=>"010100101",
  21727=>"000111001",
  21728=>"100011011",
  21729=>"100010000",
  21730=>"111010110",
  21731=>"110111111",
  21732=>"101001101",
  21733=>"111101011",
  21734=>"100011111",
  21735=>"000010001",
  21736=>"011110000",
  21737=>"010100000",
  21738=>"001110001",
  21739=>"100010110",
  21740=>"011110100",
  21741=>"010010010",
  21742=>"110111110",
  21743=>"101100011",
  21744=>"110011001",
  21745=>"111100111",
  21746=>"000000001",
  21747=>"101010100",
  21748=>"000011110",
  21749=>"000110100",
  21750=>"010111011",
  21751=>"000110000",
  21752=>"010011111",
  21753=>"100001111",
  21754=>"100001111",
  21755=>"001101110",
  21756=>"110000000",
  21757=>"010011101",
  21758=>"101011010",
  21759=>"101010101",
  21760=>"011110000",
  21761=>"100110110",
  21762=>"001011001",
  21763=>"011010111",
  21764=>"111011100",
  21765=>"110000110",
  21766=>"110100111",
  21767=>"000011001",
  21768=>"010001111",
  21769=>"000100010",
  21770=>"101111111",
  21771=>"101000011",
  21772=>"010011110",
  21773=>"110011011",
  21774=>"100101001",
  21775=>"111100000",
  21776=>"011011111",
  21777=>"110110000",
  21778=>"001101101",
  21779=>"110000011",
  21780=>"101101101",
  21781=>"010110111",
  21782=>"000010100",
  21783=>"101101110",
  21784=>"011110011",
  21785=>"000010100",
  21786=>"100110111",
  21787=>"111110000",
  21788=>"011001001",
  21789=>"100100111",
  21790=>"011100001",
  21791=>"010101000",
  21792=>"001111110",
  21793=>"101100101",
  21794=>"110001111",
  21795=>"110010110",
  21796=>"011100001",
  21797=>"110111100",
  21798=>"011010010",
  21799=>"100111110",
  21800=>"110000011",
  21801=>"101001000",
  21802=>"110000000",
  21803=>"100110001",
  21804=>"110001011",
  21805=>"110000010",
  21806=>"110110010",
  21807=>"111110011",
  21808=>"100110101",
  21809=>"000111111",
  21810=>"010000010",
  21811=>"000010000",
  21812=>"111011001",
  21813=>"000111101",
  21814=>"000010110",
  21815=>"000111010",
  21816=>"001000001",
  21817=>"001100111",
  21818=>"000000000",
  21819=>"011100111",
  21820=>"111001010",
  21821=>"011001111",
  21822=>"010001000",
  21823=>"111100110",
  21824=>"010011011",
  21825=>"111110100",
  21826=>"010101010",
  21827=>"101101010",
  21828=>"111010101",
  21829=>"010111101",
  21830=>"100011110",
  21831=>"110110100",
  21832=>"001001000",
  21833=>"010111000",
  21834=>"010101110",
  21835=>"111110011",
  21836=>"001101000",
  21837=>"111100111",
  21838=>"010101011",
  21839=>"101001000",
  21840=>"001000111",
  21841=>"101100101",
  21842=>"100001010",
  21843=>"011001101",
  21844=>"000010001",
  21845=>"000010101",
  21846=>"110110010",
  21847=>"111110000",
  21848=>"101111000",
  21849=>"101010111",
  21850=>"111011110",
  21851=>"010001100",
  21852=>"001101111",
  21853=>"110101111",
  21854=>"100101010",
  21855=>"001000111",
  21856=>"100001100",
  21857=>"111000111",
  21858=>"011100101",
  21859=>"000001111",
  21860=>"000111101",
  21861=>"110000011",
  21862=>"100010111",
  21863=>"101101101",
  21864=>"010001110",
  21865=>"000111100",
  21866=>"000010010",
  21867=>"100111000",
  21868=>"000001110",
  21869=>"111000000",
  21870=>"111110001",
  21871=>"110010110",
  21872=>"010010011",
  21873=>"000010111",
  21874=>"110111011",
  21875=>"001101100",
  21876=>"101001011",
  21877=>"111100001",
  21878=>"000111101",
  21879=>"000011010",
  21880=>"101000101",
  21881=>"101010100",
  21882=>"101001000",
  21883=>"100000111",
  21884=>"001100111",
  21885=>"110000000",
  21886=>"011000110",
  21887=>"110111011",
  21888=>"010010000",
  21889=>"100000110",
  21890=>"000101111",
  21891=>"100101111",
  21892=>"101011100",
  21893=>"001100111",
  21894=>"101001011",
  21895=>"000101110",
  21896=>"001101101",
  21897=>"111001101",
  21898=>"010000110",
  21899=>"001110101",
  21900=>"010010110",
  21901=>"000110000",
  21902=>"010110100",
  21903=>"110010001",
  21904=>"110100000",
  21905=>"000010000",
  21906=>"001001001",
  21907=>"111011100",
  21908=>"100010101",
  21909=>"110111001",
  21910=>"100111111",
  21911=>"101110111",
  21912=>"100110001",
  21913=>"100111100",
  21914=>"100111010",
  21915=>"001111011",
  21916=>"010111100",
  21917=>"000101111",
  21918=>"011011011",
  21919=>"110111111",
  21920=>"010001001",
  21921=>"100010010",
  21922=>"111111100",
  21923=>"111011101",
  21924=>"101100000",
  21925=>"001011000",
  21926=>"110100111",
  21927=>"100101010",
  21928=>"011000101",
  21929=>"111101101",
  21930=>"101111001",
  21931=>"111111001",
  21932=>"101000011",
  21933=>"011110011",
  21934=>"000000100",
  21935=>"101011100",
  21936=>"001110100",
  21937=>"111110001",
  21938=>"000000101",
  21939=>"111100111",
  21940=>"110111111",
  21941=>"111001000",
  21942=>"011001011",
  21943=>"010100100",
  21944=>"111000111",
  21945=>"100001100",
  21946=>"000111000",
  21947=>"101110001",
  21948=>"101011001",
  21949=>"110010101",
  21950=>"000101010",
  21951=>"111011111",
  21952=>"101001110",
  21953=>"000010000",
  21954=>"101001100",
  21955=>"101010011",
  21956=>"110011110",
  21957=>"011010010",
  21958=>"011001010",
  21959=>"000101000",
  21960=>"111011000",
  21961=>"110110111",
  21962=>"011001000",
  21963=>"000111101",
  21964=>"001110011",
  21965=>"000111001",
  21966=>"010000100",
  21967=>"111001001",
  21968=>"001000101",
  21969=>"011111110",
  21970=>"101010100",
  21971=>"111011010",
  21972=>"010000110",
  21973=>"110000100",
  21974=>"100011100",
  21975=>"000110111",
  21976=>"011011110",
  21977=>"111001001",
  21978=>"001000100",
  21979=>"010100001",
  21980=>"111011110",
  21981=>"101001010",
  21982=>"010110010",
  21983=>"111011110",
  21984=>"110011101",
  21985=>"001111100",
  21986=>"100011010",
  21987=>"110010000",
  21988=>"101111101",
  21989=>"111010001",
  21990=>"001001100",
  21991=>"010000110",
  21992=>"100110000",
  21993=>"001011110",
  21994=>"010101100",
  21995=>"001000111",
  21996=>"100011110",
  21997=>"110111001",
  21998=>"100100001",
  21999=>"000010100",
  22000=>"011001001",
  22001=>"010000000",
  22002=>"101011111",
  22003=>"001000111",
  22004=>"101101110",
  22005=>"110001010",
  22006=>"110000101",
  22007=>"101001010",
  22008=>"001110101",
  22009=>"111001101",
  22010=>"000110100",
  22011=>"010000110",
  22012=>"000000010",
  22013=>"001100101",
  22014=>"010110100",
  22015=>"100000010",
  22016=>"101100111",
  22017=>"111100010",
  22018=>"000000111",
  22019=>"101011011",
  22020=>"011101011",
  22021=>"000000001",
  22022=>"000010100",
  22023=>"001000001",
  22024=>"111001011",
  22025=>"010100001",
  22026=>"000110111",
  22027=>"011100011",
  22028=>"101100110",
  22029=>"111111101",
  22030=>"000010101",
  22031=>"110000101",
  22032=>"101011111",
  22033=>"101111110",
  22034=>"100110101",
  22035=>"011111011",
  22036=>"110111100",
  22037=>"001101011",
  22038=>"010111111",
  22039=>"101110110",
  22040=>"110010100",
  22041=>"101010000",
  22042=>"101111101",
  22043=>"111110010",
  22044=>"101000001",
  22045=>"110100000",
  22046=>"010000101",
  22047=>"110001101",
  22048=>"010101011",
  22049=>"101100011",
  22050=>"111100001",
  22051=>"000101100",
  22052=>"100100101",
  22053=>"001111110",
  22054=>"010010011",
  22055=>"000001000",
  22056=>"110101000",
  22057=>"001011111",
  22058=>"000101000",
  22059=>"011010100",
  22060=>"010110001",
  22061=>"010100010",
  22062=>"010001011",
  22063=>"101110110",
  22064=>"110100000",
  22065=>"000110100",
  22066=>"111101111",
  22067=>"100000101",
  22068=>"101010000",
  22069=>"001100110",
  22070=>"100100000",
  22071=>"010001111",
  22072=>"000001101",
  22073=>"010011111",
  22074=>"111000101",
  22075=>"111001100",
  22076=>"100100011",
  22077=>"001111000",
  22078=>"111000100",
  22079=>"011010110",
  22080=>"100100100",
  22081=>"100010001",
  22082=>"110001011",
  22083=>"011100010",
  22084=>"110110010",
  22085=>"010110110",
  22086=>"010111001",
  22087=>"011110001",
  22088=>"000010111",
  22089=>"101001111",
  22090=>"000011110",
  22091=>"001010100",
  22092=>"111111100",
  22093=>"011000001",
  22094=>"111111000",
  22095=>"111111100",
  22096=>"000110010",
  22097=>"001000100",
  22098=>"100001100",
  22099=>"010001110",
  22100=>"110011011",
  22101=>"111010010",
  22102=>"101000101",
  22103=>"011110101",
  22104=>"011100101",
  22105=>"001100011",
  22106=>"111100000",
  22107=>"000000100",
  22108=>"011001110",
  22109=>"000001011",
  22110=>"111001100",
  22111=>"100000000",
  22112=>"100111001",
  22113=>"100110110",
  22114=>"001111010",
  22115=>"010110010",
  22116=>"111000001",
  22117=>"010100100",
  22118=>"001011111",
  22119=>"000011100",
  22120=>"100110011",
  22121=>"101110111",
  22122=>"000100011",
  22123=>"100000000",
  22124=>"101010000",
  22125=>"010001000",
  22126=>"101000100",
  22127=>"010000101",
  22128=>"101010110",
  22129=>"001111001",
  22130=>"011101001",
  22131=>"101110001",
  22132=>"101111001",
  22133=>"101111001",
  22134=>"101111011",
  22135=>"100010100",
  22136=>"101000011",
  22137=>"101001111",
  22138=>"110101100",
  22139=>"011000010",
  22140=>"000101111",
  22141=>"100100010",
  22142=>"111000000",
  22143=>"110111101",
  22144=>"010100000",
  22145=>"000110000",
  22146=>"101101100",
  22147=>"001101111",
  22148=>"001110000",
  22149=>"010010101",
  22150=>"111010011",
  22151=>"101101100",
  22152=>"100100111",
  22153=>"000001010",
  22154=>"110001101",
  22155=>"110010000",
  22156=>"001001010",
  22157=>"001011010",
  22158=>"010101100",
  22159=>"011011011",
  22160=>"101101101",
  22161=>"010010010",
  22162=>"010111000",
  22163=>"000100001",
  22164=>"111001110",
  22165=>"111100110",
  22166=>"110011111",
  22167=>"100011001",
  22168=>"100110110",
  22169=>"011101011",
  22170=>"101111101",
  22171=>"101110010",
  22172=>"011011000",
  22173=>"000000001",
  22174=>"101110110",
  22175=>"010100100",
  22176=>"001100000",
  22177=>"000001001",
  22178=>"000110100",
  22179=>"101010010",
  22180=>"011100001",
  22181=>"001110110",
  22182=>"101001011",
  22183=>"010000000",
  22184=>"111111010",
  22185=>"011010000",
  22186=>"011111010",
  22187=>"010011100",
  22188=>"101011101",
  22189=>"011011011",
  22190=>"110000011",
  22191=>"111101111",
  22192=>"001010010",
  22193=>"111011011",
  22194=>"011110111",
  22195=>"100011110",
  22196=>"010000101",
  22197=>"111111010",
  22198=>"111100001",
  22199=>"011000000",
  22200=>"100111001",
  22201=>"001101011",
  22202=>"000000110",
  22203=>"111001010",
  22204=>"000101011",
  22205=>"000010011",
  22206=>"011011110",
  22207=>"110111111",
  22208=>"000010010",
  22209=>"010100100",
  22210=>"100001001",
  22211=>"000010110",
  22212=>"101111011",
  22213=>"000100100",
  22214=>"100100001",
  22215=>"001000001",
  22216=>"011000110",
  22217=>"011001001",
  22218=>"101110001",
  22219=>"001111011",
  22220=>"100100011",
  22221=>"010100111",
  22222=>"100001000",
  22223=>"110011100",
  22224=>"111010101",
  22225=>"111101010",
  22226=>"110000101",
  22227=>"000111010",
  22228=>"111111010",
  22229=>"010111010",
  22230=>"111000110",
  22231=>"001101101",
  22232=>"100110101",
  22233=>"100101110",
  22234=>"001010000",
  22235=>"101110100",
  22236=>"011111011",
  22237=>"010011010",
  22238=>"111011100",
  22239=>"001101010",
  22240=>"011101100",
  22241=>"001010000",
  22242=>"000100111",
  22243=>"000010000",
  22244=>"000011001",
  22245=>"111111100",
  22246=>"001000100",
  22247=>"100011110",
  22248=>"001100111",
  22249=>"110100110",
  22250=>"001000101",
  22251=>"011001101",
  22252=>"011011001",
  22253=>"000011110",
  22254=>"011110110",
  22255=>"100010011",
  22256=>"000101000",
  22257=>"000010110",
  22258=>"101010101",
  22259=>"111011111",
  22260=>"010111101",
  22261=>"111011110",
  22262=>"110100111",
  22263=>"100110100",
  22264=>"100010001",
  22265=>"111110110",
  22266=>"100110001",
  22267=>"000000101",
  22268=>"010000111",
  22269=>"011100101",
  22270=>"000011001",
  22271=>"010001000",
  22272=>"101000101",
  22273=>"010000001",
  22274=>"001011010",
  22275=>"010001001",
  22276=>"001001010",
  22277=>"110101101",
  22278=>"111101111",
  22279=>"110001010",
  22280=>"001000011",
  22281=>"100100010",
  22282=>"110001010",
  22283=>"110110100",
  22284=>"000001010",
  22285=>"101011000",
  22286=>"001100100",
  22287=>"110000001",
  22288=>"010001000",
  22289=>"111111100",
  22290=>"111000100",
  22291=>"011110000",
  22292=>"101000101",
  22293=>"111110011",
  22294=>"001101001",
  22295=>"101000010",
  22296=>"000101000",
  22297=>"110000011",
  22298=>"111100000",
  22299=>"111111101",
  22300=>"111100110",
  22301=>"010110000",
  22302=>"011100101",
  22303=>"111111111",
  22304=>"010010101",
  22305=>"011111000",
  22306=>"110000011",
  22307=>"110111001",
  22308=>"000101111",
  22309=>"100111101",
  22310=>"110110011",
  22311=>"010110110",
  22312=>"001110000",
  22313=>"000000001",
  22314=>"000101010",
  22315=>"010010010",
  22316=>"110111001",
  22317=>"001000000",
  22318=>"110111001",
  22319=>"010001110",
  22320=>"011000000",
  22321=>"011010111",
  22322=>"010100111",
  22323=>"000011001",
  22324=>"000101010",
  22325=>"101000001",
  22326=>"110000110",
  22327=>"110111001",
  22328=>"000111001",
  22329=>"000010000",
  22330=>"101011001",
  22331=>"100110100",
  22332=>"000010110",
  22333=>"101111110",
  22334=>"000011100",
  22335=>"110101100",
  22336=>"010010010",
  22337=>"100010010",
  22338=>"000010010",
  22339=>"101011011",
  22340=>"000101101",
  22341=>"111111001",
  22342=>"010111110",
  22343=>"110100111",
  22344=>"010101001",
  22345=>"001000111",
  22346=>"011110001",
  22347=>"010001000",
  22348=>"011110110",
  22349=>"000010111",
  22350=>"111101101",
  22351=>"111010100",
  22352=>"001110011",
  22353=>"000110111",
  22354=>"011110110",
  22355=>"011000010",
  22356=>"000001111",
  22357=>"101011011",
  22358=>"001100111",
  22359=>"011001111",
  22360=>"101110100",
  22361=>"101010111",
  22362=>"001110001",
  22363=>"000100110",
  22364=>"000000100",
  22365=>"011110010",
  22366=>"100001001",
  22367=>"010111101",
  22368=>"001001010",
  22369=>"000110110",
  22370=>"110010000",
  22371=>"010110100",
  22372=>"000110111",
  22373=>"111001011",
  22374=>"100101001",
  22375=>"111110000",
  22376=>"011111111",
  22377=>"101110000",
  22378=>"111000011",
  22379=>"000101111",
  22380=>"000101111",
  22381=>"110110000",
  22382=>"100010001",
  22383=>"000101000",
  22384=>"111010101",
  22385=>"111000011",
  22386=>"000011111",
  22387=>"111111010",
  22388=>"011010110",
  22389=>"000110011",
  22390=>"000011100",
  22391=>"010110000",
  22392=>"111011010",
  22393=>"111001101",
  22394=>"101001110",
  22395=>"110111011",
  22396=>"000010100",
  22397=>"110011011",
  22398=>"101100010",
  22399=>"111100100",
  22400=>"010110101",
  22401=>"001010010",
  22402=>"111111111",
  22403=>"101101011",
  22404=>"011010101",
  22405=>"111000110",
  22406=>"100101000",
  22407=>"001110110",
  22408=>"101101111",
  22409=>"101100000",
  22410=>"111101100",
  22411=>"111011111",
  22412=>"000010101",
  22413=>"011110111",
  22414=>"101101110",
  22415=>"001010011",
  22416=>"100100111",
  22417=>"111001110",
  22418=>"000000111",
  22419=>"001010111",
  22420=>"011001110",
  22421=>"111000111",
  22422=>"100111101",
  22423=>"100001000",
  22424=>"111111110",
  22425=>"111110000",
  22426=>"101001000",
  22427=>"010100110",
  22428=>"110101110",
  22429=>"011111010",
  22430=>"011111111",
  22431=>"100001000",
  22432=>"101011110",
  22433=>"010101000",
  22434=>"101000100",
  22435=>"101101011",
  22436=>"000101101",
  22437=>"110101111",
  22438=>"110001011",
  22439=>"000111110",
  22440=>"110001110",
  22441=>"010010010",
  22442=>"100001101",
  22443=>"111011001",
  22444=>"111100001",
  22445=>"101001000",
  22446=>"100110111",
  22447=>"110000000",
  22448=>"011100100",
  22449=>"111111010",
  22450=>"111100101",
  22451=>"110011000",
  22452=>"001101101",
  22453=>"110101111",
  22454=>"110011111",
  22455=>"010000011",
  22456=>"101010010",
  22457=>"011000011",
  22458=>"001001011",
  22459=>"110111011",
  22460=>"001000000",
  22461=>"000010001",
  22462=>"000000101",
  22463=>"000000000",
  22464=>"011110100",
  22465=>"000011110",
  22466=>"000000001",
  22467=>"001110010",
  22468=>"010010111",
  22469=>"010111111",
  22470=>"110111111",
  22471=>"100101001",
  22472=>"011000111",
  22473=>"101111100",
  22474=>"001111001",
  22475=>"100010000",
  22476=>"111010110",
  22477=>"000110111",
  22478=>"110011100",
  22479=>"111001111",
  22480=>"000011010",
  22481=>"100111100",
  22482=>"010111111",
  22483=>"110011011",
  22484=>"000110111",
  22485=>"001101101",
  22486=>"100110010",
  22487=>"110100010",
  22488=>"111011001",
  22489=>"000100011",
  22490=>"001011110",
  22491=>"100101001",
  22492=>"010111001",
  22493=>"001011101",
  22494=>"000101001",
  22495=>"111110010",
  22496=>"110101001",
  22497=>"010001100",
  22498=>"001000100",
  22499=>"000010110",
  22500=>"001111000",
  22501=>"000111010",
  22502=>"110011000",
  22503=>"001101000",
  22504=>"011000101",
  22505=>"111000000",
  22506=>"111100000",
  22507=>"000000111",
  22508=>"110101111",
  22509=>"110010101",
  22510=>"101010101",
  22511=>"011010001",
  22512=>"110110010",
  22513=>"010011101",
  22514=>"110100001",
  22515=>"110011100",
  22516=>"100010010",
  22517=>"000101111",
  22518=>"010100011",
  22519=>"001000101",
  22520=>"111110110",
  22521=>"111111110",
  22522=>"011100001",
  22523=>"000010111",
  22524=>"101000010",
  22525=>"101111100",
  22526=>"001011001",
  22527=>"100001001",
  22528=>"100101100",
  22529=>"011001001",
  22530=>"000110000",
  22531=>"000100010",
  22532=>"011101001",
  22533=>"010111001",
  22534=>"001010100",
  22535=>"110001111",
  22536=>"010011010",
  22537=>"001101110",
  22538=>"111001100",
  22539=>"001011101",
  22540=>"111111100",
  22541=>"011010001",
  22542=>"010001010",
  22543=>"001110011",
  22544=>"010010000",
  22545=>"110010000",
  22546=>"100010000",
  22547=>"010001001",
  22548=>"001011101",
  22549=>"011100111",
  22550=>"010100000",
  22551=>"000101100",
  22552=>"111010000",
  22553=>"000010110",
  22554=>"110110010",
  22555=>"111111010",
  22556=>"010100101",
  22557=>"100011101",
  22558=>"001100011",
  22559=>"101100010",
  22560=>"111001000",
  22561=>"011100111",
  22562=>"111111101",
  22563=>"101110111",
  22564=>"111111111",
  22565=>"101000001",
  22566=>"111101000",
  22567=>"011101101",
  22568=>"010011000",
  22569=>"100001110",
  22570=>"100110101",
  22571=>"010101001",
  22572=>"001000000",
  22573=>"000011101",
  22574=>"110100110",
  22575=>"101000000",
  22576=>"111011110",
  22577=>"001001011",
  22578=>"111100010",
  22579=>"111111110",
  22580=>"110110110",
  22581=>"100111010",
  22582=>"101110111",
  22583=>"100001011",
  22584=>"100001101",
  22585=>"100110000",
  22586=>"011011110",
  22587=>"101010101",
  22588=>"111010100",
  22589=>"100000100",
  22590=>"001111101",
  22591=>"110101101",
  22592=>"011001101",
  22593=>"001000010",
  22594=>"010100111",
  22595=>"110010000",
  22596=>"111101000",
  22597=>"101100101",
  22598=>"101000010",
  22599=>"100010100",
  22600=>"111100100",
  22601=>"010111011",
  22602=>"000110010",
  22603=>"001100011",
  22604=>"010111001",
  22605=>"010011111",
  22606=>"010011110",
  22607=>"010001001",
  22608=>"010110001",
  22609=>"110110110",
  22610=>"111001011",
  22611=>"001111000",
  22612=>"000011100",
  22613=>"100101000",
  22614=>"001011000",
  22615=>"110110111",
  22616=>"010100001",
  22617=>"110101100",
  22618=>"001010110",
  22619=>"000110010",
  22620=>"110010110",
  22621=>"000101111",
  22622=>"110111111",
  22623=>"010110001",
  22624=>"110100110",
  22625=>"000000111",
  22626=>"111111001",
  22627=>"001100001",
  22628=>"110001111",
  22629=>"100100111",
  22630=>"010110111",
  22631=>"001011100",
  22632=>"100001110",
  22633=>"011000010",
  22634=>"000011001",
  22635=>"001111111",
  22636=>"111100100",
  22637=>"010100110",
  22638=>"111011110",
  22639=>"100100101",
  22640=>"011110001",
  22641=>"001110000",
  22642=>"001110111",
  22643=>"100001001",
  22644=>"100100000",
  22645=>"100010000",
  22646=>"111110101",
  22647=>"111010011",
  22648=>"011110011",
  22649=>"101111101",
  22650=>"100001010",
  22651=>"001101011",
  22652=>"110100100",
  22653=>"001011000",
  22654=>"011000010",
  22655=>"100000110",
  22656=>"011100000",
  22657=>"010110000",
  22658=>"100001110",
  22659=>"000001101",
  22660=>"010010110",
  22661=>"110011011",
  22662=>"010001000",
  22663=>"010110011",
  22664=>"111111110",
  22665=>"010010000",
  22666=>"101100001",
  22667=>"011000101",
  22668=>"010011011",
  22669=>"101000101",
  22670=>"000011100",
  22671=>"010100011",
  22672=>"110111001",
  22673=>"000001000",
  22674=>"011011011",
  22675=>"111010100",
  22676=>"010101000",
  22677=>"101000011",
  22678=>"101110000",
  22679=>"001100010",
  22680=>"110011100",
  22681=>"101100010",
  22682=>"110000101",
  22683=>"111100001",
  22684=>"110100000",
  22685=>"000101000",
  22686=>"110010111",
  22687=>"110010001",
  22688=>"101011010",
  22689=>"010110110",
  22690=>"011001110",
  22691=>"000000110",
  22692=>"001111011",
  22693=>"100111110",
  22694=>"000111110",
  22695=>"001000011",
  22696=>"110001100",
  22697=>"110001011",
  22698=>"010010010",
  22699=>"011010111",
  22700=>"000101011",
  22701=>"111010001",
  22702=>"101011010",
  22703=>"101110100",
  22704=>"101001001",
  22705=>"101010111",
  22706=>"000111111",
  22707=>"101010000",
  22708=>"000100110",
  22709=>"010100000",
  22710=>"111010001",
  22711=>"110111110",
  22712=>"010011000",
  22713=>"100000110",
  22714=>"011110000",
  22715=>"011011100",
  22716=>"100000110",
  22717=>"010111011",
  22718=>"111101110",
  22719=>"011000101",
  22720=>"000000001",
  22721=>"010100101",
  22722=>"010110110",
  22723=>"101101110",
  22724=>"100101000",
  22725=>"100000110",
  22726=>"100111100",
  22727=>"101000111",
  22728=>"000110111",
  22729=>"100100000",
  22730=>"001000001",
  22731=>"010100110",
  22732=>"011111010",
  22733=>"111011101",
  22734=>"101011100",
  22735=>"101001110",
  22736=>"001101101",
  22737=>"001100111",
  22738=>"100100100",
  22739=>"010100101",
  22740=>"100000001",
  22741=>"000011001",
  22742=>"010001100",
  22743=>"010101101",
  22744=>"010000101",
  22745=>"000010000",
  22746=>"010010111",
  22747=>"110000100",
  22748=>"111100110",
  22749=>"100000110",
  22750=>"001000101",
  22751=>"111111000",
  22752=>"101101110",
  22753=>"001100100",
  22754=>"011111100",
  22755=>"000110000",
  22756=>"011000001",
  22757=>"111000110",
  22758=>"010111100",
  22759=>"011100101",
  22760=>"111101001",
  22761=>"100101001",
  22762=>"000001101",
  22763=>"110010010",
  22764=>"001011010",
  22765=>"000010011",
  22766=>"001001010",
  22767=>"111100000",
  22768=>"110001001",
  22769=>"011111010",
  22770=>"100101100",
  22771=>"000100000",
  22772=>"110001110",
  22773=>"110011011",
  22774=>"011000111",
  22775=>"110111001",
  22776=>"111010110",
  22777=>"000000110",
  22778=>"000110011",
  22779=>"101101000",
  22780=>"010010101",
  22781=>"111100110",
  22782=>"111110100",
  22783=>"001100110",
  22784=>"010101100",
  22785=>"100100111",
  22786=>"100111011",
  22787=>"001000000",
  22788=>"011001111",
  22789=>"010000101",
  22790=>"100001010",
  22791=>"000111000",
  22792=>"010101010",
  22793=>"000001111",
  22794=>"110101001",
  22795=>"011010101",
  22796=>"000110000",
  22797=>"011001000",
  22798=>"100001100",
  22799=>"001100001",
  22800=>"001111100",
  22801=>"000101101",
  22802=>"000111110",
  22803=>"101111001",
  22804=>"011010100",
  22805=>"011101011",
  22806=>"110110010",
  22807=>"001100110",
  22808=>"100010111",
  22809=>"010001000",
  22810=>"110001001",
  22811=>"011011110",
  22812=>"001010111",
  22813=>"110011000",
  22814=>"100110011",
  22815=>"010011001",
  22816=>"001110100",
  22817=>"100101010",
  22818=>"000001111",
  22819=>"110100000",
  22820=>"110111011",
  22821=>"111001000",
  22822=>"001111000",
  22823=>"010000001",
  22824=>"101101001",
  22825=>"110110111",
  22826=>"110101100",
  22827=>"110111110",
  22828=>"011110110",
  22829=>"101011111",
  22830=>"110100001",
  22831=>"010001011",
  22832=>"110110110",
  22833=>"001011111",
  22834=>"110000000",
  22835=>"110000001",
  22836=>"000111101",
  22837=>"000000111",
  22838=>"111011011",
  22839=>"001010110",
  22840=>"111100000",
  22841=>"100101000",
  22842=>"110100111",
  22843=>"100010000",
  22844=>"111110100",
  22845=>"111111001",
  22846=>"010111000",
  22847=>"001111110",
  22848=>"101110110",
  22849=>"111100100",
  22850=>"100011011",
  22851=>"100000010",
  22852=>"110011100",
  22853=>"000001000",
  22854=>"111010000",
  22855=>"100011101",
  22856=>"001101001",
  22857=>"100100101",
  22858=>"010010101",
  22859=>"110000100",
  22860=>"100011101",
  22861=>"100100110",
  22862=>"010100011",
  22863=>"011110100",
  22864=>"011010111",
  22865=>"111111000",
  22866=>"111011000",
  22867=>"000110110",
  22868=>"001110111",
  22869=>"011000000",
  22870=>"110101000",
  22871=>"010110010",
  22872=>"000100010",
  22873=>"111101001",
  22874=>"111110110",
  22875=>"011010111",
  22876=>"110100101",
  22877=>"001110110",
  22878=>"001000000",
  22879=>"111011111",
  22880=>"101011111",
  22881=>"000111011",
  22882=>"110000010",
  22883=>"100010000",
  22884=>"101101110",
  22885=>"000110000",
  22886=>"001100110",
  22887=>"111111100",
  22888=>"110010010",
  22889=>"110010001",
  22890=>"000111010",
  22891=>"010110111",
  22892=>"011011111",
  22893=>"001100011",
  22894=>"111011101",
  22895=>"100100011",
  22896=>"011111000",
  22897=>"111101001",
  22898=>"101000000",
  22899=>"011010100",
  22900=>"011000101",
  22901=>"000000101",
  22902=>"100001101",
  22903=>"101011001",
  22904=>"110100101",
  22905=>"000101001",
  22906=>"000001110",
  22907=>"101001011",
  22908=>"100001110",
  22909=>"011011110",
  22910=>"010100000",
  22911=>"011010001",
  22912=>"010000110",
  22913=>"110000010",
  22914=>"000111111",
  22915=>"101101000",
  22916=>"001011111",
  22917=>"100111101",
  22918=>"111111011",
  22919=>"010000010",
  22920=>"110100101",
  22921=>"101001111",
  22922=>"000101010",
  22923=>"011101110",
  22924=>"010101011",
  22925=>"001101100",
  22926=>"101010101",
  22927=>"011011111",
  22928=>"000000101",
  22929=>"001010011",
  22930=>"111101001",
  22931=>"100101110",
  22932=>"010000110",
  22933=>"100110000",
  22934=>"000100001",
  22935=>"101111010",
  22936=>"100010001",
  22937=>"000000000",
  22938=>"111000001",
  22939=>"010000100",
  22940=>"110100011",
  22941=>"000100011",
  22942=>"100001111",
  22943=>"001001001",
  22944=>"111111110",
  22945=>"010110101",
  22946=>"010111100",
  22947=>"001010000",
  22948=>"110010010",
  22949=>"110011111",
  22950=>"111010000",
  22951=>"101100100",
  22952=>"000101011",
  22953=>"111110000",
  22954=>"110101001",
  22955=>"100011110",
  22956=>"110111101",
  22957=>"011001001",
  22958=>"000100110",
  22959=>"111100110",
  22960=>"110111100",
  22961=>"000001000",
  22962=>"000010010",
  22963=>"110110100",
  22964=>"100001110",
  22965=>"111001101",
  22966=>"110000101",
  22967=>"000000001",
  22968=>"000110010",
  22969=>"101100000",
  22970=>"000100100",
  22971=>"010101000",
  22972=>"011111001",
  22973=>"110000010",
  22974=>"001101001",
  22975=>"010100011",
  22976=>"100101100",
  22977=>"001010011",
  22978=>"000111001",
  22979=>"001001001",
  22980=>"101000001",
  22981=>"001011000",
  22982=>"011100000",
  22983=>"111111010",
  22984=>"010001100",
  22985=>"001001100",
  22986=>"110011000",
  22987=>"000001001",
  22988=>"000111110",
  22989=>"011000110",
  22990=>"100000011",
  22991=>"001011001",
  22992=>"000001011",
  22993=>"110110101",
  22994=>"000111110",
  22995=>"101001010",
  22996=>"100110111",
  22997=>"100011100",
  22998=>"110000111",
  22999=>"100101001",
  23000=>"011001001",
  23001=>"100010010",
  23002=>"110000001",
  23003=>"100011010",
  23004=>"100010100",
  23005=>"101001011",
  23006=>"010001010",
  23007=>"100000110",
  23008=>"100110101",
  23009=>"001110011",
  23010=>"100001010",
  23011=>"010010110",
  23012=>"100001000",
  23013=>"101001000",
  23014=>"110000010",
  23015=>"101111100",
  23016=>"100011100",
  23017=>"101110000",
  23018=>"100110110",
  23019=>"111100110",
  23020=>"100100000",
  23021=>"000001111",
  23022=>"000111100",
  23023=>"100100010",
  23024=>"000011101",
  23025=>"101111111",
  23026=>"100110010",
  23027=>"010101110",
  23028=>"110010101",
  23029=>"100010010",
  23030=>"100000011",
  23031=>"010000111",
  23032=>"010010000",
  23033=>"111011110",
  23034=>"100000101",
  23035=>"110100101",
  23036=>"011000100",
  23037=>"111110101",
  23038=>"111011101",
  23039=>"010101110",
  23040=>"101100011",
  23041=>"111011001",
  23042=>"100111110",
  23043=>"111010000",
  23044=>"111010000",
  23045=>"000001100",
  23046=>"111110111",
  23047=>"100010111",
  23048=>"001000110",
  23049=>"110000001",
  23050=>"010011110",
  23051=>"110110000",
  23052=>"111110101",
  23053=>"111110101",
  23054=>"101100110",
  23055=>"000111011",
  23056=>"000010011",
  23057=>"011001111",
  23058=>"001001001",
  23059=>"001100010",
  23060=>"100000010",
  23061=>"101100111",
  23062=>"101111010",
  23063=>"010110010",
  23064=>"111010011",
  23065=>"110000111",
  23066=>"101011000",
  23067=>"000101010",
  23068=>"100011101",
  23069=>"111101100",
  23070=>"111101000",
  23071=>"000100010",
  23072=>"111110101",
  23073=>"110001100",
  23074=>"100001100",
  23075=>"011001001",
  23076=>"010000010",
  23077=>"001100111",
  23078=>"100101010",
  23079=>"111111010",
  23080=>"001100100",
  23081=>"110000101",
  23082=>"110100101",
  23083=>"010101010",
  23084=>"100000001",
  23085=>"001110011",
  23086=>"100000010",
  23087=>"100111000",
  23088=>"001111110",
  23089=>"011110000",
  23090=>"101101101",
  23091=>"111110111",
  23092=>"100100101",
  23093=>"110010000",
  23094=>"001011100",
  23095=>"001110100",
  23096=>"110101001",
  23097=>"100001110",
  23098=>"101001000",
  23099=>"011011110",
  23100=>"101101000",
  23101=>"011100011",
  23102=>"000100100",
  23103=>"111110101",
  23104=>"011110000",
  23105=>"001011100",
  23106=>"000010000",
  23107=>"001111100",
  23108=>"011000101",
  23109=>"101001111",
  23110=>"000100001",
  23111=>"110000111",
  23112=>"100010011",
  23113=>"010111101",
  23114=>"010011110",
  23115=>"100000100",
  23116=>"110111111",
  23117=>"010010001",
  23118=>"000011101",
  23119=>"111111101",
  23120=>"010001010",
  23121=>"000010101",
  23122=>"100110100",
  23123=>"010000101",
  23124=>"101011011",
  23125=>"000011100",
  23126=>"001110001",
  23127=>"101010100",
  23128=>"100101111",
  23129=>"100110010",
  23130=>"111000001",
  23131=>"111010101",
  23132=>"000101001",
  23133=>"110110110",
  23134=>"000001110",
  23135=>"101111000",
  23136=>"110101000",
  23137=>"010111000",
  23138=>"111010100",
  23139=>"101101111",
  23140=>"101001001",
  23141=>"111011110",
  23142=>"111000000",
  23143=>"110111110",
  23144=>"110010101",
  23145=>"011110001",
  23146=>"111011111",
  23147=>"000010000",
  23148=>"110101001",
  23149=>"110011011",
  23150=>"100011011",
  23151=>"000011010",
  23152=>"010010001",
  23153=>"001111000",
  23154=>"100010100",
  23155=>"000000100",
  23156=>"100110010",
  23157=>"011111111",
  23158=>"001010101",
  23159=>"001000100",
  23160=>"001100001",
  23161=>"001100100",
  23162=>"101111100",
  23163=>"100001100",
  23164=>"000000100",
  23165=>"001011001",
  23166=>"011011010",
  23167=>"111110010",
  23168=>"111111100",
  23169=>"101001111",
  23170=>"100110011",
  23171=>"001001001",
  23172=>"101010010",
  23173=>"110010100",
  23174=>"100100111",
  23175=>"010111100",
  23176=>"110001101",
  23177=>"010111101",
  23178=>"010000000",
  23179=>"110011000",
  23180=>"001010001",
  23181=>"111001001",
  23182=>"111101000",
  23183=>"011010110",
  23184=>"101111010",
  23185=>"101110110",
  23186=>"010111111",
  23187=>"100011110",
  23188=>"000000110",
  23189=>"110000100",
  23190=>"011111110",
  23191=>"000001111",
  23192=>"011110111",
  23193=>"111011110",
  23194=>"100100011",
  23195=>"111010101",
  23196=>"001100100",
  23197=>"001110111",
  23198=>"111100001",
  23199=>"101101010",
  23200=>"110110101",
  23201=>"110010011",
  23202=>"001100110",
  23203=>"100101101",
  23204=>"011101000",
  23205=>"100000000",
  23206=>"010111001",
  23207=>"001101000",
  23208=>"000100111",
  23209=>"011001100",
  23210=>"001001000",
  23211=>"000000101",
  23212=>"000100111",
  23213=>"111000100",
  23214=>"111011000",
  23215=>"100000000",
  23216=>"100011010",
  23217=>"011000010",
  23218=>"001001110",
  23219=>"100110010",
  23220=>"000001110",
  23221=>"110110101",
  23222=>"100011110",
  23223=>"110010000",
  23224=>"011001101",
  23225=>"101001101",
  23226=>"100100011",
  23227=>"110001010",
  23228=>"101110000",
  23229=>"000110110",
  23230=>"101111101",
  23231=>"101001010",
  23232=>"001001000",
  23233=>"000000100",
  23234=>"010010000",
  23235=>"100000111",
  23236=>"001101000",
  23237=>"000110101",
  23238=>"010111010",
  23239=>"000010011",
  23240=>"010001010",
  23241=>"010001000",
  23242=>"000001101",
  23243=>"010010011",
  23244=>"101000111",
  23245=>"001011000",
  23246=>"011101000",
  23247=>"010110001",
  23248=>"111111000",
  23249=>"110011111",
  23250=>"110100011",
  23251=>"100001110",
  23252=>"111011111",
  23253=>"010000100",
  23254=>"100010101",
  23255=>"000101100",
  23256=>"110010000",
  23257=>"111101111",
  23258=>"010010110",
  23259=>"011100101",
  23260=>"111000101",
  23261=>"101010011",
  23262=>"000100110",
  23263=>"110110111",
  23264=>"011001100",
  23265=>"111101000",
  23266=>"000111000",
  23267=>"100101001",
  23268=>"110111000",
  23269=>"011101101",
  23270=>"011100110",
  23271=>"111101110",
  23272=>"000010001",
  23273=>"111100101",
  23274=>"111000100",
  23275=>"111100010",
  23276=>"000000101",
  23277=>"101011100",
  23278=>"100001001",
  23279=>"111100111",
  23280=>"011111001",
  23281=>"101001000",
  23282=>"001010001",
  23283=>"100001111",
  23284=>"001000110",
  23285=>"110011100",
  23286=>"011001001",
  23287=>"001110110",
  23288=>"111011010",
  23289=>"010110010",
  23290=>"001000011",
  23291=>"011101110",
  23292=>"000111001",
  23293=>"010100101",
  23294=>"001110101",
  23295=>"100101110",
  23296=>"101011111",
  23297=>"001100001",
  23298=>"100010111",
  23299=>"101111011",
  23300=>"111010001",
  23301=>"010000110",
  23302=>"100011100",
  23303=>"111101111",
  23304=>"110100111",
  23305=>"010101110",
  23306=>"001100001",
  23307=>"010110101",
  23308=>"000110110",
  23309=>"011111111",
  23310=>"111001110",
  23311=>"111010111",
  23312=>"001110110",
  23313=>"000000100",
  23314=>"011101001",
  23315=>"110101001",
  23316=>"011100110",
  23317=>"100100111",
  23318=>"100000111",
  23319=>"111101010",
  23320=>"110111101",
  23321=>"001100010",
  23322=>"010101100",
  23323=>"001111100",
  23324=>"100100101",
  23325=>"011111110",
  23326=>"100110110",
  23327=>"000000111",
  23328=>"100000000",
  23329=>"000001010",
  23330=>"001010110",
  23331=>"001100011",
  23332=>"100101101",
  23333=>"111101000",
  23334=>"000010011",
  23335=>"100101010",
  23336=>"010000010",
  23337=>"011111111",
  23338=>"011110001",
  23339=>"111100000",
  23340=>"011010001",
  23341=>"110000011",
  23342=>"100011110",
  23343=>"101010111",
  23344=>"110011000",
  23345=>"110110010",
  23346=>"001001000",
  23347=>"100110100",
  23348=>"000100111",
  23349=>"111100010",
  23350=>"000101000",
  23351=>"111100011",
  23352=>"000000010",
  23353=>"101000101",
  23354=>"110100111",
  23355=>"110011000",
  23356=>"011110001",
  23357=>"000101101",
  23358=>"101010101",
  23359=>"100111101",
  23360=>"110101101",
  23361=>"100100010",
  23362=>"111101100",
  23363=>"011010001",
  23364=>"101110000",
  23365=>"111000110",
  23366=>"111010101",
  23367=>"110010010",
  23368=>"000010010",
  23369=>"010101001",
  23370=>"110100111",
  23371=>"001001111",
  23372=>"011000100",
  23373=>"001001000",
  23374=>"010000111",
  23375=>"111111001",
  23376=>"111110100",
  23377=>"010000101",
  23378=>"010101000",
  23379=>"111100001",
  23380=>"011101010",
  23381=>"111011101",
  23382=>"010110110",
  23383=>"100000001",
  23384=>"110101000",
  23385=>"001010101",
  23386=>"101010011",
  23387=>"101010011",
  23388=>"000111010",
  23389=>"101001000",
  23390=>"011110110",
  23391=>"010110000",
  23392=>"101110111",
  23393=>"011101000",
  23394=>"010101110",
  23395=>"010001001",
  23396=>"000101100",
  23397=>"010100010",
  23398=>"010101011",
  23399=>"010100111",
  23400=>"101111111",
  23401=>"110110010",
  23402=>"010110110",
  23403=>"110000000",
  23404=>"011100010",
  23405=>"101101011",
  23406=>"011101110",
  23407=>"010011111",
  23408=>"011001011",
  23409=>"011010100",
  23410=>"001001100",
  23411=>"101001011",
  23412=>"001110010",
  23413=>"100011101",
  23414=>"100110100",
  23415=>"111110011",
  23416=>"101100001",
  23417=>"100111011",
  23418=>"111000100",
  23419=>"110101111",
  23420=>"010011010",
  23421=>"001110101",
  23422=>"001000010",
  23423=>"100010100",
  23424=>"101000111",
  23425=>"101000000",
  23426=>"110010101",
  23427=>"111111101",
  23428=>"111011001",
  23429=>"111111100",
  23430=>"010110110",
  23431=>"110010000",
  23432=>"111111000",
  23433=>"001111111",
  23434=>"000011001",
  23435=>"111011110",
  23436=>"101000111",
  23437=>"100011010",
  23438=>"001110101",
  23439=>"110000000",
  23440=>"001010010",
  23441=>"110100000",
  23442=>"100111100",
  23443=>"000110110",
  23444=>"111011011",
  23445=>"000110100",
  23446=>"100101001",
  23447=>"111101100",
  23448=>"011001110",
  23449=>"111001100",
  23450=>"110001101",
  23451=>"011001111",
  23452=>"000101000",
  23453=>"010001111",
  23454=>"011111101",
  23455=>"010001101",
  23456=>"111111100",
  23457=>"000101110",
  23458=>"001011100",
  23459=>"010001011",
  23460=>"011010010",
  23461=>"110111101",
  23462=>"000010010",
  23463=>"010001111",
  23464=>"000101101",
  23465=>"110100111",
  23466=>"111000001",
  23467=>"011101110",
  23468=>"101001001",
  23469=>"000011000",
  23470=>"110010000",
  23471=>"011011010",
  23472=>"100001001",
  23473=>"001010111",
  23474=>"100000001",
  23475=>"111001111",
  23476=>"010000111",
  23477=>"101001101",
  23478=>"001000000",
  23479=>"011101100",
  23480=>"111111000",
  23481=>"001001110",
  23482=>"111010101",
  23483=>"101111011",
  23484=>"001110101",
  23485=>"100100001",
  23486=>"000110110",
  23487=>"000000011",
  23488=>"010000000",
  23489=>"000001000",
  23490=>"100110001",
  23491=>"111101100",
  23492=>"111001110",
  23493=>"101111000",
  23494=>"011000110",
  23495=>"001000001",
  23496=>"000000000",
  23497=>"100010110",
  23498=>"111000111",
  23499=>"011000011",
  23500=>"111111000",
  23501=>"010011001",
  23502=>"100000010",
  23503=>"000111011",
  23504=>"011101110",
  23505=>"100100001",
  23506=>"111010010",
  23507=>"010101010",
  23508=>"011000100",
  23509=>"011100011",
  23510=>"110100000",
  23511=>"111010001",
  23512=>"011100010",
  23513=>"101010111",
  23514=>"111110000",
  23515=>"100100010",
  23516=>"000100000",
  23517=>"111100100",
  23518=>"110011101",
  23519=>"001011100",
  23520=>"010011111",
  23521=>"100001010",
  23522=>"110101011",
  23523=>"011010100",
  23524=>"110011010",
  23525=>"101100111",
  23526=>"011100111",
  23527=>"010111100",
  23528=>"010010110",
  23529=>"001001110",
  23530=>"011010000",
  23531=>"111000000",
  23532=>"101001110",
  23533=>"110011110",
  23534=>"101100010",
  23535=>"111101110",
  23536=>"111110111",
  23537=>"011111000",
  23538=>"110110000",
  23539=>"001000010",
  23540=>"111110011",
  23541=>"000010010",
  23542=>"100100010",
  23543=>"100111001",
  23544=>"111001110",
  23545=>"111000011",
  23546=>"100000000",
  23547=>"010100010",
  23548=>"001000001",
  23549=>"011101110",
  23550=>"000001000",
  23551=>"011110000",
  23552=>"001100101",
  23553=>"011101101",
  23554=>"110101110",
  23555=>"001001100",
  23556=>"010000100",
  23557=>"001010011",
  23558=>"011111110",
  23559=>"110100011",
  23560=>"101011101",
  23561=>"000110111",
  23562=>"011001001",
  23563=>"011101111",
  23564=>"001100011",
  23565=>"001101001",
  23566=>"000000110",
  23567=>"001101010",
  23568=>"111000010",
  23569=>"110110110",
  23570=>"100010001",
  23571=>"001010000",
  23572=>"000001110",
  23573=>"011010111",
  23574=>"001000100",
  23575=>"011111100",
  23576=>"111110111",
  23577=>"001100110",
  23578=>"011010100",
  23579=>"001100000",
  23580=>"111100101",
  23581=>"110111101",
  23582=>"010101010",
  23583=>"000100010",
  23584=>"110111011",
  23585=>"100111000",
  23586=>"110000110",
  23587=>"000010110",
  23588=>"101000000",
  23589=>"111000001",
  23590=>"100000011",
  23591=>"100011011",
  23592=>"111111001",
  23593=>"010100110",
  23594=>"111101110",
  23595=>"000001100",
  23596=>"101110101",
  23597=>"100001111",
  23598=>"011101010",
  23599=>"100111010",
  23600=>"001001101",
  23601=>"111100001",
  23602=>"110100110",
  23603=>"110001101",
  23604=>"111111001",
  23605=>"110111100",
  23606=>"000000110",
  23607=>"111010000",
  23608=>"111010101",
  23609=>"111000001",
  23610=>"101111110",
  23611=>"010010101",
  23612=>"100010000",
  23613=>"000010110",
  23614=>"010111011",
  23615=>"111101111",
  23616=>"101111010",
  23617=>"110001010",
  23618=>"000010001",
  23619=>"001011110",
  23620=>"100100100",
  23621=>"001101111",
  23622=>"001101111",
  23623=>"000111001",
  23624=>"000010000",
  23625=>"000100101",
  23626=>"110101010",
  23627=>"011011001",
  23628=>"001110101",
  23629=>"001011001",
  23630=>"111010000",
  23631=>"000111110",
  23632=>"111011011",
  23633=>"101100110",
  23634=>"010001111",
  23635=>"010101011",
  23636=>"111000110",
  23637=>"011001000",
  23638=>"001111000",
  23639=>"111111110",
  23640=>"110010010",
  23641=>"001010011",
  23642=>"100100101",
  23643=>"000010101",
  23644=>"111111011",
  23645=>"010101010",
  23646=>"011110000",
  23647=>"100001000",
  23648=>"000000010",
  23649=>"010000000",
  23650=>"101101000",
  23651=>"000011011",
  23652=>"000100100",
  23653=>"000100000",
  23654=>"011001101",
  23655=>"111001110",
  23656=>"001010001",
  23657=>"010100110",
  23658=>"101111000",
  23659=>"001100000",
  23660=>"111011100",
  23661=>"111011011",
  23662=>"111001111",
  23663=>"000110111",
  23664=>"000001101",
  23665=>"010010110",
  23666=>"101111001",
  23667=>"000000000",
  23668=>"001010010",
  23669=>"111100100",
  23670=>"011100000",
  23671=>"010101110",
  23672=>"011011101",
  23673=>"100110010",
  23674=>"011101010",
  23675=>"111111110",
  23676=>"011001011",
  23677=>"011111111",
  23678=>"101111111",
  23679=>"110111011",
  23680=>"101111111",
  23681=>"101000110",
  23682=>"101011011",
  23683=>"011101001",
  23684=>"011111111",
  23685=>"111100110",
  23686=>"101001100",
  23687=>"100100000",
  23688=>"110110001",
  23689=>"111001001",
  23690=>"100010100",
  23691=>"100100100",
  23692=>"111110011",
  23693=>"101111111",
  23694=>"000111111",
  23695=>"010001100",
  23696=>"000110110",
  23697=>"111010100",
  23698=>"000000001",
  23699=>"101000001",
  23700=>"000100010",
  23701=>"110010111",
  23702=>"101100001",
  23703=>"010100001",
  23704=>"111110010",
  23705=>"101000010",
  23706=>"011111010",
  23707=>"000111111",
  23708=>"100111110",
  23709=>"111001100",
  23710=>"000010100",
  23711=>"011110011",
  23712=>"001000101",
  23713=>"000110111",
  23714=>"010010011",
  23715=>"010010110",
  23716=>"011000011",
  23717=>"111100100",
  23718=>"111001001",
  23719=>"001101111",
  23720=>"101110000",
  23721=>"110101100",
  23722=>"110111111",
  23723=>"011101000",
  23724=>"000101101",
  23725=>"100111011",
  23726=>"101101000",
  23727=>"100001011",
  23728=>"111010101",
  23729=>"000011000",
  23730=>"011010110",
  23731=>"000000010",
  23732=>"000011101",
  23733=>"100011011",
  23734=>"000010011",
  23735=>"100001111",
  23736=>"101100001",
  23737=>"100001111",
  23738=>"101101000",
  23739=>"000101111",
  23740=>"111110001",
  23741=>"010111101",
  23742=>"110010000",
  23743=>"110111111",
  23744=>"111000000",
  23745=>"010101101",
  23746=>"011101011",
  23747=>"001110101",
  23748=>"100110111",
  23749=>"001111111",
  23750=>"111110001",
  23751=>"111101100",
  23752=>"111010111",
  23753=>"010111110",
  23754=>"010001000",
  23755=>"100001101",
  23756=>"101001110",
  23757=>"101100100",
  23758=>"111111100",
  23759=>"110010001",
  23760=>"001110000",
  23761=>"111001111",
  23762=>"111111111",
  23763=>"011001111",
  23764=>"001010101",
  23765=>"110000100",
  23766=>"101110101",
  23767=>"101101001",
  23768=>"111101000",
  23769=>"100111000",
  23770=>"100011111",
  23771=>"000101111",
  23772=>"011011101",
  23773=>"101101111",
  23774=>"000101100",
  23775=>"010011101",
  23776=>"111000000",
  23777=>"001110101",
  23778=>"000110111",
  23779=>"101000111",
  23780=>"001001010",
  23781=>"110001110",
  23782=>"111010011",
  23783=>"111101000",
  23784=>"011011011",
  23785=>"101111111",
  23786=>"000000111",
  23787=>"110111100",
  23788=>"011011010",
  23789=>"000000011",
  23790=>"111000001",
  23791=>"010000011",
  23792=>"001100111",
  23793=>"111010110",
  23794=>"010110101",
  23795=>"100100011",
  23796=>"111100111",
  23797=>"111110111",
  23798=>"111111000",
  23799=>"110010000",
  23800=>"010101001",
  23801=>"000001100",
  23802=>"101011011",
  23803=>"001111111",
  23804=>"111000100",
  23805=>"000111100",
  23806=>"000111100",
  23807=>"000001000",
  23808=>"100110010",
  23809=>"100011011",
  23810=>"001110110",
  23811=>"111111000",
  23812=>"110010110",
  23813=>"011110111",
  23814=>"100001110",
  23815=>"100010011",
  23816=>"100111101",
  23817=>"000001101",
  23818=>"001010101",
  23819=>"101100111",
  23820=>"001010100",
  23821=>"001001001",
  23822=>"101100010",
  23823=>"000100110",
  23824=>"111001110",
  23825=>"101011000",
  23826=>"110000010",
  23827=>"110111001",
  23828=>"011001110",
  23829=>"011101001",
  23830=>"110110100",
  23831=>"010011110",
  23832=>"000010001",
  23833=>"110000001",
  23834=>"010101010",
  23835=>"001000111",
  23836=>"000010011",
  23837=>"001001100",
  23838=>"001011010",
  23839=>"100110010",
  23840=>"111000000",
  23841=>"010001110",
  23842=>"010011100",
  23843=>"111101110",
  23844=>"100001101",
  23845=>"100000010",
  23846=>"100100011",
  23847=>"100001011",
  23848=>"010010111",
  23849=>"101011100",
  23850=>"111111011",
  23851=>"011001101",
  23852=>"111011111",
  23853=>"101100010",
  23854=>"011011111",
  23855=>"000011101",
  23856=>"010111000",
  23857=>"110110101",
  23858=>"011000100",
  23859=>"010010110",
  23860=>"001100010",
  23861=>"010001110",
  23862=>"100110010",
  23863=>"000101011",
  23864=>"010100101",
  23865=>"111111011",
  23866=>"011110000",
  23867=>"110011001",
  23868=>"010010101",
  23869=>"000011011",
  23870=>"111111100",
  23871=>"111111100",
  23872=>"110101110",
  23873=>"101011000",
  23874=>"101110000",
  23875=>"011000011",
  23876=>"011110001",
  23877=>"001101101",
  23878=>"110011010",
  23879=>"100101111",
  23880=>"111010110",
  23881=>"001000100",
  23882=>"011010010",
  23883=>"001000010",
  23884=>"100001111",
  23885=>"000000100",
  23886=>"111000111",
  23887=>"001000001",
  23888=>"000100001",
  23889=>"000011011",
  23890=>"111100000",
  23891=>"111001100",
  23892=>"000010000",
  23893=>"001001011",
  23894=>"001100111",
  23895=>"110101101",
  23896=>"011010010",
  23897=>"111100010",
  23898=>"111111011",
  23899=>"001000110",
  23900=>"000001010",
  23901=>"000111101",
  23902=>"000110111",
  23903=>"010011000",
  23904=>"001010010",
  23905=>"001100101",
  23906=>"000000010",
  23907=>"010001011",
  23908=>"010111000",
  23909=>"101000101",
  23910=>"010000110",
  23911=>"111011111",
  23912=>"000000110",
  23913=>"000010111",
  23914=>"101001101",
  23915=>"110111101",
  23916=>"011000111",
  23917=>"001100100",
  23918=>"001000010",
  23919=>"100110010",
  23920=>"011000100",
  23921=>"011000100",
  23922=>"011011111",
  23923=>"000010100",
  23924=>"011100001",
  23925=>"001011010",
  23926=>"001010010",
  23927=>"010100010",
  23928=>"111111001",
  23929=>"101101011",
  23930=>"111101011",
  23931=>"000011110",
  23932=>"111000101",
  23933=>"110010110",
  23934=>"111111100",
  23935=>"110011000",
  23936=>"001111111",
  23937=>"010100001",
  23938=>"101011001",
  23939=>"001101111",
  23940=>"010110000",
  23941=>"001001000",
  23942=>"010001101",
  23943=>"111010010",
  23944=>"101110000",
  23945=>"011111011",
  23946=>"110111001",
  23947=>"100011000",
  23948=>"011100011",
  23949=>"111101100",
  23950=>"111110101",
  23951=>"100000000",
  23952=>"101101011",
  23953=>"011111100",
  23954=>"100111010",
  23955=>"000000110",
  23956=>"000100100",
  23957=>"011101011",
  23958=>"110100100",
  23959=>"011000000",
  23960=>"011110001",
  23961=>"000100111",
  23962=>"101111101",
  23963=>"101000000",
  23964=>"011101011",
  23965=>"111100010",
  23966=>"010001110",
  23967=>"001001101",
  23968=>"111100110",
  23969=>"010111010",
  23970=>"111010001",
  23971=>"101101110",
  23972=>"101000101",
  23973=>"100010111",
  23974=>"100000010",
  23975=>"000000111",
  23976=>"001100000",
  23977=>"110010100",
  23978=>"000100111",
  23979=>"010111111",
  23980=>"110101111",
  23981=>"110011000",
  23982=>"100111100",
  23983=>"100010000",
  23984=>"000011100",
  23985=>"001111100",
  23986=>"111011111",
  23987=>"100000100",
  23988=>"101001110",
  23989=>"110010101",
  23990=>"111010100",
  23991=>"101011010",
  23992=>"100001000",
  23993=>"010100010",
  23994=>"000100101",
  23995=>"001000100",
  23996=>"001111011",
  23997=>"100111001",
  23998=>"011000000",
  23999=>"001110000",
  24000=>"001101001",
  24001=>"101010001",
  24002=>"001110111",
  24003=>"000000000",
  24004=>"111101000",
  24005=>"111010001",
  24006=>"010100010",
  24007=>"111011101",
  24008=>"110011110",
  24009=>"110110110",
  24010=>"000010111",
  24011=>"111001101",
  24012=>"000000111",
  24013=>"111001000",
  24014=>"000010110",
  24015=>"101011111",
  24016=>"111000001",
  24017=>"001010111",
  24018=>"010001110",
  24019=>"110101011",
  24020=>"100001010",
  24021=>"011110101",
  24022=>"000111100",
  24023=>"011011001",
  24024=>"111010110",
  24025=>"000110000",
  24026=>"001010010",
  24027=>"100101111",
  24028=>"011011000",
  24029=>"111100100",
  24030=>"000001101",
  24031=>"010111001",
  24032=>"010110101",
  24033=>"111010000",
  24034=>"111010110",
  24035=>"100000110",
  24036=>"001001000",
  24037=>"011100110",
  24038=>"010110101",
  24039=>"001000010",
  24040=>"110001110",
  24041=>"010000011",
  24042=>"110111100",
  24043=>"111011101",
  24044=>"011001100",
  24045=>"110111111",
  24046=>"111110000",
  24047=>"010010100",
  24048=>"011101100",
  24049=>"101011000",
  24050=>"011001100",
  24051=>"111101110",
  24052=>"010100001",
  24053=>"100110010",
  24054=>"001110011",
  24055=>"111010100",
  24056=>"010011001",
  24057=>"100010100",
  24058=>"000110001",
  24059=>"100000111",
  24060=>"101011010",
  24061=>"110011110",
  24062=>"101111101",
  24063=>"111111111",
  24064=>"001110110",
  24065=>"111001011",
  24066=>"111111001",
  24067=>"110110000",
  24068=>"000010001",
  24069=>"110001010",
  24070=>"001100111",
  24071=>"010000000",
  24072=>"100000111",
  24073=>"000100001",
  24074=>"111000100",
  24075=>"101011100",
  24076=>"011000001",
  24077=>"111000000",
  24078=>"101101111",
  24079=>"100101100",
  24080=>"100101010",
  24081=>"111001110",
  24082=>"111101101",
  24083=>"111111000",
  24084=>"011001100",
  24085=>"110110001",
  24086=>"011110010",
  24087=>"011000000",
  24088=>"101011110",
  24089=>"110000010",
  24090=>"111001101",
  24091=>"000111000",
  24092=>"101001001",
  24093=>"110010111",
  24094=>"101111101",
  24095=>"101100101",
  24096=>"111101100",
  24097=>"001100011",
  24098=>"011000000",
  24099=>"111101010",
  24100=>"111100111",
  24101=>"110011110",
  24102=>"001010001",
  24103=>"010110110",
  24104=>"000111011",
  24105=>"011011101",
  24106=>"111010110",
  24107=>"100011000",
  24108=>"011011110",
  24109=>"000101101",
  24110=>"001000101",
  24111=>"110111001",
  24112=>"110101001",
  24113=>"000000110",
  24114=>"001100010",
  24115=>"010110111",
  24116=>"100100111",
  24117=>"011010010",
  24118=>"010101110",
  24119=>"011111100",
  24120=>"001001110",
  24121=>"011101111",
  24122=>"101011111",
  24123=>"101010011",
  24124=>"110010101",
  24125=>"000101111",
  24126=>"011100001",
  24127=>"011110011",
  24128=>"100000100",
  24129=>"111011101",
  24130=>"111111010",
  24131=>"001011011",
  24132=>"001000000",
  24133=>"010011111",
  24134=>"111101111",
  24135=>"110100000",
  24136=>"011001011",
  24137=>"010000110",
  24138=>"001111111",
  24139=>"100001100",
  24140=>"111100101",
  24141=>"010111000",
  24142=>"101011111",
  24143=>"000101010",
  24144=>"000011101",
  24145=>"000010001",
  24146=>"110101010",
  24147=>"101011000",
  24148=>"110010101",
  24149=>"100100011",
  24150=>"110010110",
  24151=>"000110011",
  24152=>"100000111",
  24153=>"011111011",
  24154=>"111001111",
  24155=>"100110110",
  24156=>"000010111",
  24157=>"111111011",
  24158=>"101011100",
  24159=>"110000101",
  24160=>"010000111",
  24161=>"100110111",
  24162=>"011111100",
  24163=>"110100010",
  24164=>"000011010",
  24165=>"001001010",
  24166=>"111100000",
  24167=>"111011001",
  24168=>"100010010",
  24169=>"110111010",
  24170=>"000011011",
  24171=>"001100101",
  24172=>"111011000",
  24173=>"110110001",
  24174=>"101100010",
  24175=>"100101101",
  24176=>"111000001",
  24177=>"001001011",
  24178=>"001111100",
  24179=>"111010010",
  24180=>"000000111",
  24181=>"110110011",
  24182=>"001001000",
  24183=>"010101101",
  24184=>"000110010",
  24185=>"000100111",
  24186=>"001001011",
  24187=>"110111110",
  24188=>"010000101",
  24189=>"110011011",
  24190=>"010111101",
  24191=>"000100100",
  24192=>"110010101",
  24193=>"010110001",
  24194=>"100110101",
  24195=>"111011011",
  24196=>"101100000",
  24197=>"001000111",
  24198=>"100001000",
  24199=>"111110001",
  24200=>"011010010",
  24201=>"000010001",
  24202=>"100010000",
  24203=>"111010001",
  24204=>"100111011",
  24205=>"111111011",
  24206=>"000010000",
  24207=>"001111110",
  24208=>"011000100",
  24209=>"100110110",
  24210=>"000000100",
  24211=>"011100100",
  24212=>"000100111",
  24213=>"111111001",
  24214=>"000011000",
  24215=>"111011011",
  24216=>"001000100",
  24217=>"101111111",
  24218=>"110111011",
  24219=>"010100010",
  24220=>"111101110",
  24221=>"011110111",
  24222=>"001110000",
  24223=>"000111111",
  24224=>"001101000",
  24225=>"011000101",
  24226=>"001000111",
  24227=>"011001000",
  24228=>"100111100",
  24229=>"110111110",
  24230=>"110111000",
  24231=>"111000000",
  24232=>"010010110",
  24233=>"101110100",
  24234=>"110011111",
  24235=>"111101001",
  24236=>"000111011",
  24237=>"010111010",
  24238=>"110101101",
  24239=>"111011111",
  24240=>"110100111",
  24241=>"000101110",
  24242=>"100110000",
  24243=>"100100010",
  24244=>"000110011",
  24245=>"001110010",
  24246=>"010101011",
  24247=>"010101100",
  24248=>"001101011",
  24249=>"010001010",
  24250=>"111001110",
  24251=>"100010101",
  24252=>"111110111",
  24253=>"010000011",
  24254=>"011000001",
  24255=>"110010101",
  24256=>"111010101",
  24257=>"010011011",
  24258=>"001011001",
  24259=>"111100010",
  24260=>"011001001",
  24261=>"000101101",
  24262=>"111000111",
  24263=>"100010010",
  24264=>"101010110",
  24265=>"010000000",
  24266=>"000001100",
  24267=>"111101100",
  24268=>"000111011",
  24269=>"100101011",
  24270=>"101100101",
  24271=>"110100101",
  24272=>"111101110",
  24273=>"001101111",
  24274=>"110101101",
  24275=>"111100010",
  24276=>"110110000",
  24277=>"010010010",
  24278=>"100010100",
  24279=>"000101100",
  24280=>"001101001",
  24281=>"000101010",
  24282=>"001001100",
  24283=>"010000000",
  24284=>"100010010",
  24285=>"111110111",
  24286=>"101111011",
  24287=>"000001110",
  24288=>"101010010",
  24289=>"001010110",
  24290=>"110010100",
  24291=>"010010011",
  24292=>"110001001",
  24293=>"000011101",
  24294=>"111100001",
  24295=>"011110000",
  24296=>"111011001",
  24297=>"010111101",
  24298=>"010010110",
  24299=>"100111010",
  24300=>"001010010",
  24301=>"001111010",
  24302=>"101100010",
  24303=>"101010100",
  24304=>"101100101",
  24305=>"011011011",
  24306=>"011011110",
  24307=>"101100101",
  24308=>"111111100",
  24309=>"011101011",
  24310=>"100000001",
  24311=>"011001101",
  24312=>"010011001",
  24313=>"000101101",
  24314=>"000011100",
  24315=>"110000001",
  24316=>"011110010",
  24317=>"001010010",
  24318=>"110000110",
  24319=>"101111101",
  24320=>"000110110",
  24321=>"111010000",
  24322=>"111100010",
  24323=>"011111110",
  24324=>"000000001",
  24325=>"111100111",
  24326=>"111110011",
  24327=>"111010000",
  24328=>"101010011",
  24329=>"100010000",
  24330=>"011011110",
  24331=>"101010100",
  24332=>"011101011",
  24333=>"010001000",
  24334=>"110011111",
  24335=>"111110000",
  24336=>"011001001",
  24337=>"001101101",
  24338=>"010010110",
  24339=>"001101011",
  24340=>"111010011",
  24341=>"100010110",
  24342=>"111001110",
  24343=>"001101100",
  24344=>"100001111",
  24345=>"111000100",
  24346=>"100101001",
  24347=>"010011001",
  24348=>"101010101",
  24349=>"010000001",
  24350=>"111010000",
  24351=>"000111101",
  24352=>"101100101",
  24353=>"110001001",
  24354=>"011011111",
  24355=>"100101011",
  24356=>"100100110",
  24357=>"110011110",
  24358=>"111111000",
  24359=>"111111100",
  24360=>"001010000",
  24361=>"001011010",
  24362=>"011011110",
  24363=>"110101100",
  24364=>"011011000",
  24365=>"000101000",
  24366=>"101011111",
  24367=>"000011011",
  24368=>"100000011",
  24369=>"100100100",
  24370=>"110011000",
  24371=>"100100100",
  24372=>"001100000",
  24373=>"110100101",
  24374=>"101100100",
  24375=>"011001000",
  24376=>"000010111",
  24377=>"111100010",
  24378=>"110110001",
  24379=>"001001011",
  24380=>"000101001",
  24381=>"110010100",
  24382=>"010100000",
  24383=>"011000010",
  24384=>"000111011",
  24385=>"100110010",
  24386=>"000110110",
  24387=>"101000011",
  24388=>"000101011",
  24389=>"001000111",
  24390=>"111111111",
  24391=>"000111010",
  24392=>"010110100",
  24393=>"110011111",
  24394=>"000011101",
  24395=>"110100111",
  24396=>"101001110",
  24397=>"111010101",
  24398=>"010010110",
  24399=>"001000000",
  24400=>"001010111",
  24401=>"111100100",
  24402=>"110000111",
  24403=>"000000000",
  24404=>"100001110",
  24405=>"000000001",
  24406=>"000111101",
  24407=>"000001001",
  24408=>"010010101",
  24409=>"010011110",
  24410=>"010011101",
  24411=>"011100000",
  24412=>"001100100",
  24413=>"101111100",
  24414=>"011011000",
  24415=>"111010011",
  24416=>"110111110",
  24417=>"010011111",
  24418=>"111110100",
  24419=>"101000000",
  24420=>"011000111",
  24421=>"100001000",
  24422=>"111100110",
  24423=>"000010011",
  24424=>"111000011",
  24425=>"011100101",
  24426=>"110001010",
  24427=>"110001010",
  24428=>"000110111",
  24429=>"101111101",
  24430=>"110110001",
  24431=>"001111111",
  24432=>"100000010",
  24433=>"111101101",
  24434=>"001100011",
  24435=>"110100010",
  24436=>"000101011",
  24437=>"011110111",
  24438=>"010110101",
  24439=>"001111100",
  24440=>"010011011",
  24441=>"010110111",
  24442=>"101110000",
  24443=>"001101101",
  24444=>"000010000",
  24445=>"111000010",
  24446=>"101101111",
  24447=>"010111010",
  24448=>"100111101",
  24449=>"011010111",
  24450=>"011000001",
  24451=>"001100010",
  24452=>"111011101",
  24453=>"000010111",
  24454=>"000111100",
  24455=>"100000100",
  24456=>"000010101",
  24457=>"111010001",
  24458=>"001010100",
  24459=>"011000100",
  24460=>"110100101",
  24461=>"101001001",
  24462=>"101001011",
  24463=>"000110010",
  24464=>"101111101",
  24465=>"110010110",
  24466=>"111001111",
  24467=>"010110010",
  24468=>"001011000",
  24469=>"001111010",
  24470=>"001111000",
  24471=>"110011010",
  24472=>"100011100",
  24473=>"111100100",
  24474=>"011100110",
  24475=>"000000100",
  24476=>"000111011",
  24477=>"001111000",
  24478=>"100111111",
  24479=>"100010110",
  24480=>"111100101",
  24481=>"100110010",
  24482=>"111101100",
  24483=>"000010010",
  24484=>"111011001",
  24485=>"111110100",
  24486=>"010101100",
  24487=>"111100101",
  24488=>"100111000",
  24489=>"010010100",
  24490=>"101000010",
  24491=>"010011001",
  24492=>"101100000",
  24493=>"001010111",
  24494=>"010110011",
  24495=>"111011110",
  24496=>"110110111",
  24497=>"110110111",
  24498=>"011111110",
  24499=>"110111111",
  24500=>"001100011",
  24501=>"110011010",
  24502=>"110101111",
  24503=>"110111011",
  24504=>"101100111",
  24505=>"011110100",
  24506=>"000111001",
  24507=>"101000110",
  24508=>"101101001",
  24509=>"110100010",
  24510=>"011111110",
  24511=>"100011010",
  24512=>"110110100",
  24513=>"011011110",
  24514=>"101100010",
  24515=>"011011110",
  24516=>"101111100",
  24517=>"011111101",
  24518=>"001010101",
  24519=>"010101000",
  24520=>"101011010",
  24521=>"100111011",
  24522=>"000010000",
  24523=>"011111001",
  24524=>"100111011",
  24525=>"111011111",
  24526=>"010010100",
  24527=>"110110110",
  24528=>"011000101",
  24529=>"011000101",
  24530=>"000000000",
  24531=>"100000101",
  24532=>"000100010",
  24533=>"000011101",
  24534=>"111011010",
  24535=>"011001000",
  24536=>"110101001",
  24537=>"000011101",
  24538=>"111111011",
  24539=>"000110100",
  24540=>"001001000",
  24541=>"011100001",
  24542=>"101101000",
  24543=>"000011111",
  24544=>"100010101",
  24545=>"000010100",
  24546=>"110110111",
  24547=>"011001010",
  24548=>"111100111",
  24549=>"100010001",
  24550=>"101111010",
  24551=>"101000111",
  24552=>"100000001",
  24553=>"010000000",
  24554=>"111111100",
  24555=>"101111111",
  24556=>"000011011",
  24557=>"110111010",
  24558=>"000000110",
  24559=>"110110111",
  24560=>"110100101",
  24561=>"100111000",
  24562=>"100101011",
  24563=>"011010101",
  24564=>"001010100",
  24565=>"010111111",
  24566=>"011111010",
  24567=>"111111000",
  24568=>"111101000",
  24569=>"011000110",
  24570=>"000110000",
  24571=>"100000100",
  24572=>"111111111",
  24573=>"011101111",
  24574=>"001011110",
  24575=>"111100110",
  24576=>"101001101",
  24577=>"100001110",
  24578=>"000011011",
  24579=>"001010011",
  24580=>"110000100",
  24581=>"011101111",
  24582=>"011000000",
  24583=>"000111001",
  24584=>"011011100",
  24585=>"100111111",
  24586=>"001011100",
  24587=>"001100011",
  24588=>"110010001",
  24589=>"010111100",
  24590=>"111001100",
  24591=>"110111100",
  24592=>"111110010",
  24593=>"111011110",
  24594=>"000100111",
  24595=>"101100011",
  24596=>"010010100",
  24597=>"010101111",
  24598=>"011100000",
  24599=>"100110010",
  24600=>"110001010",
  24601=>"100001000",
  24602=>"110110100",
  24603=>"000001100",
  24604=>"011000011",
  24605=>"011001110",
  24606=>"110011000",
  24607=>"000011110",
  24608=>"001101111",
  24609=>"001001100",
  24610=>"111110101",
  24611=>"111101010",
  24612=>"001100110",
  24613=>"010111101",
  24614=>"111001011",
  24615=>"000001000",
  24616=>"001100101",
  24617=>"100110010",
  24618=>"101101010",
  24619=>"110101010",
  24620=>"011010000",
  24621=>"110010100",
  24622=>"001011111",
  24623=>"001001000",
  24624=>"101100001",
  24625=>"001111001",
  24626=>"100100111",
  24627=>"001110111",
  24628=>"111101011",
  24629=>"001101010",
  24630=>"000110011",
  24631=>"100100110",
  24632=>"101000000",
  24633=>"100111111",
  24634=>"000111010",
  24635=>"010100110",
  24636=>"111111111",
  24637=>"100001101",
  24638=>"100011000",
  24639=>"000011010",
  24640=>"011010101",
  24641=>"001000111",
  24642=>"000100000",
  24643=>"111011000",
  24644=>"111000110",
  24645=>"101111011",
  24646=>"010011011",
  24647=>"101010001",
  24648=>"010110111",
  24649=>"111111101",
  24650=>"000101111",
  24651=>"011101001",
  24652=>"110111101",
  24653=>"110000101",
  24654=>"010111010",
  24655=>"000110101",
  24656=>"101111100",
  24657=>"110000100",
  24658=>"010110111",
  24659=>"011100111",
  24660=>"110101110",
  24661=>"010010000",
  24662=>"101100101",
  24663=>"101111000",
  24664=>"100001110",
  24665=>"101100110",
  24666=>"101011100",
  24667=>"111101010",
  24668=>"010100101",
  24669=>"110001011",
  24670=>"011101000",
  24671=>"001000010",
  24672=>"101100101",
  24673=>"101000010",
  24674=>"000001101",
  24675=>"011111000",
  24676=>"100100011",
  24677=>"111111111",
  24678=>"000010000",
  24679=>"001100110",
  24680=>"001011110",
  24681=>"110101110",
  24682=>"010101010",
  24683=>"001010110",
  24684=>"111100011",
  24685=>"111101011",
  24686=>"101111110",
  24687=>"000000001",
  24688=>"101010110",
  24689=>"010010111",
  24690=>"010001111",
  24691=>"110110011",
  24692=>"011100100",
  24693=>"100110110",
  24694=>"100100111",
  24695=>"111100101",
  24696=>"010110011",
  24697=>"011001000",
  24698=>"010010110",
  24699=>"000100100",
  24700=>"000011111",
  24701=>"111101011",
  24702=>"000110011",
  24703=>"111001001",
  24704=>"110110111",
  24705=>"110010000",
  24706=>"001001101",
  24707=>"110000101",
  24708=>"011100000",
  24709=>"001010000",
  24710=>"001011001",
  24711=>"101101101",
  24712=>"101010100",
  24713=>"001111101",
  24714=>"001000010",
  24715=>"110111111",
  24716=>"110010001",
  24717=>"010011001",
  24718=>"000000110",
  24719=>"111010110",
  24720=>"101100100",
  24721=>"000101011",
  24722=>"110100000",
  24723=>"111011001",
  24724=>"101110010",
  24725=>"000011010",
  24726=>"100100101",
  24727=>"000011111",
  24728=>"000000000",
  24729=>"011001100",
  24730=>"100101111",
  24731=>"000111010",
  24732=>"000010001",
  24733=>"011011111",
  24734=>"011101010",
  24735=>"111100010",
  24736=>"010110110",
  24737=>"101001001",
  24738=>"100100010",
  24739=>"001001100",
  24740=>"000001101",
  24741=>"101010110",
  24742=>"100000100",
  24743=>"101100000",
  24744=>"100111111",
  24745=>"000110110",
  24746=>"011000000",
  24747=>"011100111",
  24748=>"001011011",
  24749=>"010110100",
  24750=>"111010100",
  24751=>"100110010",
  24752=>"110001101",
  24753=>"100011011",
  24754=>"010110100",
  24755=>"001100101",
  24756=>"000010100",
  24757=>"001001000",
  24758=>"000101011",
  24759=>"110100010",
  24760=>"000011010",
  24761=>"100011000",
  24762=>"010011110",
  24763=>"111100000",
  24764=>"110100011",
  24765=>"000000010",
  24766=>"001001011",
  24767=>"100111110",
  24768=>"101101001",
  24769=>"000001011",
  24770=>"011101001",
  24771=>"111011111",
  24772=>"111010111",
  24773=>"010000000",
  24774=>"000100001",
  24775=>"010111101",
  24776=>"011011111",
  24777=>"100011111",
  24778=>"011011010",
  24779=>"010010111",
  24780=>"001100010",
  24781=>"101111111",
  24782=>"000101011",
  24783=>"111010010",
  24784=>"011110101",
  24785=>"001101100",
  24786=>"110001111",
  24787=>"101010010",
  24788=>"101001110",
  24789=>"010000000",
  24790=>"000000011",
  24791=>"110100011",
  24792=>"000010100",
  24793=>"111110111",
  24794=>"000110011",
  24795=>"111011100",
  24796=>"110111111",
  24797=>"100111011",
  24798=>"110000000",
  24799=>"010010111",
  24800=>"000101010",
  24801=>"011100100",
  24802=>"010011111",
  24803=>"000010011",
  24804=>"100000110",
  24805=>"010010101",
  24806=>"111000100",
  24807=>"011010000",
  24808=>"010100010",
  24809=>"110101010",
  24810=>"001111110",
  24811=>"100010111",
  24812=>"110111011",
  24813=>"010001110",
  24814=>"000111001",
  24815=>"110101001",
  24816=>"100101011",
  24817=>"100010000",
  24818=>"100010111",
  24819=>"011110110",
  24820=>"010010000",
  24821=>"111001100",
  24822=>"010100010",
  24823=>"111011010",
  24824=>"100101010",
  24825=>"100010111",
  24826=>"000010111",
  24827=>"011100100",
  24828=>"101100010",
  24829=>"101001110",
  24830=>"110101111",
  24831=>"000110100",
  24832=>"010100000",
  24833=>"001111111",
  24834=>"100011111",
  24835=>"000110100",
  24836=>"010000000",
  24837=>"111010101",
  24838=>"000011001",
  24839=>"100000110",
  24840=>"111011010",
  24841=>"010000101",
  24842=>"000001100",
  24843=>"111101000",
  24844=>"011011111",
  24845=>"100111001",
  24846=>"010001011",
  24847=>"100011111",
  24848=>"011000001",
  24849=>"110011101",
  24850=>"001111001",
  24851=>"010101100",
  24852=>"000100110",
  24853=>"000110110",
  24854=>"010000001",
  24855=>"101000110",
  24856=>"110011111",
  24857=>"100000010",
  24858=>"110011010",
  24859=>"110011011",
  24860=>"100000001",
  24861=>"010110111",
  24862=>"101100000",
  24863=>"101010100",
  24864=>"000000001",
  24865=>"110110110",
  24866=>"010001011",
  24867=>"001111011",
  24868=>"011001000",
  24869=>"111010101",
  24870=>"011001111",
  24871=>"101010110",
  24872=>"000100000",
  24873=>"100100010",
  24874=>"010000110",
  24875=>"110001111",
  24876=>"000010111",
  24877=>"101110011",
  24878=>"010100110",
  24879=>"000000010",
  24880=>"110101000",
  24881=>"001000101",
  24882=>"111010011",
  24883=>"110011001",
  24884=>"100110111",
  24885=>"001001100",
  24886=>"011000010",
  24887=>"100101000",
  24888=>"000100111",
  24889=>"011011110",
  24890=>"010111111",
  24891=>"010110111",
  24892=>"001100110",
  24893=>"011001100",
  24894=>"111101100",
  24895=>"000011100",
  24896=>"001101100",
  24897=>"110100111",
  24898=>"011111110",
  24899=>"011001100",
  24900=>"100111001",
  24901=>"010001110",
  24902=>"110000111",
  24903=>"000010001",
  24904=>"010000100",
  24905=>"010010110",
  24906=>"100001111",
  24907=>"100111011",
  24908=>"011101100",
  24909=>"111000101",
  24910=>"000100001",
  24911=>"001000101",
  24912=>"110011000",
  24913=>"010101000",
  24914=>"100101000",
  24915=>"110100100",
  24916=>"000100000",
  24917=>"010001110",
  24918=>"101110000",
  24919=>"010101101",
  24920=>"000001010",
  24921=>"011001101",
  24922=>"111111110",
  24923=>"010011010",
  24924=>"100101110",
  24925=>"000100100",
  24926=>"011100001",
  24927=>"000001110",
  24928=>"101110110",
  24929=>"100100110",
  24930=>"100001001",
  24931=>"011000001",
  24932=>"110001101",
  24933=>"101000111",
  24934=>"011010001",
  24935=>"111001101",
  24936=>"010010110",
  24937=>"000111000",
  24938=>"101000010",
  24939=>"100110110",
  24940=>"011100111",
  24941=>"101110011",
  24942=>"000111001",
  24943=>"001100000",
  24944=>"000000101",
  24945=>"111001010",
  24946=>"010100001",
  24947=>"101010011",
  24948=>"011000011",
  24949=>"000100100",
  24950=>"000101101",
  24951=>"101000011",
  24952=>"100101101",
  24953=>"100001100",
  24954=>"101000110",
  24955=>"111011110",
  24956=>"100110001",
  24957=>"011100110",
  24958=>"111101111",
  24959=>"100100101",
  24960=>"001111100",
  24961=>"101010011",
  24962=>"000000011",
  24963=>"111111010",
  24964=>"111010110",
  24965=>"001100000",
  24966=>"100001011",
  24967=>"100000001",
  24968=>"000100101",
  24969=>"101000000",
  24970=>"000000111",
  24971=>"100001100",
  24972=>"011101010",
  24973=>"100111010",
  24974=>"110100011",
  24975=>"100111000",
  24976=>"011000101",
  24977=>"101000011",
  24978=>"000000001",
  24979=>"110001110",
  24980=>"001001100",
  24981=>"001100101",
  24982=>"111111001",
  24983=>"110111010",
  24984=>"011010100",
  24985=>"011100100",
  24986=>"111100001",
  24987=>"101010101",
  24988=>"001100101",
  24989=>"001011100",
  24990=>"100101110",
  24991=>"101101101",
  24992=>"011111101",
  24993=>"111111010",
  24994=>"100001100",
  24995=>"011110110",
  24996=>"111000100",
  24997=>"111110011",
  24998=>"001000001",
  24999=>"111000111",
  25000=>"010000000",
  25001=>"000101001",
  25002=>"000111000",
  25003=>"001010001",
  25004=>"100111000",
  25005=>"010001011",
  25006=>"100000110",
  25007=>"010011010",
  25008=>"101001110",
  25009=>"010100110",
  25010=>"110100101",
  25011=>"101111011",
  25012=>"010011111",
  25013=>"110000010",
  25014=>"000010100",
  25015=>"010111000",
  25016=>"010101110",
  25017=>"111100011",
  25018=>"001001001",
  25019=>"100001000",
  25020=>"011010011",
  25021=>"010101111",
  25022=>"010011000",
  25023=>"111011110",
  25024=>"000001101",
  25025=>"010000001",
  25026=>"011010010",
  25027=>"111100111",
  25028=>"101111010",
  25029=>"001000010",
  25030=>"010000100",
  25031=>"100110110",
  25032=>"111100101",
  25033=>"001111010",
  25034=>"010110100",
  25035=>"010000010",
  25036=>"000011100",
  25037=>"000110111",
  25038=>"000010000",
  25039=>"000111001",
  25040=>"110100000",
  25041=>"001000001",
  25042=>"011100010",
  25043=>"110110101",
  25044=>"001011011",
  25045=>"001001101",
  25046=>"001000110",
  25047=>"011111110",
  25048=>"011110110",
  25049=>"011001100",
  25050=>"000000111",
  25051=>"001010000",
  25052=>"001111111",
  25053=>"011111110",
  25054=>"000011000",
  25055=>"111110110",
  25056=>"001011011",
  25057=>"100011111",
  25058=>"101110110",
  25059=>"111100110",
  25060=>"111010011",
  25061=>"011101101",
  25062=>"110111111",
  25063=>"011000001",
  25064=>"011001101",
  25065=>"011001100",
  25066=>"000001100",
  25067=>"011000011",
  25068=>"101101000",
  25069=>"011101011",
  25070=>"010010100",
  25071=>"001110000",
  25072=>"011011110",
  25073=>"011011101",
  25074=>"111011000",
  25075=>"101000100",
  25076=>"110100000",
  25077=>"110010100",
  25078=>"111011011",
  25079=>"010101110",
  25080=>"001000000",
  25081=>"001101011",
  25082=>"100110111",
  25083=>"100111011",
  25084=>"000111101",
  25085=>"110111001",
  25086=>"000001101",
  25087=>"000001110",
  25088=>"011000010",
  25089=>"000101011",
  25090=>"001110010",
  25091=>"100001010",
  25092=>"101101000",
  25093=>"101100101",
  25094=>"111000011",
  25095=>"110110101",
  25096=>"001100111",
  25097=>"111110011",
  25098=>"000010101",
  25099=>"011110010",
  25100=>"101100111",
  25101=>"101101100",
  25102=>"001100010",
  25103=>"001110111",
  25104=>"000110101",
  25105=>"000100111",
  25106=>"100110111",
  25107=>"001101001",
  25108=>"110000111",
  25109=>"001100111",
  25110=>"010000000",
  25111=>"001110100",
  25112=>"000000011",
  25113=>"101110111",
  25114=>"001100100",
  25115=>"100111011",
  25116=>"101110001",
  25117=>"100010011",
  25118=>"000010111",
  25119=>"101011101",
  25120=>"001100010",
  25121=>"111101111",
  25122=>"011001000",
  25123=>"001000000",
  25124=>"110111110",
  25125=>"110011111",
  25126=>"100011100",
  25127=>"011101101",
  25128=>"010100011",
  25129=>"111100001",
  25130=>"101000011",
  25131=>"001111110",
  25132=>"111010011",
  25133=>"000100111",
  25134=>"110101100",
  25135=>"010100011",
  25136=>"110111110",
  25137=>"000100000",
  25138=>"110001110",
  25139=>"101100010",
  25140=>"000010101",
  25141=>"100100010",
  25142=>"000000111",
  25143=>"000001110",
  25144=>"001000000",
  25145=>"001000110",
  25146=>"010110010",
  25147=>"110110010",
  25148=>"110001010",
  25149=>"010010110",
  25150=>"110111100",
  25151=>"111001101",
  25152=>"111010000",
  25153=>"111110000",
  25154=>"100100110",
  25155=>"111010111",
  25156=>"010001100",
  25157=>"011100101",
  25158=>"110000010",
  25159=>"011011000",
  25160=>"001100010",
  25161=>"010110101",
  25162=>"000100111",
  25163=>"010110001",
  25164=>"111100100",
  25165=>"101011100",
  25166=>"011101011",
  25167=>"000111101",
  25168=>"011100111",
  25169=>"010010010",
  25170=>"010110100",
  25171=>"101010011",
  25172=>"011001011",
  25173=>"011110100",
  25174=>"101010001",
  25175=>"100110110",
  25176=>"001101001",
  25177=>"110100010",
  25178=>"110101000",
  25179=>"110001000",
  25180=>"100001010",
  25181=>"111001010",
  25182=>"001110000",
  25183=>"100101111",
  25184=>"111110111",
  25185=>"101101000",
  25186=>"000101011",
  25187=>"110100101",
  25188=>"001100001",
  25189=>"101111110",
  25190=>"010011000",
  25191=>"001001010",
  25192=>"001110100",
  25193=>"011000100",
  25194=>"111010101",
  25195=>"111001101",
  25196=>"100100111",
  25197=>"001011110",
  25198=>"010100010",
  25199=>"000001110",
  25200=>"011111111",
  25201=>"111011111",
  25202=>"101111000",
  25203=>"000001100",
  25204=>"110111011",
  25205=>"101100001",
  25206=>"001111110",
  25207=>"011110100",
  25208=>"111110011",
  25209=>"001011001",
  25210=>"011000111",
  25211=>"010000001",
  25212=>"001111000",
  25213=>"001000111",
  25214=>"100011110",
  25215=>"110101001",
  25216=>"110000101",
  25217=>"011100011",
  25218=>"101001110",
  25219=>"110010100",
  25220=>"000001100",
  25221=>"000001001",
  25222=>"100000110",
  25223=>"101000001",
  25224=>"101110011",
  25225=>"110110100",
  25226=>"110110111",
  25227=>"100010000",
  25228=>"101001011",
  25229=>"100011011",
  25230=>"111000001",
  25231=>"110101101",
  25232=>"110001111",
  25233=>"101011000",
  25234=>"011000101",
  25235=>"000110001",
  25236=>"010100010",
  25237=>"010000100",
  25238=>"011001111",
  25239=>"101001010",
  25240=>"000100000",
  25241=>"001111111",
  25242=>"101011000",
  25243=>"010110011",
  25244=>"110101101",
  25245=>"010011011",
  25246=>"000001011",
  25247=>"110000100",
  25248=>"101001110",
  25249=>"110000101",
  25250=>"011010000",
  25251=>"110001111",
  25252=>"100110100",
  25253=>"011101110",
  25254=>"000010111",
  25255=>"010100000",
  25256=>"011101100",
  25257=>"011011110",
  25258=>"100000001",
  25259=>"101011011",
  25260=>"000001010",
  25261=>"101010100",
  25262=>"001101001",
  25263=>"000110100",
  25264=>"001110100",
  25265=>"110000110",
  25266=>"101001100",
  25267=>"100010010",
  25268=>"000000100",
  25269=>"110010010",
  25270=>"101001110",
  25271=>"111000110",
  25272=>"000110100",
  25273=>"011110011",
  25274=>"000101110",
  25275=>"101010100",
  25276=>"000001000",
  25277=>"000011010",
  25278=>"001000100",
  25279=>"101000011",
  25280=>"011101000",
  25281=>"110011011",
  25282=>"110100111",
  25283=>"111001011",
  25284=>"100001000",
  25285=>"100110101",
  25286=>"110000110",
  25287=>"010110001",
  25288=>"111011101",
  25289=>"010111000",
  25290=>"010110111",
  25291=>"111000010",
  25292=>"100110100",
  25293=>"001110010",
  25294=>"001101011",
  25295=>"011010010",
  25296=>"001111011",
  25297=>"011111001",
  25298=>"100100001",
  25299=>"111001111",
  25300=>"100010101",
  25301=>"110110011",
  25302=>"001111011",
  25303=>"000110000",
  25304=>"000000011",
  25305=>"110000011",
  25306=>"111011011",
  25307=>"000001101",
  25308=>"110110001",
  25309=>"110100000",
  25310=>"011111000",
  25311=>"111011111",
  25312=>"011110000",
  25313=>"001100000",
  25314=>"000110010",
  25315=>"011101100",
  25316=>"100010110",
  25317=>"000100100",
  25318=>"011011111",
  25319=>"101000000",
  25320=>"101001110",
  25321=>"111110100",
  25322=>"011000110",
  25323=>"001011111",
  25324=>"101101001",
  25325=>"101111110",
  25326=>"111011111",
  25327=>"000001000",
  25328=>"110100100",
  25329=>"001011000",
  25330=>"111110001",
  25331=>"101000011",
  25332=>"101011101",
  25333=>"001001010",
  25334=>"111011111",
  25335=>"101100011",
  25336=>"001000010",
  25337=>"110110110",
  25338=>"000000111",
  25339=>"100111100",
  25340=>"101011010",
  25341=>"001000001",
  25342=>"101110011",
  25343=>"101110101",
  25344=>"101111100",
  25345=>"010100000",
  25346=>"010000000",
  25347=>"000011110",
  25348=>"101100101",
  25349=>"000111100",
  25350=>"001011010",
  25351=>"001000110",
  25352=>"000001010",
  25353=>"011111000",
  25354=>"010111101",
  25355=>"000101111",
  25356=>"111001111",
  25357=>"101110100",
  25358=>"001011000",
  25359=>"001001101",
  25360=>"010001110",
  25361=>"010101001",
  25362=>"011010110",
  25363=>"010000100",
  25364=>"100010100",
  25365=>"110011111",
  25366=>"011100011",
  25367=>"000100000",
  25368=>"010000111",
  25369=>"101010001",
  25370=>"100011001",
  25371=>"110111000",
  25372=>"011010101",
  25373=>"001100011",
  25374=>"110100000",
  25375=>"100110111",
  25376=>"101001000",
  25377=>"110001010",
  25378=>"110011011",
  25379=>"001101110",
  25380=>"111010011",
  25381=>"001001001",
  25382=>"111110110",
  25383=>"011100001",
  25384=>"011010110",
  25385=>"101110010",
  25386=>"101101011",
  25387=>"111111110",
  25388=>"001100110",
  25389=>"011000010",
  25390=>"100111100",
  25391=>"010010000",
  25392=>"000101000",
  25393=>"100111110",
  25394=>"100011010",
  25395=>"101011001",
  25396=>"010000110",
  25397=>"011001010",
  25398=>"001010001",
  25399=>"001000010",
  25400=>"110100101",
  25401=>"001001011",
  25402=>"001101110",
  25403=>"110011100",
  25404=>"000100010",
  25405=>"000011101",
  25406=>"100100101",
  25407=>"101111101",
  25408=>"010001000",
  25409=>"101111011",
  25410=>"010000101",
  25411=>"010010111",
  25412=>"011010111",
  25413=>"010010001",
  25414=>"000010111",
  25415=>"000110101",
  25416=>"110001011",
  25417=>"011111100",
  25418=>"010101110",
  25419=>"100100011",
  25420=>"010100111",
  25421=>"011011101",
  25422=>"001100101",
  25423=>"001110000",
  25424=>"000110101",
  25425=>"010111110",
  25426=>"110111010",
  25427=>"101101000",
  25428=>"011011111",
  25429=>"001101111",
  25430=>"100111111",
  25431=>"000110000",
  25432=>"011100111",
  25433=>"111011100",
  25434=>"010001010",
  25435=>"101111100",
  25436=>"101111010",
  25437=>"111000110",
  25438=>"110111111",
  25439=>"100100011",
  25440=>"001100001",
  25441=>"011001101",
  25442=>"000010000",
  25443=>"010000010",
  25444=>"100100111",
  25445=>"110000001",
  25446=>"101001110",
  25447=>"100000111",
  25448=>"000110010",
  25449=>"001101110",
  25450=>"111111000",
  25451=>"011000001",
  25452=>"101000100",
  25453=>"111110000",
  25454=>"010000001",
  25455=>"111010010",
  25456=>"001110001",
  25457=>"111100110",
  25458=>"101010001",
  25459=>"001101011",
  25460=>"110010100",
  25461=>"010001100",
  25462=>"011011111",
  25463=>"110100111",
  25464=>"110011100",
  25465=>"000011101",
  25466=>"000111000",
  25467=>"111110110",
  25468=>"000101000",
  25469=>"011101101",
  25470=>"111101110",
  25471=>"100011001",
  25472=>"010011110",
  25473=>"000101100",
  25474=>"011111110",
  25475=>"101101100",
  25476=>"010100111",
  25477=>"111010100",
  25478=>"101001010",
  25479=>"100000000",
  25480=>"101100000",
  25481=>"101100100",
  25482=>"110101011",
  25483=>"000011010",
  25484=>"111010110",
  25485=>"011000110",
  25486=>"110000100",
  25487=>"001100000",
  25488=>"110001111",
  25489=>"101010011",
  25490=>"101110000",
  25491=>"010010010",
  25492=>"101100001",
  25493=>"011101101",
  25494=>"110111010",
  25495=>"000101111",
  25496=>"110101000",
  25497=>"010101100",
  25498=>"100011101",
  25499=>"000011001",
  25500=>"010111110",
  25501=>"111000010",
  25502=>"001011010",
  25503=>"101010010",
  25504=>"011000011",
  25505=>"000011111",
  25506=>"001101110",
  25507=>"011011101",
  25508=>"000100010",
  25509=>"011100000",
  25510=>"011000000",
  25511=>"111111110",
  25512=>"110101110",
  25513=>"100010110",
  25514=>"001111101",
  25515=>"100111001",
  25516=>"101100101",
  25517=>"001001011",
  25518=>"011110110",
  25519=>"111100100",
  25520=>"101101110",
  25521=>"111001010",
  25522=>"001000101",
  25523=>"011011110",
  25524=>"000011010",
  25525=>"011101100",
  25526=>"000101111",
  25527=>"100110101",
  25528=>"111010010",
  25529=>"101101110",
  25530=>"111000101",
  25531=>"000100001",
  25532=>"101111011",
  25533=>"011111001",
  25534=>"010011011",
  25535=>"000010111",
  25536=>"110011101",
  25537=>"000000000",
  25538=>"110100010",
  25539=>"111011010",
  25540=>"011110000",
  25541=>"101001001",
  25542=>"100011010",
  25543=>"011101110",
  25544=>"100001000",
  25545=>"100000000",
  25546=>"011001011",
  25547=>"101010110",
  25548=>"000011100",
  25549=>"101100000",
  25550=>"010100100",
  25551=>"110010010",
  25552=>"000110001",
  25553=>"001100100",
  25554=>"001010100",
  25555=>"011011100",
  25556=>"111011010",
  25557=>"111011101",
  25558=>"111000100",
  25559=>"111010110",
  25560=>"101110101",
  25561=>"011111011",
  25562=>"101111110",
  25563=>"110100010",
  25564=>"000100101",
  25565=>"010101100",
  25566=>"100100110",
  25567=>"000100001",
  25568=>"010101001",
  25569=>"111000100",
  25570=>"110100001",
  25571=>"100100100",
  25572=>"000000101",
  25573=>"011111111",
  25574=>"011010000",
  25575=>"000101101",
  25576=>"001101010",
  25577=>"110111110",
  25578=>"101001011",
  25579=>"010110000",
  25580=>"010111101",
  25581=>"111011110",
  25582=>"000001110",
  25583=>"001110011",
  25584=>"000100001",
  25585=>"001011011",
  25586=>"000111011",
  25587=>"110111111",
  25588=>"100101010",
  25589=>"110011110",
  25590=>"010111011",
  25591=>"100101011",
  25592=>"101110100",
  25593=>"011001001",
  25594=>"100100011",
  25595=>"010000110",
  25596=>"011101000",
  25597=>"000101011",
  25598=>"101010011",
  25599=>"110010010",
  25600=>"110101000",
  25601=>"101010001",
  25602=>"011101011",
  25603=>"011111011",
  25604=>"110110100",
  25605=>"101110001",
  25606=>"111101011",
  25607=>"011011000",
  25608=>"101000011",
  25609=>"000001010",
  25610=>"011100001",
  25611=>"010110111",
  25612=>"010011000",
  25613=>"101000000",
  25614=>"111000010",
  25615=>"011110110",
  25616=>"101010000",
  25617=>"000100000",
  25618=>"001000111",
  25619=>"011100110",
  25620=>"111010100",
  25621=>"111011010",
  25622=>"001011010",
  25623=>"100100101",
  25624=>"011010010",
  25625=>"000000010",
  25626=>"110000000",
  25627=>"001000110",
  25628=>"000111111",
  25629=>"111110111",
  25630=>"001110000",
  25631=>"000110011",
  25632=>"100110000",
  25633=>"000100101",
  25634=>"101110111",
  25635=>"001111000",
  25636=>"011110001",
  25637=>"101101010",
  25638=>"000100001",
  25639=>"110011100",
  25640=>"010100011",
  25641=>"010011110",
  25642=>"101100101",
  25643=>"000101110",
  25644=>"100001101",
  25645=>"101011101",
  25646=>"100110111",
  25647=>"100110100",
  25648=>"101110111",
  25649=>"110110100",
  25650=>"111000000",
  25651=>"000101110",
  25652=>"100100111",
  25653=>"101001000",
  25654=>"000001101",
  25655=>"011010110",
  25656=>"001011100",
  25657=>"110111111",
  25658=>"010001011",
  25659=>"000110000",
  25660=>"011000000",
  25661=>"011000001",
  25662=>"010011000",
  25663=>"111111100",
  25664=>"111100110",
  25665=>"100011100",
  25666=>"011110100",
  25667=>"011011010",
  25668=>"100011000",
  25669=>"110001001",
  25670=>"011001100",
  25671=>"100100000",
  25672=>"000101001",
  25673=>"001100100",
  25674=>"000010010",
  25675=>"111000001",
  25676=>"110111101",
  25677=>"101111111",
  25678=>"000010011",
  25679=>"001001000",
  25680=>"001111101",
  25681=>"010001101",
  25682=>"101010001",
  25683=>"100010101",
  25684=>"110000101",
  25685=>"001010101",
  25686=>"111110111",
  25687=>"100110010",
  25688=>"111001101",
  25689=>"100101000",
  25690=>"110110111",
  25691=>"101011010",
  25692=>"000100110",
  25693=>"000101010",
  25694=>"000000011",
  25695=>"010011010",
  25696=>"111000000",
  25697=>"100011000",
  25698=>"001001111",
  25699=>"010111111",
  25700=>"000010011",
  25701=>"001000000",
  25702=>"000101101",
  25703=>"110100111",
  25704=>"110110101",
  25705=>"111010000",
  25706=>"111001101",
  25707=>"111011111",
  25708=>"110001111",
  25709=>"010111001",
  25710=>"111011011",
  25711=>"110010001",
  25712=>"111001011",
  25713=>"110111101",
  25714=>"000101111",
  25715=>"111001001",
  25716=>"000110010",
  25717=>"010100101",
  25718=>"111000111",
  25719=>"011101011",
  25720=>"100100110",
  25721=>"010000101",
  25722=>"010111110",
  25723=>"011010000",
  25724=>"100101001",
  25725=>"000111111",
  25726=>"101101110",
  25727=>"110001001",
  25728=>"011110101",
  25729=>"111111010",
  25730=>"101101000",
  25731=>"111110001",
  25732=>"001001100",
  25733=>"000101001",
  25734=>"111001110",
  25735=>"010000000",
  25736=>"000101101",
  25737=>"000100100",
  25738=>"010000111",
  25739=>"101000110",
  25740=>"111000100",
  25741=>"011001111",
  25742=>"111011000",
  25743=>"011001101",
  25744=>"111011000",
  25745=>"101101000",
  25746=>"010000001",
  25747=>"001110101",
  25748=>"101111111",
  25749=>"010101000",
  25750=>"010010010",
  25751=>"100100100",
  25752=>"000010000",
  25753=>"001011101",
  25754=>"001010110",
  25755=>"000010010",
  25756=>"000011001",
  25757=>"101000010",
  25758=>"001010110",
  25759=>"011100100",
  25760=>"110010001",
  25761=>"100101110",
  25762=>"110100110",
  25763=>"001000110",
  25764=>"100011000",
  25765=>"111001101",
  25766=>"100000100",
  25767=>"100110100",
  25768=>"110101010",
  25769=>"101111110",
  25770=>"011001010",
  25771=>"011001010",
  25772=>"101001111",
  25773=>"101101111",
  25774=>"011010110",
  25775=>"110111111",
  25776=>"010101000",
  25777=>"111000000",
  25778=>"101011111",
  25779=>"000011101",
  25780=>"000111110",
  25781=>"100101111",
  25782=>"100011000",
  25783=>"000001011",
  25784=>"001000101",
  25785=>"000110011",
  25786=>"101101010",
  25787=>"011100101",
  25788=>"111011011",
  25789=>"110001000",
  25790=>"000010010",
  25791=>"010011111",
  25792=>"101110111",
  25793=>"111000000",
  25794=>"010000000",
  25795=>"100010100",
  25796=>"001111001",
  25797=>"100101010",
  25798=>"100000010",
  25799=>"010001011",
  25800=>"101001100",
  25801=>"010110001",
  25802=>"101001111",
  25803=>"000011101",
  25804=>"111001000",
  25805=>"000001111",
  25806=>"000100001",
  25807=>"001011011",
  25808=>"100111111",
  25809=>"100110110",
  25810=>"001000001",
  25811=>"101101100",
  25812=>"000111010",
  25813=>"000100111",
  25814=>"001000000",
  25815=>"001100100",
  25816=>"001000100",
  25817=>"000011110",
  25818=>"010110011",
  25819=>"100011000",
  25820=>"010110000",
  25821=>"101100010",
  25822=>"000001000",
  25823=>"110110110",
  25824=>"010111000",
  25825=>"000100010",
  25826=>"011110011",
  25827=>"000010100",
  25828=>"111101000",
  25829=>"010011101",
  25830=>"000111110",
  25831=>"101001101",
  25832=>"010000010",
  25833=>"010011010",
  25834=>"100000001",
  25835=>"100110100",
  25836=>"011011101",
  25837=>"000101010",
  25838=>"011100010",
  25839=>"111100110",
  25840=>"000011110",
  25841=>"001000100",
  25842=>"100011000",
  25843=>"110101000",
  25844=>"110110100",
  25845=>"110010101",
  25846=>"110001111",
  25847=>"000101101",
  25848=>"111101010",
  25849=>"010001011",
  25850=>"001101101",
  25851=>"011110001",
  25852=>"011100101",
  25853=>"110100001",
  25854=>"001011010",
  25855=>"111000010",
  25856=>"111010000",
  25857=>"110101011",
  25858=>"010111000",
  25859=>"010100101",
  25860=>"010000100",
  25861=>"110111001",
  25862=>"011111111",
  25863=>"000010011",
  25864=>"111101101",
  25865=>"100101001",
  25866=>"011000101",
  25867=>"101010011",
  25868=>"110000100",
  25869=>"000010111",
  25870=>"001110100",
  25871=>"110101011",
  25872=>"000001111",
  25873=>"010111110",
  25874=>"011110110",
  25875=>"110000110",
  25876=>"101011111",
  25877=>"111110100",
  25878=>"011001100",
  25879=>"011011011",
  25880=>"101001000",
  25881=>"000000010",
  25882=>"111101000",
  25883=>"000100010",
  25884=>"010101010",
  25885=>"101010110",
  25886=>"110011001",
  25887=>"011000110",
  25888=>"000111111",
  25889=>"000000001",
  25890=>"011010110",
  25891=>"010100101",
  25892=>"000111000",
  25893=>"110101001",
  25894=>"000000101",
  25895=>"101011100",
  25896=>"110110100",
  25897=>"000011100",
  25898=>"010100111",
  25899=>"100000111",
  25900=>"110000100",
  25901=>"000111100",
  25902=>"111110010",
  25903=>"011100110",
  25904=>"011110111",
  25905=>"001111111",
  25906=>"010111010",
  25907=>"110011001",
  25908=>"111001011",
  25909=>"101010000",
  25910=>"010010010",
  25911=>"100111011",
  25912=>"110000000",
  25913=>"110010001",
  25914=>"111001111",
  25915=>"111011111",
  25916=>"110011111",
  25917=>"111010011",
  25918=>"100000001",
  25919=>"001100110",
  25920=>"101001011",
  25921=>"010110001",
  25922=>"000011110",
  25923=>"001000011",
  25924=>"000110010",
  25925=>"110001111",
  25926=>"111111001",
  25927=>"010111000",
  25928=>"010001100",
  25929=>"100001111",
  25930=>"000001100",
  25931=>"111000011",
  25932=>"000000001",
  25933=>"001011000",
  25934=>"001111000",
  25935=>"010111111",
  25936=>"001110101",
  25937=>"000001111",
  25938=>"000101100",
  25939=>"001100100",
  25940=>"000111111",
  25941=>"110001111",
  25942=>"000010000",
  25943=>"111010010",
  25944=>"010000000",
  25945=>"111100111",
  25946=>"000100001",
  25947=>"001010000",
  25948=>"100110111",
  25949=>"110111111",
  25950=>"111111101",
  25951=>"110000011",
  25952=>"001001111",
  25953=>"010101000",
  25954=>"100100110",
  25955=>"000111001",
  25956=>"101010011",
  25957=>"001010101",
  25958=>"011101100",
  25959=>"011001000",
  25960=>"100000000",
  25961=>"000010000",
  25962=>"111000100",
  25963=>"110010000",
  25964=>"110011010",
  25965=>"100100000",
  25966=>"100010100",
  25967=>"111110101",
  25968=>"010110111",
  25969=>"001111001",
  25970=>"110100100",
  25971=>"011010000",
  25972=>"011101011",
  25973=>"001110011",
  25974=>"010100011",
  25975=>"111101111",
  25976=>"101001110",
  25977=>"001011010",
  25978=>"111011001",
  25979=>"110100111",
  25980=>"010011000",
  25981=>"000000011",
  25982=>"011111001",
  25983=>"011010000",
  25984=>"111000011",
  25985=>"010110110",
  25986=>"010000110",
  25987=>"110100111",
  25988=>"101111011",
  25989=>"101110111",
  25990=>"001001101",
  25991=>"011111110",
  25992=>"010001000",
  25993=>"011100110",
  25994=>"000011101",
  25995=>"010000100",
  25996=>"110101110",
  25997=>"100011110",
  25998=>"001001000",
  25999=>"011100110",
  26000=>"110111100",
  26001=>"000100110",
  26002=>"111101101",
  26003=>"101001001",
  26004=>"111010110",
  26005=>"000010000",
  26006=>"000001000",
  26007=>"001001010",
  26008=>"100101011",
  26009=>"000111001",
  26010=>"110001110",
  26011=>"111010111",
  26012=>"110100100",
  26013=>"000000111",
  26014=>"000111100",
  26015=>"000000000",
  26016=>"111011110",
  26017=>"111111001",
  26018=>"100110010",
  26019=>"000000000",
  26020=>"010011110",
  26021=>"111100100",
  26022=>"100101011",
  26023=>"101111011",
  26024=>"011110101",
  26025=>"011000000",
  26026=>"000000111",
  26027=>"000101000",
  26028=>"101100111",
  26029=>"101110101",
  26030=>"110010101",
  26031=>"100100001",
  26032=>"000000000",
  26033=>"010101100",
  26034=>"010100001",
  26035=>"110001000",
  26036=>"111101011",
  26037=>"010100101",
  26038=>"000011111",
  26039=>"110100010",
  26040=>"100110110",
  26041=>"101011011",
  26042=>"001110110",
  26043=>"000000111",
  26044=>"011001010",
  26045=>"100110011",
  26046=>"010100111",
  26047=>"000001010",
  26048=>"110011000",
  26049=>"000001111",
  26050=>"000111000",
  26051=>"100001001",
  26052=>"110001001",
  26053=>"100111011",
  26054=>"011010001",
  26055=>"010011000",
  26056=>"010011111",
  26057=>"110010011",
  26058=>"110000011",
  26059=>"110101100",
  26060=>"101011101",
  26061=>"001011000",
  26062=>"000100111",
  26063=>"111010111",
  26064=>"101010001",
  26065=>"101100100",
  26066=>"010110111",
  26067=>"110001000",
  26068=>"110011111",
  26069=>"101101010",
  26070=>"000110100",
  26071=>"011101100",
  26072=>"011001001",
  26073=>"001111101",
  26074=>"000011010",
  26075=>"000010101",
  26076=>"001000111",
  26077=>"111111000",
  26078=>"011011011",
  26079=>"111001000",
  26080=>"001111000",
  26081=>"111010110",
  26082=>"100111001",
  26083=>"000000000",
  26084=>"001010101",
  26085=>"000000010",
  26086=>"001001011",
  26087=>"111011110",
  26088=>"111100000",
  26089=>"010100011",
  26090=>"001000101",
  26091=>"101001011",
  26092=>"000000000",
  26093=>"111111011",
  26094=>"010000000",
  26095=>"000100001",
  26096=>"010111001",
  26097=>"100111110",
  26098=>"000100111",
  26099=>"110101010",
  26100=>"111010101",
  26101=>"100101000",
  26102=>"101100100",
  26103=>"000110101",
  26104=>"000010111",
  26105=>"000000111",
  26106=>"001010111",
  26107=>"000000110",
  26108=>"011101001",
  26109=>"011110110",
  26110=>"101110011",
  26111=>"001100000",
  26112=>"011110110",
  26113=>"111000101",
  26114=>"011110011",
  26115=>"100011111",
  26116=>"101100101",
  26117=>"000000110",
  26118=>"000100111",
  26119=>"111010110",
  26120=>"110010011",
  26121=>"010101111",
  26122=>"011100110",
  26123=>"111011000",
  26124=>"110010000",
  26125=>"100110101",
  26126=>"000010111",
  26127=>"001111100",
  26128=>"000100011",
  26129=>"000000110",
  26130=>"010010100",
  26131=>"100011000",
  26132=>"000011010",
  26133=>"101110000",
  26134=>"001111010",
  26135=>"111011011",
  26136=>"111101011",
  26137=>"111001001",
  26138=>"100110011",
  26139=>"001100010",
  26140=>"000100101",
  26141=>"101001011",
  26142=>"101100110",
  26143=>"100111111",
  26144=>"011111111",
  26145=>"101001011",
  26146=>"111101110",
  26147=>"000100000",
  26148=>"010001000",
  26149=>"100111010",
  26150=>"011010010",
  26151=>"000010101",
  26152=>"100010000",
  26153=>"110011001",
  26154=>"000001000",
  26155=>"001001011",
  26156=>"110010110",
  26157=>"100111101",
  26158=>"100001010",
  26159=>"011010100",
  26160=>"101011100",
  26161=>"001011100",
  26162=>"101101011",
  26163=>"001000011",
  26164=>"000110000",
  26165=>"000000010",
  26166=>"011100001",
  26167=>"100111100",
  26168=>"011111100",
  26169=>"110010111",
  26170=>"001110010",
  26171=>"100011011",
  26172=>"101101100",
  26173=>"100000110",
  26174=>"011010101",
  26175=>"001010010",
  26176=>"111100011",
  26177=>"100110111",
  26178=>"111110000",
  26179=>"000111010",
  26180=>"111110110",
  26181=>"001111110",
  26182=>"101011001",
  26183=>"000010110",
  26184=>"000100100",
  26185=>"000100001",
  26186=>"000101111",
  26187=>"100010111",
  26188=>"010110011",
  26189=>"011011100",
  26190=>"111011010",
  26191=>"000100001",
  26192=>"000011101",
  26193=>"100110011",
  26194=>"001010110",
  26195=>"110000001",
  26196=>"100100111",
  26197=>"111110101",
  26198=>"010011100",
  26199=>"101100110",
  26200=>"100111001",
  26201=>"010110101",
  26202=>"110010100",
  26203=>"111100110",
  26204=>"000100001",
  26205=>"000000001",
  26206=>"010001001",
  26207=>"001000000",
  26208=>"001000111",
  26209=>"000010001",
  26210=>"100111111",
  26211=>"111110111",
  26212=>"100101100",
  26213=>"100101001",
  26214=>"110011011",
  26215=>"001101111",
  26216=>"000101010",
  26217=>"011111110",
  26218=>"110101001",
  26219=>"010000010",
  26220=>"110000001",
  26221=>"111011100",
  26222=>"011101001",
  26223=>"000000101",
  26224=>"000100000",
  26225=>"011000111",
  26226=>"001101111",
  26227=>"000000010",
  26228=>"100101001",
  26229=>"011011100",
  26230=>"111111000",
  26231=>"111011010",
  26232=>"000010100",
  26233=>"001000011",
  26234=>"111100000",
  26235=>"000000110",
  26236=>"100000100",
  26237=>"111111101",
  26238=>"011011101",
  26239=>"110010010",
  26240=>"010111100",
  26241=>"001100000",
  26242=>"010110101",
  26243=>"001000001",
  26244=>"010110010",
  26245=>"000000101",
  26246=>"110100001",
  26247=>"101011001",
  26248=>"111101110",
  26249=>"100100010",
  26250=>"111001011",
  26251=>"110110000",
  26252=>"110011111",
  26253=>"010100110",
  26254=>"001001010",
  26255=>"011111001",
  26256=>"110000101",
  26257=>"000011010",
  26258=>"010100011",
  26259=>"110001110",
  26260=>"010110101",
  26261=>"110110100",
  26262=>"111110111",
  26263=>"111101100",
  26264=>"001010001",
  26265=>"111100000",
  26266=>"010000101",
  26267=>"110101100",
  26268=>"000100011",
  26269=>"000000111",
  26270=>"011111111",
  26271=>"000011101",
  26272=>"111101000",
  26273=>"010011001",
  26274=>"000001000",
  26275=>"011011101",
  26276=>"101101111",
  26277=>"011101100",
  26278=>"011010011",
  26279=>"010110000",
  26280=>"101111110",
  26281=>"000001101",
  26282=>"110000101",
  26283=>"010000000",
  26284=>"000001101",
  26285=>"001001101",
  26286=>"011011000",
  26287=>"110010001",
  26288=>"010100111",
  26289=>"101011111",
  26290=>"000011111",
  26291=>"001001000",
  26292=>"101110101",
  26293=>"011000010",
  26294=>"000100110",
  26295=>"001011010",
  26296=>"001011111",
  26297=>"000101010",
  26298=>"100001111",
  26299=>"001010001",
  26300=>"000111011",
  26301=>"011100100",
  26302=>"010111011",
  26303=>"000000000",
  26304=>"111110101",
  26305=>"010110100",
  26306=>"000010010",
  26307=>"100111111",
  26308=>"011011011",
  26309=>"001100101",
  26310=>"011111001",
  26311=>"000100100",
  26312=>"001110000",
  26313=>"101010001",
  26314=>"100100010",
  26315=>"101101111",
  26316=>"000111000",
  26317=>"101111111",
  26318=>"111101001",
  26319=>"110111111",
  26320=>"100000000",
  26321=>"010100001",
  26322=>"011100010",
  26323=>"001101000",
  26324=>"111000111",
  26325=>"101001101",
  26326=>"111001111",
  26327=>"100001110",
  26328=>"000100101",
  26329=>"100001111",
  26330=>"101000000",
  26331=>"101000000",
  26332=>"001110011",
  26333=>"111101001",
  26334=>"101110101",
  26335=>"110000001",
  26336=>"001101011",
  26337=>"010000000",
  26338=>"100100110",
  26339=>"011100000",
  26340=>"011000001",
  26341=>"100100010",
  26342=>"010101000",
  26343=>"101011011",
  26344=>"000110111",
  26345=>"000110110",
  26346=>"100110100",
  26347=>"111010011",
  26348=>"001100001",
  26349=>"000100100",
  26350=>"101101100",
  26351=>"110101100",
  26352=>"101000111",
  26353=>"011001000",
  26354=>"001100110",
  26355=>"000011000",
  26356=>"010001011",
  26357=>"101010110",
  26358=>"100011101",
  26359=>"001111101",
  26360=>"101001000",
  26361=>"100101100",
  26362=>"100111001",
  26363=>"000000101",
  26364=>"101111111",
  26365=>"000110010",
  26366=>"101111111",
  26367=>"111001000",
  26368=>"011000010",
  26369=>"111010011",
  26370=>"101100111",
  26371=>"101001001",
  26372=>"011011000",
  26373=>"000000011",
  26374=>"000001101",
  26375=>"000101111",
  26376=>"011111000",
  26377=>"100011110",
  26378=>"101000111",
  26379=>"010011000",
  26380=>"101011000",
  26381=>"001010001",
  26382=>"001101100",
  26383=>"100001101",
  26384=>"110010000",
  26385=>"000101000",
  26386=>"001010110",
  26387=>"001100100",
  26388=>"000100111",
  26389=>"100001100",
  26390=>"000101101",
  26391=>"001110000",
  26392=>"110111000",
  26393=>"001010101",
  26394=>"100000010",
  26395=>"001011110",
  26396=>"000101110",
  26397=>"101110111",
  26398=>"011010100",
  26399=>"101010101",
  26400=>"101111100",
  26401=>"011111100",
  26402=>"001101000",
  26403=>"111001100",
  26404=>"101101101",
  26405=>"000100101",
  26406=>"111100111",
  26407=>"000110111",
  26408=>"101110111",
  26409=>"000011000",
  26410=>"101110100",
  26411=>"110001100",
  26412=>"111101011",
  26413=>"010001011",
  26414=>"010000001",
  26415=>"101011111",
  26416=>"110010101",
  26417=>"000011000",
  26418=>"001011111",
  26419=>"010000110",
  26420=>"110000100",
  26421=>"110011100",
  26422=>"011110011",
  26423=>"111111000",
  26424=>"011010110",
  26425=>"010110111",
  26426=>"111000001",
  26427=>"001101111",
  26428=>"101011111",
  26429=>"100000111",
  26430=>"000100101",
  26431=>"100101111",
  26432=>"000010101",
  26433=>"110110110",
  26434=>"111111011",
  26435=>"001101110",
  26436=>"000100010",
  26437=>"110100010",
  26438=>"001101110",
  26439=>"001110010",
  26440=>"010110101",
  26441=>"011011101",
  26442=>"001010001",
  26443=>"001111000",
  26444=>"100000001",
  26445=>"010000110",
  26446=>"110010110",
  26447=>"101111001",
  26448=>"011111111",
  26449=>"000000110",
  26450=>"011101011",
  26451=>"010001011",
  26452=>"011000111",
  26453=>"100011111",
  26454=>"111111101",
  26455=>"101001111",
  26456=>"000101111",
  26457=>"111000010",
  26458=>"110101001",
  26459=>"100101100",
  26460=>"111100010",
  26461=>"100001110",
  26462=>"001000111",
  26463=>"011001000",
  26464=>"000010000",
  26465=>"010111011",
  26466=>"001101110",
  26467=>"000111001",
  26468=>"011100011",
  26469=>"111111111",
  26470=>"000111011",
  26471=>"111001111",
  26472=>"101111010",
  26473=>"111100010",
  26474=>"011110011",
  26475=>"000101001",
  26476=>"100111101",
  26477=>"011111000",
  26478=>"000001110",
  26479=>"001010110",
  26480=>"000011000",
  26481=>"101011100",
  26482=>"010100000",
  26483=>"001110000",
  26484=>"000000011",
  26485=>"000011110",
  26486=>"111001000",
  26487=>"011100000",
  26488=>"010000011",
  26489=>"000101101",
  26490=>"001111001",
  26491=>"110101110",
  26492=>"010100111",
  26493=>"101101010",
  26494=>"101010010",
  26495=>"001001000",
  26496=>"011100110",
  26497=>"010110011",
  26498=>"000101111",
  26499=>"111011000",
  26500=>"010001100",
  26501=>"100110010",
  26502=>"110001000",
  26503=>"111111101",
  26504=>"100000100",
  26505=>"111111000",
  26506=>"101011110",
  26507=>"110100000",
  26508=>"111000000",
  26509=>"000100110",
  26510=>"001000000",
  26511=>"110000111",
  26512=>"100111010",
  26513=>"110111101",
  26514=>"000000101",
  26515=>"100101101",
  26516=>"101110111",
  26517=>"111111000",
  26518=>"000111011",
  26519=>"101100000",
  26520=>"010101000",
  26521=>"001111001",
  26522=>"010001000",
  26523=>"000000101",
  26524=>"001110110",
  26525=>"011001100",
  26526=>"000001000",
  26527=>"011011111",
  26528=>"100111000",
  26529=>"011001010",
  26530=>"001010011",
  26531=>"100011010",
  26532=>"001111010",
  26533=>"101001110",
  26534=>"011110000",
  26535=>"101010111",
  26536=>"000011100",
  26537=>"011001110",
  26538=>"111010000",
  26539=>"011000100",
  26540=>"110101100",
  26541=>"011111101",
  26542=>"001001010",
  26543=>"101111011",
  26544=>"001011011",
  26545=>"101000111",
  26546=>"010101111",
  26547=>"001010001",
  26548=>"000001010",
  26549=>"001111111",
  26550=>"110100100",
  26551=>"010110011",
  26552=>"111110110",
  26553=>"011001101",
  26554=>"011000110",
  26555=>"001111111",
  26556=>"011010000",
  26557=>"010100000",
  26558=>"001100101",
  26559=>"010000000",
  26560=>"010010011",
  26561=>"000001111",
  26562=>"011001001",
  26563=>"000101100",
  26564=>"100100111",
  26565=>"111001010",
  26566=>"010100010",
  26567=>"110000100",
  26568=>"111101110",
  26569=>"011011000",
  26570=>"110110011",
  26571=>"011010100",
  26572=>"000111111",
  26573=>"001111001",
  26574=>"100001000",
  26575=>"001110111",
  26576=>"101101101",
  26577=>"111001001",
  26578=>"101011001",
  26579=>"000010111",
  26580=>"111010100",
  26581=>"101001110",
  26582=>"000110110",
  26583=>"011101111",
  26584=>"111101111",
  26585=>"111011110",
  26586=>"000111111",
  26587=>"010110000",
  26588=>"000010000",
  26589=>"100101100",
  26590=>"111010010",
  26591=>"010111101",
  26592=>"111000100",
  26593=>"101110010",
  26594=>"101011001",
  26595=>"000011110",
  26596=>"000001000",
  26597=>"010001010",
  26598=>"001110111",
  26599=>"111110010",
  26600=>"001111111",
  26601=>"001101101",
  26602=>"110001000",
  26603=>"010001111",
  26604=>"010001110",
  26605=>"000101110",
  26606=>"111101001",
  26607=>"110001111",
  26608=>"001100101",
  26609=>"110010100",
  26610=>"001101111",
  26611=>"110100000",
  26612=>"011011110",
  26613=>"100000111",
  26614=>"010001110",
  26615=>"000110110",
  26616=>"111100001",
  26617=>"111111101",
  26618=>"100000100",
  26619=>"000010001",
  26620=>"100001101",
  26621=>"000110011",
  26622=>"010000101",
  26623=>"100100110",
  26624=>"100000000",
  26625=>"010111000",
  26626=>"000001011",
  26627=>"010001111",
  26628=>"011010011",
  26629=>"110000110",
  26630=>"001010110",
  26631=>"000100111",
  26632=>"011010001",
  26633=>"011000001",
  26634=>"000101000",
  26635=>"001000100",
  26636=>"010010001",
  26637=>"000111010",
  26638=>"010001000",
  26639=>"011100000",
  26640=>"110010111",
  26641=>"111010110",
  26642=>"111101101",
  26643=>"100011101",
  26644=>"011001010",
  26645=>"110001100",
  26646=>"110010110",
  26647=>"100110100",
  26648=>"000111100",
  26649=>"111111001",
  26650=>"100010110",
  26651=>"110001011",
  26652=>"011101100",
  26653=>"011111111",
  26654=>"100010100",
  26655=>"110110010",
  26656=>"000111000",
  26657=>"010110010",
  26658=>"011100010",
  26659=>"011100100",
  26660=>"111101011",
  26661=>"110100010",
  26662=>"111101011",
  26663=>"111000000",
  26664=>"100010110",
  26665=>"110010000",
  26666=>"010000111",
  26667=>"001100001",
  26668=>"101101101",
  26669=>"110111110",
  26670=>"001000000",
  26671=>"000011111",
  26672=>"000011000",
  26673=>"001001010",
  26674=>"000011111",
  26675=>"010001000",
  26676=>"011110010",
  26677=>"000101000",
  26678=>"010011001",
  26679=>"000111111",
  26680=>"000101001",
  26681=>"101101001",
  26682=>"010001000",
  26683=>"100000110",
  26684=>"010001000",
  26685=>"011101010",
  26686=>"000110101",
  26687=>"000110001",
  26688=>"010110110",
  26689=>"000000000",
  26690=>"001101001",
  26691=>"101001111",
  26692=>"100010111",
  26693=>"011010001",
  26694=>"101001010",
  26695=>"111000001",
  26696=>"111111010",
  26697=>"010011100",
  26698=>"101100110",
  26699=>"001100110",
  26700=>"010000001",
  26701=>"000001011",
  26702=>"011010010",
  26703=>"001101100",
  26704=>"010101111",
  26705=>"111101111",
  26706=>"011101110",
  26707=>"010000110",
  26708=>"100011001",
  26709=>"111110110",
  26710=>"011001100",
  26711=>"101100010",
  26712=>"011010001",
  26713=>"010100110",
  26714=>"101010111",
  26715=>"111010100",
  26716=>"100100010",
  26717=>"100100000",
  26718=>"010010010",
  26719=>"010001111",
  26720=>"100010010",
  26721=>"011000010",
  26722=>"000001000",
  26723=>"111010001",
  26724=>"110010101",
  26725=>"010011001",
  26726=>"011111000",
  26727=>"000000110",
  26728=>"000001011",
  26729=>"110000011",
  26730=>"001010010",
  26731=>"011111010",
  26732=>"000010010",
  26733=>"111100010",
  26734=>"011000110",
  26735=>"011001001",
  26736=>"000010100",
  26737=>"010011011",
  26738=>"111101101",
  26739=>"101100010",
  26740=>"000110011",
  26741=>"101110110",
  26742=>"011101111",
  26743=>"111101001",
  26744=>"100011011",
  26745=>"001111000",
  26746=>"101110010",
  26747=>"000110000",
  26748=>"000110011",
  26749=>"010110010",
  26750=>"010000000",
  26751=>"000111101",
  26752=>"010100101",
  26753=>"010000000",
  26754=>"111101010",
  26755=>"011011011",
  26756=>"110011100",
  26757=>"001111011",
  26758=>"011010000",
  26759=>"110101111",
  26760=>"111010101",
  26761=>"000110001",
  26762=>"100001011",
  26763=>"010001101",
  26764=>"101100011",
  26765=>"010010011",
  26766=>"100000111",
  26767=>"100000011",
  26768=>"110100100",
  26769=>"001110001",
  26770=>"001010010",
  26771=>"111110011",
  26772=>"011011011",
  26773=>"101011011",
  26774=>"000110010",
  26775=>"110011100",
  26776=>"011000000",
  26777=>"100010100",
  26778=>"011000000",
  26779=>"110100110",
  26780=>"101001010",
  26781=>"111111010",
  26782=>"000010010",
  26783=>"010110010",
  26784=>"101001001",
  26785=>"010001110",
  26786=>"110000111",
  26787=>"110110110",
  26788=>"100001011",
  26789=>"100000100",
  26790=>"111010110",
  26791=>"010000101",
  26792=>"010000110",
  26793=>"101001001",
  26794=>"100111010",
  26795=>"001010010",
  26796=>"100001111",
  26797=>"110001001",
  26798=>"001100011",
  26799=>"101111100",
  26800=>"010111010",
  26801=>"010000011",
  26802=>"001001101",
  26803=>"101101011",
  26804=>"011101110",
  26805=>"000010111",
  26806=>"110110111",
  26807=>"010101111",
  26808=>"101011010",
  26809=>"110110101",
  26810=>"010100000",
  26811=>"100111101",
  26812=>"000001101",
  26813=>"101000101",
  26814=>"000100110",
  26815=>"111011000",
  26816=>"010100011",
  26817=>"011110010",
  26818=>"000101000",
  26819=>"010111110",
  26820=>"000000100",
  26821=>"101010010",
  26822=>"101000011",
  26823=>"010101101",
  26824=>"010010110",
  26825=>"000100001",
  26826=>"011010110",
  26827=>"000010110",
  26828=>"110010001",
  26829=>"110111111",
  26830=>"011101110",
  26831=>"000011101",
  26832=>"010101111",
  26833=>"111110111",
  26834=>"100010000",
  26835=>"010111010",
  26836=>"011001001",
  26837=>"000111010",
  26838=>"000000000",
  26839=>"011111011",
  26840=>"100110111",
  26841=>"011010110",
  26842=>"000011100",
  26843=>"110100011",
  26844=>"111010001",
  26845=>"001100010",
  26846=>"110011001",
  26847=>"000011100",
  26848=>"000110110",
  26849=>"111011110",
  26850=>"100011110",
  26851=>"111110010",
  26852=>"111101101",
  26853=>"011001110",
  26854=>"010100010",
  26855=>"101000101",
  26856=>"101000011",
  26857=>"100011000",
  26858=>"010110011",
  26859=>"101000010",
  26860=>"100011110",
  26861=>"101111110",
  26862=>"101001010",
  26863=>"100010101",
  26864=>"011100100",
  26865=>"001110001",
  26866=>"011011010",
  26867=>"001000000",
  26868=>"010100110",
  26869=>"101101000",
  26870=>"101010011",
  26871=>"101100010",
  26872=>"010110000",
  26873=>"000000010",
  26874=>"110000001",
  26875=>"111001000",
  26876=>"010011000",
  26877=>"111011011",
  26878=>"111111000",
  26879=>"000101001",
  26880=>"010110011",
  26881=>"100111010",
  26882=>"010000011",
  26883=>"000010100",
  26884=>"110010101",
  26885=>"000010101",
  26886=>"000011110",
  26887=>"001011001",
  26888=>"011111000",
  26889=>"000001001",
  26890=>"011000100",
  26891=>"111101011",
  26892=>"000000001",
  26893=>"011001101",
  26894=>"000011100",
  26895=>"001001000",
  26896=>"111011101",
  26897=>"000000000",
  26898=>"001000010",
  26899=>"010101001",
  26900=>"001011000",
  26901=>"111010010",
  26902=>"111111101",
  26903=>"111000100",
  26904=>"010111000",
  26905=>"000110100",
  26906=>"001100111",
  26907=>"011001010",
  26908=>"000111001",
  26909=>"000100000",
  26910=>"100100010",
  26911=>"110000110",
  26912=>"101011101",
  26913=>"110011111",
  26914=>"000000000",
  26915=>"000000111",
  26916=>"101000001",
  26917=>"101110110",
  26918=>"000101110",
  26919=>"000111101",
  26920=>"010010101",
  26921=>"100001111",
  26922=>"000010001",
  26923=>"001100001",
  26924=>"000000001",
  26925=>"100000011",
  26926=>"000000001",
  26927=>"000001111",
  26928=>"110111001",
  26929=>"011101110",
  26930=>"010000011",
  26931=>"000110000",
  26932=>"100101000",
  26933=>"001000001",
  26934=>"011000000",
  26935=>"010001011",
  26936=>"001001000",
  26937=>"101011001",
  26938=>"110111001",
  26939=>"111111101",
  26940=>"001110101",
  26941=>"110110110",
  26942=>"000111001",
  26943=>"110000100",
  26944=>"011111001",
  26945=>"101100100",
  26946=>"111100100",
  26947=>"100100100",
  26948=>"011110010",
  26949=>"101110001",
  26950=>"001001101",
  26951=>"110001000",
  26952=>"010100000",
  26953=>"100001011",
  26954=>"101111100",
  26955=>"000110100",
  26956=>"010101110",
  26957=>"011010111",
  26958=>"001110011",
  26959=>"011111000",
  26960=>"101111100",
  26961=>"111100010",
  26962=>"111010011",
  26963=>"010010110",
  26964=>"100100110",
  26965=>"001011101",
  26966=>"010011010",
  26967=>"110110111",
  26968=>"100000110",
  26969=>"001011001",
  26970=>"000010001",
  26971=>"100001000",
  26972=>"001001001",
  26973=>"101011111",
  26974=>"010111010",
  26975=>"000001011",
  26976=>"000110001",
  26977=>"111000111",
  26978=>"101100010",
  26979=>"100100100",
  26980=>"011011001",
  26981=>"111100011",
  26982=>"011111011",
  26983=>"111001101",
  26984=>"111011011",
  26985=>"011100110",
  26986=>"000110010",
  26987=>"000000000",
  26988=>"100010100",
  26989=>"000010101",
  26990=>"100000100",
  26991=>"001010001",
  26992=>"000101111",
  26993=>"110111000",
  26994=>"110001110",
  26995=>"011101011",
  26996=>"101111001",
  26997=>"111111011",
  26998=>"111010111",
  26999=>"010111000",
  27000=>"010100100",
  27001=>"011001000",
  27002=>"111011100",
  27003=>"111100011",
  27004=>"000011000",
  27005=>"101011001",
  27006=>"101011111",
  27007=>"101100010",
  27008=>"001001001",
  27009=>"000000000",
  27010=>"111110111",
  27011=>"001101111",
  27012=>"010011111",
  27013=>"110110110",
  27014=>"101011111",
  27015=>"000000110",
  27016=>"110001001",
  27017=>"010011111",
  27018=>"110000010",
  27019=>"011000001",
  27020=>"001001000",
  27021=>"100011101",
  27022=>"111101001",
  27023=>"011100100",
  27024=>"001101111",
  27025=>"101000010",
  27026=>"001001001",
  27027=>"011000011",
  27028=>"011110110",
  27029=>"010100111",
  27030=>"111111111",
  27031=>"110010001",
  27032=>"001110100",
  27033=>"001111001",
  27034=>"001110100",
  27035=>"111110001",
  27036=>"100101000",
  27037=>"011111101",
  27038=>"100000110",
  27039=>"111111011",
  27040=>"100001011",
  27041=>"001000000",
  27042=>"110110010",
  27043=>"101100001",
  27044=>"110100001",
  27045=>"111101100",
  27046=>"111010110",
  27047=>"010010111",
  27048=>"010101010",
  27049=>"111101010",
  27050=>"000111101",
  27051=>"110011001",
  27052=>"000001011",
  27053=>"111000010",
  27054=>"010101101",
  27055=>"111111000",
  27056=>"010001001",
  27057=>"111110100",
  27058=>"101011111",
  27059=>"111011000",
  27060=>"011000111",
  27061=>"010101011",
  27062=>"000101010",
  27063=>"010011110",
  27064=>"111101010",
  27065=>"001100111",
  27066=>"001101001",
  27067=>"001010010",
  27068=>"010010000",
  27069=>"000110101",
  27070=>"011101111",
  27071=>"111010000",
  27072=>"101000001",
  27073=>"010100111",
  27074=>"010001011",
  27075=>"101011000",
  27076=>"000010101",
  27077=>"010101100",
  27078=>"100100100",
  27079=>"000000000",
  27080=>"101101100",
  27081=>"000111111",
  27082=>"000011111",
  27083=>"000100111",
  27084=>"001001101",
  27085=>"110000110",
  27086=>"001011111",
  27087=>"101010001",
  27088=>"100010001",
  27089=>"110101111",
  27090=>"000011001",
  27091=>"000000110",
  27092=>"000100010",
  27093=>"011101010",
  27094=>"011100100",
  27095=>"010010010",
  27096=>"100101111",
  27097=>"011110010",
  27098=>"111010010",
  27099=>"000000110",
  27100=>"001001101",
  27101=>"111001100",
  27102=>"010011001",
  27103=>"110111100",
  27104=>"110011110",
  27105=>"111011001",
  27106=>"111100110",
  27107=>"110110001",
  27108=>"010010111",
  27109=>"001001111",
  27110=>"111101000",
  27111=>"001001000",
  27112=>"000110110",
  27113=>"000011001",
  27114=>"101101100",
  27115=>"011111110",
  27116=>"010001001",
  27117=>"010101000",
  27118=>"110100001",
  27119=>"001000110",
  27120=>"000000000",
  27121=>"111010100",
  27122=>"111010001",
  27123=>"010000101",
  27124=>"101000001",
  27125=>"110010000",
  27126=>"000000110",
  27127=>"001100110",
  27128=>"001001011",
  27129=>"111011110",
  27130=>"001100001",
  27131=>"101001010",
  27132=>"101111011",
  27133=>"010001000",
  27134=>"111110111",
  27135=>"110110001",
  27136=>"011111011",
  27137=>"001011000",
  27138=>"011101101",
  27139=>"010100000",
  27140=>"000101110",
  27141=>"111110101",
  27142=>"101001011",
  27143=>"101100101",
  27144=>"010111000",
  27145=>"010101001",
  27146=>"101100011",
  27147=>"011101110",
  27148=>"000110000",
  27149=>"111110110",
  27150=>"110000010",
  27151=>"010010111",
  27152=>"110010011",
  27153=>"000001110",
  27154=>"111000000",
  27155=>"100101011",
  27156=>"010010000",
  27157=>"100100100",
  27158=>"010111110",
  27159=>"001010010",
  27160=>"110000001",
  27161=>"001111001",
  27162=>"011001100",
  27163=>"101000001",
  27164=>"111000111",
  27165=>"001001011",
  27166=>"101100000",
  27167=>"001101010",
  27168=>"110010001",
  27169=>"101001110",
  27170=>"100010001",
  27171=>"011000010",
  27172=>"110100001",
  27173=>"001010000",
  27174=>"111101110",
  27175=>"001000000",
  27176=>"111001001",
  27177=>"110011010",
  27178=>"101010110",
  27179=>"001010001",
  27180=>"001001000",
  27181=>"000101110",
  27182=>"101100010",
  27183=>"100000001",
  27184=>"010101111",
  27185=>"000010011",
  27186=>"000000011",
  27187=>"100111111",
  27188=>"001000110",
  27189=>"001111010",
  27190=>"101100011",
  27191=>"100100111",
  27192=>"100010101",
  27193=>"111011111",
  27194=>"011110011",
  27195=>"111000101",
  27196=>"110111011",
  27197=>"000010110",
  27198=>"111010101",
  27199=>"010111100",
  27200=>"101001110",
  27201=>"111100110",
  27202=>"110110111",
  27203=>"001110001",
  27204=>"010110110",
  27205=>"000111001",
  27206=>"001000001",
  27207=>"010000111",
  27208=>"101010001",
  27209=>"110100001",
  27210=>"000011011",
  27211=>"011001011",
  27212=>"110001110",
  27213=>"100101110",
  27214=>"110111001",
  27215=>"010111110",
  27216=>"110110001",
  27217=>"101110000",
  27218=>"101111001",
  27219=>"110010010",
  27220=>"011001000",
  27221=>"001000001",
  27222=>"101001100",
  27223=>"000111100",
  27224=>"101010101",
  27225=>"111001010",
  27226=>"110011010",
  27227=>"011100101",
  27228=>"110011001",
  27229=>"001000100",
  27230=>"000111101",
  27231=>"111000000",
  27232=>"101100110",
  27233=>"001100101",
  27234=>"110000011",
  27235=>"111010110",
  27236=>"110110111",
  27237=>"101100000",
  27238=>"010100000",
  27239=>"101110011",
  27240=>"000101011",
  27241=>"110101010",
  27242=>"010010010",
  27243=>"111000000",
  27244=>"100010110",
  27245=>"110111000",
  27246=>"101111011",
  27247=>"100000110",
  27248=>"110110110",
  27249=>"000000001",
  27250=>"111110101",
  27251=>"010000001",
  27252=>"101110111",
  27253=>"110100101",
  27254=>"011010101",
  27255=>"010101010",
  27256=>"111101000",
  27257=>"000101111",
  27258=>"001001101",
  27259=>"011000000",
  27260=>"100100001",
  27261=>"000100101",
  27262=>"010000100",
  27263=>"100000101",
  27264=>"000000110",
  27265=>"011001101",
  27266=>"110111111",
  27267=>"001010101",
  27268=>"000100110",
  27269=>"100000010",
  27270=>"000011001",
  27271=>"010101100",
  27272=>"000000010",
  27273=>"011111110",
  27274=>"111111111",
  27275=>"000000011",
  27276=>"111000001",
  27277=>"101110110",
  27278=>"011100001",
  27279=>"010000001",
  27280=>"011001110",
  27281=>"001000000",
  27282=>"111000101",
  27283=>"100111011",
  27284=>"001100001",
  27285=>"100011101",
  27286=>"010011000",
  27287=>"111111100",
  27288=>"010110010",
  27289=>"010111110",
  27290=>"010011110",
  27291=>"101100101",
  27292=>"011010001",
  27293=>"011011100",
  27294=>"111010101",
  27295=>"001001110",
  27296=>"101100011",
  27297=>"110100111",
  27298=>"100010011",
  27299=>"100100101",
  27300=>"000011110",
  27301=>"101000100",
  27302=>"001000101",
  27303=>"111000001",
  27304=>"001101111",
  27305=>"110101111",
  27306=>"010101101",
  27307=>"111111001",
  27308=>"000011000",
  27309=>"111111111",
  27310=>"111110000",
  27311=>"010111010",
  27312=>"101001001",
  27313=>"100010000",
  27314=>"110010010",
  27315=>"010100010",
  27316=>"010010100",
  27317=>"111100111",
  27318=>"110111000",
  27319=>"001111111",
  27320=>"010001100",
  27321=>"000100000",
  27322=>"101010001",
  27323=>"101001111",
  27324=>"010010111",
  27325=>"000010001",
  27326=>"000000001",
  27327=>"110100110",
  27328=>"110000110",
  27329=>"111101111",
  27330=>"110010100",
  27331=>"000110100",
  27332=>"101001110",
  27333=>"001001000",
  27334=>"001000111",
  27335=>"011010010",
  27336=>"000000000",
  27337=>"011110000",
  27338=>"000000011",
  27339=>"000101110",
  27340=>"000100011",
  27341=>"000011000",
  27342=>"101000101",
  27343=>"110011111",
  27344=>"111101101",
  27345=>"111100000",
  27346=>"110110010",
  27347=>"001011000",
  27348=>"001010101",
  27349=>"110000100",
  27350=>"000010100",
  27351=>"010111000",
  27352=>"110110000",
  27353=>"101101111",
  27354=>"000010100",
  27355=>"010000011",
  27356=>"000010010",
  27357=>"001001001",
  27358=>"100001010",
  27359=>"001000011",
  27360=>"100100101",
  27361=>"000010110",
  27362=>"000111100",
  27363=>"010100000",
  27364=>"001001001",
  27365=>"101000001",
  27366=>"001000000",
  27367=>"101010010",
  27368=>"001011111",
  27369=>"000010111",
  27370=>"001100001",
  27371=>"100111111",
  27372=>"010101100",
  27373=>"010100100",
  27374=>"111000000",
  27375=>"110000110",
  27376=>"110100101",
  27377=>"011110001",
  27378=>"101100000",
  27379=>"000010000",
  27380=>"100000110",
  27381=>"100010111",
  27382=>"111110001",
  27383=>"011101000",
  27384=>"101111111",
  27385=>"110110110",
  27386=>"110001010",
  27387=>"001011010",
  27388=>"010101101",
  27389=>"010011000",
  27390=>"010010100",
  27391=>"111010000",
  27392=>"000100110",
  27393=>"110011001",
  27394=>"110111110",
  27395=>"001100001",
  27396=>"100101001",
  27397=>"101101110",
  27398=>"010100011",
  27399=>"000000000",
  27400=>"000101111",
  27401=>"101011011",
  27402=>"101100110",
  27403=>"010010110",
  27404=>"110101000",
  27405=>"110110001",
  27406=>"000100111",
  27407=>"011111110",
  27408=>"101000011",
  27409=>"100001100",
  27410=>"011111011",
  27411=>"000001001",
  27412=>"000011000",
  27413=>"100101101",
  27414=>"010001010",
  27415=>"010100000",
  27416=>"111001110",
  27417=>"100010000",
  27418=>"000100000",
  27419=>"110001100",
  27420=>"101000001",
  27421=>"100011001",
  27422=>"000101011",
  27423=>"010111001",
  27424=>"010010110",
  27425=>"000011000",
  27426=>"001000111",
  27427=>"100100111",
  27428=>"010100101",
  27429=>"100000111",
  27430=>"011111000",
  27431=>"011001011",
  27432=>"111110011",
  27433=>"000010010",
  27434=>"111001101",
  27435=>"000001100",
  27436=>"001110001",
  27437=>"000100100",
  27438=>"011100011",
  27439=>"001111111",
  27440=>"101100000",
  27441=>"101000111",
  27442=>"100101010",
  27443=>"000101110",
  27444=>"100000000",
  27445=>"100100111",
  27446=>"010001111",
  27447=>"001100100",
  27448=>"011011100",
  27449=>"001111101",
  27450=>"011001000",
  27451=>"000101011",
  27452=>"000011110",
  27453=>"110100001",
  27454=>"001000000",
  27455=>"001000011",
  27456=>"110100010",
  27457=>"001000000",
  27458=>"011101010",
  27459=>"111011011",
  27460=>"111001110",
  27461=>"101011100",
  27462=>"101011010",
  27463=>"101111000",
  27464=>"010110011",
  27465=>"011110000",
  27466=>"101010000",
  27467=>"000010101",
  27468=>"001111101",
  27469=>"011011011",
  27470=>"000100011",
  27471=>"001101000",
  27472=>"111100010",
  27473=>"000110101",
  27474=>"000000001",
  27475=>"001001101",
  27476=>"011000011",
  27477=>"010000101",
  27478=>"000100011",
  27479=>"010111111",
  27480=>"001010001",
  27481=>"111000010",
  27482=>"000101001",
  27483=>"110101000",
  27484=>"011111110",
  27485=>"100011110",
  27486=>"110110110",
  27487=>"101011100",
  27488=>"000100000",
  27489=>"011000111",
  27490=>"000000000",
  27491=>"101011001",
  27492=>"101101010",
  27493=>"100000100",
  27494=>"001001000",
  27495=>"010010111",
  27496=>"110100010",
  27497=>"000111010",
  27498=>"001111110",
  27499=>"011101100",
  27500=>"110101010",
  27501=>"000000100",
  27502=>"000101000",
  27503=>"010001110",
  27504=>"011100000",
  27505=>"101100100",
  27506=>"111110110",
  27507=>"100110100",
  27508=>"000110110",
  27509=>"000010101",
  27510=>"101001010",
  27511=>"011011111",
  27512=>"000011000",
  27513=>"011101111",
  27514=>"011101011",
  27515=>"010011101",
  27516=>"011000001",
  27517=>"001100101",
  27518=>"010001001",
  27519=>"110000011",
  27520=>"000000011",
  27521=>"110011100",
  27522=>"000000010",
  27523=>"010010010",
  27524=>"100111001",
  27525=>"011010100",
  27526=>"101000101",
  27527=>"011111110",
  27528=>"111111111",
  27529=>"110010101",
  27530=>"110100110",
  27531=>"001000110",
  27532=>"100001001",
  27533=>"101101011",
  27534=>"000100011",
  27535=>"101011111",
  27536=>"001101001",
  27537=>"001110110",
  27538=>"101000100",
  27539=>"011000100",
  27540=>"010111110",
  27541=>"101110010",
  27542=>"111111110",
  27543=>"001010100",
  27544=>"100110111",
  27545=>"110001000",
  27546=>"000000000",
  27547=>"000111110",
  27548=>"001100000",
  27549=>"011011101",
  27550=>"100111000",
  27551=>"000100000",
  27552=>"101100010",
  27553=>"011111011",
  27554=>"001001111",
  27555=>"110000001",
  27556=>"111000011",
  27557=>"100011111",
  27558=>"100010011",
  27559=>"100110100",
  27560=>"000101000",
  27561=>"000011100",
  27562=>"110110101",
  27563=>"111010110",
  27564=>"001010001",
  27565=>"011000001",
  27566=>"011011101",
  27567=>"011111000",
  27568=>"010010111",
  27569=>"001011011",
  27570=>"101110011",
  27571=>"111000100",
  27572=>"010010111",
  27573=>"111010000",
  27574=>"000000101",
  27575=>"000000100",
  27576=>"001000100",
  27577=>"000011001",
  27578=>"111001010",
  27579=>"100101111",
  27580=>"010011011",
  27581=>"101001011",
  27582=>"001000111",
  27583=>"111111010",
  27584=>"100101001",
  27585=>"111111011",
  27586=>"001000110",
  27587=>"110010100",
  27588=>"001001111",
  27589=>"011010000",
  27590=>"110110110",
  27591=>"010101101",
  27592=>"001110100",
  27593=>"100010101",
  27594=>"111111101",
  27595=>"111100011",
  27596=>"101000111",
  27597=>"010001110",
  27598=>"001001101",
  27599=>"000111110",
  27600=>"101111011",
  27601=>"010100100",
  27602=>"001000111",
  27603=>"110110000",
  27604=>"000011111",
  27605=>"101010000",
  27606=>"010001001",
  27607=>"100110011",
  27608=>"010100111",
  27609=>"110001001",
  27610=>"011100011",
  27611=>"110111111",
  27612=>"010010000",
  27613=>"011100001",
  27614=>"101001111",
  27615=>"000000010",
  27616=>"000111000",
  27617=>"010001110",
  27618=>"001010110",
  27619=>"011110000",
  27620=>"010001110",
  27621=>"101000000",
  27622=>"001100000",
  27623=>"111110001",
  27624=>"011001010",
  27625=>"011011001",
  27626=>"111000000",
  27627=>"100010111",
  27628=>"101101010",
  27629=>"101111111",
  27630=>"000011000",
  27631=>"010010011",
  27632=>"010110000",
  27633=>"010110100",
  27634=>"000010101",
  27635=>"100100011",
  27636=>"110000011",
  27637=>"110100100",
  27638=>"010110001",
  27639=>"000000101",
  27640=>"111100101",
  27641=>"000000000",
  27642=>"100010100",
  27643=>"001100111",
  27644=>"111100100",
  27645=>"110111000",
  27646=>"001100100",
  27647=>"000101111",
  27648=>"100000011",
  27649=>"000110011",
  27650=>"001000101",
  27651=>"110101101",
  27652=>"011111101",
  27653=>"000110011",
  27654=>"010110110",
  27655=>"010110001",
  27656=>"001100010",
  27657=>"010101111",
  27658=>"010011100",
  27659=>"111111000",
  27660=>"011111010",
  27661=>"010111010",
  27662=>"011010101",
  27663=>"110101111",
  27664=>"100101000",
  27665=>"100100111",
  27666=>"110101000",
  27667=>"001111010",
  27668=>"110010101",
  27669=>"000000001",
  27670=>"001000010",
  27671=>"111111001",
  27672=>"100110110",
  27673=>"000101001",
  27674=>"001001101",
  27675=>"001100001",
  27676=>"000101011",
  27677=>"100111100",
  27678=>"011100100",
  27679=>"000111000",
  27680=>"110001100",
  27681=>"011011111",
  27682=>"001000101",
  27683=>"110011100",
  27684=>"010000000",
  27685=>"111111010",
  27686=>"001000001",
  27687=>"111111001",
  27688=>"010100111",
  27689=>"001000111",
  27690=>"001001001",
  27691=>"110111010",
  27692=>"001101000",
  27693=>"001010001",
  27694=>"100101111",
  27695=>"010000010",
  27696=>"001110011",
  27697=>"010111101",
  27698=>"100000010",
  27699=>"010101110",
  27700=>"100110100",
  27701=>"001111111",
  27702=>"000000000",
  27703=>"111010100",
  27704=>"101001100",
  27705=>"000000101",
  27706=>"000100000",
  27707=>"100100001",
  27708=>"011010100",
  27709=>"110111001",
  27710=>"110101001",
  27711=>"010010000",
  27712=>"110110010",
  27713=>"110000000",
  27714=>"100010110",
  27715=>"101010100",
  27716=>"111011100",
  27717=>"100110011",
  27718=>"111101011",
  27719=>"001101000",
  27720=>"111101000",
  27721=>"010001110",
  27722=>"101001000",
  27723=>"100001001",
  27724=>"100010011",
  27725=>"001001011",
  27726=>"001001000",
  27727=>"100101101",
  27728=>"010000010",
  27729=>"000110010",
  27730=>"010111010",
  27731=>"111001101",
  27732=>"010000001",
  27733=>"010000110",
  27734=>"111110011",
  27735=>"100100010",
  27736=>"010110000",
  27737=>"100101010",
  27738=>"000001111",
  27739=>"000100001",
  27740=>"000001101",
  27741=>"101011100",
  27742=>"000000010",
  27743=>"001011110",
  27744=>"000000001",
  27745=>"010000100",
  27746=>"100011111",
  27747=>"100111001",
  27748=>"001001111",
  27749=>"001010101",
  27750=>"111011011",
  27751=>"011100111",
  27752=>"010010110",
  27753=>"010111011",
  27754=>"100000101",
  27755=>"010100001",
  27756=>"001011000",
  27757=>"010100001",
  27758=>"010001100",
  27759=>"101001011",
  27760=>"111101100",
  27761=>"001000001",
  27762=>"001000000",
  27763=>"110000010",
  27764=>"011110101",
  27765=>"101000010",
  27766=>"110011010",
  27767=>"001111101",
  27768=>"101001110",
  27769=>"110000000",
  27770=>"011001000",
  27771=>"010110011",
  27772=>"000101010",
  27773=>"000000010",
  27774=>"000100100",
  27775=>"000011110",
  27776=>"111101010",
  27777=>"000010111",
  27778=>"100111101",
  27779=>"110100111",
  27780=>"011001001",
  27781=>"101111111",
  27782=>"011001111",
  27783=>"101001101",
  27784=>"110111001",
  27785=>"011000101",
  27786=>"010010001",
  27787=>"110011010",
  27788=>"100000000",
  27789=>"111011100",
  27790=>"110000000",
  27791=>"011011100",
  27792=>"101010000",
  27793=>"101101101",
  27794=>"110000101",
  27795=>"100000010",
  27796=>"010101011",
  27797=>"011001001",
  27798=>"100000100",
  27799=>"110001110",
  27800=>"001010111",
  27801=>"000111101",
  27802=>"010011001",
  27803=>"001011100",
  27804=>"010010101",
  27805=>"010010110",
  27806=>"110111011",
  27807=>"011101100",
  27808=>"001111010",
  27809=>"011100010",
  27810=>"001101101",
  27811=>"000000011",
  27812=>"101110011",
  27813=>"111111110",
  27814=>"000010000",
  27815=>"111111111",
  27816=>"111010110",
  27817=>"100011110",
  27818=>"010101011",
  27819=>"011111000",
  27820=>"100011011",
  27821=>"111110101",
  27822=>"110001001",
  27823=>"010000011",
  27824=>"111100011",
  27825=>"110010110",
  27826=>"100111110",
  27827=>"101110010",
  27828=>"000001111",
  27829=>"100101010",
  27830=>"110100010",
  27831=>"001010010",
  27832=>"001100010",
  27833=>"010001001",
  27834=>"110101100",
  27835=>"100011111",
  27836=>"101001000",
  27837=>"101011010",
  27838=>"011110000",
  27839=>"000000110",
  27840=>"101111111",
  27841=>"001100010",
  27842=>"101100101",
  27843=>"100111110",
  27844=>"111001011",
  27845=>"111101000",
  27846=>"101011111",
  27847=>"011100001",
  27848=>"111101000",
  27849=>"011011101",
  27850=>"011100010",
  27851=>"001110111",
  27852=>"011010110",
  27853=>"010111001",
  27854=>"011010001",
  27855=>"000100111",
  27856=>"101011000",
  27857=>"110111100",
  27858=>"101111000",
  27859=>"010110110",
  27860=>"101110110",
  27861=>"100100011",
  27862=>"011111111",
  27863=>"001111001",
  27864=>"100111001",
  27865=>"011000100",
  27866=>"110001101",
  27867=>"000000001",
  27868=>"000001100",
  27869=>"010100111",
  27870=>"001100001",
  27871=>"111001000",
  27872=>"101000011",
  27873=>"000100000",
  27874=>"110010100",
  27875=>"000100001",
  27876=>"000111011",
  27877=>"001000010",
  27878=>"011001100",
  27879=>"000001110",
  27880=>"100110111",
  27881=>"010101100",
  27882=>"000000101",
  27883=>"101101101",
  27884=>"000000000",
  27885=>"001111000",
  27886=>"100001000",
  27887=>"001001100",
  27888=>"011000101",
  27889=>"101111000",
  27890=>"011101000",
  27891=>"010100001",
  27892=>"101110010",
  27893=>"101101000",
  27894=>"110100010",
  27895=>"011100100",
  27896=>"001011000",
  27897=>"011011110",
  27898=>"100101001",
  27899=>"101100101",
  27900=>"010111000",
  27901=>"111010000",
  27902=>"110111100",
  27903=>"001000010",
  27904=>"001100101",
  27905=>"100001011",
  27906=>"111101101",
  27907=>"110001101",
  27908=>"011110011",
  27909=>"011111001",
  27910=>"000000010",
  27911=>"011110110",
  27912=>"010111000",
  27913=>"110101101",
  27914=>"111010011",
  27915=>"101111100",
  27916=>"101100110",
  27917=>"011011110",
  27918=>"111110111",
  27919=>"000010011",
  27920=>"001110111",
  27921=>"010100101",
  27922=>"100101010",
  27923=>"111001100",
  27924=>"010101110",
  27925=>"011101000",
  27926=>"101111101",
  27927=>"101111101",
  27928=>"111100100",
  27929=>"101000110",
  27930=>"000010011",
  27931=>"011101001",
  27932=>"101011110",
  27933=>"111010101",
  27934=>"111010011",
  27935=>"000001001",
  27936=>"011010111",
  27937=>"100101111",
  27938=>"111011011",
  27939=>"101001111",
  27940=>"011010010",
  27941=>"001001000",
  27942=>"100101110",
  27943=>"100111101",
  27944=>"101011011",
  27945=>"110101110",
  27946=>"001000011",
  27947=>"001000100",
  27948=>"111110101",
  27949=>"100100010",
  27950=>"110010001",
  27951=>"100111000",
  27952=>"101010001",
  27953=>"011101010",
  27954=>"100010010",
  27955=>"010100001",
  27956=>"011010111",
  27957=>"010001010",
  27958=>"110100110",
  27959=>"111101001",
  27960=>"111000110",
  27961=>"111001001",
  27962=>"011010111",
  27963=>"101111100",
  27964=>"100100111",
  27965=>"111110010",
  27966=>"101000001",
  27967=>"011001000",
  27968=>"100001111",
  27969=>"100100101",
  27970=>"110000011",
  27971=>"000101101",
  27972=>"111110110",
  27973=>"100000111",
  27974=>"111000100",
  27975=>"001010100",
  27976=>"101100000",
  27977=>"011101000",
  27978=>"100100100",
  27979=>"110011110",
  27980=>"011000001",
  27981=>"010000000",
  27982=>"110111010",
  27983=>"101011011",
  27984=>"000001011",
  27985=>"001111010",
  27986=>"010111000",
  27987=>"000010111",
  27988=>"000101110",
  27989=>"100110110",
  27990=>"000110001",
  27991=>"000101000",
  27992=>"000010101",
  27993=>"100011111",
  27994=>"101101000",
  27995=>"000010000",
  27996=>"111010110",
  27997=>"001111100",
  27998=>"110111110",
  27999=>"001000011",
  28000=>"011011100",
  28001=>"001100011",
  28002=>"000110011",
  28003=>"111100001",
  28004=>"101010010",
  28005=>"110101000",
  28006=>"110101010",
  28007=>"011101101",
  28008=>"001101011",
  28009=>"111110110",
  28010=>"001001101",
  28011=>"110000000",
  28012=>"100110111",
  28013=>"100001011",
  28014=>"110110111",
  28015=>"011110010",
  28016=>"001000111",
  28017=>"111001111",
  28018=>"010110110",
  28019=>"010011101",
  28020=>"000000111",
  28021=>"000100000",
  28022=>"101101100",
  28023=>"100000111",
  28024=>"111001101",
  28025=>"101001010",
  28026=>"111001111",
  28027=>"001001100",
  28028=>"000101101",
  28029=>"000110001",
  28030=>"101001101",
  28031=>"110110010",
  28032=>"001100000",
  28033=>"100000001",
  28034=>"101111010",
  28035=>"110001001",
  28036=>"010000110",
  28037=>"000010010",
  28038=>"100010100",
  28039=>"011011011",
  28040=>"111111001",
  28041=>"001101000",
  28042=>"000101001",
  28043=>"000011011",
  28044=>"001110010",
  28045=>"000000000",
  28046=>"111001111",
  28047=>"001000100",
  28048=>"001000100",
  28049=>"100000100",
  28050=>"111000000",
  28051=>"000000011",
  28052=>"111110010",
  28053=>"001101101",
  28054=>"000110000",
  28055=>"010001100",
  28056=>"011111111",
  28057=>"101110110",
  28058=>"111001001",
  28059=>"000000010",
  28060=>"011101000",
  28061=>"011111011",
  28062=>"110110101",
  28063=>"001000000",
  28064=>"101110101",
  28065=>"110110100",
  28066=>"101111010",
  28067=>"000010010",
  28068=>"111000100",
  28069=>"001111011",
  28070=>"100110100",
  28071=>"001010100",
  28072=>"011001011",
  28073=>"101010110",
  28074=>"110010100",
  28075=>"001000001",
  28076=>"001001100",
  28077=>"110111010",
  28078=>"110010101",
  28079=>"010000100",
  28080=>"010110100",
  28081=>"111011001",
  28082=>"111101111",
  28083=>"001001100",
  28084=>"101011101",
  28085=>"111010001",
  28086=>"100000011",
  28087=>"001101101",
  28088=>"011111010",
  28089=>"111010101",
  28090=>"110111010",
  28091=>"100011011",
  28092=>"110000110",
  28093=>"000000110",
  28094=>"001010100",
  28095=>"101010111",
  28096=>"011101010",
  28097=>"011000011",
  28098=>"010000010",
  28099=>"110010111",
  28100=>"101111110",
  28101=>"100010111",
  28102=>"101010010",
  28103=>"111000011",
  28104=>"011001110",
  28105=>"010110111",
  28106=>"101010111",
  28107=>"100101110",
  28108=>"011111001",
  28109=>"100111011",
  28110=>"101100000",
  28111=>"000011010",
  28112=>"101011101",
  28113=>"011000101",
  28114=>"101010000",
  28115=>"001000100",
  28116=>"111000101",
  28117=>"110011110",
  28118=>"100000000",
  28119=>"000010101",
  28120=>"001111100",
  28121=>"110010111",
  28122=>"000000111",
  28123=>"001111000",
  28124=>"111101100",
  28125=>"010110101",
  28126=>"010001010",
  28127=>"110011100",
  28128=>"010011111",
  28129=>"111011101",
  28130=>"001010101",
  28131=>"110101111",
  28132=>"101110010",
  28133=>"101000110",
  28134=>"101101111",
  28135=>"110110000",
  28136=>"101001010",
  28137=>"111101011",
  28138=>"010110001",
  28139=>"001011010",
  28140=>"101000010",
  28141=>"100101010",
  28142=>"010001111",
  28143=>"010111011",
  28144=>"011011001",
  28145=>"011001101",
  28146=>"000101010",
  28147=>"100100011",
  28148=>"010001001",
  28149=>"100110111",
  28150=>"110010001",
  28151=>"101010010",
  28152=>"011110011",
  28153=>"001110000",
  28154=>"001001111",
  28155=>"100000001",
  28156=>"100111101",
  28157=>"011000001",
  28158=>"000010000",
  28159=>"101010101",
  28160=>"000011101",
  28161=>"101001011",
  28162=>"100011101",
  28163=>"010100110",
  28164=>"010111111",
  28165=>"100011110",
  28166=>"011111000",
  28167=>"111110101",
  28168=>"001111011",
  28169=>"001110010",
  28170=>"110000110",
  28171=>"001111110",
  28172=>"000001110",
  28173=>"000100100",
  28174=>"000011011",
  28175=>"100000110",
  28176=>"100000101",
  28177=>"010010101",
  28178=>"100000101",
  28179=>"110001011",
  28180=>"100011001",
  28181=>"101100010",
  28182=>"010011111",
  28183=>"001010000",
  28184=>"110111001",
  28185=>"110100001",
  28186=>"101101000",
  28187=>"101111110",
  28188=>"011000110",
  28189=>"111001101",
  28190=>"011100000",
  28191=>"111101000",
  28192=>"111100001",
  28193=>"000101110",
  28194=>"100010101",
  28195=>"001111001",
  28196=>"110110110",
  28197=>"000100010",
  28198=>"001111101",
  28199=>"000010000",
  28200=>"001110010",
  28201=>"001100011",
  28202=>"010111011",
  28203=>"101100001",
  28204=>"000110101",
  28205=>"110111111",
  28206=>"001101110",
  28207=>"100011100",
  28208=>"000111011",
  28209=>"010111101",
  28210=>"000111100",
  28211=>"011011111",
  28212=>"110111111",
  28213=>"001100110",
  28214=>"011000110",
  28215=>"010001011",
  28216=>"001100110",
  28217=>"000000111",
  28218=>"010101101",
  28219=>"000011111",
  28220=>"111100001",
  28221=>"010101111",
  28222=>"000011100",
  28223=>"110001000",
  28224=>"010110000",
  28225=>"101110100",
  28226=>"100011001",
  28227=>"011000010",
  28228=>"101110010",
  28229=>"010101110",
  28230=>"100010010",
  28231=>"100010001",
  28232=>"011000111",
  28233=>"011110000",
  28234=>"110110111",
  28235=>"010001011",
  28236=>"011101100",
  28237=>"001010000",
  28238=>"111111101",
  28239=>"000000110",
  28240=>"000111000",
  28241=>"011101111",
  28242=>"110100000",
  28243=>"001110001",
  28244=>"101010101",
  28245=>"101000000",
  28246=>"101010011",
  28247=>"010011000",
  28248=>"110001110",
  28249=>"001101001",
  28250=>"100111111",
  28251=>"001100101",
  28252=>"100000111",
  28253=>"000000010",
  28254=>"010010010",
  28255=>"010101001",
  28256=>"011100100",
  28257=>"000001000",
  28258=>"110001010",
  28259=>"100100101",
  28260=>"110001000",
  28261=>"111001011",
  28262=>"001000011",
  28263=>"111111011",
  28264=>"110001110",
  28265=>"100100100",
  28266=>"111010100",
  28267=>"100001010",
  28268=>"010001011",
  28269=>"100010111",
  28270=>"110000011",
  28271=>"000100001",
  28272=>"110100110",
  28273=>"101100001",
  28274=>"111001111",
  28275=>"101010111",
  28276=>"011111000",
  28277=>"010000110",
  28278=>"111011100",
  28279=>"110001110",
  28280=>"100100000",
  28281=>"100001101",
  28282=>"101111001",
  28283=>"101111010",
  28284=>"000010101",
  28285=>"100000000",
  28286=>"011011101",
  28287=>"001011100",
  28288=>"001001110",
  28289=>"111010001",
  28290=>"111100010",
  28291=>"001001010",
  28292=>"101001101",
  28293=>"100100100",
  28294=>"101010100",
  28295=>"110100011",
  28296=>"100011010",
  28297=>"111100111",
  28298=>"010001110",
  28299=>"010110001",
  28300=>"101110001",
  28301=>"000101011",
  28302=>"101001000",
  28303=>"101000011",
  28304=>"000000001",
  28305=>"000001111",
  28306=>"011100010",
  28307=>"101011111",
  28308=>"001010010",
  28309=>"110111100",
  28310=>"110000101",
  28311=>"001110110",
  28312=>"001101111",
  28313=>"111101011",
  28314=>"110001001",
  28315=>"011000110",
  28316=>"010011000",
  28317=>"000010010",
  28318=>"110110000",
  28319=>"000111110",
  28320=>"101011001",
  28321=>"010111011",
  28322=>"001110100",
  28323=>"100110010",
  28324=>"000001110",
  28325=>"000110101",
  28326=>"100011110",
  28327=>"110000111",
  28328=>"010111100",
  28329=>"011011111",
  28330=>"101001011",
  28331=>"000000100",
  28332=>"011110101",
  28333=>"001100001",
  28334=>"000110110",
  28335=>"010110011",
  28336=>"000011011",
  28337=>"000000100",
  28338=>"010011011",
  28339=>"011010111",
  28340=>"101111101",
  28341=>"111111101",
  28342=>"000010101",
  28343=>"111111001",
  28344=>"101100110",
  28345=>"010001101",
  28346=>"101110011",
  28347=>"000000111",
  28348=>"001010110",
  28349=>"011101001",
  28350=>"101011011",
  28351=>"000011101",
  28352=>"111010010",
  28353=>"101110111",
  28354=>"011100100",
  28355=>"010011101",
  28356=>"001101010",
  28357=>"001011111",
  28358=>"011001101",
  28359=>"001000110",
  28360=>"000101000",
  28361=>"100000010",
  28362=>"001110101",
  28363=>"101001001",
  28364=>"000000011",
  28365=>"110001101",
  28366=>"111011110",
  28367=>"100101101",
  28368=>"011100010",
  28369=>"101010101",
  28370=>"101010100",
  28371=>"101101100",
  28372=>"000110000",
  28373=>"110110110",
  28374=>"111011000",
  28375=>"011111001",
  28376=>"101101101",
  28377=>"110111111",
  28378=>"010110000",
  28379=>"000100100",
  28380=>"100100011",
  28381=>"000110011",
  28382=>"100101001",
  28383=>"001100010",
  28384=>"100000111",
  28385=>"011011110",
  28386=>"010000011",
  28387=>"000111001",
  28388=>"101001111",
  28389=>"000001000",
  28390=>"001011010",
  28391=>"111101000",
  28392=>"001101100",
  28393=>"101110011",
  28394=>"011110000",
  28395=>"001101111",
  28396=>"001101110",
  28397=>"001111000",
  28398=>"110011100",
  28399=>"011100000",
  28400=>"010110001",
  28401=>"111010110",
  28402=>"001011111",
  28403=>"110011100",
  28404=>"001100101",
  28405=>"011001011",
  28406=>"101000001",
  28407=>"000001101",
  28408=>"010010100",
  28409=>"100010100",
  28410=>"011011000",
  28411=>"010100001",
  28412=>"010100110",
  28413=>"000010011",
  28414=>"001001001",
  28415=>"000010110",
  28416=>"001010101",
  28417=>"111111100",
  28418=>"111111100",
  28419=>"110011000",
  28420=>"010010010",
  28421=>"000011111",
  28422=>"001100100",
  28423=>"000110100",
  28424=>"001000000",
  28425=>"001100000",
  28426=>"101010110",
  28427=>"001100000",
  28428=>"011100010",
  28429=>"101111100",
  28430=>"001100010",
  28431=>"001111101",
  28432=>"110000100",
  28433=>"101001110",
  28434=>"000010000",
  28435=>"101110001",
  28436=>"100110110",
  28437=>"010000100",
  28438=>"010010100",
  28439=>"001011011",
  28440=>"101110100",
  28441=>"011111110",
  28442=>"110101001",
  28443=>"011011000",
  28444=>"000110101",
  28445=>"001011101",
  28446=>"010111000",
  28447=>"001110111",
  28448=>"011110111",
  28449=>"011111010",
  28450=>"101101111",
  28451=>"111010011",
  28452=>"111010001",
  28453=>"111101010",
  28454=>"010000011",
  28455=>"101111000",
  28456=>"001110110",
  28457=>"000101110",
  28458=>"110110100",
  28459=>"000100000",
  28460=>"010100010",
  28461=>"010000101",
  28462=>"111101100",
  28463=>"001010011",
  28464=>"100000011",
  28465=>"001000101",
  28466=>"000111010",
  28467=>"100010111",
  28468=>"100011010",
  28469=>"100010110",
  28470=>"000010011",
  28471=>"011000010",
  28472=>"001011111",
  28473=>"000000000",
  28474=>"010101101",
  28475=>"011011001",
  28476=>"000000100",
  28477=>"001011000",
  28478=>"110100110",
  28479=>"010101100",
  28480=>"011111101",
  28481=>"011001000",
  28482=>"001001011",
  28483=>"001101011",
  28484=>"011100110",
  28485=>"111010001",
  28486=>"110101100",
  28487=>"111000000",
  28488=>"110101111",
  28489=>"101001010",
  28490=>"111100001",
  28491=>"000010011",
  28492=>"001101110",
  28493=>"011001111",
  28494=>"110011001",
  28495=>"110011010",
  28496=>"001010011",
  28497=>"111100111",
  28498=>"011000010",
  28499=>"000001000",
  28500=>"110011000",
  28501=>"110001010",
  28502=>"000000000",
  28503=>"010011100",
  28504=>"000110111",
  28505=>"010101000",
  28506=>"011110001",
  28507=>"101000101",
  28508=>"011100001",
  28509=>"000010010",
  28510=>"110110111",
  28511=>"100100101",
  28512=>"100000100",
  28513=>"010000001",
  28514=>"111110100",
  28515=>"010100111",
  28516=>"011011000",
  28517=>"001000000",
  28518=>"101000001",
  28519=>"101111110",
  28520=>"000111100",
  28521=>"100100100",
  28522=>"101101011",
  28523=>"010110100",
  28524=>"001111111",
  28525=>"100010010",
  28526=>"111011010",
  28527=>"101011000",
  28528=>"111111101",
  28529=>"000001101",
  28530=>"110001110",
  28531=>"011010010",
  28532=>"010111001",
  28533=>"001101011",
  28534=>"001010101",
  28535=>"010011110",
  28536=>"101101100",
  28537=>"001101001",
  28538=>"111011001",
  28539=>"100111001",
  28540=>"100101101",
  28541=>"000111111",
  28542=>"001100010",
  28543=>"111111011",
  28544=>"101010110",
  28545=>"001010010",
  28546=>"111010110",
  28547=>"010000111",
  28548=>"000011010",
  28549=>"010110001",
  28550=>"010000110",
  28551=>"110010001",
  28552=>"101010100",
  28553=>"100000011",
  28554=>"110101111",
  28555=>"001010101",
  28556=>"001000111",
  28557=>"001100001",
  28558=>"000100100",
  28559=>"000100111",
  28560=>"111001000",
  28561=>"111111111",
  28562=>"011011111",
  28563=>"111010101",
  28564=>"011010100",
  28565=>"000111011",
  28566=>"100100000",
  28567=>"101000010",
  28568=>"001001000",
  28569=>"110000111",
  28570=>"111110101",
  28571=>"010111000",
  28572=>"001110111",
  28573=>"000110010",
  28574=>"000110010",
  28575=>"110011110",
  28576=>"111110111",
  28577=>"011010111",
  28578=>"011011111",
  28579=>"011100010",
  28580=>"011000100",
  28581=>"101101011",
  28582=>"111110010",
  28583=>"100111111",
  28584=>"100111110",
  28585=>"101110000",
  28586=>"010101111",
  28587=>"100001100",
  28588=>"000000011",
  28589=>"000100010",
  28590=>"110101001",
  28591=>"101110100",
  28592=>"001001000",
  28593=>"100101011",
  28594=>"011101101",
  28595=>"101001101",
  28596=>"111011011",
  28597=>"011011110",
  28598=>"111011010",
  28599=>"100100111",
  28600=>"000101111",
  28601=>"000101110",
  28602=>"001000111",
  28603=>"000110011",
  28604=>"000100001",
  28605=>"001010000",
  28606=>"001110101",
  28607=>"010110101",
  28608=>"110011001",
  28609=>"110110011",
  28610=>"110011000",
  28611=>"111100011",
  28612=>"110100100",
  28613=>"000011111",
  28614=>"110001110",
  28615=>"010110000",
  28616=>"100100111",
  28617=>"101000001",
  28618=>"001001101",
  28619=>"011100001",
  28620=>"001110100",
  28621=>"010100010",
  28622=>"000100010",
  28623=>"110101010",
  28624=>"011010110",
  28625=>"001000011",
  28626=>"000001111",
  28627=>"101000110",
  28628=>"000110101",
  28629=>"011110010",
  28630=>"110010111",
  28631=>"001110111",
  28632=>"111110011",
  28633=>"111111011",
  28634=>"101110000",
  28635=>"010101101",
  28636=>"010000101",
  28637=>"001000111",
  28638=>"101010011",
  28639=>"010110001",
  28640=>"101100000",
  28641=>"101100100",
  28642=>"101100100",
  28643=>"000110110",
  28644=>"100010101",
  28645=>"011000101",
  28646=>"010110010",
  28647=>"011110111",
  28648=>"000111100",
  28649=>"100111001",
  28650=>"101100101",
  28651=>"111100101",
  28652=>"010010001",
  28653=>"000111110",
  28654=>"100110000",
  28655=>"001000111",
  28656=>"111001000",
  28657=>"011010100",
  28658=>"011101011",
  28659=>"010110100",
  28660=>"010111101",
  28661=>"101001111",
  28662=>"010011011",
  28663=>"111101001",
  28664=>"010110110",
  28665=>"100011011",
  28666=>"000110111",
  28667=>"001100100",
  28668=>"010101100",
  28669=>"000000110",
  28670=>"110110110",
  28671=>"001110100",
  28672=>"011001111",
  28673=>"100011001",
  28674=>"100111100",
  28675=>"111001011",
  28676=>"001101001",
  28677=>"001010011",
  28678=>"100000000",
  28679=>"001000100",
  28680=>"010101101",
  28681=>"100001111",
  28682=>"111100110",
  28683=>"111010001",
  28684=>"101010001",
  28685=>"001111100",
  28686=>"001100001",
  28687=>"110011000",
  28688=>"101101000",
  28689=>"001010001",
  28690=>"101010111",
  28691=>"011000110",
  28692=>"101001110",
  28693=>"001110000",
  28694=>"111011101",
  28695=>"100010110",
  28696=>"111101111",
  28697=>"111101111",
  28698=>"101000001",
  28699=>"001011111",
  28700=>"101100011",
  28701=>"010111111",
  28702=>"010000001",
  28703=>"000011111",
  28704=>"010010001",
  28705=>"011110010",
  28706=>"000001101",
  28707=>"100000001",
  28708=>"010010111",
  28709=>"100010111",
  28710=>"010110111",
  28711=>"100110110",
  28712=>"100100010",
  28713=>"101011110",
  28714=>"010110011",
  28715=>"010111101",
  28716=>"101000101",
  28717=>"001000101",
  28718=>"101010000",
  28719=>"111111111",
  28720=>"110100011",
  28721=>"011010110",
  28722=>"000000110",
  28723=>"111101110",
  28724=>"110001011",
  28725=>"101111011",
  28726=>"001100110",
  28727=>"011101101",
  28728=>"011101010",
  28729=>"100111001",
  28730=>"111000010",
  28731=>"111110010",
  28732=>"010010001",
  28733=>"010111100",
  28734=>"101111000",
  28735=>"110011001",
  28736=>"111011000",
  28737=>"101111111",
  28738=>"001110111",
  28739=>"100011000",
  28740=>"111111001",
  28741=>"100100000",
  28742=>"000000001",
  28743=>"110010101",
  28744=>"100000010",
  28745=>"101001010",
  28746=>"010000111",
  28747=>"101100100",
  28748=>"110000011",
  28749=>"010001110",
  28750=>"101000010",
  28751=>"111110001",
  28752=>"101100111",
  28753=>"110101110",
  28754=>"000011010",
  28755=>"111011100",
  28756=>"000111011",
  28757=>"011011111",
  28758=>"011101111",
  28759=>"001010011",
  28760=>"100001000",
  28761=>"100011011",
  28762=>"001110110",
  28763=>"111110100",
  28764=>"101000100",
  28765=>"001100001",
  28766=>"100110101",
  28767=>"101000000",
  28768=>"010101100",
  28769=>"110000100",
  28770=>"101101000",
  28771=>"010100010",
  28772=>"110000110",
  28773=>"010111101",
  28774=>"111101111",
  28775=>"001100111",
  28776=>"101001100",
  28777=>"010111100",
  28778=>"000100010",
  28779=>"100100011",
  28780=>"001000100",
  28781=>"101101101",
  28782=>"110001010",
  28783=>"100100111",
  28784=>"101010101",
  28785=>"001000100",
  28786=>"010110100",
  28787=>"010010011",
  28788=>"111001001",
  28789=>"110001001",
  28790=>"101011010",
  28791=>"010001111",
  28792=>"000110110",
  28793=>"100110111",
  28794=>"001000011",
  28795=>"111111100",
  28796=>"011000111",
  28797=>"001001000",
  28798=>"111100000",
  28799=>"100100111",
  28800=>"000110111",
  28801=>"100101100",
  28802=>"001000001",
  28803=>"100001101",
  28804=>"011000000",
  28805=>"101000010",
  28806=>"000101011",
  28807=>"011101100",
  28808=>"111111011",
  28809=>"010110010",
  28810=>"110011011",
  28811=>"010111010",
  28812=>"001111101",
  28813=>"000000010",
  28814=>"000111000",
  28815=>"110111100",
  28816=>"100000111",
  28817=>"010101111",
  28818=>"101110010",
  28819=>"100100111",
  28820=>"110010100",
  28821=>"100110011",
  28822=>"010001101",
  28823=>"111011011",
  28824=>"011110100",
  28825=>"111001111",
  28826=>"110101100",
  28827=>"111111111",
  28828=>"011100010",
  28829=>"110100110",
  28830=>"111100110",
  28831=>"100010100",
  28832=>"010011111",
  28833=>"110000101",
  28834=>"001001010",
  28835=>"101001001",
  28836=>"010110111",
  28837=>"001001101",
  28838=>"100010000",
  28839=>"100101000",
  28840=>"111010101",
  28841=>"111010011",
  28842=>"011010011",
  28843=>"010100101",
  28844=>"101000000",
  28845=>"011000000",
  28846=>"010101010",
  28847=>"000101011",
  28848=>"000010110",
  28849=>"111001001",
  28850=>"101100011",
  28851=>"100101100",
  28852=>"010000100",
  28853=>"000000001",
  28854=>"110001111",
  28855=>"110011001",
  28856=>"000110011",
  28857=>"011100101",
  28858=>"001000010",
  28859=>"001011000",
  28860=>"110100000",
  28861=>"101001100",
  28862=>"010000101",
  28863=>"110101111",
  28864=>"001110010",
  28865=>"001111111",
  28866=>"110001010",
  28867=>"111011000",
  28868=>"010111000",
  28869=>"000110100",
  28870=>"100100010",
  28871=>"000100000",
  28872=>"111011011",
  28873=>"011101100",
  28874=>"110110001",
  28875=>"111110111",
  28876=>"110000111",
  28877=>"101001000",
  28878=>"010000010",
  28879=>"101011101",
  28880=>"011110111",
  28881=>"010111011",
  28882=>"001110000",
  28883=>"000000111",
  28884=>"011110110",
  28885=>"110010000",
  28886=>"000011111",
  28887=>"110010010",
  28888=>"001101010",
  28889=>"011000101",
  28890=>"001111001",
  28891=>"000011010",
  28892=>"010000010",
  28893=>"000011110",
  28894=>"100111101",
  28895=>"110110000",
  28896=>"000001101",
  28897=>"100101111",
  28898=>"001100011",
  28899=>"100111111",
  28900=>"110111010",
  28901=>"111000110",
  28902=>"010000000",
  28903=>"100110011",
  28904=>"000010100",
  28905=>"100000111",
  28906=>"111111111",
  28907=>"100010110",
  28908=>"111101101",
  28909=>"010010011",
  28910=>"000100011",
  28911=>"001110010",
  28912=>"011011100",
  28913=>"111010111",
  28914=>"110000000",
  28915=>"111100100",
  28916=>"010111110",
  28917=>"111001001",
  28918=>"110011111",
  28919=>"100001100",
  28920=>"100101110",
  28921=>"101100100",
  28922=>"000011100",
  28923=>"000111110",
  28924=>"100000010",
  28925=>"111100011",
  28926=>"001010101",
  28927=>"101001011",
  28928=>"101110001",
  28929=>"010111100",
  28930=>"001000100",
  28931=>"000000111",
  28932=>"010101001",
  28933=>"101100000",
  28934=>"100010010",
  28935=>"111001101",
  28936=>"001010011",
  28937=>"001100100",
  28938=>"110000110",
  28939=>"000001110",
  28940=>"110001010",
  28941=>"010111011",
  28942=>"000111010",
  28943=>"110001010",
  28944=>"011000110",
  28945=>"111100001",
  28946=>"100011111",
  28947=>"110110000",
  28948=>"100110101",
  28949=>"101001001",
  28950=>"010101011",
  28951=>"001101010",
  28952=>"011100001",
  28953=>"010110000",
  28954=>"010100100",
  28955=>"101001000",
  28956=>"101011111",
  28957=>"010100000",
  28958=>"100010101",
  28959=>"101110001",
  28960=>"110111010",
  28961=>"000110010",
  28962=>"000001010",
  28963=>"100110101",
  28964=>"101011101",
  28965=>"101010001",
  28966=>"000001010",
  28967=>"000001110",
  28968=>"100100000",
  28969=>"000101001",
  28970=>"101100001",
  28971=>"000100111",
  28972=>"111100000",
  28973=>"100110111",
  28974=>"111000010",
  28975=>"111111001",
  28976=>"111100101",
  28977=>"011101111",
  28978=>"100001011",
  28979=>"100111110",
  28980=>"110110101",
  28981=>"010010111",
  28982=>"011111000",
  28983=>"101100001",
  28984=>"010101001",
  28985=>"110010011",
  28986=>"100011111",
  28987=>"010101010",
  28988=>"100011101",
  28989=>"001001001",
  28990=>"000100000",
  28991=>"100000010",
  28992=>"010101100",
  28993=>"010010111",
  28994=>"110110010",
  28995=>"001001100",
  28996=>"100110110",
  28997=>"101101101",
  28998=>"100100001",
  28999=>"001111111",
  29000=>"011011001",
  29001=>"110000110",
  29002=>"001010001",
  29003=>"001111010",
  29004=>"011110100",
  29005=>"011000001",
  29006=>"010011001",
  29007=>"011110001",
  29008=>"010111000",
  29009=>"101110110",
  29010=>"010010011",
  29011=>"010001011",
  29012=>"001110001",
  29013=>"101111101",
  29014=>"101111111",
  29015=>"101111001",
  29016=>"010000100",
  29017=>"010100111",
  29018=>"011010100",
  29019=>"111010001",
  29020=>"000111101",
  29021=>"000100111",
  29022=>"010001101",
  29023=>"101011000",
  29024=>"000101000",
  29025=>"111000100",
  29026=>"011110101",
  29027=>"010100101",
  29028=>"110000110",
  29029=>"001111011",
  29030=>"010011110",
  29031=>"001100000",
  29032=>"110000010",
  29033=>"010000111",
  29034=>"000000100",
  29035=>"000000110",
  29036=>"110001000",
  29037=>"111010001",
  29038=>"000001010",
  29039=>"000100101",
  29040=>"101101101",
  29041=>"101011000",
  29042=>"011010000",
  29043=>"101111011",
  29044=>"001000000",
  29045=>"101000000",
  29046=>"011101111",
  29047=>"001110111",
  29048=>"111011111",
  29049=>"000111100",
  29050=>"010000111",
  29051=>"101001000",
  29052=>"100111100",
  29053=>"010000110",
  29054=>"000100111",
  29055=>"011110001",
  29056=>"000010010",
  29057=>"111010010",
  29058=>"101011010",
  29059=>"000100001",
  29060=>"011010010",
  29061=>"001000001",
  29062=>"100111001",
  29063=>"110001010",
  29064=>"000001010",
  29065=>"011001100",
  29066=>"001010001",
  29067=>"101011100",
  29068=>"111101010",
  29069=>"100010011",
  29070=>"010010100",
  29071=>"111110101",
  29072=>"100100101",
  29073=>"000010010",
  29074=>"000000001",
  29075=>"100010011",
  29076=>"011010111",
  29077=>"000010101",
  29078=>"001100011",
  29079=>"001110101",
  29080=>"001000111",
  29081=>"001000101",
  29082=>"101110110",
  29083=>"111100001",
  29084=>"101001010",
  29085=>"111010101",
  29086=>"011000100",
  29087=>"110000101",
  29088=>"011100001",
  29089=>"001011000",
  29090=>"001000000",
  29091=>"001101001",
  29092=>"011100011",
  29093=>"011011100",
  29094=>"001000011",
  29095=>"100001000",
  29096=>"111010100",
  29097=>"101101110",
  29098=>"100110111",
  29099=>"111110010",
  29100=>"110001101",
  29101=>"100010010",
  29102=>"001001111",
  29103=>"001010100",
  29104=>"010110100",
  29105=>"000011011",
  29106=>"111111111",
  29107=>"001101100",
  29108=>"100001110",
  29109=>"010010100",
  29110=>"010101001",
  29111=>"111111010",
  29112=>"111101101",
  29113=>"111001010",
  29114=>"110101000",
  29115=>"010011001",
  29116=>"011111111",
  29117=>"101100110",
  29118=>"111100011",
  29119=>"000001011",
  29120=>"010001010",
  29121=>"101101001",
  29122=>"111111110",
  29123=>"100111001",
  29124=>"001010100",
  29125=>"000011001",
  29126=>"100101101",
  29127=>"101000111",
  29128=>"000001111",
  29129=>"010010111",
  29130=>"110001010",
  29131=>"010011111",
  29132=>"000100101",
  29133=>"011000111",
  29134=>"010010011",
  29135=>"101111011",
  29136=>"111010010",
  29137=>"001000110",
  29138=>"011110110",
  29139=>"111001010",
  29140=>"000110111",
  29141=>"011001010",
  29142=>"101101100",
  29143=>"001110111",
  29144=>"000101111",
  29145=>"010100001",
  29146=>"010001011",
  29147=>"010110001",
  29148=>"110111110",
  29149=>"001100011",
  29150=>"111000110",
  29151=>"000100001",
  29152=>"011001111",
  29153=>"010110000",
  29154=>"110100100",
  29155=>"101101001",
  29156=>"001100110",
  29157=>"101111011",
  29158=>"001100100",
  29159=>"001100000",
  29160=>"110001000",
  29161=>"111110100",
  29162=>"110101110",
  29163=>"001010101",
  29164=>"000111100",
  29165=>"111011010",
  29166=>"010010100",
  29167=>"000001100",
  29168=>"011011111",
  29169=>"001100000",
  29170=>"000111010",
  29171=>"000010000",
  29172=>"101101000",
  29173=>"000111011",
  29174=>"110111000",
  29175=>"101101100",
  29176=>"111100011",
  29177=>"110000100",
  29178=>"101010001",
  29179=>"001111001",
  29180=>"000000011",
  29181=>"111101011",
  29182=>"000100111",
  29183=>"101011110",
  29184=>"101010101",
  29185=>"111011100",
  29186=>"000100011",
  29187=>"101111111",
  29188=>"011000110",
  29189=>"111101011",
  29190=>"111110011",
  29191=>"101010011",
  29192=>"100111110",
  29193=>"001010000",
  29194=>"101000111",
  29195=>"000111001",
  29196=>"101011100",
  29197=>"000101100",
  29198=>"101001001",
  29199=>"100000001",
  29200=>"101110111",
  29201=>"001000011",
  29202=>"111100010",
  29203=>"011010010",
  29204=>"101001101",
  29205=>"001100101",
  29206=>"001111110",
  29207=>"101111111",
  29208=>"110111010",
  29209=>"100000101",
  29210=>"001001001",
  29211=>"000010001",
  29212=>"010001011",
  29213=>"010000110",
  29214=>"100011110",
  29215=>"101101100",
  29216=>"110100100",
  29217=>"000000000",
  29218=>"001001101",
  29219=>"000111001",
  29220=>"010111111",
  29221=>"100010001",
  29222=>"110101011",
  29223=>"100101000",
  29224=>"100101110",
  29225=>"000110010",
  29226=>"010010011",
  29227=>"011111110",
  29228=>"000100000",
  29229=>"000011101",
  29230=>"110110000",
  29231=>"001101010",
  29232=>"010101101",
  29233=>"100101111",
  29234=>"000000110",
  29235=>"110100111",
  29236=>"011010000",
  29237=>"010110100",
  29238=>"110001101",
  29239=>"011111110",
  29240=>"110110110",
  29241=>"110101110",
  29242=>"010111011",
  29243=>"100010110",
  29244=>"011000001",
  29245=>"111110100",
  29246=>"101000100",
  29247=>"011101010",
  29248=>"100100011",
  29249=>"111011000",
  29250=>"001000011",
  29251=>"110110011",
  29252=>"001101000",
  29253=>"011111001",
  29254=>"000000000",
  29255=>"000011101",
  29256=>"111110000",
  29257=>"100110111",
  29258=>"001000100",
  29259=>"000110111",
  29260=>"110000000",
  29261=>"000100111",
  29262=>"101001001",
  29263=>"010111110",
  29264=>"000111101",
  29265=>"010010101",
  29266=>"000001001",
  29267=>"001001000",
  29268=>"110000100",
  29269=>"000011011",
  29270=>"001111100",
  29271=>"000100011",
  29272=>"111100011",
  29273=>"101001001",
  29274=>"011100101",
  29275=>"000100111",
  29276=>"100010000",
  29277=>"001111100",
  29278=>"010111110",
  29279=>"100100111",
  29280=>"110001011",
  29281=>"000010100",
  29282=>"100101101",
  29283=>"001001011",
  29284=>"101011100",
  29285=>"011110100",
  29286=>"011010110",
  29287=>"110011000",
  29288=>"110000010",
  29289=>"011001000",
  29290=>"000111001",
  29291=>"111001101",
  29292=>"011010000",
  29293=>"101011000",
  29294=>"001111101",
  29295=>"010011101",
  29296=>"111000111",
  29297=>"011100110",
  29298=>"010000101",
  29299=>"110011111",
  29300=>"100010000",
  29301=>"000001111",
  29302=>"000001101",
  29303=>"110011111",
  29304=>"100100111",
  29305=>"100011001",
  29306=>"000110001",
  29307=>"110100001",
  29308=>"000110000",
  29309=>"110010110",
  29310=>"101100011",
  29311=>"111100101",
  29312=>"001100110",
  29313=>"010100000",
  29314=>"110110110",
  29315=>"100001011",
  29316=>"011100011",
  29317=>"100100000",
  29318=>"001111110",
  29319=>"000100000",
  29320=>"110100100",
  29321=>"000010101",
  29322=>"101111110",
  29323=>"010111100",
  29324=>"101100100",
  29325=>"101011011",
  29326=>"100010001",
  29327=>"000111110",
  29328=>"101001111",
  29329=>"101110100",
  29330=>"100101011",
  29331=>"000001010",
  29332=>"000000110",
  29333=>"010000101",
  29334=>"111100100",
  29335=>"100001111",
  29336=>"101110111",
  29337=>"001101111",
  29338=>"000101110",
  29339=>"001010001",
  29340=>"001000001",
  29341=>"110101111",
  29342=>"011101011",
  29343=>"110001001",
  29344=>"111001111",
  29345=>"111011111",
  29346=>"010000001",
  29347=>"010101001",
  29348=>"100100010",
  29349=>"111101011",
  29350=>"010001110",
  29351=>"000101010",
  29352=>"100101010",
  29353=>"000110000",
  29354=>"011011110",
  29355=>"101011000",
  29356=>"111100011",
  29357=>"110111111",
  29358=>"100100001",
  29359=>"100001001",
  29360=>"001010110",
  29361=>"101000111",
  29362=>"101110100",
  29363=>"110101111",
  29364=>"110101111",
  29365=>"100101000",
  29366=>"010010001",
  29367=>"011000101",
  29368=>"101000100",
  29369=>"100010111",
  29370=>"000100000",
  29371=>"111101011",
  29372=>"110001111",
  29373=>"100110000",
  29374=>"001101100",
  29375=>"111101000",
  29376=>"100111010",
  29377=>"000101100",
  29378=>"000010001",
  29379=>"100110100",
  29380=>"000110111",
  29381=>"100000111",
  29382=>"010011000",
  29383=>"110001100",
  29384=>"110010011",
  29385=>"110110111",
  29386=>"101101000",
  29387=>"110010001",
  29388=>"110110001",
  29389=>"001101110",
  29390=>"101101001",
  29391=>"110010111",
  29392=>"100100000",
  29393=>"110010010",
  29394=>"011101001",
  29395=>"001100000",
  29396=>"000000101",
  29397=>"001101101",
  29398=>"001111110",
  29399=>"000111100",
  29400=>"000011110",
  29401=>"110011100",
  29402=>"111000000",
  29403=>"000001010",
  29404=>"101011101",
  29405=>"001011011",
  29406=>"001111110",
  29407=>"100001101",
  29408=>"000100111",
  29409=>"011100011",
  29410=>"011011110",
  29411=>"110110110",
  29412=>"001111000",
  29413=>"110111001",
  29414=>"010001111",
  29415=>"001000011",
  29416=>"100010100",
  29417=>"010100111",
  29418=>"101000000",
  29419=>"001101000",
  29420=>"011001001",
  29421=>"000011111",
  29422=>"110111111",
  29423=>"010110101",
  29424=>"110010101",
  29425=>"011000000",
  29426=>"111101000",
  29427=>"111100110",
  29428=>"110111000",
  29429=>"101100101",
  29430=>"011111000",
  29431=>"000000010",
  29432=>"011011100",
  29433=>"000001110",
  29434=>"111110100",
  29435=>"100000000",
  29436=>"101100100",
  29437=>"101010010",
  29438=>"010001110",
  29439=>"100110101",
  29440=>"100100100",
  29441=>"110000011",
  29442=>"110010011",
  29443=>"010110011",
  29444=>"000101101",
  29445=>"000001101",
  29446=>"011001010",
  29447=>"100000001",
  29448=>"110101010",
  29449=>"010110100",
  29450=>"000100101",
  29451=>"001101111",
  29452=>"000000100",
  29453=>"010000010",
  29454=>"101010100",
  29455=>"010110110",
  29456=>"001110010",
  29457=>"100011010",
  29458=>"010011110",
  29459=>"001100011",
  29460=>"010100110",
  29461=>"110010000",
  29462=>"101100110",
  29463=>"110001100",
  29464=>"001011010",
  29465=>"001011011",
  29466=>"000100111",
  29467=>"111001011",
  29468=>"110101101",
  29469=>"000111010",
  29470=>"100001010",
  29471=>"111001101",
  29472=>"110010110",
  29473=>"010100000",
  29474=>"100001100",
  29475=>"100111101",
  29476=>"010010111",
  29477=>"011111111",
  29478=>"010100000",
  29479=>"011100110",
  29480=>"101011001",
  29481=>"101010001",
  29482=>"011111001",
  29483=>"000001010",
  29484=>"100111010",
  29485=>"000001111",
  29486=>"111000100",
  29487=>"010000111",
  29488=>"011101101",
  29489=>"001011101",
  29490=>"010001000",
  29491=>"000000111",
  29492=>"111001001",
  29493=>"100101010",
  29494=>"011111101",
  29495=>"011100111",
  29496=>"111011000",
  29497=>"011001011",
  29498=>"000111111",
  29499=>"000110101",
  29500=>"111000000",
  29501=>"000101011",
  29502=>"111011111",
  29503=>"100111101",
  29504=>"010001011",
  29505=>"001110000",
  29506=>"011110111",
  29507=>"010010100",
  29508=>"010010001",
  29509=>"111111110",
  29510=>"100001101",
  29511=>"101110111",
  29512=>"010111101",
  29513=>"010011001",
  29514=>"010101001",
  29515=>"001001000",
  29516=>"010110100",
  29517=>"100111100",
  29518=>"000011111",
  29519=>"101101010",
  29520=>"111101110",
  29521=>"110101100",
  29522=>"100010010",
  29523=>"011001001",
  29524=>"001110100",
  29525=>"001110101",
  29526=>"011010011",
  29527=>"111111011",
  29528=>"101100110",
  29529=>"011010000",
  29530=>"001001110",
  29531=>"111110111",
  29532=>"100010100",
  29533=>"000001101",
  29534=>"100100111",
  29535=>"000000011",
  29536=>"001000100",
  29537=>"111010111",
  29538=>"111110011",
  29539=>"010000011",
  29540=>"000111101",
  29541=>"011100000",
  29542=>"101011101",
  29543=>"010001000",
  29544=>"011110010",
  29545=>"101010000",
  29546=>"110110100",
  29547=>"001101011",
  29548=>"101011100",
  29549=>"000000010",
  29550=>"110000111",
  29551=>"000010110",
  29552=>"100000010",
  29553=>"000000000",
  29554=>"100010101",
  29555=>"011010110",
  29556=>"110000100",
  29557=>"001010000",
  29558=>"100101010",
  29559=>"001101011",
  29560=>"010110100",
  29561=>"111100111",
  29562=>"100101001",
  29563=>"001110010",
  29564=>"000000111",
  29565=>"111001001",
  29566=>"100100111",
  29567=>"110100011",
  29568=>"100000100",
  29569=>"000000011",
  29570=>"001001101",
  29571=>"101011111",
  29572=>"111000000",
  29573=>"100011101",
  29574=>"101001100",
  29575=>"100011011",
  29576=>"100011011",
  29577=>"010111000",
  29578=>"011101110",
  29579=>"100110111",
  29580=>"100000101",
  29581=>"111101010",
  29582=>"010111001",
  29583=>"100001100",
  29584=>"011000001",
  29585=>"001101000",
  29586=>"101000110",
  29587=>"100110100",
  29588=>"011111101",
  29589=>"100010101",
  29590=>"110001101",
  29591=>"111011100",
  29592=>"010010010",
  29593=>"110000000",
  29594=>"110010010",
  29595=>"111011110",
  29596=>"010000100",
  29597=>"110010100",
  29598=>"000001101",
  29599=>"000000101",
  29600=>"000011011",
  29601=>"011100100",
  29602=>"100001111",
  29603=>"000100000",
  29604=>"100001011",
  29605=>"010111000",
  29606=>"101110011",
  29607=>"010000011",
  29608=>"101110100",
  29609=>"000000100",
  29610=>"101000101",
  29611=>"011101011",
  29612=>"101100001",
  29613=>"010000010",
  29614=>"010011111",
  29615=>"100001000",
  29616=>"101100110",
  29617=>"010000000",
  29618=>"010000010",
  29619=>"001111100",
  29620=>"100111000",
  29621=>"010000101",
  29622=>"111011110",
  29623=>"100000010",
  29624=>"010001111",
  29625=>"000101111",
  29626=>"010101001",
  29627=>"111110111",
  29628=>"111010100",
  29629=>"000111010",
  29630=>"111100011",
  29631=>"111100010",
  29632=>"001111110",
  29633=>"101110001",
  29634=>"000011101",
  29635=>"001010100",
  29636=>"101010011",
  29637=>"110001110",
  29638=>"111111000",
  29639=>"000111110",
  29640=>"011000010",
  29641=>"000011100",
  29642=>"100010100",
  29643=>"011111010",
  29644=>"111011000",
  29645=>"001010101",
  29646=>"010000001",
  29647=>"011000011",
  29648=>"100010101",
  29649=>"100100010",
  29650=>"001000111",
  29651=>"001010010",
  29652=>"010000001",
  29653=>"001100111",
  29654=>"100100110",
  29655=>"101110111",
  29656=>"111101110",
  29657=>"100011100",
  29658=>"111010010",
  29659=>"101011100",
  29660=>"101111111",
  29661=>"000000100",
  29662=>"011000000",
  29663=>"001001110",
  29664=>"100101111",
  29665=>"000011011",
  29666=>"110110000",
  29667=>"100001110",
  29668=>"011110011",
  29669=>"101010100",
  29670=>"100011111",
  29671=>"100111111",
  29672=>"110100010",
  29673=>"110000111",
  29674=>"001000010",
  29675=>"000100001",
  29676=>"110100010",
  29677=>"010001001",
  29678=>"011100110",
  29679=>"111010001",
  29680=>"011110100",
  29681=>"100111011",
  29682=>"101101110",
  29683=>"110111001",
  29684=>"000011001",
  29685=>"110000001",
  29686=>"011110110",
  29687=>"110011110",
  29688=>"000000010",
  29689=>"011111000",
  29690=>"100101101",
  29691=>"101100010",
  29692=>"111111010",
  29693=>"101111000",
  29694=>"001110011",
  29695=>"001001001",
  29696=>"111101110",
  29697=>"111001011",
  29698=>"000101011",
  29699=>"010111011",
  29700=>"101001101",
  29701=>"100010001",
  29702=>"011111110",
  29703=>"011100010",
  29704=>"100011101",
  29705=>"011110010",
  29706=>"101000110",
  29707=>"111010100",
  29708=>"001100100",
  29709=>"111011110",
  29710=>"011001011",
  29711=>"101110000",
  29712=>"010111000",
  29713=>"000101000",
  29714=>"011100101",
  29715=>"110000100",
  29716=>"100000001",
  29717=>"101011100",
  29718=>"001101000",
  29719=>"010000001",
  29720=>"111000000",
  29721=>"101001001",
  29722=>"110111100",
  29723=>"011000001",
  29724=>"110101010",
  29725=>"111111100",
  29726=>"001100100",
  29727=>"101111010",
  29728=>"111011010",
  29729=>"100111111",
  29730=>"100101001",
  29731=>"000001111",
  29732=>"000010010",
  29733=>"101101110",
  29734=>"100001001",
  29735=>"000101101",
  29736=>"001011110",
  29737=>"101000000",
  29738=>"001101001",
  29739=>"100100000",
  29740=>"100101101",
  29741=>"111011110",
  29742=>"001001011",
  29743=>"110011011",
  29744=>"110000100",
  29745=>"100000000",
  29746=>"011111010",
  29747=>"110101111",
  29748=>"010011011",
  29749=>"000100001",
  29750=>"100010011",
  29751=>"000110011",
  29752=>"000100010",
  29753=>"000101111",
  29754=>"100001101",
  29755=>"001101010",
  29756=>"111000100",
  29757=>"111001100",
  29758=>"100011101",
  29759=>"100100111",
  29760=>"101010010",
  29761=>"011001100",
  29762=>"101010000",
  29763=>"011011111",
  29764=>"111110000",
  29765=>"000001110",
  29766=>"111001100",
  29767=>"111001001",
  29768=>"011000110",
  29769=>"111011111",
  29770=>"011011000",
  29771=>"001110111",
  29772=>"010000001",
  29773=>"101100111",
  29774=>"100100001",
  29775=>"010100010",
  29776=>"111010111",
  29777=>"001001000",
  29778=>"101010100",
  29779=>"111001011",
  29780=>"010100000",
  29781=>"111110010",
  29782=>"100101100",
  29783=>"100001101",
  29784=>"110000001",
  29785=>"010101100",
  29786=>"100011000",
  29787=>"100100010",
  29788=>"011000111",
  29789=>"000100110",
  29790=>"000011110",
  29791=>"101001001",
  29792=>"101110101",
  29793=>"001010001",
  29794=>"010010000",
  29795=>"000101101",
  29796=>"110100011",
  29797=>"110100011",
  29798=>"010011110",
  29799=>"000100100",
  29800=>"010001111",
  29801=>"111000101",
  29802=>"111101110",
  29803=>"110001001",
  29804=>"011000001",
  29805=>"111101101",
  29806=>"111000000",
  29807=>"001110011",
  29808=>"001111000",
  29809=>"001110000",
  29810=>"100001000",
  29811=>"110000010",
  29812=>"001011000",
  29813=>"110001010",
  29814=>"110010011",
  29815=>"100001010",
  29816=>"110010111",
  29817=>"110110001",
  29818=>"001101001",
  29819=>"111100010",
  29820=>"001111111",
  29821=>"011111010",
  29822=>"001010111",
  29823=>"011011011",
  29824=>"101001101",
  29825=>"111011110",
  29826=>"100011001",
  29827=>"000111000",
  29828=>"000110000",
  29829=>"010101100",
  29830=>"101100000",
  29831=>"101101000",
  29832=>"011000001",
  29833=>"000100010",
  29834=>"110101011",
  29835=>"010001010",
  29836=>"101111101",
  29837=>"101010011",
  29838=>"111100101",
  29839=>"111101110",
  29840=>"111000101",
  29841=>"011010111",
  29842=>"001100101",
  29843=>"111001111",
  29844=>"100101111",
  29845=>"010111011",
  29846=>"101000001",
  29847=>"000101100",
  29848=>"010011011",
  29849=>"001110110",
  29850=>"101111111",
  29851=>"001011000",
  29852=>"000010100",
  29853=>"110011100",
  29854=>"011100101",
  29855=>"000101010",
  29856=>"111000100",
  29857=>"010110010",
  29858=>"101010010",
  29859=>"001110110",
  29860=>"000010101",
  29861=>"101110000",
  29862=>"100110111",
  29863=>"011000100",
  29864=>"001001100",
  29865=>"011011010",
  29866=>"000010000",
  29867=>"101101001",
  29868=>"110100001",
  29869=>"010100100",
  29870=>"010100010",
  29871=>"110110010",
  29872=>"011011111",
  29873=>"010011101",
  29874=>"101001101",
  29875=>"101010010",
  29876=>"111010011",
  29877=>"100000001",
  29878=>"111110011",
  29879=>"111010111",
  29880=>"001011011",
  29881=>"100011001",
  29882=>"000100101",
  29883=>"101101001",
  29884=>"111100111",
  29885=>"110010111",
  29886=>"001000110",
  29887=>"011010001",
  29888=>"000001011",
  29889=>"101111110",
  29890=>"111110011",
  29891=>"010111011",
  29892=>"010110000",
  29893=>"000000000",
  29894=>"101001110",
  29895=>"010100111",
  29896=>"000010000",
  29897=>"001011011",
  29898=>"001001001",
  29899=>"111100110",
  29900=>"110001000",
  29901=>"111111100",
  29902=>"000010010",
  29903=>"010110100",
  29904=>"001000010",
  29905=>"100011001",
  29906=>"100000111",
  29907=>"111001101",
  29908=>"001000101",
  29909=>"110001101",
  29910=>"110000110",
  29911=>"101010010",
  29912=>"011001011",
  29913=>"000111000",
  29914=>"001110101",
  29915=>"101011010",
  29916=>"111100110",
  29917=>"100011010",
  29918=>"101000011",
  29919=>"010010011",
  29920=>"110001110",
  29921=>"010111101",
  29922=>"011010100",
  29923=>"011100011",
  29924=>"100110111",
  29925=>"101010110",
  29926=>"001000111",
  29927=>"000111000",
  29928=>"000111100",
  29929=>"001001110",
  29930=>"010110010",
  29931=>"101010011",
  29932=>"110011101",
  29933=>"101100000",
  29934=>"001101010",
  29935=>"000001101",
  29936=>"010110011",
  29937=>"111100111",
  29938=>"000111101",
  29939=>"101101110",
  29940=>"001011001",
  29941=>"011101111",
  29942=>"010100101",
  29943=>"001011010",
  29944=>"011000111",
  29945=>"100111101",
  29946=>"111100011",
  29947=>"100010101",
  29948=>"011111101",
  29949=>"111111000",
  29950=>"010001100",
  29951=>"001001111",
  29952=>"011011100",
  29953=>"101110111",
  29954=>"111011110",
  29955=>"011111000",
  29956=>"100011000",
  29957=>"100110011",
  29958=>"010011011",
  29959=>"111011100",
  29960=>"000001111",
  29961=>"100000110",
  29962=>"010110011",
  29963=>"100010101",
  29964=>"001101001",
  29965=>"000000101",
  29966=>"001000011",
  29967=>"000000110",
  29968=>"001101010",
  29969=>"000000101",
  29970=>"010101010",
  29971=>"001101000",
  29972=>"011010001",
  29973=>"100101001",
  29974=>"100101100",
  29975=>"111010011",
  29976=>"010010000",
  29977=>"100100001",
  29978=>"011010111",
  29979=>"111000100",
  29980=>"100000101",
  29981=>"010000010",
  29982=>"000011100",
  29983=>"000001000",
  29984=>"000010111",
  29985=>"001001011",
  29986=>"010011110",
  29987=>"101011101",
  29988=>"111111010",
  29989=>"001000011",
  29990=>"101001001",
  29991=>"101100000",
  29992=>"101111100",
  29993=>"001100001",
  29994=>"000000111",
  29995=>"000010010",
  29996=>"010101010",
  29997=>"001101101",
  29998=>"000111101",
  29999=>"110111100",
  30000=>"100001101",
  30001=>"010101110",
  30002=>"000101011",
  30003=>"010001010",
  30004=>"100000100",
  30005=>"010100000",
  30006=>"010110101",
  30007=>"111001111",
  30008=>"000100100",
  30009=>"000110010",
  30010=>"100011100",
  30011=>"110110100",
  30012=>"110001100",
  30013=>"010001011",
  30014=>"010100111",
  30015=>"111001010",
  30016=>"010011111",
  30017=>"001110001",
  30018=>"100000001",
  30019=>"010000101",
  30020=>"101101011",
  30021=>"111010100",
  30022=>"100010100",
  30023=>"101111001",
  30024=>"011111100",
  30025=>"010111101",
  30026=>"100100010",
  30027=>"101101000",
  30028=>"111110000",
  30029=>"000111111",
  30030=>"001101010",
  30031=>"011100101",
  30032=>"101000001",
  30033=>"001101001",
  30034=>"011010010",
  30035=>"000101101",
  30036=>"111110011",
  30037=>"101000010",
  30038=>"010110000",
  30039=>"001101110",
  30040=>"000000111",
  30041=>"010101000",
  30042=>"001000110",
  30043=>"010100001",
  30044=>"001110111",
  30045=>"011100100",
  30046=>"100010101",
  30047=>"010010100",
  30048=>"001100110",
  30049=>"101001110",
  30050=>"100000110",
  30051=>"001101010",
  30052=>"101000111",
  30053=>"100100011",
  30054=>"100011111",
  30055=>"100111110",
  30056=>"011100001",
  30057=>"100101111",
  30058=>"000000111",
  30059=>"000110111",
  30060=>"000111110",
  30061=>"101011001",
  30062=>"001101000",
  30063=>"110100110",
  30064=>"010100110",
  30065=>"010101000",
  30066=>"100000010",
  30067=>"110111000",
  30068=>"000000010",
  30069=>"011010111",
  30070=>"010101100",
  30071=>"111011000",
  30072=>"010111111",
  30073=>"100011001",
  30074=>"000101001",
  30075=>"111110000",
  30076=>"001100101",
  30077=>"111010000",
  30078=>"000110101",
  30079=>"001000100",
  30080=>"000110101",
  30081=>"100110010",
  30082=>"001001011",
  30083=>"010000000",
  30084=>"100111110",
  30085=>"000010000",
  30086=>"101100101",
  30087=>"010000011",
  30088=>"011100111",
  30089=>"101111010",
  30090=>"000110100",
  30091=>"010000111",
  30092=>"011100100",
  30093=>"101100001",
  30094=>"000101100",
  30095=>"000000110",
  30096=>"010001001",
  30097=>"000000010",
  30098=>"111011011",
  30099=>"001111010",
  30100=>"110101101",
  30101=>"101001101",
  30102=>"100111100",
  30103=>"000000010",
  30104=>"100111001",
  30105=>"001100111",
  30106=>"001101101",
  30107=>"111110111",
  30108=>"010111101",
  30109=>"101111011",
  30110=>"111101101",
  30111=>"100000001",
  30112=>"000100000",
  30113=>"101001101",
  30114=>"111000010",
  30115=>"001001001",
  30116=>"000001101",
  30117=>"010101111",
  30118=>"110000001",
  30119=>"010111000",
  30120=>"110110110",
  30121=>"111010001",
  30122=>"101101100",
  30123=>"001100010",
  30124=>"100011111",
  30125=>"001101111",
  30126=>"011010100",
  30127=>"001110101",
  30128=>"111000110",
  30129=>"100001111",
  30130=>"010000010",
  30131=>"000010110",
  30132=>"110001001",
  30133=>"001100001",
  30134=>"110011011",
  30135=>"111110110",
  30136=>"001001101",
  30137=>"000000101",
  30138=>"001100000",
  30139=>"100000011",
  30140=>"110101000",
  30141=>"011000100",
  30142=>"111011000",
  30143=>"100011100",
  30144=>"111111111",
  30145=>"110001101",
  30146=>"111101111",
  30147=>"110101000",
  30148=>"110101100",
  30149=>"010000100",
  30150=>"100110101",
  30151=>"111010000",
  30152=>"011000011",
  30153=>"001001011",
  30154=>"010110101",
  30155=>"111000001",
  30156=>"100000011",
  30157=>"101001100",
  30158=>"111010000",
  30159=>"111010001",
  30160=>"101100010",
  30161=>"011100011",
  30162=>"010101100",
  30163=>"011011100",
  30164=>"010000111",
  30165=>"001110110",
  30166=>"011111010",
  30167=>"001001011",
  30168=>"110111110",
  30169=>"010001010",
  30170=>"110110010",
  30171=>"000101011",
  30172=>"010110010",
  30173=>"101010010",
  30174=>"110110100",
  30175=>"111011010",
  30176=>"010010011",
  30177=>"000111110",
  30178=>"011011011",
  30179=>"110001010",
  30180=>"010101010",
  30181=>"010110101",
  30182=>"010101010",
  30183=>"011111011",
  30184=>"111010110",
  30185=>"000010011",
  30186=>"010010010",
  30187=>"110101000",
  30188=>"111101100",
  30189=>"101001110",
  30190=>"011111101",
  30191=>"011010110",
  30192=>"111011000",
  30193=>"101101010",
  30194=>"100101001",
  30195=>"100001110",
  30196=>"001101010",
  30197=>"111110100",
  30198=>"111000101",
  30199=>"101011111",
  30200=>"010010001",
  30201=>"001010001",
  30202=>"100010110",
  30203=>"000010001",
  30204=>"001100110",
  30205=>"010000010",
  30206=>"011110110",
  30207=>"000100100",
  30208=>"101011110",
  30209=>"011011001",
  30210=>"101101101",
  30211=>"000010111",
  30212=>"100100111",
  30213=>"110100001",
  30214=>"110100101",
  30215=>"011000010",
  30216=>"011001000",
  30217=>"010111010",
  30218=>"101010010",
  30219=>"000110100",
  30220=>"101111010",
  30221=>"101010000",
  30222=>"011000110",
  30223=>"100010010",
  30224=>"111010111",
  30225=>"110101110",
  30226=>"101110110",
  30227=>"011010011",
  30228=>"011001011",
  30229=>"100100010",
  30230=>"110101000",
  30231=>"110101001",
  30232=>"010101001",
  30233=>"001011001",
  30234=>"010001000",
  30235=>"011111011",
  30236=>"001000110",
  30237=>"001000111",
  30238=>"111010111",
  30239=>"000000000",
  30240=>"101111010",
  30241=>"101110000",
  30242=>"100110000",
  30243=>"000101000",
  30244=>"110001100",
  30245=>"011100101",
  30246=>"111010000",
  30247=>"100001000",
  30248=>"100001000",
  30249=>"010111111",
  30250=>"101001111",
  30251=>"010101110",
  30252=>"110100011",
  30253=>"010101111",
  30254=>"010001000",
  30255=>"101001001",
  30256=>"001010101",
  30257=>"110011000",
  30258=>"101000101",
  30259=>"111000001",
  30260=>"011001010",
  30261=>"010011110",
  30262=>"010110000",
  30263=>"000110111",
  30264=>"110010111",
  30265=>"011010010",
  30266=>"000101000",
  30267=>"101010000",
  30268=>"110111011",
  30269=>"111011010",
  30270=>"110000110",
  30271=>"101011001",
  30272=>"011011111",
  30273=>"001001000",
  30274=>"000011011",
  30275=>"101101110",
  30276=>"000010000",
  30277=>"100001000",
  30278=>"000100011",
  30279=>"000101110",
  30280=>"010011111",
  30281=>"100100010",
  30282=>"110010001",
  30283=>"111011111",
  30284=>"111110111",
  30285=>"001100011",
  30286=>"101101001",
  30287=>"100111110",
  30288=>"100110010",
  30289=>"101110100",
  30290=>"111001111",
  30291=>"001100010",
  30292=>"111100101",
  30293=>"000001010",
  30294=>"001110010",
  30295=>"010010001",
  30296=>"100001110",
  30297=>"110111111",
  30298=>"101011010",
  30299=>"101100110",
  30300=>"110000010",
  30301=>"000000000",
  30302=>"001111111",
  30303=>"110000110",
  30304=>"110101101",
  30305=>"010110101",
  30306=>"101000001",
  30307=>"000110100",
  30308=>"011000010",
  30309=>"000010110",
  30310=>"011101010",
  30311=>"001111111",
  30312=>"110101001",
  30313=>"000100000",
  30314=>"001100001",
  30315=>"010000101",
  30316=>"000010111",
  30317=>"101110101",
  30318=>"110110011",
  30319=>"110011001",
  30320=>"010100010",
  30321=>"000000111",
  30322=>"111000100",
  30323=>"000111110",
  30324=>"000111001",
  30325=>"110001110",
  30326=>"000001000",
  30327=>"101001001",
  30328=>"111011101",
  30329=>"001000101",
  30330=>"110100001",
  30331=>"011100111",
  30332=>"100110100",
  30333=>"100111100",
  30334=>"011100101",
  30335=>"111111110",
  30336=>"001001111",
  30337=>"010100000",
  30338=>"111001100",
  30339=>"001000110",
  30340=>"100110110",
  30341=>"100010100",
  30342=>"000101100",
  30343=>"111000010",
  30344=>"011111010",
  30345=>"001010010",
  30346=>"110010101",
  30347=>"011010111",
  30348=>"111100111",
  30349=>"011010110",
  30350=>"011110100",
  30351=>"111100100",
  30352=>"101101111",
  30353=>"010110000",
  30354=>"110110111",
  30355=>"000000000",
  30356=>"000101010",
  30357=>"001001101",
  30358=>"111001010",
  30359=>"101000100",
  30360=>"100001011",
  30361=>"110111010",
  30362=>"001100010",
  30363=>"001101100",
  30364=>"000000000",
  30365=>"000101110",
  30366=>"111000111",
  30367=>"111000101",
  30368=>"110000100",
  30369=>"110111001",
  30370=>"101000001",
  30371=>"101111100",
  30372=>"000010100",
  30373=>"010010101",
  30374=>"011011011",
  30375=>"010010001",
  30376=>"110100010",
  30377=>"100010000",
  30378=>"101100010",
  30379=>"000010110",
  30380=>"000000111",
  30381=>"011010111",
  30382=>"010101011",
  30383=>"000000010",
  30384=>"000111101",
  30385=>"011101001",
  30386=>"100001110",
  30387=>"001000000",
  30388=>"001001111",
  30389=>"001110000",
  30390=>"010000001",
  30391=>"110000011",
  30392=>"100001000",
  30393=>"011111101",
  30394=>"110110011",
  30395=>"001110011",
  30396=>"101010100",
  30397=>"011011110",
  30398=>"100100111",
  30399=>"101000101",
  30400=>"001111000",
  30401=>"010011101",
  30402=>"011100100",
  30403=>"100111000",
  30404=>"111011000",
  30405=>"001000101",
  30406=>"111010000",
  30407=>"011100010",
  30408=>"101011111",
  30409=>"111001000",
  30410=>"011100111",
  30411=>"001000001",
  30412=>"000010100",
  30413=>"101011111",
  30414=>"001011101",
  30415=>"001111011",
  30416=>"110001111",
  30417=>"100101011",
  30418=>"100011010",
  30419=>"011101001",
  30420=>"100001110",
  30421=>"010000010",
  30422=>"110011010",
  30423=>"111110001",
  30424=>"100111100",
  30425=>"100001001",
  30426=>"000100111",
  30427=>"011100100",
  30428=>"100001001",
  30429=>"001110010",
  30430=>"001101010",
  30431=>"111001110",
  30432=>"011111111",
  30433=>"010010011",
  30434=>"001001110",
  30435=>"001100000",
  30436=>"000111111",
  30437=>"000000010",
  30438=>"111101000",
  30439=>"001100101",
  30440=>"011001100",
  30441=>"010001001",
  30442=>"010000011",
  30443=>"111101000",
  30444=>"010101110",
  30445=>"010000010",
  30446=>"100101111",
  30447=>"110101010",
  30448=>"011001111",
  30449=>"111010000",
  30450=>"001111000",
  30451=>"100001011",
  30452=>"010000110",
  30453=>"100101100",
  30454=>"101101100",
  30455=>"110111000",
  30456=>"101101001",
  30457=>"010010100",
  30458=>"111000000",
  30459=>"101000110",
  30460=>"000000011",
  30461=>"000101000",
  30462=>"010101101",
  30463=>"001011010",
  30464=>"101110010",
  30465=>"010001110",
  30466=>"011011100",
  30467=>"110101000",
  30468=>"111100010",
  30469=>"100010111",
  30470=>"101001010",
  30471=>"100000110",
  30472=>"010000101",
  30473=>"001110110",
  30474=>"100101101",
  30475=>"000000011",
  30476=>"110110010",
  30477=>"110001111",
  30478=>"110010101",
  30479=>"010000001",
  30480=>"111010111",
  30481=>"000000011",
  30482=>"111011111",
  30483=>"100101110",
  30484=>"100101010",
  30485=>"001101110",
  30486=>"010001001",
  30487=>"010111101",
  30488=>"100001100",
  30489=>"001110011",
  30490=>"101111101",
  30491=>"001110101",
  30492=>"100110101",
  30493=>"101010001",
  30494=>"000100110",
  30495=>"010100101",
  30496=>"011000010",
  30497=>"011011011",
  30498=>"001000101",
  30499=>"100001010",
  30500=>"010010100",
  30501=>"000001010",
  30502=>"100101100",
  30503=>"111110000",
  30504=>"101111100",
  30505=>"001110010",
  30506=>"101100010",
  30507=>"111011101",
  30508=>"111100111",
  30509=>"110110000",
  30510=>"101101111",
  30511=>"111011111",
  30512=>"111111110",
  30513=>"001111111",
  30514=>"100011001",
  30515=>"100101011",
  30516=>"110000110",
  30517=>"111100000",
  30518=>"100000111",
  30519=>"111010000",
  30520=>"000001001",
  30521=>"100000000",
  30522=>"100111110",
  30523=>"111000011",
  30524=>"110111111",
  30525=>"000111110",
  30526=>"011111011",
  30527=>"100000110",
  30528=>"001000111",
  30529=>"001010000",
  30530=>"111100110",
  30531=>"001010000",
  30532=>"010101110",
  30533=>"110100101",
  30534=>"100101111",
  30535=>"111001101",
  30536=>"010100001",
  30537=>"111101001",
  30538=>"111111111",
  30539=>"001100011",
  30540=>"001100111",
  30541=>"100000011",
  30542=>"101101000",
  30543=>"000011101",
  30544=>"101000100",
  30545=>"000000110",
  30546=>"110111010",
  30547=>"111001111",
  30548=>"010010010",
  30549=>"100000101",
  30550=>"011100011",
  30551=>"011010001",
  30552=>"100011000",
  30553=>"010111110",
  30554=>"111110011",
  30555=>"000111111",
  30556=>"000000100",
  30557=>"110110010",
  30558=>"111100101",
  30559=>"100011110",
  30560=>"111110000",
  30561=>"111111111",
  30562=>"101100011",
  30563=>"101000110",
  30564=>"001010111",
  30565=>"001010001",
  30566=>"000101011",
  30567=>"101101001",
  30568=>"100000000",
  30569=>"101010001",
  30570=>"100000001",
  30571=>"010001111",
  30572=>"010101011",
  30573=>"110011100",
  30574=>"110110110",
  30575=>"101011000",
  30576=>"111101000",
  30577=>"001000011",
  30578=>"011000011",
  30579=>"100011110",
  30580=>"001101011",
  30581=>"010010110",
  30582=>"000110000",
  30583=>"101100000",
  30584=>"001000010",
  30585=>"110000000",
  30586=>"000011010",
  30587=>"001000001",
  30588=>"100100000",
  30589=>"011010100",
  30590=>"000101111",
  30591=>"100011111",
  30592=>"001110010",
  30593=>"110001010",
  30594=>"001100110",
  30595=>"000100100",
  30596=>"100110100",
  30597=>"110011001",
  30598=>"000110110",
  30599=>"110011100",
  30600=>"101111001",
  30601=>"100001110",
  30602=>"001100110",
  30603=>"001111010",
  30604=>"011111001",
  30605=>"011100000",
  30606=>"101010000",
  30607=>"101111011",
  30608=>"001000110",
  30609=>"111001011",
  30610=>"000010001",
  30611=>"011100100",
  30612=>"110010011",
  30613=>"101000011",
  30614=>"010000111",
  30615=>"101001001",
  30616=>"011101110",
  30617=>"111111111",
  30618=>"001100100",
  30619=>"111110011",
  30620=>"000000110",
  30621=>"010001001",
  30622=>"010111111",
  30623=>"000001111",
  30624=>"101011111",
  30625=>"001010000",
  30626=>"000011111",
  30627=>"000100110",
  30628=>"000000011",
  30629=>"100111110",
  30630=>"000110111",
  30631=>"000110101",
  30632=>"100101110",
  30633=>"110001011",
  30634=>"110110100",
  30635=>"010110001",
  30636=>"100110010",
  30637=>"001000000",
  30638=>"100110101",
  30639=>"001001100",
  30640=>"101101110",
  30641=>"001010011",
  30642=>"111000101",
  30643=>"100011110",
  30644=>"111110111",
  30645=>"101011011",
  30646=>"110000111",
  30647=>"111110101",
  30648=>"011011011",
  30649=>"111111111",
  30650=>"110101110",
  30651=>"100110001",
  30652=>"100100111",
  30653=>"101000000",
  30654=>"010010101",
  30655=>"001100110",
  30656=>"001010100",
  30657=>"011110101",
  30658=>"101111110",
  30659=>"110000000",
  30660=>"000101011",
  30661=>"110111011",
  30662=>"001011011",
  30663=>"100110101",
  30664=>"110100110",
  30665=>"001001101",
  30666=>"111001100",
  30667=>"100011010",
  30668=>"000110000",
  30669=>"101111010",
  30670=>"010010110",
  30671=>"111100110",
  30672=>"010010001",
  30673=>"010010000",
  30674=>"010010100",
  30675=>"101100010",
  30676=>"001001111",
  30677=>"111111000",
  30678=>"010110011",
  30679=>"101001010",
  30680=>"001100100",
  30681=>"000010000",
  30682=>"110110001",
  30683=>"111001101",
  30684=>"011000100",
  30685=>"011110100",
  30686=>"000001110",
  30687=>"000000100",
  30688=>"010101010",
  30689=>"000111111",
  30690=>"100111010",
  30691=>"011000101",
  30692=>"110001010",
  30693=>"011000100",
  30694=>"000111010",
  30695=>"000100001",
  30696=>"000110111",
  30697=>"001110111",
  30698=>"100101000",
  30699=>"100110011",
  30700=>"011111001",
  30701=>"100010101",
  30702=>"111001111",
  30703=>"101000010",
  30704=>"011101001",
  30705=>"000001001",
  30706=>"011111100",
  30707=>"100001101",
  30708=>"100000011",
  30709=>"010100111",
  30710=>"011111110",
  30711=>"010100111",
  30712=>"001000000",
  30713=>"101010101",
  30714=>"100100101",
  30715=>"011111010",
  30716=>"000110010",
  30717=>"101011110",
  30718=>"101001100",
  30719=>"110110011",
  30720=>"010011000",
  30721=>"111010101",
  30722=>"000111101",
  30723=>"100111001",
  30724=>"101001000",
  30725=>"101010000",
  30726=>"001001011",
  30727=>"000011000",
  30728=>"111000111",
  30729=>"000000000",
  30730=>"010100000",
  30731=>"100000100",
  30732=>"011101010",
  30733=>"011111111",
  30734=>"111001100",
  30735=>"000000000",
  30736=>"000101001",
  30737=>"010101010",
  30738=>"011010101",
  30739=>"111010111",
  30740=>"011110101",
  30741=>"110100110",
  30742=>"100001001",
  30743=>"010011101",
  30744=>"010000100",
  30745=>"111110010",
  30746=>"111000000",
  30747=>"000011011",
  30748=>"100011110",
  30749=>"010001010",
  30750=>"000110111",
  30751=>"100110110",
  30752=>"111110001",
  30753=>"000010000",
  30754=>"111101011",
  30755=>"110000100",
  30756=>"000101000",
  30757=>"110011101",
  30758=>"111000100",
  30759=>"000000001",
  30760=>"011000000",
  30761=>"010101010",
  30762=>"101100110",
  30763=>"011000100",
  30764=>"010010110",
  30765=>"101110100",
  30766=>"101001110",
  30767=>"100110010",
  30768=>"000000111",
  30769=>"101011000",
  30770=>"101110100",
  30771=>"001110110",
  30772=>"111010000",
  30773=>"010100011",
  30774=>"010110011",
  30775=>"011000010",
  30776=>"010110000",
  30777=>"101110101",
  30778=>"000011100",
  30779=>"000111011",
  30780=>"000011000",
  30781=>"001000011",
  30782=>"010111101",
  30783=>"000000000",
  30784=>"001010011",
  30785=>"000001011",
  30786=>"100011000",
  30787=>"110011000",
  30788=>"010110010",
  30789=>"100001000",
  30790=>"111011111",
  30791=>"000001000",
  30792=>"100001011",
  30793=>"101000000",
  30794=>"010100011",
  30795=>"101010110",
  30796=>"101011001",
  30797=>"110000000",
  30798=>"101011000",
  30799=>"010100000",
  30800=>"001000001",
  30801=>"011001001",
  30802=>"010111000",
  30803=>"001000001",
  30804=>"111001011",
  30805=>"001110001",
  30806=>"101010101",
  30807=>"000111001",
  30808=>"111011110",
  30809=>"011111110",
  30810=>"010111110",
  30811=>"101010000",
  30812=>"011100010",
  30813=>"010011101",
  30814=>"010100110",
  30815=>"000010000",
  30816=>"010010011",
  30817=>"100010110",
  30818=>"000010011",
  30819=>"110101101",
  30820=>"100111001",
  30821=>"110110100",
  30822=>"111101011",
  30823=>"011010011",
  30824=>"001110001",
  30825=>"010110010",
  30826=>"110011001",
  30827=>"011011111",
  30828=>"010001111",
  30829=>"010000010",
  30830=>"010001100",
  30831=>"010000010",
  30832=>"010101010",
  30833=>"000011111",
  30834=>"000100100",
  30835=>"111010111",
  30836=>"000111100",
  30837=>"110101101",
  30838=>"110111001",
  30839=>"100011000",
  30840=>"011001010",
  30841=>"110110101",
  30842=>"111111110",
  30843=>"010111001",
  30844=>"001001110",
  30845=>"111111001",
  30846=>"110000010",
  30847=>"000111100",
  30848=>"011001000",
  30849=>"101101011",
  30850=>"000000101",
  30851=>"000000011",
  30852=>"001110001",
  30853=>"111110101",
  30854=>"110111000",
  30855=>"110000011",
  30856=>"000010001",
  30857=>"100001110",
  30858=>"101111111",
  30859=>"111001010",
  30860=>"100100111",
  30861=>"111001110",
  30862=>"010000111",
  30863=>"011110000",
  30864=>"110101010",
  30865=>"100011100",
  30866=>"110101010",
  30867=>"101110100",
  30868=>"101110110",
  30869=>"100100101",
  30870=>"000110001",
  30871=>"001110011",
  30872=>"011001111",
  30873=>"100010101",
  30874=>"100000110",
  30875=>"011010011",
  30876=>"000001110",
  30877=>"100000100",
  30878=>"000110011",
  30879=>"101011101",
  30880=>"110010100",
  30881=>"000100110",
  30882=>"000110100",
  30883=>"011001110",
  30884=>"101101011",
  30885=>"111001000",
  30886=>"001000111",
  30887=>"000100000",
  30888=>"101100000",
  30889=>"001111000",
  30890=>"001010000",
  30891=>"101101010",
  30892=>"001000101",
  30893=>"100111110",
  30894=>"000011101",
  30895=>"111011100",
  30896=>"100111110",
  30897=>"010111000",
  30898=>"100100100",
  30899=>"000101011",
  30900=>"111000011",
  30901=>"011011111",
  30902=>"100000100",
  30903=>"110011100",
  30904=>"111010000",
  30905=>"111111100",
  30906=>"111000001",
  30907=>"101011001",
  30908=>"101001110",
  30909=>"111110011",
  30910=>"100111110",
  30911=>"010111010",
  30912=>"010101011",
  30913=>"100010101",
  30914=>"011111110",
  30915=>"101101101",
  30916=>"111101111",
  30917=>"011111001",
  30918=>"110101110",
  30919=>"010101011",
  30920=>"011110111",
  30921=>"001111010",
  30922=>"100011111",
  30923=>"001010100",
  30924=>"010000110",
  30925=>"100101100",
  30926=>"010010001",
  30927=>"111100100",
  30928=>"010000100",
  30929=>"000100101",
  30930=>"111111001",
  30931=>"101011100",
  30932=>"111101010",
  30933=>"001100110",
  30934=>"100100011",
  30935=>"001101011",
  30936=>"111001110",
  30937=>"110111101",
  30938=>"100011001",
  30939=>"001101001",
  30940=>"111111100",
  30941=>"000011110",
  30942=>"001001000",
  30943=>"000110111",
  30944=>"111101011",
  30945=>"001011010",
  30946=>"100001101",
  30947=>"110111010",
  30948=>"111001110",
  30949=>"110110110",
  30950=>"010110001",
  30951=>"111001101",
  30952=>"100110101",
  30953=>"100000001",
  30954=>"101101000",
  30955=>"101001101",
  30956=>"010110000",
  30957=>"111001010",
  30958=>"000000010",
  30959=>"100010110",
  30960=>"000100001",
  30961=>"011001001",
  30962=>"011110100",
  30963=>"101101010",
  30964=>"111011111",
  30965=>"110101010",
  30966=>"110111000",
  30967=>"000011000",
  30968=>"100100110",
  30969=>"101100111",
  30970=>"000110101",
  30971=>"101000000",
  30972=>"111100110",
  30973=>"011100010",
  30974=>"110001010",
  30975=>"010010001",
  30976=>"001000001",
  30977=>"101101111",
  30978=>"110000101",
  30979=>"001111000",
  30980=>"110101010",
  30981=>"111111000",
  30982=>"010100000",
  30983=>"100000110",
  30984=>"010110100",
  30985=>"000010110",
  30986=>"001000111",
  30987=>"110010001",
  30988=>"111100111",
  30989=>"100011111",
  30990=>"010101111",
  30991=>"100010010",
  30992=>"001000001",
  30993=>"011111101",
  30994=>"110011101",
  30995=>"110001110",
  30996=>"001100101",
  30997=>"000000101",
  30998=>"111011010",
  30999=>"111110101",
  31000=>"101110011",
  31001=>"011110110",
  31002=>"111101010",
  31003=>"111011000",
  31004=>"000110011",
  31005=>"111001011",
  31006=>"001100001",
  31007=>"001001110",
  31008=>"101010111",
  31009=>"111111100",
  31010=>"100100010",
  31011=>"101100101",
  31012=>"011101010",
  31013=>"010010111",
  31014=>"111001010",
  31015=>"010011111",
  31016=>"111100101",
  31017=>"001100000",
  31018=>"100111111",
  31019=>"000000010",
  31020=>"111111001",
  31021=>"110101000",
  31022=>"101100000",
  31023=>"000011100",
  31024=>"010010001",
  31025=>"111011101",
  31026=>"001101111",
  31027=>"010010101",
  31028=>"001101000",
  31029=>"000101100",
  31030=>"111110100",
  31031=>"000101011",
  31032=>"000000101",
  31033=>"101110000",
  31034=>"110101111",
  31035=>"000000011",
  31036=>"110010111",
  31037=>"000110000",
  31038=>"110000000",
  31039=>"110100101",
  31040=>"000010001",
  31041=>"000001000",
  31042=>"110111001",
  31043=>"010100100",
  31044=>"001001010",
  31045=>"010011111",
  31046=>"000010010",
  31047=>"110101000",
  31048=>"001001100",
  31049=>"111110000",
  31050=>"101011111",
  31051=>"001001111",
  31052=>"000101001",
  31053=>"011100000",
  31054=>"111110001",
  31055=>"011000000",
  31056=>"101111010",
  31057=>"101100110",
  31058=>"110000101",
  31059=>"000001110",
  31060=>"100010000",
  31061=>"110110010",
  31062=>"010110101",
  31063=>"000111010",
  31064=>"001101100",
  31065=>"100000000",
  31066=>"110000111",
  31067=>"011100100",
  31068=>"100001101",
  31069=>"100000111",
  31070=>"001111011",
  31071=>"010000100",
  31072=>"000001101",
  31073=>"110010110",
  31074=>"101001001",
  31075=>"010101011",
  31076=>"000000011",
  31077=>"111101100",
  31078=>"010100000",
  31079=>"000011001",
  31080=>"011001101",
  31081=>"011000001",
  31082=>"001010011",
  31083=>"111101011",
  31084=>"100010000",
  31085=>"110101001",
  31086=>"000000011",
  31087=>"100100101",
  31088=>"011011101",
  31089=>"110001111",
  31090=>"101101111",
  31091=>"110110100",
  31092=>"011000011",
  31093=>"101101010",
  31094=>"001101010",
  31095=>"011110111",
  31096=>"000000011",
  31097=>"010010110",
  31098=>"100111011",
  31099=>"100011111",
  31100=>"100100100",
  31101=>"000110111",
  31102=>"101111000",
  31103=>"110110000",
  31104=>"010011101",
  31105=>"100111111",
  31106=>"011011010",
  31107=>"000110001",
  31108=>"000110000",
  31109=>"101101010",
  31110=>"101111010",
  31111=>"011011011",
  31112=>"111110101",
  31113=>"000101110",
  31114=>"001101101",
  31115=>"110010101",
  31116=>"001110000",
  31117=>"000100101",
  31118=>"010110101",
  31119=>"010110111",
  31120=>"010100101",
  31121=>"011000000",
  31122=>"100101111",
  31123=>"111011101",
  31124=>"100101010",
  31125=>"100110100",
  31126=>"110010001",
  31127=>"110110011",
  31128=>"110110000",
  31129=>"001110000",
  31130=>"011001011",
  31131=>"000011000",
  31132=>"111110110",
  31133=>"010101001",
  31134=>"100010010",
  31135=>"101110110",
  31136=>"011011111",
  31137=>"010111010",
  31138=>"101111111",
  31139=>"110011010",
  31140=>"001101000",
  31141=>"100000100",
  31142=>"010111010",
  31143=>"100101000",
  31144=>"000011000",
  31145=>"110000000",
  31146=>"000100010",
  31147=>"000001111",
  31148=>"101101110",
  31149=>"000001010",
  31150=>"011001110",
  31151=>"101010111",
  31152=>"100100011",
  31153=>"010010011",
  31154=>"000011111",
  31155=>"111000001",
  31156=>"010010101",
  31157=>"000111110",
  31158=>"010100111",
  31159=>"010111011",
  31160=>"101000101",
  31161=>"000101000",
  31162=>"001100001",
  31163=>"111011000",
  31164=>"000010001",
  31165=>"010000101",
  31166=>"101110000",
  31167=>"111010011",
  31168=>"100010000",
  31169=>"100000010",
  31170=>"110011111",
  31171=>"001111110",
  31172=>"000011101",
  31173=>"111001100",
  31174=>"111101100",
  31175=>"101100000",
  31176=>"111111001",
  31177=>"110011111",
  31178=>"010010000",
  31179=>"000000110",
  31180=>"000010101",
  31181=>"011010001",
  31182=>"000101111",
  31183=>"001011101",
  31184=>"111100000",
  31185=>"100110001",
  31186=>"101101001",
  31187=>"011111111",
  31188=>"010111010",
  31189=>"111110111",
  31190=>"101000100",
  31191=>"111011010",
  31192=>"100000001",
  31193=>"011101001",
  31194=>"101111001",
  31195=>"100000011",
  31196=>"011010100",
  31197=>"001001011",
  31198=>"111000111",
  31199=>"010010101",
  31200=>"010101001",
  31201=>"100000011",
  31202=>"110011111",
  31203=>"111011001",
  31204=>"000001010",
  31205=>"110000010",
  31206=>"100000011",
  31207=>"100110010",
  31208=>"000011001",
  31209=>"110001101",
  31210=>"110011000",
  31211=>"110010110",
  31212=>"100001101",
  31213=>"000011000",
  31214=>"111010000",
  31215=>"001110111",
  31216=>"111010111",
  31217=>"000100000",
  31218=>"000010001",
  31219=>"011100111",
  31220=>"101110111",
  31221=>"001001011",
  31222=>"111001100",
  31223=>"010011001",
  31224=>"001101010",
  31225=>"111001011",
  31226=>"111011010",
  31227=>"010100011",
  31228=>"101011001",
  31229=>"101110111",
  31230=>"001100111",
  31231=>"000001001",
  31232=>"101101101",
  31233=>"110001011",
  31234=>"011100100",
  31235=>"111001010",
  31236=>"000110100",
  31237=>"100000000",
  31238=>"101110010",
  31239=>"110010001",
  31240=>"101011000",
  31241=>"111111101",
  31242=>"101001001",
  31243=>"011101101",
  31244=>"111011110",
  31245=>"101001000",
  31246=>"111010001",
  31247=>"100010001",
  31248=>"000111001",
  31249=>"000000110",
  31250=>"010111001",
  31251=>"010010001",
  31252=>"000110000",
  31253=>"101100001",
  31254=>"000011011",
  31255=>"010001011",
  31256=>"010000001",
  31257=>"001010011",
  31258=>"010010010",
  31259=>"000000001",
  31260=>"011100001",
  31261=>"110000000",
  31262=>"000110011",
  31263=>"100101100",
  31264=>"011100011",
  31265=>"011101001",
  31266=>"111111111",
  31267=>"111011011",
  31268=>"110010000",
  31269=>"111010110",
  31270=>"010001011",
  31271=>"110110001",
  31272=>"101011000",
  31273=>"110111111",
  31274=>"100101011",
  31275=>"101111101",
  31276=>"001011000",
  31277=>"101000100",
  31278=>"100010101",
  31279=>"011100100",
  31280=>"011010100",
  31281=>"110001000",
  31282=>"001011011",
  31283=>"000000101",
  31284=>"100000100",
  31285=>"011111010",
  31286=>"011001111",
  31287=>"111100110",
  31288=>"100011101",
  31289=>"011101001",
  31290=>"001101111",
  31291=>"111100011",
  31292=>"011100111",
  31293=>"000000100",
  31294=>"110011110",
  31295=>"011101101",
  31296=>"000000001",
  31297=>"100111111",
  31298=>"110101100",
  31299=>"010011111",
  31300=>"010000000",
  31301=>"101001001",
  31302=>"011001100",
  31303=>"101001100",
  31304=>"001000010",
  31305=>"000110101",
  31306=>"101111111",
  31307=>"000111111",
  31308=>"101000000",
  31309=>"011001101",
  31310=>"010101100",
  31311=>"100100000",
  31312=>"111111011",
  31313=>"111011110",
  31314=>"011101111",
  31315=>"010111000",
  31316=>"011100110",
  31317=>"001010000",
  31318=>"100100111",
  31319=>"100111100",
  31320=>"110001110",
  31321=>"001100010",
  31322=>"010110001",
  31323=>"010010110",
  31324=>"010000100",
  31325=>"000000000",
  31326=>"101000110",
  31327=>"100111000",
  31328=>"000100110",
  31329=>"111001010",
  31330=>"101110011",
  31331=>"111000010",
  31332=>"011111001",
  31333=>"001000000",
  31334=>"001001000",
  31335=>"011011100",
  31336=>"000011001",
  31337=>"001100110",
  31338=>"000011010",
  31339=>"011000111",
  31340=>"111000011",
  31341=>"001110000",
  31342=>"000111010",
  31343=>"001001101",
  31344=>"011001000",
  31345=>"111001010",
  31346=>"110101101",
  31347=>"000000110",
  31348=>"111011110",
  31349=>"111011010",
  31350=>"011111011",
  31351=>"111110110",
  31352=>"010010011",
  31353=>"111110010",
  31354=>"100111010",
  31355=>"100100011",
  31356=>"100000010",
  31357=>"111110111",
  31358=>"010101011",
  31359=>"101110011",
  31360=>"010000000",
  31361=>"110001100",
  31362=>"000011101",
  31363=>"101001100",
  31364=>"000000011",
  31365=>"001100101",
  31366=>"000101110",
  31367=>"101101110",
  31368=>"101000101",
  31369=>"111101111",
  31370=>"100111001",
  31371=>"110011111",
  31372=>"010111011",
  31373=>"110101011",
  31374=>"111011110",
  31375=>"010010010",
  31376=>"011110101",
  31377=>"000110101",
  31378=>"001001111",
  31379=>"100100101",
  31380=>"110001000",
  31381=>"111111110",
  31382=>"110000100",
  31383=>"101100011",
  31384=>"101011110",
  31385=>"100001011",
  31386=>"101001110",
  31387=>"111010110",
  31388=>"101001000",
  31389=>"001010010",
  31390=>"011001100",
  31391=>"011001001",
  31392=>"100001010",
  31393=>"000001010",
  31394=>"101110110",
  31395=>"011011001",
  31396=>"101001001",
  31397=>"000000011",
  31398=>"011111100",
  31399=>"000010111",
  31400=>"100001001",
  31401=>"101110001",
  31402=>"000111001",
  31403=>"110000111",
  31404=>"000001101",
  31405=>"111101110",
  31406=>"110010100",
  31407=>"011100101",
  31408=>"110011010",
  31409=>"011101010",
  31410=>"101100101",
  31411=>"011111101",
  31412=>"100111110",
  31413=>"011101000",
  31414=>"100010010",
  31415=>"000101101",
  31416=>"110101011",
  31417=>"000110101",
  31418=>"000001000",
  31419=>"000010000",
  31420=>"000100100",
  31421=>"000001011",
  31422=>"001011011",
  31423=>"110000011",
  31424=>"101111010",
  31425=>"100000011",
  31426=>"011011001",
  31427=>"010001010",
  31428=>"011100111",
  31429=>"100100111",
  31430=>"010110001",
  31431=>"000101101",
  31432=>"011111010",
  31433=>"101011101",
  31434=>"000101000",
  31435=>"110100010",
  31436=>"001010001",
  31437=>"000100001",
  31438=>"100000110",
  31439=>"000000010",
  31440=>"101001011",
  31441=>"100010100",
  31442=>"010100001",
  31443=>"001011100",
  31444=>"000000010",
  31445=>"111111010",
  31446=>"011000010",
  31447=>"000011111",
  31448=>"101010111",
  31449=>"011000011",
  31450=>"010111100",
  31451=>"010010110",
  31452=>"111111000",
  31453=>"011101111",
  31454=>"001111100",
  31455=>"010110011",
  31456=>"000001011",
  31457=>"110111011",
  31458=>"100000100",
  31459=>"111110111",
  31460=>"101010100",
  31461=>"011010101",
  31462=>"111010001",
  31463=>"101011101",
  31464=>"000101001",
  31465=>"011111011",
  31466=>"100010110",
  31467=>"111000000",
  31468=>"010100011",
  31469=>"101010011",
  31470=>"011100001",
  31471=>"000110010",
  31472=>"100111000",
  31473=>"000001101",
  31474=>"000010000",
  31475=>"001110110",
  31476=>"010100001",
  31477=>"001111011",
  31478=>"111100111",
  31479=>"110111110",
  31480=>"010111110",
  31481=>"110100100",
  31482=>"110101101",
  31483=>"100110011",
  31484=>"011110010",
  31485=>"011111000",
  31486=>"101000101",
  31487=>"100100010",
  31488=>"000001100",
  31489=>"111111010",
  31490=>"110111101",
  31491=>"001101101",
  31492=>"000111001",
  31493=>"011000001",
  31494=>"111101010",
  31495=>"011110110",
  31496=>"010000000",
  31497=>"101111011",
  31498=>"001000001",
  31499=>"101111001",
  31500=>"010100011",
  31501=>"111101010",
  31502=>"010000110",
  31503=>"010101100",
  31504=>"101101011",
  31505=>"101010011",
  31506=>"110011101",
  31507=>"100111101",
  31508=>"111110111",
  31509=>"011000100",
  31510=>"010001000",
  31511=>"001110100",
  31512=>"101111010",
  31513=>"110110101",
  31514=>"011010011",
  31515=>"110100000",
  31516=>"011000100",
  31517=>"110010000",
  31518=>"000010000",
  31519=>"010001100",
  31520=>"100111000",
  31521=>"010101100",
  31522=>"101011111",
  31523=>"110100100",
  31524=>"000110010",
  31525=>"111001000",
  31526=>"110100010",
  31527=>"111011111",
  31528=>"110001111",
  31529=>"010011110",
  31530=>"111000100",
  31531=>"011010010",
  31532=>"111010001",
  31533=>"010001010",
  31534=>"110000101",
  31535=>"101010000",
  31536=>"010011000",
  31537=>"100100100",
  31538=>"101110100",
  31539=>"100110100",
  31540=>"110111000",
  31541=>"010110010",
  31542=>"000011101",
  31543=>"000010011",
  31544=>"101011101",
  31545=>"000010000",
  31546=>"000110010",
  31547=>"011111000",
  31548=>"010001000",
  31549=>"001100001",
  31550=>"000000000",
  31551=>"010001100",
  31552=>"100011011",
  31553=>"110100111",
  31554=>"011001010",
  31555=>"011110011",
  31556=>"100110100",
  31557=>"001111110",
  31558=>"001111000",
  31559=>"000001110",
  31560=>"011110111",
  31561=>"101111111",
  31562=>"001100010",
  31563=>"110011011",
  31564=>"010100110",
  31565=>"101111110",
  31566=>"110001001",
  31567=>"110010010",
  31568=>"000100100",
  31569=>"111010011",
  31570=>"010111011",
  31571=>"000110011",
  31572=>"010101010",
  31573=>"100101100",
  31574=>"000110000",
  31575=>"010001000",
  31576=>"111110101",
  31577=>"011110111",
  31578=>"010011011",
  31579=>"010011000",
  31580=>"011110011",
  31581=>"000001110",
  31582=>"000100111",
  31583=>"010001111",
  31584=>"000111010",
  31585=>"111001111",
  31586=>"000000100",
  31587=>"011000001",
  31588=>"101110110",
  31589=>"000001010",
  31590=>"110100100",
  31591=>"101100010",
  31592=>"111111110",
  31593=>"101001001",
  31594=>"111011000",
  31595=>"011000101",
  31596=>"001000000",
  31597=>"111001000",
  31598=>"001001011",
  31599=>"000000000",
  31600=>"011110001",
  31601=>"100000011",
  31602=>"110100100",
  31603=>"110111010",
  31604=>"000010110",
  31605=>"011000001",
  31606=>"110110100",
  31607=>"100010100",
  31608=>"110110001",
  31609=>"111101101",
  31610=>"000110111",
  31611=>"111100110",
  31612=>"010010001",
  31613=>"110110100",
  31614=>"011010100",
  31615=>"001001011",
  31616=>"011111000",
  31617=>"100000001",
  31618=>"000100111",
  31619=>"100000101",
  31620=>"000010000",
  31621=>"011111101",
  31622=>"011000110",
  31623=>"111011111",
  31624=>"111010000",
  31625=>"100100011",
  31626=>"100101001",
  31627=>"010110001",
  31628=>"000111001",
  31629=>"111100110",
  31630=>"111000110",
  31631=>"100110000",
  31632=>"111101110",
  31633=>"100000110",
  31634=>"000000000",
  31635=>"100011110",
  31636=>"001100100",
  31637=>"010111100",
  31638=>"001001101",
  31639=>"100101111",
  31640=>"011010100",
  31641=>"100000001",
  31642=>"010110001",
  31643=>"110000011",
  31644=>"000100110",
  31645=>"000001101",
  31646=>"011001110",
  31647=>"111111100",
  31648=>"001010010",
  31649=>"101010010",
  31650=>"100110001",
  31651=>"001010110",
  31652=>"001110011",
  31653=>"111111111",
  31654=>"101000001",
  31655=>"111111100",
  31656=>"110001111",
  31657=>"110111011",
  31658=>"100111011",
  31659=>"000111100",
  31660=>"001000001",
  31661=>"110011010",
  31662=>"100111110",
  31663=>"111111110",
  31664=>"100110101",
  31665=>"011111110",
  31666=>"011100010",
  31667=>"101100010",
  31668=>"111111010",
  31669=>"001000010",
  31670=>"011111110",
  31671=>"100101011",
  31672=>"100100101",
  31673=>"011110101",
  31674=>"111010110",
  31675=>"001011011",
  31676=>"110011100",
  31677=>"101111000",
  31678=>"001011011",
  31679=>"001000010",
  31680=>"110000100",
  31681=>"000111101",
  31682=>"111110010",
  31683=>"101100000",
  31684=>"010000110",
  31685=>"100001110",
  31686=>"111111001",
  31687=>"111111100",
  31688=>"010011011",
  31689=>"110001110",
  31690=>"011100111",
  31691=>"101111111",
  31692=>"110010010",
  31693=>"010111010",
  31694=>"000101110",
  31695=>"111101110",
  31696=>"000100110",
  31697=>"101000001",
  31698=>"100101100",
  31699=>"011011000",
  31700=>"000110110",
  31701=>"001011010",
  31702=>"000101000",
  31703=>"111101101",
  31704=>"111011001",
  31705=>"010000111",
  31706=>"101110101",
  31707=>"111010010",
  31708=>"010111101",
  31709=>"011101110",
  31710=>"010000000",
  31711=>"011011001",
  31712=>"111111111",
  31713=>"000110000",
  31714=>"111100100",
  31715=>"001000011",
  31716=>"111101010",
  31717=>"000101010",
  31718=>"010000000",
  31719=>"010111001",
  31720=>"000101000",
  31721=>"111110001",
  31722=>"010000001",
  31723=>"010011110",
  31724=>"110111111",
  31725=>"010111101",
  31726=>"010111011",
  31727=>"111000001",
  31728=>"000101001",
  31729=>"101100010",
  31730=>"101011111",
  31731=>"000100000",
  31732=>"000101001",
  31733=>"101111101",
  31734=>"111011110",
  31735=>"110001111",
  31736=>"011001111",
  31737=>"110111000",
  31738=>"000000000",
  31739=>"000111111",
  31740=>"111101010",
  31741=>"110100000",
  31742=>"011111110",
  31743=>"010011001",
  31744=>"111101011",
  31745=>"010101011",
  31746=>"011111101",
  31747=>"001010110",
  31748=>"000011000",
  31749=>"011000000",
  31750=>"111011011",
  31751=>"001111101",
  31752=>"101100111",
  31753=>"010011100",
  31754=>"110101010",
  31755=>"110011110",
  31756=>"001001011",
  31757=>"110011001",
  31758=>"111001100",
  31759=>"110110111",
  31760=>"000010001",
  31761=>"000100111",
  31762=>"000111100",
  31763=>"000110001",
  31764=>"001000100",
  31765=>"101000101",
  31766=>"110110111",
  31767=>"111100101",
  31768=>"010000001",
  31769=>"011000000",
  31770=>"111011001",
  31771=>"001001110",
  31772=>"100110010",
  31773=>"100010101",
  31774=>"110000001",
  31775=>"100101110",
  31776=>"001011111",
  31777=>"111101110",
  31778=>"010101000",
  31779=>"101000111",
  31780=>"111101010",
  31781=>"011011010",
  31782=>"000101001",
  31783=>"100011001",
  31784=>"011011011",
  31785=>"011011101",
  31786=>"011011111",
  31787=>"010111000",
  31788=>"111011111",
  31789=>"010111111",
  31790=>"110011011",
  31791=>"100101110",
  31792=>"010001111",
  31793=>"101010101",
  31794=>"101000101",
  31795=>"110110110",
  31796=>"100001100",
  31797=>"001111011",
  31798=>"110101111",
  31799=>"101100000",
  31800=>"101000100",
  31801=>"100100111",
  31802=>"000101101",
  31803=>"100110000",
  31804=>"110111000",
  31805=>"111000110",
  31806=>"000010110",
  31807=>"000010011",
  31808=>"000100100",
  31809=>"100010010",
  31810=>"101000000",
  31811=>"111100100",
  31812=>"111011011",
  31813=>"100101101",
  31814=>"111111100",
  31815=>"100101000",
  31816=>"010101011",
  31817=>"101011010",
  31818=>"000011011",
  31819=>"000111110",
  31820=>"011000000",
  31821=>"110110110",
  31822=>"100000110",
  31823=>"111101111",
  31824=>"000110111",
  31825=>"111001011",
  31826=>"101100010",
  31827=>"111110101",
  31828=>"011010010",
  31829=>"100110111",
  31830=>"000110011",
  31831=>"010100011",
  31832=>"000101100",
  31833=>"101011111",
  31834=>"001110000",
  31835=>"001100000",
  31836=>"100001101",
  31837=>"111111011",
  31838=>"101010100",
  31839=>"011110011",
  31840=>"111101001",
  31841=>"011101110",
  31842=>"111011100",
  31843=>"000100101",
  31844=>"000001100",
  31845=>"111101110",
  31846=>"110011001",
  31847=>"101110111",
  31848=>"101011010",
  31849=>"111110011",
  31850=>"100100111",
  31851=>"100101000",
  31852=>"001010100",
  31853=>"010001011",
  31854=>"100101001",
  31855=>"001000111",
  31856=>"011001000",
  31857=>"110101110",
  31858=>"100011010",
  31859=>"110010100",
  31860=>"110001010",
  31861=>"110000011",
  31862=>"111001110",
  31863=>"110001010",
  31864=>"010110110",
  31865=>"011111100",
  31866=>"111011010",
  31867=>"101111000",
  31868=>"010000001",
  31869=>"010010011",
  31870=>"101011000",
  31871=>"011111101",
  31872=>"111110100",
  31873=>"001100100",
  31874=>"001000100",
  31875=>"010011101",
  31876=>"001000000",
  31877=>"111100101",
  31878=>"001111110",
  31879=>"111001001",
  31880=>"111001011",
  31881=>"000110011",
  31882=>"111101001",
  31883=>"110101001",
  31884=>"101100111",
  31885=>"000001101",
  31886=>"010011001",
  31887=>"011001100",
  31888=>"110001101",
  31889=>"010111110",
  31890=>"100001000",
  31891=>"001011101",
  31892=>"011111100",
  31893=>"001100000",
  31894=>"110010100",
  31895=>"010111001",
  31896=>"100011001",
  31897=>"000100111",
  31898=>"001011000",
  31899=>"011111011",
  31900=>"111101011",
  31901=>"010111100",
  31902=>"001000100",
  31903=>"000111101",
  31904=>"011111001",
  31905=>"001001000",
  31906=>"111101111",
  31907=>"110000010",
  31908=>"001101111",
  31909=>"010100000",
  31910=>"010001101",
  31911=>"001111010",
  31912=>"101111011",
  31913=>"001101010",
  31914=>"000111000",
  31915=>"110101100",
  31916=>"000000001",
  31917=>"111101001",
  31918=>"111011111",
  31919=>"101000111",
  31920=>"011110011",
  31921=>"001100111",
  31922=>"010110101",
  31923=>"100001001",
  31924=>"010001110",
  31925=>"011111111",
  31926=>"000110100",
  31927=>"111111111",
  31928=>"110100101",
  31929=>"111001011",
  31930=>"001100011",
  31931=>"111001011",
  31932=>"111001111",
  31933=>"111110010",
  31934=>"010011110",
  31935=>"100011010",
  31936=>"011110100",
  31937=>"001101010",
  31938=>"010000011",
  31939=>"011011110",
  31940=>"100010111",
  31941=>"101001010",
  31942=>"001100110",
  31943=>"010000000",
  31944=>"101101000",
  31945=>"100110001",
  31946=>"000100111",
  31947=>"000001001",
  31948=>"000010101",
  31949=>"100111001",
  31950=>"000100000",
  31951=>"000001011",
  31952=>"110101111",
  31953=>"000000001",
  31954=>"000011110",
  31955=>"100110101",
  31956=>"101111111",
  31957=>"001101100",
  31958=>"000010101",
  31959=>"100101110",
  31960=>"000101101",
  31961=>"110000000",
  31962=>"010011001",
  31963=>"000101000",
  31964=>"010010010",
  31965=>"101101010",
  31966=>"001000101",
  31967=>"101100100",
  31968=>"011001000",
  31969=>"111010011",
  31970=>"001110011",
  31971=>"000110101",
  31972=>"000111101",
  31973=>"101010000",
  31974=>"001000010",
  31975=>"000110100",
  31976=>"100111101",
  31977=>"101010110",
  31978=>"011000001",
  31979=>"100010110",
  31980=>"000101001",
  31981=>"000100111",
  31982=>"111111011",
  31983=>"100110010",
  31984=>"001111110",
  31985=>"001111010",
  31986=>"111000111",
  31987=>"111011011",
  31988=>"000110001",
  31989=>"111010100",
  31990=>"010010100",
  31991=>"111010001",
  31992=>"011011110",
  31993=>"010010111",
  31994=>"010101000",
  31995=>"000010110",
  31996=>"001111001",
  31997=>"000000010",
  31998=>"001010000",
  31999=>"000001000",
  32000=>"100010001",
  32001=>"011111000",
  32002=>"101011010",
  32003=>"100001100",
  32004=>"011111100",
  32005=>"010011110",
  32006=>"101010010",
  32007=>"011110111",
  32008=>"000110001",
  32009=>"010010010",
  32010=>"100100001",
  32011=>"110000110",
  32012=>"110110001",
  32013=>"111011000",
  32014=>"111010111",
  32015=>"100010011",
  32016=>"000000101",
  32017=>"110110011",
  32018=>"110001101",
  32019=>"110101101",
  32020=>"101111110",
  32021=>"100011110",
  32022=>"001000000",
  32023=>"101001011",
  32024=>"011101100",
  32025=>"110101001",
  32026=>"110000110",
  32027=>"110011110",
  32028=>"010000000",
  32029=>"111100111",
  32030=>"001111111",
  32031=>"010011011",
  32032=>"100101100",
  32033=>"001000111",
  32034=>"101000010",
  32035=>"100110001",
  32036=>"101001110",
  32037=>"010100101",
  32038=>"011011111",
  32039=>"010100001",
  32040=>"111110111",
  32041=>"010010001",
  32042=>"011110011",
  32043=>"100111010",
  32044=>"110101111",
  32045=>"001111011",
  32046=>"000111101",
  32047=>"110101110",
  32048=>"111110111",
  32049=>"000101101",
  32050=>"001110011",
  32051=>"000000101",
  32052=>"110010001",
  32053=>"010100101",
  32054=>"100011110",
  32055=>"110001110",
  32056=>"101010001",
  32057=>"110110101",
  32058=>"111110110",
  32059=>"010100010",
  32060=>"101111100",
  32061=>"110100000",
  32062=>"110000011",
  32063=>"011000111",
  32064=>"101001010",
  32065=>"000101000",
  32066=>"111110111",
  32067=>"111000000",
  32068=>"111111010",
  32069=>"101110111",
  32070=>"001010001",
  32071=>"010101001",
  32072=>"001001101",
  32073=>"110101101",
  32074=>"010111000",
  32075=>"010011110",
  32076=>"100010111",
  32077=>"001100001",
  32078=>"100110011",
  32079=>"000011011",
  32080=>"111111100",
  32081=>"110111000",
  32082=>"111010101",
  32083=>"111001000",
  32084=>"111111010",
  32085=>"101011010",
  32086=>"010001011",
  32087=>"110111111",
  32088=>"100110011",
  32089=>"111000001",
  32090=>"000010001",
  32091=>"011110011",
  32092=>"001000100",
  32093=>"011100011",
  32094=>"000000001",
  32095=>"001011010",
  32096=>"110010110",
  32097=>"010000101",
  32098=>"110100010",
  32099=>"010111111",
  32100=>"110010010",
  32101=>"001010011",
  32102=>"000100111",
  32103=>"111100001",
  32104=>"010111001",
  32105=>"000010111",
  32106=>"011100000",
  32107=>"111011101",
  32108=>"100011100",
  32109=>"110111010",
  32110=>"010001000",
  32111=>"111010100",
  32112=>"010111010",
  32113=>"000000111",
  32114=>"111101101",
  32115=>"100101111",
  32116=>"000001011",
  32117=>"010100011",
  32118=>"010000001",
  32119=>"011110010",
  32120=>"111110100",
  32121=>"010111010",
  32122=>"100000101",
  32123=>"100001100",
  32124=>"101000101",
  32125=>"001011110",
  32126=>"111110011",
  32127=>"111110010",
  32128=>"010101100",
  32129=>"000110011",
  32130=>"110011000",
  32131=>"001001111",
  32132=>"000110010",
  32133=>"001101011",
  32134=>"100001010",
  32135=>"011101011",
  32136=>"010100110",
  32137=>"111011000",
  32138=>"100111011",
  32139=>"011001111",
  32140=>"000010010",
  32141=>"001111100",
  32142=>"010001101",
  32143=>"011010001",
  32144=>"111011101",
  32145=>"111001101",
  32146=>"011001100",
  32147=>"111110011",
  32148=>"010100100",
  32149=>"010001000",
  32150=>"000010101",
  32151=>"101100001",
  32152=>"010001000",
  32153=>"000010110",
  32154=>"011011100",
  32155=>"010111111",
  32156=>"100100001",
  32157=>"011000000",
  32158=>"000010001",
  32159=>"010010001",
  32160=>"000011010",
  32161=>"101100000",
  32162=>"011111010",
  32163=>"100001110",
  32164=>"011100000",
  32165=>"000010110",
  32166=>"100100011",
  32167=>"110000011",
  32168=>"010011111",
  32169=>"111101001",
  32170=>"000100000",
  32171=>"010111110",
  32172=>"110001111",
  32173=>"100011000",
  32174=>"011110111",
  32175=>"111000001",
  32176=>"100100110",
  32177=>"111110011",
  32178=>"111100000",
  32179=>"111001001",
  32180=>"101010100",
  32181=>"011010101",
  32182=>"101100101",
  32183=>"001001101",
  32184=>"100000111",
  32185=>"000101101",
  32186=>"110110000",
  32187=>"111011010",
  32188=>"011100111",
  32189=>"111000100",
  32190=>"111100001",
  32191=>"011010010",
  32192=>"110001100",
  32193=>"011110011",
  32194=>"010001111",
  32195=>"010101101",
  32196=>"100000110",
  32197=>"010000100",
  32198=>"001100111",
  32199=>"111101110",
  32200=>"101111110",
  32201=>"100001101",
  32202=>"010011111",
  32203=>"111110101",
  32204=>"110111001",
  32205=>"111001101",
  32206=>"000101111",
  32207=>"011111000",
  32208=>"100100111",
  32209=>"100110110",
  32210=>"100110001",
  32211=>"111001001",
  32212=>"101111111",
  32213=>"101000111",
  32214=>"110011010",
  32215=>"101001110",
  32216=>"111000011",
  32217=>"110110111",
  32218=>"011101010",
  32219=>"001000101",
  32220=>"010100011",
  32221=>"000000100",
  32222=>"100111111",
  32223=>"110011001",
  32224=>"110010001",
  32225=>"011110101",
  32226=>"101000110",
  32227=>"001010000",
  32228=>"111100010",
  32229=>"111011111",
  32230=>"000111010",
  32231=>"100001110",
  32232=>"000011111",
  32233=>"110011101",
  32234=>"001001101",
  32235=>"101101111",
  32236=>"110001110",
  32237=>"000101001",
  32238=>"000010111",
  32239=>"111100010",
  32240=>"101000100",
  32241=>"011001011",
  32242=>"011110000",
  32243=>"010100110",
  32244=>"101111010",
  32245=>"111101001",
  32246=>"010101110",
  32247=>"110000000",
  32248=>"101101100",
  32249=>"011010010",
  32250=>"000101110",
  32251=>"010011001",
  32252=>"100001000",
  32253=>"111000011",
  32254=>"000011101",
  32255=>"000100001",
  32256=>"110011110",
  32257=>"001100010",
  32258=>"100101101",
  32259=>"111111110",
  32260=>"011000011",
  32261=>"101110001",
  32262=>"110110100",
  32263=>"110100110",
  32264=>"000000100",
  32265=>"001001011",
  32266=>"101101000",
  32267=>"010100001",
  32268=>"101100101",
  32269=>"110001001",
  32270=>"111101001",
  32271=>"100000000",
  32272=>"010001010",
  32273=>"110101110",
  32274=>"110101111",
  32275=>"111001000",
  32276=>"010010000",
  32277=>"001011111",
  32278=>"111000011",
  32279=>"100101000",
  32280=>"111000011",
  32281=>"111100011",
  32282=>"000001001",
  32283=>"110001000",
  32284=>"001100010",
  32285=>"111000101",
  32286=>"001100100",
  32287=>"101110101",
  32288=>"010000010",
  32289=>"101001100",
  32290=>"000001010",
  32291=>"010110000",
  32292=>"100110101",
  32293=>"101100110",
  32294=>"100101000",
  32295=>"010001001",
  32296=>"011100110",
  32297=>"110010011",
  32298=>"110010110",
  32299=>"011110111",
  32300=>"111010011",
  32301=>"101111100",
  32302=>"111000010",
  32303=>"110011111",
  32304=>"101100010",
  32305=>"111100000",
  32306=>"110110111",
  32307=>"111000100",
  32308=>"010101001",
  32309=>"111111000",
  32310=>"001010001",
  32311=>"111100111",
  32312=>"101110111",
  32313=>"001011011",
  32314=>"001001000",
  32315=>"000110100",
  32316=>"101110011",
  32317=>"000110101",
  32318=>"100100101",
  32319=>"000001010",
  32320=>"010100010",
  32321=>"110100101",
  32322=>"011000000",
  32323=>"101100110",
  32324=>"000010111",
  32325=>"111011111",
  32326=>"100000110",
  32327=>"010100000",
  32328=>"110110110",
  32329=>"010010010",
  32330=>"110010110",
  32331=>"001101110",
  32332=>"100110101",
  32333=>"001100100",
  32334=>"110001101",
  32335=>"010011101",
  32336=>"101101011",
  32337=>"110110011",
  32338=>"101101000",
  32339=>"100011111",
  32340=>"101110001",
  32341=>"110110111",
  32342=>"000010101",
  32343=>"001011010",
  32344=>"110111110",
  32345=>"010110101",
  32346=>"010110010",
  32347=>"000000000",
  32348=>"000011010",
  32349=>"011111110",
  32350=>"000000110",
  32351=>"001111001",
  32352=>"110000100",
  32353=>"011011000",
  32354=>"101010000",
  32355=>"100000101",
  32356=>"001011001",
  32357=>"011000000",
  32358=>"111100010",
  32359=>"111111001",
  32360=>"001101110",
  32361=>"101011010",
  32362=>"001110000",
  32363=>"010100111",
  32364=>"011011001",
  32365=>"010101011",
  32366=>"111111111",
  32367=>"001001101",
  32368=>"101000010",
  32369=>"100000010",
  32370=>"011101101",
  32371=>"101111101",
  32372=>"010101111",
  32373=>"111111111",
  32374=>"000000000",
  32375=>"011111011",
  32376=>"100101000",
  32377=>"001110101",
  32378=>"010111101",
  32379=>"110101101",
  32380=>"001101100",
  32381=>"101110101",
  32382=>"011010101",
  32383=>"101010001",
  32384=>"111010101",
  32385=>"110001011",
  32386=>"100010000",
  32387=>"001001010",
  32388=>"001101000",
  32389=>"111100110",
  32390=>"100010010",
  32391=>"110001101",
  32392=>"100101010",
  32393=>"101101110",
  32394=>"111000010",
  32395=>"100110111",
  32396=>"110000001",
  32397=>"110001011",
  32398=>"110111001",
  32399=>"110000001",
  32400=>"010101110",
  32401=>"111001100",
  32402=>"000000010",
  32403=>"101000101",
  32404=>"111100000",
  32405=>"000101010",
  32406=>"001110001",
  32407=>"111101111",
  32408=>"100010101",
  32409=>"011001010",
  32410=>"101000000",
  32411=>"111110010",
  32412=>"111110001",
  32413=>"110001101",
  32414=>"110111100",
  32415=>"011010001",
  32416=>"110101011",
  32417=>"000110101",
  32418=>"100001110",
  32419=>"010101000",
  32420=>"101101000",
  32421=>"001101100",
  32422=>"101110111",
  32423=>"110111000",
  32424=>"111010111",
  32425=>"000101010",
  32426=>"111010110",
  32427=>"011110010",
  32428=>"110011001",
  32429=>"011011010",
  32430=>"001010010",
  32431=>"001101111",
  32432=>"001001100",
  32433=>"000011000",
  32434=>"000010001",
  32435=>"010100101",
  32436=>"000111110",
  32437=>"011100001",
  32438=>"011001011",
  32439=>"100011001",
  32440=>"100011011",
  32441=>"010100100",
  32442=>"110010000",
  32443=>"010011000",
  32444=>"001001101",
  32445=>"100100010",
  32446=>"000100111",
  32447=>"000000001",
  32448=>"110000000",
  32449=>"110100011",
  32450=>"000011001",
  32451=>"111111100",
  32452=>"111010000",
  32453=>"101010110",
  32454=>"001010100",
  32455=>"000010101",
  32456=>"100100010",
  32457=>"110110010",
  32458=>"101101001",
  32459=>"011011010",
  32460=>"110101110",
  32461=>"000111111",
  32462=>"110000011",
  32463=>"100101000",
  32464=>"100010100",
  32465=>"001001000",
  32466=>"111110101",
  32467=>"101000010",
  32468=>"000000000",
  32469=>"011010101",
  32470=>"100001000",
  32471=>"001101010",
  32472=>"000101100",
  32473=>"011011000",
  32474=>"000101011",
  32475=>"001011011",
  32476=>"000110001",
  32477=>"011010100",
  32478=>"000111101",
  32479=>"001010100",
  32480=>"100111010",
  32481=>"000111010",
  32482=>"010100011",
  32483=>"001000111",
  32484=>"011000101",
  32485=>"111010010",
  32486=>"011100111",
  32487=>"001101110",
  32488=>"111011110",
  32489=>"101101001",
  32490=>"110011011",
  32491=>"000011000",
  32492=>"100110101",
  32493=>"011001001",
  32494=>"111110101",
  32495=>"100000010",
  32496=>"110001000",
  32497=>"001000110",
  32498=>"110111011",
  32499=>"111100110",
  32500=>"100001101",
  32501=>"001001011",
  32502=>"100001111",
  32503=>"110000001",
  32504=>"100111111",
  32505=>"001101000",
  32506=>"101110001",
  32507=>"100001100",
  32508=>"011100100",
  32509=>"000100110",
  32510=>"110101110",
  32511=>"100101110",
  32512=>"000010100",
  32513=>"000101000",
  32514=>"101111000",
  32515=>"101010000",
  32516=>"000101101",
  32517=>"101011010",
  32518=>"110111111",
  32519=>"001001000",
  32520=>"010110100",
  32521=>"101100000",
  32522=>"000100111",
  32523=>"101100100",
  32524=>"011101101",
  32525=>"011011000",
  32526=>"100010100",
  32527=>"000110100",
  32528=>"001100111",
  32529=>"110011010",
  32530=>"011111011",
  32531=>"001101001",
  32532=>"010010011",
  32533=>"110001111",
  32534=>"000101101",
  32535=>"001001101",
  32536=>"010110110",
  32537=>"000011110",
  32538=>"000010100",
  32539=>"111101000",
  32540=>"000010100",
  32541=>"010111000",
  32542=>"101110011",
  32543=>"111000001",
  32544=>"100001011",
  32545=>"101011111",
  32546=>"010110010",
  32547=>"011000000",
  32548=>"110010011",
  32549=>"111111110",
  32550=>"001001001",
  32551=>"100010011",
  32552=>"010010001",
  32553=>"111000010",
  32554=>"000100101",
  32555=>"101111110",
  32556=>"001101101",
  32557=>"000111101",
  32558=>"001001111",
  32559=>"000101100",
  32560=>"010100011",
  32561=>"111101001",
  32562=>"000111001",
  32563=>"110100110",
  32564=>"100000111",
  32565=>"111011100",
  32566=>"001000001",
  32567=>"011101101",
  32568=>"101010101",
  32569=>"110001101",
  32570=>"010001110",
  32571=>"110110011",
  32572=>"010101111",
  32573=>"000010110",
  32574=>"110101010",
  32575=>"100101110",
  32576=>"111011101",
  32577=>"001010111",
  32578=>"101111101",
  32579=>"111101010",
  32580=>"011011111",
  32581=>"000110000",
  32582=>"010000111",
  32583=>"001110010",
  32584=>"011111111",
  32585=>"010001101",
  32586=>"111110001",
  32587=>"110111001",
  32588=>"001011000",
  32589=>"010010100",
  32590=>"101110100",
  32591=>"111000001",
  32592=>"011011000",
  32593=>"100011111",
  32594=>"111101001",
  32595=>"010011001",
  32596=>"101001001",
  32597=>"000111000",
  32598=>"011100000",
  32599=>"100100000",
  32600=>"010011000",
  32601=>"011010011",
  32602=>"010111001",
  32603=>"110100001",
  32604=>"010100100",
  32605=>"001101110",
  32606=>"001011110",
  32607=>"100100110",
  32608=>"011010100",
  32609=>"110100110",
  32610=>"100101011",
  32611=>"011010011",
  32612=>"011001010",
  32613=>"001100010",
  32614=>"101111110",
  32615=>"010100111",
  32616=>"111100110",
  32617=>"000000011",
  32618=>"101110001",
  32619=>"000111110",
  32620=>"110010100",
  32621=>"000010010",
  32622=>"110011010",
  32623=>"000000101",
  32624=>"110011001",
  32625=>"010000010",
  32626=>"111001101",
  32627=>"100110101",
  32628=>"000110110",
  32629=>"101011001",
  32630=>"010000010",
  32631=>"000000101",
  32632=>"100001100",
  32633=>"111100001",
  32634=>"011110001",
  32635=>"000111011",
  32636=>"110010000",
  32637=>"111010110",
  32638=>"100110010",
  32639=>"101101110",
  32640=>"111010101",
  32641=>"010101100",
  32642=>"000000010",
  32643=>"111010110",
  32644=>"000110001",
  32645=>"100011101",
  32646=>"101000011",
  32647=>"111011101",
  32648=>"110100110",
  32649=>"100000101",
  32650=>"000011110",
  32651=>"111010001",
  32652=>"101111011",
  32653=>"110111100",
  32654=>"110101000",
  32655=>"110101100",
  32656=>"110101111",
  32657=>"011111010",
  32658=>"000110001",
  32659=>"100011011",
  32660=>"111111110",
  32661=>"001001101",
  32662=>"000100100",
  32663=>"011000000",
  32664=>"111010100",
  32665=>"101001000",
  32666=>"101011110",
  32667=>"000000000",
  32668=>"001111001",
  32669=>"011011010",
  32670=>"000000011",
  32671=>"001011101",
  32672=>"101011010",
  32673=>"000111000",
  32674=>"100000011",
  32675=>"100101110",
  32676=>"000100101",
  32677=>"001110101",
  32678=>"000100010",
  32679=>"001011110",
  32680=>"000011001",
  32681=>"001100100",
  32682=>"100001110",
  32683=>"111110010",
  32684=>"000101101",
  32685=>"111010011",
  32686=>"111100100",
  32687=>"010110010",
  32688=>"011100100",
  32689=>"010101000",
  32690=>"111100110",
  32691=>"100101000",
  32692=>"111101111",
  32693=>"001011010",
  32694=>"001100110",
  32695=>"110100010",
  32696=>"010110110",
  32697=>"001010011",
  32698=>"000000110",
  32699=>"100101100",
  32700=>"011110101",
  32701=>"111011101",
  32702=>"111100000",
  32703=>"101010100",
  32704=>"011000111",
  32705=>"000011010",
  32706=>"011110011",
  32707=>"111110010",
  32708=>"011010001",
  32709=>"101110100",
  32710=>"111001110",
  32711=>"101000010",
  32712=>"010001100",
  32713=>"010011111",
  32714=>"000001001",
  32715=>"110110111",
  32716=>"101101010",
  32717=>"111100000",
  32718=>"011001111",
  32719=>"011110101",
  32720=>"000001001",
  32721=>"011111111",
  32722=>"001111000",
  32723=>"011100000",
  32724=>"111100110",
  32725=>"110011000",
  32726=>"011011011",
  32727=>"011101011",
  32728=>"000110101",
  32729=>"100001111",
  32730=>"010001111",
  32731=>"111110100",
  32732=>"000101000",
  32733=>"111001001",
  32734=>"010110101",
  32735=>"000001110",
  32736=>"110111100",
  32737=>"010111011",
  32738=>"101111001",
  32739=>"001011000",
  32740=>"011010111",
  32741=>"000100010",
  32742=>"100100001",
  32743=>"000101011",
  32744=>"001100100",
  32745=>"000010110",
  32746=>"100101110",
  32747=>"101100000",
  32748=>"101011010",
  32749=>"110100001",
  32750=>"001000011",
  32751=>"001101111",
  32752=>"010100101",
  32753=>"111010000",
  32754=>"101000100",
  32755=>"111011110",
  32756=>"100010001",
  32757=>"011010011",
  32758=>"110001011",
  32759=>"100001001",
  32760=>"110010000",
  32761=>"101110101",
  32762=>"100101001",
  32763=>"110101101",
  32764=>"110001001",
  32765=>"111010100",
  32766=>"001100110",
  32767=>"111001110",
  32768=>"110001010",
  32769=>"111111000",
  32770=>"101000101",
  32771=>"101011000",
  32772=>"010101100",
  32773=>"111100000",
  32774=>"101001111",
  32775=>"101110111",
  32776=>"001110100",
  32777=>"100100111",
  32778=>"111100111",
  32779=>"011111011",
  32780=>"101010011",
  32781=>"011000011",
  32782=>"010001111",
  32783=>"010011011",
  32784=>"111100011",
  32785=>"010110000",
  32786=>"110100000",
  32787=>"000110100",
  32788=>"000011111",
  32789=>"011110110",
  32790=>"111001101",
  32791=>"010001001",
  32792=>"111110000",
  32793=>"000100000",
  32794=>"010011111",
  32795=>"111010100",
  32796=>"001100110",
  32797=>"101100011",
  32798=>"100100000",
  32799=>"000110000",
  32800=>"001100101",
  32801=>"100100010",
  32802=>"011110101",
  32803=>"100011011",
  32804=>"011001101",
  32805=>"001000001",
  32806=>"010010010",
  32807=>"110010101",
  32808=>"100010001",
  32809=>"000010110",
  32810=>"001010110",
  32811=>"011001011",
  32812=>"001001111",
  32813=>"100110100",
  32814=>"001011010",
  32815=>"100010011",
  32816=>"100000100",
  32817=>"011011100",
  32818=>"101101110",
  32819=>"111110000",
  32820=>"111110010",
  32821=>"011110001",
  32822=>"000110110",
  32823=>"000100010",
  32824=>"111001111",
  32825=>"111111001",
  32826=>"000011011",
  32827=>"101010111",
  32828=>"110111100",
  32829=>"000001011",
  32830=>"001111111",
  32831=>"011001100",
  32832=>"110001100",
  32833=>"110010010",
  32834=>"001101110",
  32835=>"010000111",
  32836=>"110101111",
  32837=>"001100101",
  32838=>"110111000",
  32839=>"111000000",
  32840=>"000010001",
  32841=>"010111111",
  32842=>"010001010",
  32843=>"000011100",
  32844=>"000000011",
  32845=>"011100100",
  32846=>"101010100",
  32847=>"010101000",
  32848=>"001001101",
  32849=>"000011000",
  32850=>"110000110",
  32851=>"010001010",
  32852=>"110110110",
  32853=>"000010010",
  32854=>"000110000",
  32855=>"110101110",
  32856=>"010011110",
  32857=>"100011001",
  32858=>"001110111",
  32859=>"011110101",
  32860=>"000110100",
  32861=>"100101110",
  32862=>"100111001",
  32863=>"010110000",
  32864=>"100001001",
  32865=>"111100111",
  32866=>"101001100",
  32867=>"010011110",
  32868=>"010001100",
  32869=>"001100110",
  32870=>"010110001",
  32871=>"100100111",
  32872=>"110111010",
  32873=>"110101000",
  32874=>"101011100",
  32875=>"010000010",
  32876=>"110101101",
  32877=>"011101001",
  32878=>"011110000",
  32879=>"010101110",
  32880=>"110111010",
  32881=>"101110010",
  32882=>"000011011",
  32883=>"001000000",
  32884=>"000001100",
  32885=>"010001000",
  32886=>"011000100",
  32887=>"010100101",
  32888=>"000100010",
  32889=>"111100101",
  32890=>"000011000",
  32891=>"000000101",
  32892=>"110000100",
  32893=>"111001000",
  32894=>"011000111",
  32895=>"000000011",
  32896=>"101001000",
  32897=>"010000000",
  32898=>"101110111",
  32899=>"000011111",
  32900=>"100100010",
  32901=>"001100111",
  32902=>"100111111",
  32903=>"110111110",
  32904=>"100111111",
  32905=>"101101010",
  32906=>"110000110",
  32907=>"110111110",
  32908=>"101101111",
  32909=>"101000011",
  32910=>"111001000",
  32911=>"101101110",
  32912=>"100010001",
  32913=>"110110000",
  32914=>"100010111",
  32915=>"101111101",
  32916=>"001101011",
  32917=>"001111011",
  32918=>"101001011",
  32919=>"011110110",
  32920=>"101100000",
  32921=>"110001111",
  32922=>"000010110",
  32923=>"101001010",
  32924=>"101010011",
  32925=>"001110111",
  32926=>"110101010",
  32927=>"001100011",
  32928=>"101000101",
  32929=>"100100111",
  32930=>"000000011",
  32931=>"000101111",
  32932=>"001110000",
  32933=>"000111011",
  32934=>"111011011",
  32935=>"001101101",
  32936=>"110000001",
  32937=>"101010111",
  32938=>"100011000",
  32939=>"111111011",
  32940=>"001011011",
  32941=>"010000111",
  32942=>"010101000",
  32943=>"010101010",
  32944=>"110001101",
  32945=>"111100100",
  32946=>"111010110",
  32947=>"000001111",
  32948=>"001001001",
  32949=>"000001001",
  32950=>"111001011",
  32951=>"000110101",
  32952=>"111101111",
  32953=>"110000100",
  32954=>"111010010",
  32955=>"111100110",
  32956=>"010111100",
  32957=>"101000100",
  32958=>"001110001",
  32959=>"110011001",
  32960=>"001000100",
  32961=>"000011000",
  32962=>"001101011",
  32963=>"110111001",
  32964=>"100101110",
  32965=>"110011110",
  32966=>"011110000",
  32967=>"100000111",
  32968=>"110111011",
  32969=>"100010110",
  32970=>"011110010",
  32971=>"100101100",
  32972=>"001001101",
  32973=>"100010011",
  32974=>"111111101",
  32975=>"111100100",
  32976=>"110011010",
  32977=>"101111010",
  32978=>"111100010",
  32979=>"001111001",
  32980=>"110011001",
  32981=>"100001111",
  32982=>"001110010",
  32983=>"000000111",
  32984=>"010011001",
  32985=>"111111001",
  32986=>"110111000",
  32987=>"000000100",
  32988=>"010011101",
  32989=>"110000110",
  32990=>"101010110",
  32991=>"001000001",
  32992=>"001011111",
  32993=>"100011111",
  32994=>"011011110",
  32995=>"000100110",
  32996=>"100000100",
  32997=>"001001100",
  32998=>"000011100",
  32999=>"001001110",
  33000=>"100111111",
  33001=>"010100011",
  33002=>"110100000",
  33003=>"011000101",
  33004=>"001010111",
  33005=>"100011111",
  33006=>"110000001",
  33007=>"000000110",
  33008=>"000111001",
  33009=>"110110010",
  33010=>"001001111",
  33011=>"010010110",
  33012=>"111111010",
  33013=>"001111111",
  33014=>"111110010",
  33015=>"010110110",
  33016=>"011101100",
  33017=>"010001000",
  33018=>"000010010",
  33019=>"100000010",
  33020=>"111001001",
  33021=>"010111000",
  33022=>"011010110",
  33023=>"110010101",
  33024=>"110011011",
  33025=>"101010000",
  33026=>"001001000",
  33027=>"000111001",
  33028=>"110001011",
  33029=>"000000010",
  33030=>"101011111",
  33031=>"011010111",
  33032=>"001001001",
  33033=>"100101000",
  33034=>"010111111",
  33035=>"110101011",
  33036=>"111001111",
  33037=>"101001000",
  33038=>"010011100",
  33039=>"111111001",
  33040=>"110110111",
  33041=>"111111001",
  33042=>"001111111",
  33043=>"011111000",
  33044=>"101010010",
  33045=>"111000000",
  33046=>"110000111",
  33047=>"010110000",
  33048=>"101001011",
  33049=>"010110010",
  33050=>"111111110",
  33051=>"100111101",
  33052=>"111010011",
  33053=>"101111000",
  33054=>"010111111",
  33055=>"001000110",
  33056=>"100110101",
  33057=>"111000000",
  33058=>"100011100",
  33059=>"010011010",
  33060=>"111001101",
  33061=>"011101000",
  33062=>"000001110",
  33063=>"011110111",
  33064=>"101111111",
  33065=>"000101001",
  33066=>"110101110",
  33067=>"001100110",
  33068=>"111011100",
  33069=>"000100000",
  33070=>"110101000",
  33071=>"000111110",
  33072=>"011110010",
  33073=>"011110001",
  33074=>"110100111",
  33075=>"001100100",
  33076=>"101011111",
  33077=>"001000011",
  33078=>"110001110",
  33079=>"000000001",
  33080=>"000111000",
  33081=>"010111101",
  33082=>"111110000",
  33083=>"000010011",
  33084=>"001100110",
  33085=>"110111011",
  33086=>"010101110",
  33087=>"110000101",
  33088=>"001011000",
  33089=>"000011010",
  33090=>"011000101",
  33091=>"000100100",
  33092=>"010010100",
  33093=>"101101100",
  33094=>"010010001",
  33095=>"100101011",
  33096=>"001000001",
  33097=>"111100000",
  33098=>"111100100",
  33099=>"000011110",
  33100=>"010010010",
  33101=>"111011000",
  33102=>"010000100",
  33103=>"101001110",
  33104=>"100010001",
  33105=>"110101010",
  33106=>"111111110",
  33107=>"001100110",
  33108=>"010110110",
  33109=>"111100010",
  33110=>"001000000",
  33111=>"011001110",
  33112=>"001100111",
  33113=>"110010101",
  33114=>"101001011",
  33115=>"000110111",
  33116=>"000011111",
  33117=>"001110110",
  33118=>"111000101",
  33119=>"010111110",
  33120=>"100111100",
  33121=>"110010001",
  33122=>"001100010",
  33123=>"110101100",
  33124=>"111100001",
  33125=>"000110111",
  33126=>"010000001",
  33127=>"111110011",
  33128=>"111010001",
  33129=>"100110111",
  33130=>"001001110",
  33131=>"001110101",
  33132=>"001001000",
  33133=>"100011011",
  33134=>"111011111",
  33135=>"011010110",
  33136=>"100101001",
  33137=>"111111110",
  33138=>"010010110",
  33139=>"010110110",
  33140=>"111110001",
  33141=>"011100111",
  33142=>"011110001",
  33143=>"100000010",
  33144=>"110001010",
  33145=>"111110000",
  33146=>"001000111",
  33147=>"111110000",
  33148=>"110001001",
  33149=>"000100110",
  33150=>"011110010",
  33151=>"000101110",
  33152=>"110101101",
  33153=>"000001010",
  33154=>"100101110",
  33155=>"110110000",
  33156=>"101001110",
  33157=>"000000110",
  33158=>"110101011",
  33159=>"011111110",
  33160=>"000010000",
  33161=>"100010010",
  33162=>"010101000",
  33163=>"110101110",
  33164=>"111001101",
  33165=>"000011000",
  33166=>"010110110",
  33167=>"010111001",
  33168=>"110001000",
  33169=>"011010100",
  33170=>"101000011",
  33171=>"011011011",
  33172=>"100001010",
  33173=>"000000000",
  33174=>"000000011",
  33175=>"100111110",
  33176=>"110001010",
  33177=>"011101010",
  33178=>"011111001",
  33179=>"100001001",
  33180=>"111110011",
  33181=>"010000011",
  33182=>"100111111",
  33183=>"001000010",
  33184=>"110110100",
  33185=>"001111001",
  33186=>"101001001",
  33187=>"101100110",
  33188=>"110010100",
  33189=>"110001001",
  33190=>"100110100",
  33191=>"010001110",
  33192=>"111110000",
  33193=>"000001000",
  33194=>"100000110",
  33195=>"001100100",
  33196=>"100001110",
  33197=>"100001010",
  33198=>"101010110",
  33199=>"100100011",
  33200=>"100000001",
  33201=>"011001001",
  33202=>"000101010",
  33203=>"001010000",
  33204=>"011100101",
  33205=>"010000111",
  33206=>"000010010",
  33207=>"000100100",
  33208=>"111111100",
  33209=>"111111111",
  33210=>"110000111",
  33211=>"101001100",
  33212=>"011111101",
  33213=>"010111110",
  33214=>"000101101",
  33215=>"101111000",
  33216=>"010000010",
  33217=>"011101101",
  33218=>"010110001",
  33219=>"010101001",
  33220=>"011000011",
  33221=>"101001000",
  33222=>"101010101",
  33223=>"001001011",
  33224=>"101111000",
  33225=>"010101110",
  33226=>"000110101",
  33227=>"001001111",
  33228=>"001111001",
  33229=>"001001110",
  33230=>"100111010",
  33231=>"001100011",
  33232=>"000100001",
  33233=>"001110010",
  33234=>"011000011",
  33235=>"111011100",
  33236=>"100111011",
  33237=>"000000010",
  33238=>"101000111",
  33239=>"101101010",
  33240=>"110110101",
  33241=>"111001110",
  33242=>"001100010",
  33243=>"101000010",
  33244=>"101000101",
  33245=>"000100100",
  33246=>"110110100",
  33247=>"001010001",
  33248=>"001100001",
  33249=>"010111001",
  33250=>"101100110",
  33251=>"000101101",
  33252=>"100111010",
  33253=>"101110010",
  33254=>"000010001",
  33255=>"100101001",
  33256=>"100010000",
  33257=>"011110001",
  33258=>"010010001",
  33259=>"101001111",
  33260=>"110101001",
  33261=>"111010111",
  33262=>"010111111",
  33263=>"000000100",
  33264=>"110001010",
  33265=>"001010010",
  33266=>"010001101",
  33267=>"100010111",
  33268=>"010001101",
  33269=>"001100100",
  33270=>"111101110",
  33271=>"101000101",
  33272=>"100000100",
  33273=>"101010101",
  33274=>"100010000",
  33275=>"111001111",
  33276=>"101100011",
  33277=>"110000000",
  33278=>"011100111",
  33279=>"101010010",
  33280=>"010010010",
  33281=>"111100001",
  33282=>"010000000",
  33283=>"101001010",
  33284=>"110011111",
  33285=>"000111111",
  33286=>"010010011",
  33287=>"100000001",
  33288=>"010001110",
  33289=>"001101110",
  33290=>"010101011",
  33291=>"011001101",
  33292=>"100010000",
  33293=>"101011100",
  33294=>"001001101",
  33295=>"100111000",
  33296=>"001110100",
  33297=>"111100000",
  33298=>"011110100",
  33299=>"000110111",
  33300=>"110000110",
  33301=>"001100100",
  33302=>"000011101",
  33303=>"011000111",
  33304=>"001010011",
  33305=>"000000111",
  33306=>"000001110",
  33307=>"010111101",
  33308=>"100011101",
  33309=>"000011010",
  33310=>"001101101",
  33311=>"111111110",
  33312=>"011111010",
  33313=>"100101100",
  33314=>"010010011",
  33315=>"001110010",
  33316=>"111110110",
  33317=>"011001100",
  33318=>"101010001",
  33319=>"110100001",
  33320=>"010100000",
  33321=>"001011111",
  33322=>"111101011",
  33323=>"000000111",
  33324=>"100000111",
  33325=>"000101110",
  33326=>"010001111",
  33327=>"100100001",
  33328=>"110001010",
  33329=>"011011000",
  33330=>"101110000",
  33331=>"001101001",
  33332=>"001010110",
  33333=>"101100111",
  33334=>"110001101",
  33335=>"101000101",
  33336=>"001111010",
  33337=>"001101001",
  33338=>"101010010",
  33339=>"111100011",
  33340=>"011000000",
  33341=>"100100000",
  33342=>"100011100",
  33343=>"110100110",
  33344=>"110111001",
  33345=>"110010010",
  33346=>"011010010",
  33347=>"000011111",
  33348=>"001101101",
  33349=>"000001111",
  33350=>"100111101",
  33351=>"010101111",
  33352=>"111011110",
  33353=>"101010111",
  33354=>"000110110",
  33355=>"011100010",
  33356=>"001000111",
  33357=>"100001111",
  33358=>"111000101",
  33359=>"000010000",
  33360=>"010001111",
  33361=>"111011111",
  33362=>"101010010",
  33363=>"000101100",
  33364=>"001011100",
  33365=>"101000010",
  33366=>"110110110",
  33367=>"110100100",
  33368=>"001111011",
  33369=>"101000110",
  33370=>"101001101",
  33371=>"011001010",
  33372=>"000110000",
  33373=>"010011000",
  33374=>"010000110",
  33375=>"011011111",
  33376=>"001101110",
  33377=>"110000000",
  33378=>"001111001",
  33379=>"111101011",
  33380=>"111010111",
  33381=>"011100111",
  33382=>"101000110",
  33383=>"010011000",
  33384=>"101001000",
  33385=>"110000110",
  33386=>"011111111",
  33387=>"001100011",
  33388=>"010000101",
  33389=>"101000011",
  33390=>"001110100",
  33391=>"111011100",
  33392=>"010111111",
  33393=>"100000100",
  33394=>"110001111",
  33395=>"001111010",
  33396=>"100010010",
  33397=>"100101100",
  33398=>"100111110",
  33399=>"000000101",
  33400=>"100001110",
  33401=>"111001001",
  33402=>"101000000",
  33403=>"011100010",
  33404=>"010000101",
  33405=>"100100011",
  33406=>"001100100",
  33407=>"111011011",
  33408=>"011011011",
  33409=>"000000011",
  33410=>"010001000",
  33411=>"001101100",
  33412=>"000110000",
  33413=>"000011001",
  33414=>"011101010",
  33415=>"111110001",
  33416=>"000010101",
  33417=>"000000100",
  33418=>"110101111",
  33419=>"100101111",
  33420=>"011101000",
  33421=>"000011110",
  33422=>"000000000",
  33423=>"110100010",
  33424=>"111000000",
  33425=>"111100100",
  33426=>"100000110",
  33427=>"010010010",
  33428=>"000000011",
  33429=>"011000011",
  33430=>"110000111",
  33431=>"110111001",
  33432=>"101000011",
  33433=>"101001101",
  33434=>"110001010",
  33435=>"010001101",
  33436=>"010101001",
  33437=>"111111111",
  33438=>"000101010",
  33439=>"001100001",
  33440=>"110000011",
  33441=>"110011010",
  33442=>"011010011",
  33443=>"101010101",
  33444=>"101100000",
  33445=>"111111111",
  33446=>"011101111",
  33447=>"001000111",
  33448=>"001010111",
  33449=>"111010011",
  33450=>"111111010",
  33451=>"110110000",
  33452=>"011000110",
  33453=>"011010100",
  33454=>"101111011",
  33455=>"001110001",
  33456=>"000001000",
  33457=>"110111111",
  33458=>"000001111",
  33459=>"001011101",
  33460=>"000110111",
  33461=>"000111010",
  33462=>"100110101",
  33463=>"001010110",
  33464=>"111101010",
  33465=>"011000001",
  33466=>"010000010",
  33467=>"011011011",
  33468=>"011111010",
  33469=>"000100110",
  33470=>"000001011",
  33471=>"100100111",
  33472=>"001011110",
  33473=>"100110101",
  33474=>"111001101",
  33475=>"101111010",
  33476=>"001100110",
  33477=>"000101000",
  33478=>"001010111",
  33479=>"111001110",
  33480=>"000011101",
  33481=>"111010100",
  33482=>"111101011",
  33483=>"010011000",
  33484=>"001111111",
  33485=>"111101011",
  33486=>"110000101",
  33487=>"110110010",
  33488=>"000011100",
  33489=>"011011001",
  33490=>"111100100",
  33491=>"111111100",
  33492=>"101101100",
  33493=>"100110000",
  33494=>"000101001",
  33495=>"001001000",
  33496=>"111011010",
  33497=>"111101010",
  33498=>"001101011",
  33499=>"000001101",
  33500=>"100100111",
  33501=>"001001001",
  33502=>"101111111",
  33503=>"100101111",
  33504=>"001101010",
  33505=>"110101001",
  33506=>"001000010",
  33507=>"110100011",
  33508=>"010011100",
  33509=>"111000101",
  33510=>"111001011",
  33511=>"100001110",
  33512=>"001101101",
  33513=>"101101000",
  33514=>"000100100",
  33515=>"111010101",
  33516=>"101110110",
  33517=>"000010110",
  33518=>"111000010",
  33519=>"111111111",
  33520=>"110101011",
  33521=>"001100001",
  33522=>"101100000",
  33523=>"011011010",
  33524=>"001110000",
  33525=>"100010101",
  33526=>"000110111",
  33527=>"100100101",
  33528=>"101000011",
  33529=>"101001110",
  33530=>"111001101",
  33531=>"010110101",
  33532=>"100100010",
  33533=>"101110101",
  33534=>"010000001",
  33535=>"111110111",
  33536=>"000010010",
  33537=>"111011101",
  33538=>"001001000",
  33539=>"110000110",
  33540=>"010101000",
  33541=>"111001000",
  33542=>"110010011",
  33543=>"000111100",
  33544=>"111000010",
  33545=>"100111000",
  33546=>"000001011",
  33547=>"010001100",
  33548=>"000110111",
  33549=>"111000100",
  33550=>"110010000",
  33551=>"000110101",
  33552=>"000110010",
  33553=>"001100100",
  33554=>"111001000",
  33555=>"001010111",
  33556=>"111100010",
  33557=>"111011111",
  33558=>"100010000",
  33559=>"111001001",
  33560=>"011001010",
  33561=>"010111110",
  33562=>"100000110",
  33563=>"110011000",
  33564=>"110111000",
  33565=>"100011111",
  33566=>"110011011",
  33567=>"000001100",
  33568=>"001110010",
  33569=>"100011110",
  33570=>"111011001",
  33571=>"010101010",
  33572=>"110110110",
  33573=>"110001000",
  33574=>"110010100",
  33575=>"010110101",
  33576=>"001110000",
  33577=>"111101111",
  33578=>"001101110",
  33579=>"011101111",
  33580=>"001110111",
  33581=>"000011001",
  33582=>"101000011",
  33583=>"001011111",
  33584=>"100000111",
  33585=>"110000101",
  33586=>"000100000",
  33587=>"100101011",
  33588=>"100001100",
  33589=>"001101000",
  33590=>"101001000",
  33591=>"001000011",
  33592=>"010101011",
  33593=>"011110010",
  33594=>"010000001",
  33595=>"010100111",
  33596=>"110000011",
  33597=>"100110111",
  33598=>"010111001",
  33599=>"000111001",
  33600=>"001111000",
  33601=>"001011000",
  33602=>"101110000",
  33603=>"110011010",
  33604=>"111000001",
  33605=>"111101101",
  33606=>"100101011",
  33607=>"110000011",
  33608=>"011100001",
  33609=>"011010010",
  33610=>"011010001",
  33611=>"101000001",
  33612=>"100010001",
  33613=>"001011110",
  33614=>"000110001",
  33615=>"111110110",
  33616=>"110101011",
  33617=>"100001000",
  33618=>"111011000",
  33619=>"001001111",
  33620=>"100100001",
  33621=>"111001011",
  33622=>"100100111",
  33623=>"101010110",
  33624=>"101100111",
  33625=>"011111110",
  33626=>"011000110",
  33627=>"101000100",
  33628=>"001100100",
  33629=>"100111111",
  33630=>"110000110",
  33631=>"100010111",
  33632=>"101011000",
  33633=>"100101000",
  33634=>"100001000",
  33635=>"111011111",
  33636=>"000101111",
  33637=>"101010000",
  33638=>"111111001",
  33639=>"000011111",
  33640=>"011101101",
  33641=>"110001010",
  33642=>"000101000",
  33643=>"101100000",
  33644=>"001001000",
  33645=>"111010001",
  33646=>"000000011",
  33647=>"001101000",
  33648=>"000001000",
  33649=>"010010100",
  33650=>"001111100",
  33651=>"100111110",
  33652=>"100110110",
  33653=>"111010111",
  33654=>"100011110",
  33655=>"010010111",
  33656=>"101101000",
  33657=>"100001001",
  33658=>"110111111",
  33659=>"000001100",
  33660=>"011000000",
  33661=>"111100000",
  33662=>"000101111",
  33663=>"111111001",
  33664=>"010101101",
  33665=>"100001100",
  33666=>"011000000",
  33667=>"011000111",
  33668=>"001101000",
  33669=>"100000100",
  33670=>"000011001",
  33671=>"011100001",
  33672=>"000000100",
  33673=>"001111011",
  33674=>"000001000",
  33675=>"010110001",
  33676=>"000101010",
  33677=>"000100001",
  33678=>"101000110",
  33679=>"110001110",
  33680=>"010110100",
  33681=>"001110111",
  33682=>"110010000",
  33683=>"010001010",
  33684=>"111110111",
  33685=>"101010110",
  33686=>"100000111",
  33687=>"000110110",
  33688=>"101111101",
  33689=>"001101101",
  33690=>"000011100",
  33691=>"110110110",
  33692=>"010111111",
  33693=>"111000111",
  33694=>"000111111",
  33695=>"001010110",
  33696=>"000110111",
  33697=>"001101101",
  33698=>"100101010",
  33699=>"011111000",
  33700=>"110110011",
  33701=>"001000000",
  33702=>"101110100",
  33703=>"000101101",
  33704=>"001110110",
  33705=>"110011010",
  33706=>"000100000",
  33707=>"101100000",
  33708=>"011111001",
  33709=>"000101010",
  33710=>"010111011",
  33711=>"111101101",
  33712=>"110000111",
  33713=>"011010000",
  33714=>"100001000",
  33715=>"010000010",
  33716=>"101010100",
  33717=>"000011000",
  33718=>"110101000",
  33719=>"001010111",
  33720=>"001010100",
  33721=>"111101101",
  33722=>"101101110",
  33723=>"110011001",
  33724=>"111111000",
  33725=>"110000001",
  33726=>"111111111",
  33727=>"100010001",
  33728=>"011011101",
  33729=>"000001000",
  33730=>"000111000",
  33731=>"110010011",
  33732=>"100100101",
  33733=>"100001101",
  33734=>"001000000",
  33735=>"111010100",
  33736=>"000000001",
  33737=>"111010000",
  33738=>"110100111",
  33739=>"110011111",
  33740=>"100101001",
  33741=>"001000001",
  33742=>"011000011",
  33743=>"001111101",
  33744=>"100111001",
  33745=>"101101000",
  33746=>"010000010",
  33747=>"110111100",
  33748=>"010011010",
  33749=>"111111111",
  33750=>"001010110",
  33751=>"010100011",
  33752=>"100000101",
  33753=>"101001101",
  33754=>"010111100",
  33755=>"011110011",
  33756=>"001001111",
  33757=>"000010100",
  33758=>"101101001",
  33759=>"101111100",
  33760=>"000011100",
  33761=>"011001010",
  33762=>"110000111",
  33763=>"100100000",
  33764=>"010011000",
  33765=>"101001101",
  33766=>"000101101",
  33767=>"000001011",
  33768=>"100111000",
  33769=>"100110110",
  33770=>"100011100",
  33771=>"110010100",
  33772=>"110000010",
  33773=>"111100010",
  33774=>"000011001",
  33775=>"110111010",
  33776=>"110111000",
  33777=>"110110101",
  33778=>"110111100",
  33779=>"001011111",
  33780=>"001111110",
  33781=>"111100100",
  33782=>"111111101",
  33783=>"011111101",
  33784=>"000111010",
  33785=>"110000110",
  33786=>"100111001",
  33787=>"110101110",
  33788=>"101010101",
  33789=>"110011000",
  33790=>"011100101",
  33791=>"010011011",
  33792=>"111001100",
  33793=>"110111010",
  33794=>"010110001",
  33795=>"001110101",
  33796=>"000100000",
  33797=>"101100100",
  33798=>"110010000",
  33799=>"101110011",
  33800=>"111101110",
  33801=>"010011101",
  33802=>"010011100",
  33803=>"001111011",
  33804=>"001110110",
  33805=>"100010011",
  33806=>"110011111",
  33807=>"110001001",
  33808=>"110111000",
  33809=>"100110110",
  33810=>"011011111",
  33811=>"011011111",
  33812=>"010101001",
  33813=>"101101110",
  33814=>"101011010",
  33815=>"011110011",
  33816=>"000010011",
  33817=>"110010001",
  33818=>"111000111",
  33819=>"001001000",
  33820=>"001001000",
  33821=>"100101000",
  33822=>"111011010",
  33823=>"110001101",
  33824=>"011000100",
  33825=>"100000011",
  33826=>"111001111",
  33827=>"000010011",
  33828=>"000110000",
  33829=>"111000111",
  33830=>"101011101",
  33831=>"100010001",
  33832=>"011001111",
  33833=>"000111000",
  33834=>"101001001",
  33835=>"010011011",
  33836=>"100011000",
  33837=>"001101010",
  33838=>"111000011",
  33839=>"011010101",
  33840=>"010100011",
  33841=>"110110100",
  33842=>"111111001",
  33843=>"101111101",
  33844=>"000100001",
  33845=>"000101101",
  33846=>"111001011",
  33847=>"101101011",
  33848=>"111000000",
  33849=>"000001000",
  33850=>"110011100",
  33851=>"001001001",
  33852=>"110101001",
  33853=>"000011101",
  33854=>"111001101",
  33855=>"000001110",
  33856=>"100001101",
  33857=>"101010010",
  33858=>"011100110",
  33859=>"110110111",
  33860=>"011101010",
  33861=>"100000011",
  33862=>"010101101",
  33863=>"110011111",
  33864=>"101001010",
  33865=>"010111100",
  33866=>"010110110",
  33867=>"011000100",
  33868=>"001111100",
  33869=>"000100001",
  33870=>"010001010",
  33871=>"110111110",
  33872=>"100010111",
  33873=>"111111100",
  33874=>"100110101",
  33875=>"001100100",
  33876=>"111000010",
  33877=>"100001000",
  33878=>"001110101",
  33879=>"101000110",
  33880=>"011011111",
  33881=>"000010001",
  33882=>"010110111",
  33883=>"110010000",
  33884=>"010001110",
  33885=>"111000010",
  33886=>"100111011",
  33887=>"110000010",
  33888=>"101111001",
  33889=>"101101010",
  33890=>"001101000",
  33891=>"010001001",
  33892=>"111110100",
  33893=>"010011010",
  33894=>"011110101",
  33895=>"000100010",
  33896=>"000011000",
  33897=>"010000111",
  33898=>"000000000",
  33899=>"010111011",
  33900=>"010111100",
  33901=>"101100101",
  33902=>"010011010",
  33903=>"000100110",
  33904=>"100001111",
  33905=>"010010000",
  33906=>"111111110",
  33907=>"111010110",
  33908=>"010010101",
  33909=>"101100100",
  33910=>"111111010",
  33911=>"111111000",
  33912=>"010111111",
  33913=>"000001010",
  33914=>"101111110",
  33915=>"110010011",
  33916=>"000010011",
  33917=>"001011001",
  33918=>"110101101",
  33919=>"110001110",
  33920=>"000100100",
  33921=>"010001011",
  33922=>"010000001",
  33923=>"000010111",
  33924=>"000001100",
  33925=>"011101000",
  33926=>"010101001",
  33927=>"110001100",
  33928=>"111110111",
  33929=>"010010111",
  33930=>"011001111",
  33931=>"111101101",
  33932=>"111000000",
  33933=>"000111110",
  33934=>"011100101",
  33935=>"111011001",
  33936=>"110110010",
  33937=>"100110111",
  33938=>"001000110",
  33939=>"010101101",
  33940=>"000110010",
  33941=>"011000100",
  33942=>"110111011",
  33943=>"110010100",
  33944=>"011111000",
  33945=>"001110100",
  33946=>"110101111",
  33947=>"110000100",
  33948=>"011000111",
  33949=>"010011110",
  33950=>"000000000",
  33951=>"101110111",
  33952=>"100100111",
  33953=>"100000100",
  33954=>"101111111",
  33955=>"110000010",
  33956=>"010010001",
  33957=>"000010010",
  33958=>"110010011",
  33959=>"101100101",
  33960=>"011011000",
  33961=>"101011100",
  33962=>"110100011",
  33963=>"111011000",
  33964=>"110100010",
  33965=>"000101111",
  33966=>"101100000",
  33967=>"011000111",
  33968=>"100010101",
  33969=>"000000000",
  33970=>"100001111",
  33971=>"001100001",
  33972=>"011000101",
  33973=>"100000000",
  33974=>"010100110",
  33975=>"001110110",
  33976=>"011111001",
  33977=>"010011111",
  33978=>"011111000",
  33979=>"101000100",
  33980=>"100100101",
  33981=>"101100011",
  33982=>"010001001",
  33983=>"100111011",
  33984=>"001001100",
  33985=>"101100110",
  33986=>"111101110",
  33987=>"011000101",
  33988=>"100110000",
  33989=>"111011111",
  33990=>"010000000",
  33991=>"001101000",
  33992=>"011101011",
  33993=>"101010000",
  33994=>"111011111",
  33995=>"011010101",
  33996=>"111011001",
  33997=>"011110010",
  33998=>"001110110",
  33999=>"011111111",
  34000=>"101000001",
  34001=>"010011111",
  34002=>"001101000",
  34003=>"010001000",
  34004=>"101100001",
  34005=>"110100000",
  34006=>"110110010",
  34007=>"101011111",
  34008=>"111111001",
  34009=>"101111010",
  34010=>"010111011",
  34011=>"100011100",
  34012=>"011000000",
  34013=>"111001000",
  34014=>"000000100",
  34015=>"000010001",
  34016=>"001101100",
  34017=>"111111001",
  34018=>"001010100",
  34019=>"110000001",
  34020=>"111100000",
  34021=>"111111001",
  34022=>"110110101",
  34023=>"001101000",
  34024=>"101000011",
  34025=>"000011001",
  34026=>"000001000",
  34027=>"010100010",
  34028=>"010011010",
  34029=>"001100000",
  34030=>"000010001",
  34031=>"110110000",
  34032=>"000110111",
  34033=>"101010000",
  34034=>"000001100",
  34035=>"001010110",
  34036=>"001110111",
  34037=>"011000010",
  34038=>"000101010",
  34039=>"101100111",
  34040=>"101010011",
  34041=>"000101000",
  34042=>"111100100",
  34043=>"110111100",
  34044=>"100000100",
  34045=>"001110010",
  34046=>"111110001",
  34047=>"010110111",
  34048=>"100010001",
  34049=>"010000101",
  34050=>"100110101",
  34051=>"010010000",
  34052=>"110011001",
  34053=>"011010011",
  34054=>"100000110",
  34055=>"000011011",
  34056=>"101010010",
  34057=>"101101110",
  34058=>"101111011",
  34059=>"111011111",
  34060=>"000110111",
  34061=>"000001000",
  34062=>"110011111",
  34063=>"000100101",
  34064=>"111001101",
  34065=>"110000010",
  34066=>"010100101",
  34067=>"000000011",
  34068=>"000000010",
  34069=>"100001100",
  34070=>"101001101",
  34071=>"110000001",
  34072=>"111001001",
  34073=>"001001000",
  34074=>"110100000",
  34075=>"000101000",
  34076=>"110111001",
  34077=>"011110101",
  34078=>"101110001",
  34079=>"110111001",
  34080=>"000001110",
  34081=>"100011111",
  34082=>"010011000",
  34083=>"000000110",
  34084=>"001101111",
  34085=>"000010001",
  34086=>"000010100",
  34087=>"110000101",
  34088=>"010101000",
  34089=>"001100111",
  34090=>"010111110",
  34091=>"000001101",
  34092=>"110010111",
  34093=>"011010010",
  34094=>"001000011",
  34095=>"010001011",
  34096=>"100010010",
  34097=>"111100001",
  34098=>"111011010",
  34099=>"001110000",
  34100=>"111001111",
  34101=>"000001001",
  34102=>"100111100",
  34103=>"011010010",
  34104=>"110000011",
  34105=>"000011010",
  34106=>"111011000",
  34107=>"110010010",
  34108=>"001000000",
  34109=>"101110100",
  34110=>"010111011",
  34111=>"101111110",
  34112=>"110100000",
  34113=>"001000100",
  34114=>"110101001",
  34115=>"111000101",
  34116=>"010110101",
  34117=>"100111100",
  34118=>"000000111",
  34119=>"001111101",
  34120=>"011001001",
  34121=>"101100000",
  34122=>"001100111",
  34123=>"001000001",
  34124=>"110000010",
  34125=>"101011011",
  34126=>"001100110",
  34127=>"010010100",
  34128=>"011100001",
  34129=>"000110011",
  34130=>"010100001",
  34131=>"010000111",
  34132=>"000001001",
  34133=>"100010110",
  34134=>"100110100",
  34135=>"010010111",
  34136=>"001011011",
  34137=>"001100011",
  34138=>"010000001",
  34139=>"000001100",
  34140=>"110101100",
  34141=>"100101011",
  34142=>"010000111",
  34143=>"010100100",
  34144=>"111111101",
  34145=>"111110111",
  34146=>"110111110",
  34147=>"100011110",
  34148=>"000001111",
  34149=>"000000011",
  34150=>"000100100",
  34151=>"101010101",
  34152=>"110000100",
  34153=>"100111101",
  34154=>"001100100",
  34155=>"001111101",
  34156=>"110010101",
  34157=>"000110101",
  34158=>"111111111",
  34159=>"101000100",
  34160=>"011001010",
  34161=>"111011011",
  34162=>"010100110",
  34163=>"011011011",
  34164=>"100000010",
  34165=>"010011010",
  34166=>"000100010",
  34167=>"111011100",
  34168=>"000011111",
  34169=>"101111000",
  34170=>"110110101",
  34171=>"101000001",
  34172=>"001000101",
  34173=>"100110011",
  34174=>"010100111",
  34175=>"111111101",
  34176=>"001000101",
  34177=>"100101101",
  34178=>"010010110",
  34179=>"000011000",
  34180=>"000011110",
  34181=>"010000100",
  34182=>"111101101",
  34183=>"111001101",
  34184=>"011000100",
  34185=>"111110000",
  34186=>"001010111",
  34187=>"101111011",
  34188=>"011101101",
  34189=>"011011011",
  34190=>"111010001",
  34191=>"101010100",
  34192=>"001100111",
  34193=>"111101111",
  34194=>"001000011",
  34195=>"010100001",
  34196=>"010000000",
  34197=>"101010100",
  34198=>"001011101",
  34199=>"101011110",
  34200=>"000111101",
  34201=>"000101001",
  34202=>"110000010",
  34203=>"010000110",
  34204=>"011101001",
  34205=>"010111110",
  34206=>"000100110",
  34207=>"001001111",
  34208=>"110011000",
  34209=>"100000010",
  34210=>"011011000",
  34211=>"111001000",
  34212=>"111101111",
  34213=>"011000010",
  34214=>"011010001",
  34215=>"011000101",
  34216=>"000000010",
  34217=>"101011101",
  34218=>"110010000",
  34219=>"101111100",
  34220=>"001000011",
  34221=>"000001000",
  34222=>"011101010",
  34223=>"111111100",
  34224=>"101111110",
  34225=>"010111010",
  34226=>"111000100",
  34227=>"110111000",
  34228=>"011001000",
  34229=>"010011011",
  34230=>"111111000",
  34231=>"111010001",
  34232=>"111001001",
  34233=>"011101000",
  34234=>"010010110",
  34235=>"010101100",
  34236=>"111010111",
  34237=>"100101010",
  34238=>"001001101",
  34239=>"110110010",
  34240=>"111001011",
  34241=>"000000011",
  34242=>"101101010",
  34243=>"000011010",
  34244=>"000100000",
  34245=>"100001000",
  34246=>"111110101",
  34247=>"100001000",
  34248=>"011101010",
  34249=>"011011001",
  34250=>"001100000",
  34251=>"001000100",
  34252=>"100010111",
  34253=>"111010000",
  34254=>"011111000",
  34255=>"001110011",
  34256=>"010101111",
  34257=>"010001011",
  34258=>"101001101",
  34259=>"000110000",
  34260=>"000100110",
  34261=>"110110001",
  34262=>"000000011",
  34263=>"100000111",
  34264=>"010111000",
  34265=>"011011111",
  34266=>"101101111",
  34267=>"101001010",
  34268=>"001111011",
  34269=>"110101010",
  34270=>"101110110",
  34271=>"000010101",
  34272=>"111010100",
  34273=>"000101010",
  34274=>"101101110",
  34275=>"101110000",
  34276=>"110101101",
  34277=>"010011111",
  34278=>"100101010",
  34279=>"100110001",
  34280=>"101011110",
  34281=>"000011011",
  34282=>"001011110",
  34283=>"011000111",
  34284=>"100010100",
  34285=>"000010010",
  34286=>"010001000",
  34287=>"001010010",
  34288=>"100011100",
  34289=>"100000010",
  34290=>"011111000",
  34291=>"110100110",
  34292=>"000101111",
  34293=>"010000000",
  34294=>"010101100",
  34295=>"100010100",
  34296=>"101101111",
  34297=>"100010001",
  34298=>"001110001",
  34299=>"010100001",
  34300=>"101001000",
  34301=>"001011011",
  34302=>"011101001",
  34303=>"110001111",
  34304=>"001100010",
  34305=>"011101100",
  34306=>"000010010",
  34307=>"010110111",
  34308=>"010010010",
  34309=>"000010110",
  34310=>"100011111",
  34311=>"100001111",
  34312=>"001001001",
  34313=>"101010001",
  34314=>"110000110",
  34315=>"110010110",
  34316=>"101001001",
  34317=>"000101110",
  34318=>"101010000",
  34319=>"011110100",
  34320=>"000011001",
  34321=>"001001011",
  34322=>"110100000",
  34323=>"110101000",
  34324=>"000110101",
  34325=>"100000111",
  34326=>"100101000",
  34327=>"111110011",
  34328=>"111100100",
  34329=>"000101100",
  34330=>"101000110",
  34331=>"101110100",
  34332=>"101001000",
  34333=>"100100000",
  34334=>"110110110",
  34335=>"101001000",
  34336=>"100100010",
  34337=>"000110110",
  34338=>"111011101",
  34339=>"000011111",
  34340=>"111110000",
  34341=>"001000001",
  34342=>"110101111",
  34343=>"100111110",
  34344=>"111101110",
  34345=>"010010010",
  34346=>"000100000",
  34347=>"111000101",
  34348=>"101100000",
  34349=>"010001000",
  34350=>"110101000",
  34351=>"010010100",
  34352=>"111011001",
  34353=>"010001001",
  34354=>"101111011",
  34355=>"010001100",
  34356=>"111111111",
  34357=>"010011111",
  34358=>"000100000",
  34359=>"101010011",
  34360=>"000000101",
  34361=>"010000100",
  34362=>"101000110",
  34363=>"111000100",
  34364=>"100000111",
  34365=>"101100011",
  34366=>"000101011",
  34367=>"100000111",
  34368=>"001110111",
  34369=>"001110110",
  34370=>"100100011",
  34371=>"100101101",
  34372=>"100000100",
  34373=>"100011110",
  34374=>"110011101",
  34375=>"000110100",
  34376=>"010001011",
  34377=>"000001100",
  34378=>"101110101",
  34379=>"000101010",
  34380=>"001010000",
  34381=>"000110010",
  34382=>"001011010",
  34383=>"010011011",
  34384=>"010011111",
  34385=>"010110011",
  34386=>"001001100",
  34387=>"101001101",
  34388=>"000111001",
  34389=>"111111001",
  34390=>"111111110",
  34391=>"111010011",
  34392=>"000110000",
  34393=>"111000001",
  34394=>"001010101",
  34395=>"000010110",
  34396=>"100100010",
  34397=>"101000010",
  34398=>"000101011",
  34399=>"111101000",
  34400=>"111110010",
  34401=>"101011110",
  34402=>"000001010",
  34403=>"101110011",
  34404=>"001111000",
  34405=>"111110110",
  34406=>"100101011",
  34407=>"110001000",
  34408=>"101100100",
  34409=>"100011001",
  34410=>"011111001",
  34411=>"101010111",
  34412=>"011001000",
  34413=>"110110011",
  34414=>"111101101",
  34415=>"011011010",
  34416=>"110010001",
  34417=>"011010110",
  34418=>"101010111",
  34419=>"110110011",
  34420=>"000010101",
  34421=>"000011000",
  34422=>"000110111",
  34423=>"010110010",
  34424=>"011111101",
  34425=>"100100100",
  34426=>"111101100",
  34427=>"000101000",
  34428=>"001101110",
  34429=>"000000011",
  34430=>"111101011",
  34431=>"110011111",
  34432=>"111010000",
  34433=>"111111111",
  34434=>"000001001",
  34435=>"000011000",
  34436=>"101101100",
  34437=>"000001001",
  34438=>"110101101",
  34439=>"111101101",
  34440=>"000001100",
  34441=>"111111101",
  34442=>"011100001",
  34443=>"001011100",
  34444=>"001101110",
  34445=>"011001011",
  34446=>"110110100",
  34447=>"100111101",
  34448=>"100010100",
  34449=>"010001011",
  34450=>"100110011",
  34451=>"110001000",
  34452=>"001101100",
  34453=>"110110100",
  34454=>"010001000",
  34455=>"111011100",
  34456=>"111110101",
  34457=>"000001000",
  34458=>"011111110",
  34459=>"101111010",
  34460=>"000000111",
  34461=>"000111010",
  34462=>"001000101",
  34463=>"000010000",
  34464=>"110100110",
  34465=>"110011011",
  34466=>"011010100",
  34467=>"110010100",
  34468=>"000101110",
  34469=>"010000110",
  34470=>"110111000",
  34471=>"011000011",
  34472=>"010100101",
  34473=>"000010011",
  34474=>"010110100",
  34475=>"110001001",
  34476=>"001101001",
  34477=>"000101000",
  34478=>"001001010",
  34479=>"100100001",
  34480=>"101010011",
  34481=>"011110000",
  34482=>"111100101",
  34483=>"000000011",
  34484=>"000000010",
  34485=>"100101100",
  34486=>"010001100",
  34487=>"110000000",
  34488=>"011000000",
  34489=>"000010111",
  34490=>"111001011",
  34491=>"010011000",
  34492=>"010101011",
  34493=>"110001101",
  34494=>"101100010",
  34495=>"010100011",
  34496=>"000110100",
  34497=>"101100000",
  34498=>"010010000",
  34499=>"001000011",
  34500=>"110111100",
  34501=>"000010001",
  34502=>"000110111",
  34503=>"100010101",
  34504=>"111110111",
  34505=>"010100111",
  34506=>"001101110",
  34507=>"101111100",
  34508=>"001001000",
  34509=>"001000100",
  34510=>"100010110",
  34511=>"111010011",
  34512=>"111100111",
  34513=>"010000110",
  34514=>"001100000",
  34515=>"100000110",
  34516=>"010011000",
  34517=>"111110111",
  34518=>"101011010",
  34519=>"010111000",
  34520=>"110010000",
  34521=>"001101000",
  34522=>"010000000",
  34523=>"001001100",
  34524=>"000111010",
  34525=>"001111011",
  34526=>"101000100",
  34527=>"110000110",
  34528=>"101111111",
  34529=>"000001000",
  34530=>"000000101",
  34531=>"110100100",
  34532=>"111101010",
  34533=>"100011010",
  34534=>"010100111",
  34535=>"000110111",
  34536=>"100010000",
  34537=>"100111011",
  34538=>"110111101",
  34539=>"101101001",
  34540=>"000001101",
  34541=>"000011011",
  34542=>"101010110",
  34543=>"010110000",
  34544=>"011101111",
  34545=>"100100101",
  34546=>"100000111",
  34547=>"010011111",
  34548=>"111010100",
  34549=>"111101001",
  34550=>"111011010",
  34551=>"010101010",
  34552=>"010111000",
  34553=>"100110001",
  34554=>"100010000",
  34555=>"001001000",
  34556=>"001000010",
  34557=>"100000010",
  34558=>"000001010",
  34559=>"000000011",
  34560=>"001010111",
  34561=>"011101111",
  34562=>"100101111",
  34563=>"010001111",
  34564=>"100001110",
  34565=>"011001111",
  34566=>"010000101",
  34567=>"001001010",
  34568=>"000011100",
  34569=>"100101010",
  34570=>"101011110",
  34571=>"111100100",
  34572=>"101101010",
  34573=>"001010101",
  34574=>"101011101",
  34575=>"000010111",
  34576=>"111111101",
  34577=>"101100000",
  34578=>"011100101",
  34579=>"101001101",
  34580=>"000000000",
  34581=>"000110100",
  34582=>"001011000",
  34583=>"000000001",
  34584=>"000100010",
  34585=>"100110100",
  34586=>"000110010",
  34587=>"001101000",
  34588=>"100111111",
  34589=>"000101011",
  34590=>"010001010",
  34591=>"110001010",
  34592=>"110001001",
  34593=>"001100110",
  34594=>"010110111",
  34595=>"110111000",
  34596=>"111001101",
  34597=>"000010000",
  34598=>"101011111",
  34599=>"111111001",
  34600=>"101111000",
  34601=>"011000011",
  34602=>"111001001",
  34603=>"101100111",
  34604=>"110000011",
  34605=>"000000011",
  34606=>"101110111",
  34607=>"101001000",
  34608=>"000100101",
  34609=>"100000000",
  34610=>"010100000",
  34611=>"001100001",
  34612=>"001110001",
  34613=>"100001010",
  34614=>"111101101",
  34615=>"111100011",
  34616=>"101100100",
  34617=>"010101010",
  34618=>"111011000",
  34619=>"100011101",
  34620=>"000011000",
  34621=>"001000010",
  34622=>"101010001",
  34623=>"011101100",
  34624=>"110011101",
  34625=>"011101000",
  34626=>"111110011",
  34627=>"111101111",
  34628=>"100111010",
  34629=>"001110000",
  34630=>"100010011",
  34631=>"010101110",
  34632=>"100100000",
  34633=>"101000000",
  34634=>"111100011",
  34635=>"110011100",
  34636=>"010000010",
  34637=>"011001001",
  34638=>"100000111",
  34639=>"100000001",
  34640=>"000010100",
  34641=>"001101011",
  34642=>"000011000",
  34643=>"100101100",
  34644=>"100001110",
  34645=>"111101001",
  34646=>"001010100",
  34647=>"001111001",
  34648=>"011001100",
  34649=>"001000110",
  34650=>"010101000",
  34651=>"001011111",
  34652=>"111100101",
  34653=>"100101001",
  34654=>"100010111",
  34655=>"001000000",
  34656=>"011111111",
  34657=>"010011000",
  34658=>"101100000",
  34659=>"100010101",
  34660=>"100000110",
  34661=>"100000001",
  34662=>"010111010",
  34663=>"110110001",
  34664=>"001110101",
  34665=>"101101110",
  34666=>"000000110",
  34667=>"111100000",
  34668=>"111010010",
  34669=>"100000110",
  34670=>"100010011",
  34671=>"100010101",
  34672=>"010010001",
  34673=>"110000110",
  34674=>"101011001",
  34675=>"000001001",
  34676=>"111101110",
  34677=>"101011111",
  34678=>"111111111",
  34679=>"100000011",
  34680=>"110110010",
  34681=>"011100011",
  34682=>"010101011",
  34683=>"111010000",
  34684=>"011010000",
  34685=>"111011110",
  34686=>"011001010",
  34687=>"011100010",
  34688=>"100111101",
  34689=>"110101100",
  34690=>"111111111",
  34691=>"110110000",
  34692=>"000110111",
  34693=>"100111001",
  34694=>"011001001",
  34695=>"000000110",
  34696=>"011110101",
  34697=>"011111101",
  34698=>"111111100",
  34699=>"100010011",
  34700=>"001100100",
  34701=>"011010100",
  34702=>"101000101",
  34703=>"000101101",
  34704=>"101111111",
  34705=>"110010010",
  34706=>"000011011",
  34707=>"000000101",
  34708=>"110000011",
  34709=>"001101100",
  34710=>"010001001",
  34711=>"101110000",
  34712=>"111010101",
  34713=>"100000010",
  34714=>"100010110",
  34715=>"010111001",
  34716=>"110010111",
  34717=>"001111001",
  34718=>"110101011",
  34719=>"111101100",
  34720=>"010100011",
  34721=>"111111101",
  34722=>"000100111",
  34723=>"111111110",
  34724=>"110111001",
  34725=>"001010110",
  34726=>"010011111",
  34727=>"111011000",
  34728=>"010101001",
  34729=>"110111111",
  34730=>"101101001",
  34731=>"000001110",
  34732=>"100000110",
  34733=>"011011101",
  34734=>"011010011",
  34735=>"011111111",
  34736=>"111000000",
  34737=>"001001001",
  34738=>"011100001",
  34739=>"110111011",
  34740=>"100010110",
  34741=>"001110000",
  34742=>"011111000",
  34743=>"010001011",
  34744=>"111101100",
  34745=>"011111010",
  34746=>"101000010",
  34747=>"001011110",
  34748=>"101101011",
  34749=>"000011100",
  34750=>"001000001",
  34751=>"111100011",
  34752=>"101100000",
  34753=>"101110101",
  34754=>"001000100",
  34755=>"000101011",
  34756=>"110011010",
  34757=>"000111011",
  34758=>"111010000",
  34759=>"110010101",
  34760=>"001111000",
  34761=>"110100000",
  34762=>"110010011",
  34763=>"001010111",
  34764=>"111111100",
  34765=>"111100100",
  34766=>"110101111",
  34767=>"111001000",
  34768=>"000010101",
  34769=>"001101111",
  34770=>"010110110",
  34771=>"101101001",
  34772=>"001010010",
  34773=>"000011010",
  34774=>"001111000",
  34775=>"111001111",
  34776=>"010000000",
  34777=>"101010101",
  34778=>"110101000",
  34779=>"001000111",
  34780=>"111110100",
  34781=>"111111101",
  34782=>"100111000",
  34783=>"101011001",
  34784=>"100111111",
  34785=>"001010010",
  34786=>"000100111",
  34787=>"000010010",
  34788=>"100001111",
  34789=>"000010001",
  34790=>"001011101",
  34791=>"100111010",
  34792=>"001110000",
  34793=>"111101100",
  34794=>"101001100",
  34795=>"011111110",
  34796=>"101101101",
  34797=>"011100110",
  34798=>"100010000",
  34799=>"111000100",
  34800=>"001110100",
  34801=>"100001110",
  34802=>"101010011",
  34803=>"110000100",
  34804=>"111011010",
  34805=>"000010000",
  34806=>"000011000",
  34807=>"110111010",
  34808=>"001100110",
  34809=>"111101100",
  34810=>"101100000",
  34811=>"010100111",
  34812=>"110010100",
  34813=>"100001110",
  34814=>"001110100",
  34815=>"000101000",
  34816=>"101100000",
  34817=>"000110010",
  34818=>"101001111",
  34819=>"101001101",
  34820=>"100001011",
  34821=>"000010100",
  34822=>"000110111",
  34823=>"101100111",
  34824=>"110001010",
  34825=>"111001001",
  34826=>"111000110",
  34827=>"011001110",
  34828=>"001101001",
  34829=>"001000000",
  34830=>"100001110",
  34831=>"100110100",
  34832=>"101110010",
  34833=>"100100101",
  34834=>"100001010",
  34835=>"111101110",
  34836=>"101100010",
  34837=>"110010011",
  34838=>"110100001",
  34839=>"000001000",
  34840=>"001000000",
  34841=>"000110010",
  34842=>"101000110",
  34843=>"111001001",
  34844=>"100010110",
  34845=>"001010110",
  34846=>"001100011",
  34847=>"011110101",
  34848=>"111011100",
  34849=>"100001001",
  34850=>"101011000",
  34851=>"010010110",
  34852=>"011101010",
  34853=>"100110111",
  34854=>"000100100",
  34855=>"011010100",
  34856=>"001101001",
  34857=>"111001110",
  34858=>"010010001",
  34859=>"011100101",
  34860=>"011001100",
  34861=>"001000110",
  34862=>"010100111",
  34863=>"100010011",
  34864=>"011001110",
  34865=>"011111010",
  34866=>"000000110",
  34867=>"000101000",
  34868=>"101110000",
  34869=>"011100000",
  34870=>"100000000",
  34871=>"001011101",
  34872=>"000101011",
  34873=>"100000001",
  34874=>"001110011",
  34875=>"000100110",
  34876=>"100010111",
  34877=>"101100111",
  34878=>"100100000",
  34879=>"001100110",
  34880=>"000100100",
  34881=>"110010001",
  34882=>"111101110",
  34883=>"110000011",
  34884=>"001011101",
  34885=>"010100100",
  34886=>"100100000",
  34887=>"100000000",
  34888=>"010100011",
  34889=>"111100111",
  34890=>"000101100",
  34891=>"010010110",
  34892=>"110001000",
  34893=>"000111000",
  34894=>"101001101",
  34895=>"110010011",
  34896=>"001110001",
  34897=>"000000110",
  34898=>"101011100",
  34899=>"110010000",
  34900=>"001101010",
  34901=>"111111011",
  34902=>"101010010",
  34903=>"101100001",
  34904=>"011111011",
  34905=>"111111011",
  34906=>"011100001",
  34907=>"110111011",
  34908=>"100110001",
  34909=>"101101100",
  34910=>"101010101",
  34911=>"001101011",
  34912=>"001010100",
  34913=>"100110010",
  34914=>"100111111",
  34915=>"011001001",
  34916=>"100000010",
  34917=>"011010001",
  34918=>"011100111",
  34919=>"111010010",
  34920=>"100001100",
  34921=>"001100010",
  34922=>"011001100",
  34923=>"011000101",
  34924=>"001101101",
  34925=>"101000000",
  34926=>"100000011",
  34927=>"111110001",
  34928=>"101000100",
  34929=>"001000100",
  34930=>"100001000",
  34931=>"111001001",
  34932=>"101000011",
  34933=>"010101111",
  34934=>"000011101",
  34935=>"010100011",
  34936=>"101111100",
  34937=>"101100101",
  34938=>"110101110",
  34939=>"100000111",
  34940=>"100100101",
  34941=>"101111101",
  34942=>"011001000",
  34943=>"011111010",
  34944=>"000000010",
  34945=>"111100011",
  34946=>"001011000",
  34947=>"101100100",
  34948=>"110110110",
  34949=>"000101010",
  34950=>"001011011",
  34951=>"000111000",
  34952=>"001000000",
  34953=>"010001010",
  34954=>"111000000",
  34955=>"100011001",
  34956=>"000100010",
  34957=>"101111110",
  34958=>"110111000",
  34959=>"100111011",
  34960=>"010000001",
  34961=>"111111011",
  34962=>"111010010",
  34963=>"011101000",
  34964=>"001000001",
  34965=>"101010000",
  34966=>"100011100",
  34967=>"110110000",
  34968=>"000011111",
  34969=>"011000110",
  34970=>"111100000",
  34971=>"000111001",
  34972=>"000100110",
  34973=>"010001111",
  34974=>"101110000",
  34975=>"011011010",
  34976=>"011111011",
  34977=>"111100101",
  34978=>"110011101",
  34979=>"011010010",
  34980=>"100111110",
  34981=>"001000000",
  34982=>"011000100",
  34983=>"010100100",
  34984=>"111001010",
  34985=>"110011101",
  34986=>"001001000",
  34987=>"110110000",
  34988=>"000111010",
  34989=>"110110101",
  34990=>"101101000",
  34991=>"011101111",
  34992=>"001100111",
  34993=>"010101101",
  34994=>"001110000",
  34995=>"111110001",
  34996=>"000000001",
  34997=>"111100011",
  34998=>"110011011",
  34999=>"111000101",
  35000=>"010101111",
  35001=>"101100101",
  35002=>"101011001",
  35003=>"010111100",
  35004=>"100101001",
  35005=>"111010010",
  35006=>"000101000",
  35007=>"001001101",
  35008=>"010100011",
  35009=>"101100101",
  35010=>"100010011",
  35011=>"011111001",
  35012=>"111111100",
  35013=>"100001000",
  35014=>"100000000",
  35015=>"101001010",
  35016=>"001000100",
  35017=>"110001111",
  35018=>"110011110",
  35019=>"111110100",
  35020=>"111100111",
  35021=>"000010101",
  35022=>"001011001",
  35023=>"011101100",
  35024=>"001101111",
  35025=>"101101010",
  35026=>"110100001",
  35027=>"011011110",
  35028=>"000001111",
  35029=>"101101011",
  35030=>"001001001",
  35031=>"010101100",
  35032=>"001101101",
  35033=>"101111100",
  35034=>"000010101",
  35035=>"101100001",
  35036=>"011011101",
  35037=>"100100010",
  35038=>"000101111",
  35039=>"100111011",
  35040=>"000101101",
  35041=>"101111111",
  35042=>"101101110",
  35043=>"110100110",
  35044=>"110100011",
  35045=>"110110100",
  35046=>"000111110",
  35047=>"101100110",
  35048=>"010111111",
  35049=>"001110110",
  35050=>"011101100",
  35051=>"001101101",
  35052=>"110001010",
  35053=>"110101110",
  35054=>"100100101",
  35055=>"101101001",
  35056=>"011110000",
  35057=>"100001101",
  35058=>"110111111",
  35059=>"011110010",
  35060=>"111110011",
  35061=>"101100110",
  35062=>"000000001",
  35063=>"110000001",
  35064=>"001111010",
  35065=>"101000100",
  35066=>"100101010",
  35067=>"110000100",
  35068=>"111001000",
  35069=>"001011100",
  35070=>"111011100",
  35071=>"110011110",
  35072=>"111000000",
  35073=>"001010000",
  35074=>"110110010",
  35075=>"100001101",
  35076=>"011111000",
  35077=>"001000100",
  35078=>"000001001",
  35079=>"111001100",
  35080=>"011101010",
  35081=>"000011000",
  35082=>"011011001",
  35083=>"111100011",
  35084=>"000000010",
  35085=>"000001101",
  35086=>"001001010",
  35087=>"110010111",
  35088=>"101111000",
  35089=>"011110100",
  35090=>"000010000",
  35091=>"011110001",
  35092=>"001001001",
  35093=>"011100100",
  35094=>"010000110",
  35095=>"000101101",
  35096=>"111111000",
  35097=>"111101001",
  35098=>"000100001",
  35099=>"001100100",
  35100=>"110000100",
  35101=>"011100110",
  35102=>"101000100",
  35103=>"101100001",
  35104=>"110111110",
  35105=>"001010000",
  35106=>"011011010",
  35107=>"010011111",
  35108=>"100110110",
  35109=>"110000111",
  35110=>"111101010",
  35111=>"001111001",
  35112=>"101111001",
  35113=>"001000100",
  35114=>"100100100",
  35115=>"011001100",
  35116=>"001001111",
  35117=>"011110000",
  35118=>"001100111",
  35119=>"011101010",
  35120=>"000000111",
  35121=>"100000001",
  35122=>"010111010",
  35123=>"001101100",
  35124=>"000101100",
  35125=>"010111011",
  35126=>"001001110",
  35127=>"111011111",
  35128=>"000000110",
  35129=>"101100011",
  35130=>"010000100",
  35131=>"001011101",
  35132=>"000000101",
  35133=>"000111111",
  35134=>"000011000",
  35135=>"011100110",
  35136=>"000001010",
  35137=>"111101010",
  35138=>"001101010",
  35139=>"011110101",
  35140=>"000101101",
  35141=>"010010010",
  35142=>"011000011",
  35143=>"011101010",
  35144=>"011010000",
  35145=>"101000101",
  35146=>"111011101",
  35147=>"000100001",
  35148=>"111100100",
  35149=>"001010001",
  35150=>"010001101",
  35151=>"010011010",
  35152=>"000011001",
  35153=>"001011100",
  35154=>"000100001",
  35155=>"100110010",
  35156=>"010101100",
  35157=>"010000101",
  35158=>"100110111",
  35159=>"011001010",
  35160=>"100100010",
  35161=>"100001010",
  35162=>"100100100",
  35163=>"010100001",
  35164=>"111111111",
  35165=>"111101000",
  35166=>"011001010",
  35167=>"110100001",
  35168=>"010101110",
  35169=>"110000010",
  35170=>"000001100",
  35171=>"100000100",
  35172=>"101111000",
  35173=>"010011110",
  35174=>"101101010",
  35175=>"011000001",
  35176=>"001111100",
  35177=>"100101101",
  35178=>"011011000",
  35179=>"001101101",
  35180=>"000110111",
  35181=>"101001100",
  35182=>"100101000",
  35183=>"111101101",
  35184=>"110000010",
  35185=>"101110011",
  35186=>"011111000",
  35187=>"010010001",
  35188=>"000101111",
  35189=>"100111000",
  35190=>"011011010",
  35191=>"100011110",
  35192=>"010101010",
  35193=>"100001101",
  35194=>"011110101",
  35195=>"110101001",
  35196=>"100011111",
  35197=>"110110101",
  35198=>"001010011",
  35199=>"111001111",
  35200=>"101001001",
  35201=>"001111111",
  35202=>"100011100",
  35203=>"011101000",
  35204=>"011110100",
  35205=>"110010111",
  35206=>"111111110",
  35207=>"000101010",
  35208=>"101111110",
  35209=>"011000100",
  35210=>"110100000",
  35211=>"010101111",
  35212=>"101101100",
  35213=>"000000101",
  35214=>"111111101",
  35215=>"110111010",
  35216=>"011010100",
  35217=>"101100110",
  35218=>"011011011",
  35219=>"000000101",
  35220=>"100000000",
  35221=>"010110111",
  35222=>"000000101",
  35223=>"100101100",
  35224=>"000011111",
  35225=>"101001100",
  35226=>"001001100",
  35227=>"011000110",
  35228=>"111000110",
  35229=>"100101000",
  35230=>"000010110",
  35231=>"110110000",
  35232=>"101110001",
  35233=>"000011101",
  35234=>"011110011",
  35235=>"000000000",
  35236=>"111011101",
  35237=>"001111101",
  35238=>"100001111",
  35239=>"101111100",
  35240=>"010011111",
  35241=>"001011010",
  35242=>"101110101",
  35243=>"000100010",
  35244=>"010101000",
  35245=>"000001101",
  35246=>"000111100",
  35247=>"101100110",
  35248=>"001100000",
  35249=>"111001100",
  35250=>"000111011",
  35251=>"111010011",
  35252=>"011110111",
  35253=>"100011011",
  35254=>"010111101",
  35255=>"101001000",
  35256=>"011011010",
  35257=>"001100000",
  35258=>"000000010",
  35259=>"011001000",
  35260=>"111101101",
  35261=>"001011010",
  35262=>"100110010",
  35263=>"101011111",
  35264=>"100101111",
  35265=>"000100100",
  35266=>"111000000",
  35267=>"111101110",
  35268=>"001001101",
  35269=>"010010100",
  35270=>"100110111",
  35271=>"001001000",
  35272=>"101111001",
  35273=>"011101101",
  35274=>"011111001",
  35275=>"000101000",
  35276=>"001110001",
  35277=>"000101000",
  35278=>"101110001",
  35279=>"110010100",
  35280=>"110110101",
  35281=>"001000001",
  35282=>"100011001",
  35283=>"100101011",
  35284=>"101001011",
  35285=>"010000010",
  35286=>"010100101",
  35287=>"111011100",
  35288=>"001001110",
  35289=>"101001010",
  35290=>"111110000",
  35291=>"111101110",
  35292=>"101101101",
  35293=>"111010100",
  35294=>"000000101",
  35295=>"001110011",
  35296=>"001001001",
  35297=>"001010110",
  35298=>"011101010",
  35299=>"101000010",
  35300=>"110111001",
  35301=>"001000101",
  35302=>"110000110",
  35303=>"010000000",
  35304=>"011000000",
  35305=>"011001100",
  35306=>"101100110",
  35307=>"000101000",
  35308=>"000101001",
  35309=>"010010000",
  35310=>"001001110",
  35311=>"101011101",
  35312=>"110000001",
  35313=>"000011000",
  35314=>"010000010",
  35315=>"111000101",
  35316=>"100100010",
  35317=>"100100111",
  35318=>"011010100",
  35319=>"110000011",
  35320=>"001111011",
  35321=>"100010100",
  35322=>"101000101",
  35323=>"101000111",
  35324=>"100011001",
  35325=>"101101100",
  35326=>"011010010",
  35327=>"010110010",
  35328=>"100001101",
  35329=>"100110111",
  35330=>"111010010",
  35331=>"110100011",
  35332=>"100100011",
  35333=>"100000011",
  35334=>"001011000",
  35335=>"111000100",
  35336=>"000111001",
  35337=>"111011101",
  35338=>"111011010",
  35339=>"010011011",
  35340=>"000010000",
  35341=>"000111100",
  35342=>"101101111",
  35343=>"111111110",
  35344=>"101101010",
  35345=>"110010001",
  35346=>"101100011",
  35347=>"110100001",
  35348=>"101000000",
  35349=>"010001101",
  35350=>"001111011",
  35351=>"010011101",
  35352=>"010001100",
  35353=>"100101110",
  35354=>"011101001",
  35355=>"101001011",
  35356=>"111101001",
  35357=>"111111111",
  35358=>"110001010",
  35359=>"100010101",
  35360=>"101111011",
  35361=>"000110000",
  35362=>"100010011",
  35363=>"011100101",
  35364=>"111011011",
  35365=>"110010000",
  35366=>"100011011",
  35367=>"011001101",
  35368=>"100110100",
  35369=>"000001011",
  35370=>"000100110",
  35371=>"111000111",
  35372=>"010011101",
  35373=>"001011111",
  35374=>"100010001",
  35375=>"010010001",
  35376=>"101110101",
  35377=>"111001111",
  35378=>"101001110",
  35379=>"101111110",
  35380=>"101010010",
  35381=>"111000000",
  35382=>"110010100",
  35383=>"111110001",
  35384=>"000101101",
  35385=>"000011000",
  35386=>"110001101",
  35387=>"110111000",
  35388=>"100000110",
  35389=>"100001000",
  35390=>"000101110",
  35391=>"111111000",
  35392=>"111100101",
  35393=>"110111011",
  35394=>"111001110",
  35395=>"101110000",
  35396=>"101011101",
  35397=>"100100110",
  35398=>"100111000",
  35399=>"100010001",
  35400=>"110010000",
  35401=>"110100010",
  35402=>"101111101",
  35403=>"101101000",
  35404=>"010100100",
  35405=>"100100000",
  35406=>"000101111",
  35407=>"000111110",
  35408=>"110011001",
  35409=>"001101000",
  35410=>"011001000",
  35411=>"100111001",
  35412=>"101110011",
  35413=>"111010000",
  35414=>"001001101",
  35415=>"001000111",
  35416=>"100010101",
  35417=>"101110100",
  35418=>"111001000",
  35419=>"000011000",
  35420=>"000011011",
  35421=>"000101000",
  35422=>"011101101",
  35423=>"001110111",
  35424=>"101111110",
  35425=>"111101010",
  35426=>"100001010",
  35427=>"000001010",
  35428=>"101110001",
  35429=>"000000101",
  35430=>"010111011",
  35431=>"101011100",
  35432=>"011110110",
  35433=>"101010111",
  35434=>"010011010",
  35435=>"011111101",
  35436=>"000101011",
  35437=>"000010010",
  35438=>"111011110",
  35439=>"100101111",
  35440=>"100000101",
  35441=>"100100111",
  35442=>"000011100",
  35443=>"000110100",
  35444=>"011111110",
  35445=>"010010000",
  35446=>"111101111",
  35447=>"110011011",
  35448=>"110011001",
  35449=>"101111101",
  35450=>"001011001",
  35451=>"010100001",
  35452=>"110101000",
  35453=>"001011111",
  35454=>"110001110",
  35455=>"111111111",
  35456=>"011100000",
  35457=>"101011110",
  35458=>"011001110",
  35459=>"001011111",
  35460=>"100100111",
  35461=>"100100000",
  35462=>"000011001",
  35463=>"000100011",
  35464=>"010111111",
  35465=>"011100011",
  35466=>"011010110",
  35467=>"010101011",
  35468=>"101011011",
  35469=>"010000101",
  35470=>"111011000",
  35471=>"011111100",
  35472=>"110010110",
  35473=>"110101111",
  35474=>"010000100",
  35475=>"010111001",
  35476=>"010010100",
  35477=>"000001000",
  35478=>"110100101",
  35479=>"101001101",
  35480=>"110000001",
  35481=>"010000110",
  35482=>"011100110",
  35483=>"111001010",
  35484=>"101001010",
  35485=>"001111110",
  35486=>"100101100",
  35487=>"101100001",
  35488=>"110000111",
  35489=>"100101101",
  35490=>"111110100",
  35491=>"101000110",
  35492=>"111111111",
  35493=>"111001010",
  35494=>"100001100",
  35495=>"000111111",
  35496=>"111011001",
  35497=>"100011111",
  35498=>"110000110",
  35499=>"111000111",
  35500=>"111010101",
  35501=>"001001101",
  35502=>"001100111",
  35503=>"100000000",
  35504=>"000111011",
  35505=>"110110110",
  35506=>"100010101",
  35507=>"010001110",
  35508=>"010011100",
  35509=>"111010111",
  35510=>"000101010",
  35511=>"011101110",
  35512=>"101100100",
  35513=>"101100101",
  35514=>"101110000",
  35515=>"101111111",
  35516=>"011001001",
  35517=>"001010011",
  35518=>"101101100",
  35519=>"110111010",
  35520=>"110001001",
  35521=>"110011110",
  35522=>"011101101",
  35523=>"011000111",
  35524=>"011100010",
  35525=>"000101010",
  35526=>"110010010",
  35527=>"100010010",
  35528=>"111100011",
  35529=>"110101011",
  35530=>"100010011",
  35531=>"001000001",
  35532=>"110001001",
  35533=>"000110010",
  35534=>"010010101",
  35535=>"010001000",
  35536=>"011011010",
  35537=>"000000011",
  35538=>"000000010",
  35539=>"001000110",
  35540=>"100100010",
  35541=>"000000001",
  35542=>"111111001",
  35543=>"110001001",
  35544=>"000110010",
  35545=>"001010100",
  35546=>"111000011",
  35547=>"110100000",
  35548=>"100101111",
  35549=>"010010111",
  35550=>"001010001",
  35551=>"100110111",
  35552=>"001001010",
  35553=>"110110111",
  35554=>"001110000",
  35555=>"000001010",
  35556=>"101011011",
  35557=>"101001000",
  35558=>"001000100",
  35559=>"000000010",
  35560=>"101110010",
  35561=>"100010010",
  35562=>"000111100",
  35563=>"001101010",
  35564=>"110011010",
  35565=>"111000110",
  35566=>"110101001",
  35567=>"001000110",
  35568=>"010110110",
  35569=>"110000010",
  35570=>"101100100",
  35571=>"111101010",
  35572=>"000101110",
  35573=>"010001100",
  35574=>"110001111",
  35575=>"011101110",
  35576=>"111010001",
  35577=>"100010000",
  35578=>"000010000",
  35579=>"100101001",
  35580=>"011010010",
  35581=>"100000010",
  35582=>"011101000",
  35583=>"011110100",
  35584=>"110100000",
  35585=>"111101001",
  35586=>"001100000",
  35587=>"101010111",
  35588=>"000011001",
  35589=>"110000000",
  35590=>"001101011",
  35591=>"001011010",
  35592=>"101111100",
  35593=>"100011000",
  35594=>"110111010",
  35595=>"111011001",
  35596=>"000110000",
  35597=>"011100111",
  35598=>"011010000",
  35599=>"000110100",
  35600=>"001000010",
  35601=>"000010111",
  35602=>"001000111",
  35603=>"011101110",
  35604=>"111000001",
  35605=>"011001110",
  35606=>"000111110",
  35607=>"001000000",
  35608=>"111101001",
  35609=>"000000010",
  35610=>"001010000",
  35611=>"110000110",
  35612=>"011100110",
  35613=>"010101010",
  35614=>"111100010",
  35615=>"111011010",
  35616=>"011111111",
  35617=>"110110011",
  35618=>"100011101",
  35619=>"100100011",
  35620=>"111101000",
  35621=>"001101001",
  35622=>"011101001",
  35623=>"010011100",
  35624=>"111011110",
  35625=>"111010000",
  35626=>"111010001",
  35627=>"010001111",
  35628=>"010100101",
  35629=>"000010110",
  35630=>"000100010",
  35631=>"001110000",
  35632=>"010001000",
  35633=>"101101000",
  35634=>"011111111",
  35635=>"011110011",
  35636=>"000101111",
  35637=>"001001110",
  35638=>"111000100",
  35639=>"000010100",
  35640=>"110110110",
  35641=>"010010110",
  35642=>"111000101",
  35643=>"110101110",
  35644=>"000100111",
  35645=>"100000110",
  35646=>"110100101",
  35647=>"000001110",
  35648=>"110001011",
  35649=>"000100010",
  35650=>"101011001",
  35651=>"111100110",
  35652=>"010000111",
  35653=>"101010110",
  35654=>"101001100",
  35655=>"011001011",
  35656=>"101101101",
  35657=>"100011100",
  35658=>"100100110",
  35659=>"101000010",
  35660=>"111010111",
  35661=>"010000000",
  35662=>"010100110",
  35663=>"110011101",
  35664=>"110100001",
  35665=>"101001000",
  35666=>"000110001",
  35667=>"110001100",
  35668=>"001101101",
  35669=>"001011001",
  35670=>"001001110",
  35671=>"001001001",
  35672=>"110100110",
  35673=>"000011100",
  35674=>"011000011",
  35675=>"000110010",
  35676=>"110010000",
  35677=>"110110110",
  35678=>"010011011",
  35679=>"010101111",
  35680=>"001001101",
  35681=>"110001000",
  35682=>"000101000",
  35683=>"111101101",
  35684=>"001011000",
  35685=>"011000100",
  35686=>"000100000",
  35687=>"011101101",
  35688=>"111010101",
  35689=>"110001101",
  35690=>"001100001",
  35691=>"100101001",
  35692=>"111110101",
  35693=>"011100011",
  35694=>"111010100",
  35695=>"010100010",
  35696=>"110010000",
  35697=>"011111001",
  35698=>"110101010",
  35699=>"000101100",
  35700=>"100000000",
  35701=>"100011110",
  35702=>"111101111",
  35703=>"111101111",
  35704=>"011111111",
  35705=>"100110100",
  35706=>"111100110",
  35707=>"100011101",
  35708=>"000000101",
  35709=>"111001110",
  35710=>"110000011",
  35711=>"000110101",
  35712=>"001110111",
  35713=>"011110100",
  35714=>"101010110",
  35715=>"010110000",
  35716=>"100001000",
  35717=>"111000000",
  35718=>"010011111",
  35719=>"000010000",
  35720=>"011110011",
  35721=>"111001111",
  35722=>"000000010",
  35723=>"101000110",
  35724=>"001010111",
  35725=>"000101000",
  35726=>"001101110",
  35727=>"010100000",
  35728=>"101111111",
  35729=>"111111110",
  35730=>"111001101",
  35731=>"111001011",
  35732=>"011100001",
  35733=>"000001000",
  35734=>"110001000",
  35735=>"011100101",
  35736=>"010010011",
  35737=>"100011000",
  35738=>"010001010",
  35739=>"110001001",
  35740=>"001111010",
  35741=>"111000100",
  35742=>"010001111",
  35743=>"000101001",
  35744=>"000100000",
  35745=>"001100111",
  35746=>"100101011",
  35747=>"100000101",
  35748=>"000000000",
  35749=>"100101110",
  35750=>"000001110",
  35751=>"010110101",
  35752=>"100000110",
  35753=>"010000111",
  35754=>"101110111",
  35755=>"011011110",
  35756=>"111011111",
  35757=>"100001110",
  35758=>"100111010",
  35759=>"010011001",
  35760=>"111110000",
  35761=>"100101010",
  35762=>"111011101",
  35763=>"001000111",
  35764=>"011111111",
  35765=>"011110000",
  35766=>"010101111",
  35767=>"100000100",
  35768=>"101111101",
  35769=>"010010110",
  35770=>"001100011",
  35771=>"110100101",
  35772=>"000101001",
  35773=>"111111110",
  35774=>"000011011",
  35775=>"110101110",
  35776=>"101010110",
  35777=>"100010010",
  35778=>"010001101",
  35779=>"011110110",
  35780=>"010010010",
  35781=>"100101001",
  35782=>"111111111",
  35783=>"010010111",
  35784=>"000011111",
  35785=>"010011001",
  35786=>"111110111",
  35787=>"101111001",
  35788=>"001011011",
  35789=>"100101100",
  35790=>"110111001",
  35791=>"010010011",
  35792=>"111100101",
  35793=>"111011000",
  35794=>"111110101",
  35795=>"100010101",
  35796=>"101110110",
  35797=>"001100011",
  35798=>"000010000",
  35799=>"000100110",
  35800=>"110010000",
  35801=>"100100110",
  35802=>"111111111",
  35803=>"010111101",
  35804=>"011100111",
  35805=>"000101000",
  35806=>"101011111",
  35807=>"111001111",
  35808=>"111100010",
  35809=>"110001011",
  35810=>"010000011",
  35811=>"100100010",
  35812=>"010011100",
  35813=>"011001101",
  35814=>"100001010",
  35815=>"101001011",
  35816=>"100100100",
  35817=>"011010010",
  35818=>"001010011",
  35819=>"011000000",
  35820=>"110111111",
  35821=>"101001011",
  35822=>"010110000",
  35823=>"101101011",
  35824=>"001011000",
  35825=>"010111011",
  35826=>"001100110",
  35827=>"000001110",
  35828=>"101000000",
  35829=>"011000100",
  35830=>"010100110",
  35831=>"000100110",
  35832=>"001001001",
  35833=>"101001000",
  35834=>"110001001",
  35835=>"000100111",
  35836=>"001010011",
  35837=>"101011110",
  35838=>"000111010",
  35839=>"011011001",
  35840=>"000101000",
  35841=>"001011101",
  35842=>"010001011",
  35843=>"011100110",
  35844=>"001111010",
  35845=>"111101111",
  35846=>"010111111",
  35847=>"101000100",
  35848=>"100000001",
  35849=>"100011011",
  35850=>"101110101",
  35851=>"001010000",
  35852=>"111100101",
  35853=>"110110000",
  35854=>"010010100",
  35855=>"101000010",
  35856=>"001110001",
  35857=>"001001101",
  35858=>"001010100",
  35859=>"001110001",
  35860=>"000111101",
  35861=>"110010000",
  35862=>"000101110",
  35863=>"110011110",
  35864=>"100110100",
  35865=>"011001110",
  35866=>"000011101",
  35867=>"101101001",
  35868=>"100001111",
  35869=>"101011001",
  35870=>"010001100",
  35871=>"110011101",
  35872=>"011111000",
  35873=>"000010111",
  35874=>"111000110",
  35875=>"010010110",
  35876=>"000111000",
  35877=>"100111010",
  35878=>"000111110",
  35879=>"101100001",
  35880=>"111001001",
  35881=>"011100101",
  35882=>"010111110",
  35883=>"000010011",
  35884=>"000111100",
  35885=>"100000111",
  35886=>"001011101",
  35887=>"111111111",
  35888=>"101111100",
  35889=>"100100110",
  35890=>"101000111",
  35891=>"111011011",
  35892=>"101000000",
  35893=>"111110110",
  35894=>"000000101",
  35895=>"110111101",
  35896=>"001111001",
  35897=>"010101010",
  35898=>"010111010",
  35899=>"001011011",
  35900=>"010110101",
  35901=>"100111000",
  35902=>"000011100",
  35903=>"101011100",
  35904=>"101001010",
  35905=>"001000000",
  35906=>"010101101",
  35907=>"100110010",
  35908=>"000100011",
  35909=>"000000101",
  35910=>"010011000",
  35911=>"000110000",
  35912=>"111011000",
  35913=>"101100101",
  35914=>"010101100",
  35915=>"100010100",
  35916=>"100101001",
  35917=>"110101111",
  35918=>"011100000",
  35919=>"000111010",
  35920=>"100000011",
  35921=>"000101100",
  35922=>"000001100",
  35923=>"101010000",
  35924=>"110011111",
  35925=>"100101110",
  35926=>"010010010",
  35927=>"101111100",
  35928=>"001010011",
  35929=>"011011110",
  35930=>"101010011",
  35931=>"100010110",
  35932=>"000111110",
  35933=>"110110011",
  35934=>"111111110",
  35935=>"010110110",
  35936=>"111110101",
  35937=>"100100010",
  35938=>"101100000",
  35939=>"010001001",
  35940=>"010010111",
  35941=>"011010101",
  35942=>"011001001",
  35943=>"000001111",
  35944=>"100000110",
  35945=>"010110100",
  35946=>"001010011",
  35947=>"011100000",
  35948=>"110111011",
  35949=>"000110011",
  35950=>"100001000",
  35951=>"011101000",
  35952=>"001100101",
  35953=>"011110110",
  35954=>"101000001",
  35955=>"111111111",
  35956=>"000000001",
  35957=>"001101000",
  35958=>"101010011",
  35959=>"010001100",
  35960=>"010110000",
  35961=>"111010100",
  35962=>"100101011",
  35963=>"110011010",
  35964=>"101011110",
  35965=>"110001000",
  35966=>"110110001",
  35967=>"111001111",
  35968=>"001000101",
  35969=>"101100111",
  35970=>"100110111",
  35971=>"010100111",
  35972=>"011110110",
  35973=>"001110000",
  35974=>"011101101",
  35975=>"010110111",
  35976=>"000101101",
  35977=>"110110110",
  35978=>"010010110",
  35979=>"101111100",
  35980=>"000011000",
  35981=>"001110010",
  35982=>"001110000",
  35983=>"001011001",
  35984=>"000010001",
  35985=>"111111101",
  35986=>"010011111",
  35987=>"001100010",
  35988=>"000010110",
  35989=>"101100001",
  35990=>"101001000",
  35991=>"110100000",
  35992=>"111100101",
  35993=>"100110011",
  35994=>"010111100",
  35995=>"111000101",
  35996=>"010000101",
  35997=>"110110100",
  35998=>"101011101",
  35999=>"111011100",
  36000=>"000101010",
  36001=>"010110110",
  36002=>"010101111",
  36003=>"000111111",
  36004=>"011001010",
  36005=>"000001000",
  36006=>"010001110",
  36007=>"010000000",
  36008=>"100010001",
  36009=>"001111100",
  36010=>"010101010",
  36011=>"010101111",
  36012=>"011000011",
  36013=>"100111100",
  36014=>"111111010",
  36015=>"011101000",
  36016=>"101101101",
  36017=>"011110110",
  36018=>"011111111",
  36019=>"101110000",
  36020=>"100010010",
  36021=>"111100111",
  36022=>"010010110",
  36023=>"001010110",
  36024=>"101100000",
  36025=>"110010111",
  36026=>"110010000",
  36027=>"110110011",
  36028=>"100100010",
  36029=>"001111001",
  36030=>"111001011",
  36031=>"011000000",
  36032=>"001001001",
  36033=>"000101101",
  36034=>"011011111",
  36035=>"111000100",
  36036=>"110111110",
  36037=>"000000001",
  36038=>"101101100",
  36039=>"100000111",
  36040=>"010100001",
  36041=>"010011001",
  36042=>"101000000",
  36043=>"010001110",
  36044=>"101110111",
  36045=>"001010010",
  36046=>"000010100",
  36047=>"000100000",
  36048=>"110000111",
  36049=>"001110110",
  36050=>"110011010",
  36051=>"100110101",
  36052=>"100111101",
  36053=>"001001000",
  36054=>"101000101",
  36055=>"110110110",
  36056=>"011111111",
  36057=>"001100101",
  36058=>"101111111",
  36059=>"000011101",
  36060=>"111000010",
  36061=>"011111111",
  36062=>"110011101",
  36063=>"100010010",
  36064=>"101101110",
  36065=>"011011101",
  36066=>"111101010",
  36067=>"000110101",
  36068=>"000110011",
  36069=>"000111000",
  36070=>"101010000",
  36071=>"110101111",
  36072=>"101100110",
  36073=>"011110111",
  36074=>"101000011",
  36075=>"110000111",
  36076=>"100000010",
  36077=>"001100000",
  36078=>"111100101",
  36079=>"101000111",
  36080=>"010000000",
  36081=>"011000001",
  36082=>"110001101",
  36083=>"100000010",
  36084=>"110011100",
  36085=>"000010011",
  36086=>"101001000",
  36087=>"000100000",
  36088=>"000111110",
  36089=>"010101001",
  36090=>"010001001",
  36091=>"000110001",
  36092=>"100000110",
  36093=>"001101110",
  36094=>"100011000",
  36095=>"001001000",
  36096=>"110000011",
  36097=>"111100001",
  36098=>"001110000",
  36099=>"011001011",
  36100=>"111100100",
  36101=>"111100010",
  36102=>"000001010",
  36103=>"101001111",
  36104=>"010110000",
  36105=>"100110001",
  36106=>"101100110",
  36107=>"100101000",
  36108=>"000101110",
  36109=>"010011010",
  36110=>"001100101",
  36111=>"001110010",
  36112=>"000110001",
  36113=>"001011000",
  36114=>"010001000",
  36115=>"011110101",
  36116=>"110110011",
  36117=>"010001110",
  36118=>"111110110",
  36119=>"101100111",
  36120=>"001101001",
  36121=>"100011101",
  36122=>"001101011",
  36123=>"111011010",
  36124=>"111100011",
  36125=>"011011001",
  36126=>"001010111",
  36127=>"110110001",
  36128=>"111111001",
  36129=>"000011001",
  36130=>"110011101",
  36131=>"011101011",
  36132=>"011100000",
  36133=>"100000111",
  36134=>"101100101",
  36135=>"010100110",
  36136=>"101001110",
  36137=>"111111111",
  36138=>"010100000",
  36139=>"010100010",
  36140=>"100101111",
  36141=>"000000000",
  36142=>"110010011",
  36143=>"111001000",
  36144=>"101000100",
  36145=>"111000100",
  36146=>"111100001",
  36147=>"100110100",
  36148=>"011011111",
  36149=>"010011101",
  36150=>"000000000",
  36151=>"110000001",
  36152=>"100111111",
  36153=>"101111111",
  36154=>"000011110",
  36155=>"110011110",
  36156=>"101100010",
  36157=>"011010001",
  36158=>"001001100",
  36159=>"110111001",
  36160=>"100110110",
  36161=>"101101101",
  36162=>"010100111",
  36163=>"010101001",
  36164=>"111101101",
  36165=>"111101111",
  36166=>"010011000",
  36167=>"010110001",
  36168=>"011111101",
  36169=>"010100101",
  36170=>"111110001",
  36171=>"010010110",
  36172=>"001111001",
  36173=>"000001100",
  36174=>"001111100",
  36175=>"000101001",
  36176=>"100110110",
  36177=>"001111001",
  36178=>"100000000",
  36179=>"100111100",
  36180=>"000111000",
  36181=>"111011011",
  36182=>"000111011",
  36183=>"110111010",
  36184=>"001111000",
  36185=>"001111000",
  36186=>"111001101",
  36187=>"000011011",
  36188=>"111100101",
  36189=>"111101000",
  36190=>"100001111",
  36191=>"100011011",
  36192=>"111010110",
  36193=>"101101011",
  36194=>"010000110",
  36195=>"111100011",
  36196=>"111100000",
  36197=>"110111111",
  36198=>"001000001",
  36199=>"111100111",
  36200=>"010111100",
  36201=>"000000111",
  36202=>"101111010",
  36203=>"010100111",
  36204=>"110100010",
  36205=>"100010000",
  36206=>"001000001",
  36207=>"110100100",
  36208=>"011100110",
  36209=>"000001000",
  36210=>"100010100",
  36211=>"101100000",
  36212=>"000010101",
  36213=>"100110011",
  36214=>"000110001",
  36215=>"111101111",
  36216=>"011100111",
  36217=>"111100010",
  36218=>"101011011",
  36219=>"111010010",
  36220=>"000000010",
  36221=>"010100011",
  36222=>"111110101",
  36223=>"100011001",
  36224=>"111111101",
  36225=>"001001100",
  36226=>"111110000",
  36227=>"010101100",
  36228=>"011000100",
  36229=>"100100001",
  36230=>"110111111",
  36231=>"111011110",
  36232=>"110001100",
  36233=>"110001001",
  36234=>"000011010",
  36235=>"000000111",
  36236=>"101101100",
  36237=>"110011110",
  36238=>"010011101",
  36239=>"110011001",
  36240=>"100001100",
  36241=>"010110100",
  36242=>"110010010",
  36243=>"110110100",
  36244=>"011101011",
  36245=>"000100001",
  36246=>"000000000",
  36247=>"010100100",
  36248=>"000010000",
  36249=>"001011110",
  36250=>"000010110",
  36251=>"000001100",
  36252=>"011100100",
  36253=>"001001001",
  36254=>"100101010",
  36255=>"001000010",
  36256=>"001011111",
  36257=>"101011111",
  36258=>"111001101",
  36259=>"011010000",
  36260=>"001011100",
  36261=>"010100110",
  36262=>"010010100",
  36263=>"010010010",
  36264=>"000101100",
  36265=>"011010110",
  36266=>"010001000",
  36267=>"111110011",
  36268=>"100010011",
  36269=>"111110101",
  36270=>"011101100",
  36271=>"101100000",
  36272=>"100110000",
  36273=>"110001010",
  36274=>"110110110",
  36275=>"101011101",
  36276=>"111101110",
  36277=>"111100110",
  36278=>"001100001",
  36279=>"110011100",
  36280=>"101100110",
  36281=>"110001011",
  36282=>"000100111",
  36283=>"100101011",
  36284=>"001101001",
  36285=>"111111100",
  36286=>"001110010",
  36287=>"111100010",
  36288=>"111010111",
  36289=>"110101001",
  36290=>"110101110",
  36291=>"101111100",
  36292=>"101010001",
  36293=>"011100110",
  36294=>"100110111",
  36295=>"101011011",
  36296=>"001100101",
  36297=>"011111111",
  36298=>"010101010",
  36299=>"110000011",
  36300=>"101011001",
  36301=>"011000111",
  36302=>"010011001",
  36303=>"101101110",
  36304=>"010010111",
  36305=>"000110111",
  36306=>"101100010",
  36307=>"000011101",
  36308=>"101000111",
  36309=>"011001001",
  36310=>"110011001",
  36311=>"101110010",
  36312=>"100011101",
  36313=>"111000101",
  36314=>"111010101",
  36315=>"011001110",
  36316=>"101010110",
  36317=>"111011010",
  36318=>"111010101",
  36319=>"010111011",
  36320=>"000110101",
  36321=>"001011110",
  36322=>"001001000",
  36323=>"001110011",
  36324=>"001000111",
  36325=>"000101101",
  36326=>"011111110",
  36327=>"111011010",
  36328=>"011100000",
  36329=>"011110001",
  36330=>"010111101",
  36331=>"101101101",
  36332=>"011111011",
  36333=>"010000001",
  36334=>"010010111",
  36335=>"001101110",
  36336=>"010100000",
  36337=>"110010010",
  36338=>"111111100",
  36339=>"010010110",
  36340=>"011100010",
  36341=>"101111000",
  36342=>"110111001",
  36343=>"010100000",
  36344=>"001101101",
  36345=>"010000000",
  36346=>"000010001",
  36347=>"110101111",
  36348=>"101101100",
  36349=>"100101010",
  36350=>"101111111",
  36351=>"011111110",
  36352=>"101101000",
  36353=>"101101011",
  36354=>"011000101",
  36355=>"100110010",
  36356=>"111100000",
  36357=>"000001010",
  36358=>"100101111",
  36359=>"010001000",
  36360=>"010100100",
  36361=>"111110010",
  36362=>"100101100",
  36363=>"000100000",
  36364=>"101110000",
  36365=>"111000011",
  36366=>"011000101",
  36367=>"101011100",
  36368=>"001110001",
  36369=>"001000111",
  36370=>"110111111",
  36371=>"010100110",
  36372=>"010101000",
  36373=>"001101010",
  36374=>"101010111",
  36375=>"100100001",
  36376=>"110000111",
  36377=>"110111100",
  36378=>"111001111",
  36379=>"010111110",
  36380=>"111001100",
  36381=>"111101110",
  36382=>"001101101",
  36383=>"101110111",
  36384=>"011001111",
  36385=>"001101110",
  36386=>"000110011",
  36387=>"001010011",
  36388=>"110001011",
  36389=>"101100001",
  36390=>"101111001",
  36391=>"001011001",
  36392=>"101101000",
  36393=>"100111000",
  36394=>"010001111",
  36395=>"111010110",
  36396=>"101111111",
  36397=>"010101000",
  36398=>"101011000",
  36399=>"000111010",
  36400=>"010110010",
  36401=>"001111001",
  36402=>"001100011",
  36403=>"110011011",
  36404=>"001101011",
  36405=>"101101101",
  36406=>"101110010",
  36407=>"100111111",
  36408=>"010110001",
  36409=>"101111001",
  36410=>"101001100",
  36411=>"011101011",
  36412=>"100000010",
  36413=>"000011100",
  36414=>"010000010",
  36415=>"001100010",
  36416=>"001001111",
  36417=>"100110010",
  36418=>"000100000",
  36419=>"000010001",
  36420=>"000110100",
  36421=>"011000010",
  36422=>"111011011",
  36423=>"001101011",
  36424=>"110110100",
  36425=>"111001000",
  36426=>"110110110",
  36427=>"010011101",
  36428=>"110011011",
  36429=>"000010010",
  36430=>"100111111",
  36431=>"111101110",
  36432=>"010010101",
  36433=>"011001111",
  36434=>"011110101",
  36435=>"010100001",
  36436=>"000001011",
  36437=>"010100011",
  36438=>"101010101",
  36439=>"010110011",
  36440=>"100000110",
  36441=>"101010001",
  36442=>"100001000",
  36443=>"100011001",
  36444=>"010011000",
  36445=>"001111110",
  36446=>"100111010",
  36447=>"110000001",
  36448=>"110110000",
  36449=>"010010111",
  36450=>"010011111",
  36451=>"100101111",
  36452=>"111111100",
  36453=>"101001110",
  36454=>"000000110",
  36455=>"101010010",
  36456=>"100001010",
  36457=>"000011101",
  36458=>"101001000",
  36459=>"110011011",
  36460=>"001100110",
  36461=>"111101001",
  36462=>"000011101",
  36463=>"101101111",
  36464=>"111110111",
  36465=>"011111001",
  36466=>"111000000",
  36467=>"110111011",
  36468=>"011101101",
  36469=>"101011100",
  36470=>"100110001",
  36471=>"110010010",
  36472=>"110101100",
  36473=>"000001101",
  36474=>"001110000",
  36475=>"000100011",
  36476=>"101000010",
  36477=>"000000000",
  36478=>"111001000",
  36479=>"001101101",
  36480=>"110111000",
  36481=>"111000101",
  36482=>"111000010",
  36483=>"001110110",
  36484=>"010101110",
  36485=>"010100010",
  36486=>"110100010",
  36487=>"101101011",
  36488=>"110000101",
  36489=>"011100101",
  36490=>"010101100",
  36491=>"110100111",
  36492=>"100000100",
  36493=>"001100101",
  36494=>"111101000",
  36495=>"011111010",
  36496=>"000100001",
  36497=>"100010010",
  36498=>"011001110",
  36499=>"011100011",
  36500=>"111101011",
  36501=>"010001000",
  36502=>"101111111",
  36503=>"000100111",
  36504=>"100000011",
  36505=>"001010011",
  36506=>"111111000",
  36507=>"001110010",
  36508=>"110010010",
  36509=>"010011001",
  36510=>"101111100",
  36511=>"111011010",
  36512=>"010111101",
  36513=>"000100101",
  36514=>"110010001",
  36515=>"101111101",
  36516=>"101111111",
  36517=>"101101001",
  36518=>"001111111",
  36519=>"001101010",
  36520=>"011110100",
  36521=>"000011111",
  36522=>"000010010",
  36523=>"111011010",
  36524=>"000011011",
  36525=>"100011000",
  36526=>"101101100",
  36527=>"110101111",
  36528=>"110011111",
  36529=>"011111001",
  36530=>"010111101",
  36531=>"011100100",
  36532=>"001101010",
  36533=>"111110111",
  36534=>"111111010",
  36535=>"101111111",
  36536=>"111110100",
  36537=>"111100010",
  36538=>"011010101",
  36539=>"000011010",
  36540=>"111001111",
  36541=>"011001000",
  36542=>"110000011",
  36543=>"111010010",
  36544=>"110110110",
  36545=>"010101101",
  36546=>"100100000",
  36547=>"101000010",
  36548=>"111111001",
  36549=>"101011100",
  36550=>"011010000",
  36551=>"010101000",
  36552=>"011001010",
  36553=>"110111001",
  36554=>"101111011",
  36555=>"110111010",
  36556=>"101000010",
  36557=>"000010010",
  36558=>"110111100",
  36559=>"000010000",
  36560=>"110011111",
  36561=>"010110100",
  36562=>"110100000",
  36563=>"100001010",
  36564=>"000110001",
  36565=>"100100111",
  36566=>"101110010",
  36567=>"101000100",
  36568=>"000101101",
  36569=>"111010001",
  36570=>"111100111",
  36571=>"010001110",
  36572=>"101001010",
  36573=>"001010010",
  36574=>"011110110",
  36575=>"011101010",
  36576=>"101100111",
  36577=>"100001111",
  36578=>"010100010",
  36579=>"010110101",
  36580=>"110110111",
  36581=>"110000100",
  36582=>"110011000",
  36583=>"101011100",
  36584=>"101110001",
  36585=>"111110110",
  36586=>"100010010",
  36587=>"111111101",
  36588=>"100110110",
  36589=>"111100011",
  36590=>"110111001",
  36591=>"011100010",
  36592=>"100101110",
  36593=>"100101101",
  36594=>"101010011",
  36595=>"101011011",
  36596=>"011010110",
  36597=>"010111111",
  36598=>"000010100",
  36599=>"000001110",
  36600=>"000001100",
  36601=>"010100000",
  36602=>"110001001",
  36603=>"100100011",
  36604=>"100000000",
  36605=>"101001100",
  36606=>"001001101",
  36607=>"000001100",
  36608=>"110011111",
  36609=>"001110010",
  36610=>"010110100",
  36611=>"011100100",
  36612=>"101010000",
  36613=>"001000110",
  36614=>"111101111",
  36615=>"001010001",
  36616=>"101110100",
  36617=>"000111111",
  36618=>"101001001",
  36619=>"011001111",
  36620=>"000001110",
  36621=>"101101011",
  36622=>"100011111",
  36623=>"010111000",
  36624=>"111000111",
  36625=>"010010110",
  36626=>"110101000",
  36627=>"110000000",
  36628=>"110111101",
  36629=>"101010101",
  36630=>"001000111",
  36631=>"110011111",
  36632=>"001101111",
  36633=>"100001110",
  36634=>"010110101",
  36635=>"100111110",
  36636=>"100110111",
  36637=>"011111011",
  36638=>"010000101",
  36639=>"101011000",
  36640=>"100111101",
  36641=>"001110010",
  36642=>"111101001",
  36643=>"110000011",
  36644=>"010011110",
  36645=>"000111000",
  36646=>"001100101",
  36647=>"011110000",
  36648=>"111000010",
  36649=>"011111000",
  36650=>"100100110",
  36651=>"111101101",
  36652=>"110110000",
  36653=>"010010000",
  36654=>"001100001",
  36655=>"111010110",
  36656=>"000000011",
  36657=>"000111011",
  36658=>"001011101",
  36659=>"010011111",
  36660=>"111111001",
  36661=>"111101101",
  36662=>"010111011",
  36663=>"100001011",
  36664=>"011000110",
  36665=>"000010101",
  36666=>"111101110",
  36667=>"100001001",
  36668=>"111110001",
  36669=>"000001010",
  36670=>"010100101",
  36671=>"001011000",
  36672=>"011110110",
  36673=>"100100101",
  36674=>"001110111",
  36675=>"100011010",
  36676=>"000100111",
  36677=>"110000011",
  36678=>"011011001",
  36679=>"101010100",
  36680=>"000100010",
  36681=>"001101101",
  36682=>"010010001",
  36683=>"110100000",
  36684=>"001101100",
  36685=>"001011111",
  36686=>"111001101",
  36687=>"101111100",
  36688=>"010101000",
  36689=>"000100111",
  36690=>"101110010",
  36691=>"000010011",
  36692=>"110000110",
  36693=>"101100111",
  36694=>"001000101",
  36695=>"100110110",
  36696=>"010110100",
  36697=>"010010000",
  36698=>"010011100",
  36699=>"100001010",
  36700=>"110100100",
  36701=>"010110101",
  36702=>"001101100",
  36703=>"000010010",
  36704=>"111110000",
  36705=>"010101010",
  36706=>"111100000",
  36707=>"001011000",
  36708=>"110111001",
  36709=>"111000101",
  36710=>"101110100",
  36711=>"001010111",
  36712=>"110110111",
  36713=>"100110110",
  36714=>"110101010",
  36715=>"110001100",
  36716=>"101001001",
  36717=>"101100001",
  36718=>"110001001",
  36719=>"110011111",
  36720=>"100000111",
  36721=>"101010110",
  36722=>"001001000",
  36723=>"011100110",
  36724=>"000100110",
  36725=>"110100000",
  36726=>"101110101",
  36727=>"011001011",
  36728=>"100100100",
  36729=>"110010110",
  36730=>"001000110",
  36731=>"110001101",
  36732=>"011011110",
  36733=>"011000101",
  36734=>"000000011",
  36735=>"011011010",
  36736=>"110101101",
  36737=>"100000111",
  36738=>"100101011",
  36739=>"110000000",
  36740=>"001111100",
  36741=>"110010001",
  36742=>"001100010",
  36743=>"110100010",
  36744=>"111100111",
  36745=>"000011110",
  36746=>"001011111",
  36747=>"000110010",
  36748=>"110010000",
  36749=>"101111101",
  36750=>"100011101",
  36751=>"101010000",
  36752=>"111101111",
  36753=>"001111110",
  36754=>"000111111",
  36755=>"101010101",
  36756=>"011101000",
  36757=>"010011110",
  36758=>"001111011",
  36759=>"110011011",
  36760=>"101100100",
  36761=>"101101101",
  36762=>"000001011",
  36763=>"010110101",
  36764=>"000000111",
  36765=>"001010001",
  36766=>"000001111",
  36767=>"011010000",
  36768=>"000111111",
  36769=>"011110011",
  36770=>"010111001",
  36771=>"101110010",
  36772=>"101000001",
  36773=>"011010001",
  36774=>"000111110",
  36775=>"111110101",
  36776=>"101110101",
  36777=>"010010011",
  36778=>"100000011",
  36779=>"011110010",
  36780=>"000010011",
  36781=>"101010100",
  36782=>"100101101",
  36783=>"110000001",
  36784=>"111011001",
  36785=>"001010000",
  36786=>"001101001",
  36787=>"001011001",
  36788=>"101100111",
  36789=>"100001101",
  36790=>"001110110",
  36791=>"110010111",
  36792=>"000011111",
  36793=>"010000000",
  36794=>"110111111",
  36795=>"000000010",
  36796=>"111101100",
  36797=>"010100111",
  36798=>"111011111",
  36799=>"000001001",
  36800=>"010001010",
  36801=>"001000101",
  36802=>"101100010",
  36803=>"110110101",
  36804=>"100110010",
  36805=>"111101000",
  36806=>"101111001",
  36807=>"001000010",
  36808=>"000010011",
  36809=>"001011111",
  36810=>"110001111",
  36811=>"111011011",
  36812=>"111111010",
  36813=>"111110111",
  36814=>"001100000",
  36815=>"001100010",
  36816=>"100011111",
  36817=>"010000101",
  36818=>"101010010",
  36819=>"010011110",
  36820=>"101011000",
  36821=>"110011000",
  36822=>"100000001",
  36823=>"000110100",
  36824=>"111110001",
  36825=>"101001001",
  36826=>"011001101",
  36827=>"011110110",
  36828=>"100101111",
  36829=>"010001100",
  36830=>"100100011",
  36831=>"110111010",
  36832=>"101111110",
  36833=>"110101000",
  36834=>"010000011",
  36835=>"010010001",
  36836=>"101110111",
  36837=>"011010110",
  36838=>"100101111",
  36839=>"001011110",
  36840=>"000111011",
  36841=>"011001000",
  36842=>"100000010",
  36843=>"010111101",
  36844=>"111111000",
  36845=>"100000011",
  36846=>"101100101",
  36847=>"011011101",
  36848=>"001100011",
  36849=>"011001101",
  36850=>"101101101",
  36851=>"000110101",
  36852=>"100010001",
  36853=>"100110100",
  36854=>"100000111",
  36855=>"110000110",
  36856=>"010101101",
  36857=>"111000110",
  36858=>"110111011",
  36859=>"111110010",
  36860=>"000100101",
  36861=>"111010011",
  36862=>"000010110",
  36863=>"111000100",
  36864=>"111100000",
  36865=>"110000100",
  36866=>"101010101",
  36867=>"111010101",
  36868=>"010000000",
  36869=>"101001101",
  36870=>"001100000",
  36871=>"111101010",
  36872=>"001100101",
  36873=>"111010100",
  36874=>"010110001",
  36875=>"111110110",
  36876=>"101000000",
  36877=>"001011110",
  36878=>"101010111",
  36879=>"001110010",
  36880=>"010000101",
  36881=>"111101001",
  36882=>"000000110",
  36883=>"100100010",
  36884=>"111100000",
  36885=>"000010010",
  36886=>"110011111",
  36887=>"011101001",
  36888=>"111110111",
  36889=>"001101100",
  36890=>"010000111",
  36891=>"001010101",
  36892=>"101101011",
  36893=>"110010110",
  36894=>"010100101",
  36895=>"100100010",
  36896=>"011010101",
  36897=>"101101001",
  36898=>"010010011",
  36899=>"101101110",
  36900=>"101111011",
  36901=>"010000000",
  36902=>"111101001",
  36903=>"110010100",
  36904=>"110001001",
  36905=>"100101010",
  36906=>"010010011",
  36907=>"110000011",
  36908=>"101110111",
  36909=>"101110010",
  36910=>"010001111",
  36911=>"010110010",
  36912=>"111001100",
  36913=>"000010001",
  36914=>"100100010",
  36915=>"011010001",
  36916=>"111000010",
  36917=>"001111000",
  36918=>"110110000",
  36919=>"110100011",
  36920=>"001101001",
  36921=>"000001011",
  36922=>"101100011",
  36923=>"000000100",
  36924=>"110011101",
  36925=>"001101110",
  36926=>"001001010",
  36927=>"001100110",
  36928=>"100010100",
  36929=>"110100101",
  36930=>"110011010",
  36931=>"101001100",
  36932=>"000110110",
  36933=>"010111001",
  36934=>"000011001",
  36935=>"010001111",
  36936=>"111001010",
  36937=>"110010000",
  36938=>"000000110",
  36939=>"111100000",
  36940=>"110100000",
  36941=>"110010100",
  36942=>"110001011",
  36943=>"100100110",
  36944=>"000111111",
  36945=>"000100100",
  36946=>"010011101",
  36947=>"101110100",
  36948=>"111000111",
  36949=>"000011000",
  36950=>"111000111",
  36951=>"001001001",
  36952=>"110011001",
  36953=>"001110111",
  36954=>"100110110",
  36955=>"100010101",
  36956=>"101011000",
  36957=>"101000011",
  36958=>"001111011",
  36959=>"010001010",
  36960=>"110100000",
  36961=>"110001110",
  36962=>"001111111",
  36963=>"011001101",
  36964=>"010000010",
  36965=>"000001000",
  36966=>"000000011",
  36967=>"111111000",
  36968=>"011110000",
  36969=>"100011000",
  36970=>"111010010",
  36971=>"111000110",
  36972=>"000101010",
  36973=>"001101000",
  36974=>"011100011",
  36975=>"101011100",
  36976=>"000111101",
  36977=>"000111101",
  36978=>"110111010",
  36979=>"100011110",
  36980=>"000010101",
  36981=>"111011000",
  36982=>"101100001",
  36983=>"011011100",
  36984=>"011100101",
  36985=>"001000000",
  36986=>"000001011",
  36987=>"000000100",
  36988=>"011100110",
  36989=>"110011010",
  36990=>"000000000",
  36991=>"111101101",
  36992=>"110010010",
  36993=>"100011111",
  36994=>"101011011",
  36995=>"001100010",
  36996=>"011000011",
  36997=>"110010100",
  36998=>"001110000",
  36999=>"000110101",
  37000=>"100100000",
  37001=>"111011011",
  37002=>"000001111",
  37003=>"101111011",
  37004=>"111100101",
  37005=>"011011001",
  37006=>"111010101",
  37007=>"111000010",
  37008=>"100110110",
  37009=>"101101011",
  37010=>"111001101",
  37011=>"111000110",
  37012=>"110000010",
  37013=>"100000011",
  37014=>"000101000",
  37015=>"111101011",
  37016=>"011111100",
  37017=>"010110101",
  37018=>"111101100",
  37019=>"011011101",
  37020=>"101011010",
  37021=>"001001000",
  37022=>"010111010",
  37023=>"010010000",
  37024=>"111010101",
  37025=>"101100010",
  37026=>"100000111",
  37027=>"111011110",
  37028=>"011101111",
  37029=>"111110111",
  37030=>"010010011",
  37031=>"000010000",
  37032=>"001001000",
  37033=>"011001101",
  37034=>"010001111",
  37035=>"100010101",
  37036=>"110001000",
  37037=>"001000110",
  37038=>"110010011",
  37039=>"110101111",
  37040=>"010010001",
  37041=>"001010100",
  37042=>"100111000",
  37043=>"111101111",
  37044=>"000000110",
  37045=>"000100101",
  37046=>"101111110",
  37047=>"110010100",
  37048=>"000101000",
  37049=>"010101100",
  37050=>"110001101",
  37051=>"111001110",
  37052=>"000110111",
  37053=>"001111100",
  37054=>"000000100",
  37055=>"110110011",
  37056=>"010101110",
  37057=>"000011000",
  37058=>"111100001",
  37059=>"001011011",
  37060=>"000011101",
  37061=>"010101000",
  37062=>"101100101",
  37063=>"011110001",
  37064=>"000011011",
  37065=>"000101011",
  37066=>"000011011",
  37067=>"000000011",
  37068=>"010100110",
  37069=>"100111101",
  37070=>"011011111",
  37071=>"010100011",
  37072=>"110100110",
  37073=>"111000111",
  37074=>"001001001",
  37075=>"010111100",
  37076=>"100101010",
  37077=>"010011100",
  37078=>"010110001",
  37079=>"000011101",
  37080=>"111100100",
  37081=>"100011011",
  37082=>"000010000",
  37083=>"000010111",
  37084=>"010110011",
  37085=>"010110100",
  37086=>"011001100",
  37087=>"000101110",
  37088=>"011101011",
  37089=>"011110000",
  37090=>"001000010",
  37091=>"011111111",
  37092=>"111111001",
  37093=>"001011011",
  37094=>"100100111",
  37095=>"010110001",
  37096=>"111000010",
  37097=>"101110010",
  37098=>"101011101",
  37099=>"110111100",
  37100=>"101100110",
  37101=>"001010010",
  37102=>"011100101",
  37103=>"010110111",
  37104=>"010010011",
  37105=>"001000100",
  37106=>"000011011",
  37107=>"000101010",
  37108=>"111100111",
  37109=>"100101010",
  37110=>"010100101",
  37111=>"000100110",
  37112=>"101000111",
  37113=>"100000111",
  37114=>"110001101",
  37115=>"111101010",
  37116=>"111101011",
  37117=>"001001110",
  37118=>"110000111",
  37119=>"011000101",
  37120=>"011010000",
  37121=>"010000100",
  37122=>"100110011",
  37123=>"001000111",
  37124=>"101000111",
  37125=>"100010110",
  37126=>"111000001",
  37127=>"101100000",
  37128=>"100000010",
  37129=>"110001111",
  37130=>"011001101",
  37131=>"100001110",
  37132=>"000011011",
  37133=>"110100100",
  37134=>"010111100",
  37135=>"111001001",
  37136=>"001001111",
  37137=>"101011000",
  37138=>"001000000",
  37139=>"110010000",
  37140=>"110101000",
  37141=>"111000110",
  37142=>"001100010",
  37143=>"000101110",
  37144=>"011110111",
  37145=>"000100000",
  37146=>"101010110",
  37147=>"001110001",
  37148=>"111001000",
  37149=>"011011010",
  37150=>"000011010",
  37151=>"101101001",
  37152=>"010111000",
  37153=>"000101110",
  37154=>"101001011",
  37155=>"101100100",
  37156=>"000100111",
  37157=>"011111010",
  37158=>"001101000",
  37159=>"110111010",
  37160=>"000001101",
  37161=>"100011111",
  37162=>"110011010",
  37163=>"010011010",
  37164=>"010111111",
  37165=>"000000111",
  37166=>"001001000",
  37167=>"101011100",
  37168=>"001010011",
  37169=>"000010010",
  37170=>"101111100",
  37171=>"011000000",
  37172=>"101010110",
  37173=>"011111001",
  37174=>"000101010",
  37175=>"111100111",
  37176=>"011011000",
  37177=>"001111000",
  37178=>"111001001",
  37179=>"001100110",
  37180=>"011110010",
  37181=>"011010011",
  37182=>"000100001",
  37183=>"111100011",
  37184=>"111111100",
  37185=>"000010001",
  37186=>"110000100",
  37187=>"101100000",
  37188=>"110011010",
  37189=>"101100101",
  37190=>"001100111",
  37191=>"101101000",
  37192=>"110011111",
  37193=>"100111011",
  37194=>"100011110",
  37195=>"000010110",
  37196=>"011011000",
  37197=>"110100011",
  37198=>"101001101",
  37199=>"001110011",
  37200=>"000101110",
  37201=>"100000000",
  37202=>"010111100",
  37203=>"100100101",
  37204=>"111101111",
  37205=>"001000100",
  37206=>"111110011",
  37207=>"111001011",
  37208=>"001001000",
  37209=>"111100011",
  37210=>"010001010",
  37211=>"110110100",
  37212=>"100110011",
  37213=>"010000111",
  37214=>"011011010",
  37215=>"100001110",
  37216=>"111101110",
  37217=>"001011001",
  37218=>"110001011",
  37219=>"101001011",
  37220=>"010000011",
  37221=>"101000101",
  37222=>"011110100",
  37223=>"100011110",
  37224=>"100110000",
  37225=>"111101010",
  37226=>"100101011",
  37227=>"011000000",
  37228=>"111101111",
  37229=>"001101001",
  37230=>"000001100",
  37231=>"010101001",
  37232=>"111000100",
  37233=>"100011101",
  37234=>"100101000",
  37235=>"100110000",
  37236=>"111000111",
  37237=>"010001000",
  37238=>"000011000",
  37239=>"111000101",
  37240=>"000000010",
  37241=>"110111110",
  37242=>"001110010",
  37243=>"111111010",
  37244=>"001111110",
  37245=>"010101010",
  37246=>"000001111",
  37247=>"101100111",
  37248=>"001110100",
  37249=>"010011101",
  37250=>"111111010",
  37251=>"001010100",
  37252=>"001000010",
  37253=>"101110101",
  37254=>"110111100",
  37255=>"001001101",
  37256=>"010111000",
  37257=>"101110111",
  37258=>"110110010",
  37259=>"011101011",
  37260=>"100011101",
  37261=>"101110111",
  37262=>"001101001",
  37263=>"100101101",
  37264=>"010011111",
  37265=>"100001100",
  37266=>"010101011",
  37267=>"001101000",
  37268=>"011100011",
  37269=>"000011010",
  37270=>"101000001",
  37271=>"111011111",
  37272=>"000000000",
  37273=>"001001000",
  37274=>"100001001",
  37275=>"101001010",
  37276=>"101111100",
  37277=>"010110000",
  37278=>"010001010",
  37279=>"111000100",
  37280=>"111000000",
  37281=>"010100011",
  37282=>"111010010",
  37283=>"111010001",
  37284=>"010100011",
  37285=>"010000111",
  37286=>"010001011",
  37287=>"010000111",
  37288=>"110011100",
  37289=>"110001101",
  37290=>"000010000",
  37291=>"111100010",
  37292=>"110000110",
  37293=>"001110110",
  37294=>"100100101",
  37295=>"100011000",
  37296=>"001001011",
  37297=>"111010110",
  37298=>"100100000",
  37299=>"101011100",
  37300=>"110011111",
  37301=>"000100100",
  37302=>"001001001",
  37303=>"110000101",
  37304=>"111100101",
  37305=>"001101011",
  37306=>"000101001",
  37307=>"110101010",
  37308=>"110000111",
  37309=>"101101100",
  37310=>"000110000",
  37311=>"001011111",
  37312=>"111001111",
  37313=>"010001111",
  37314=>"100111100",
  37315=>"010001110",
  37316=>"100000111",
  37317=>"111001100",
  37318=>"011000011",
  37319=>"001101000",
  37320=>"010001110",
  37321=>"100000001",
  37322=>"110101011",
  37323=>"011000100",
  37324=>"100000001",
  37325=>"000110100",
  37326=>"111011001",
  37327=>"000111111",
  37328=>"010110100",
  37329=>"101011100",
  37330=>"001010001",
  37331=>"001011010",
  37332=>"111101111",
  37333=>"010100100",
  37334=>"111101100",
  37335=>"101100001",
  37336=>"010101101",
  37337=>"010110100",
  37338=>"010011011",
  37339=>"000100100",
  37340=>"111100101",
  37341=>"110000011",
  37342=>"011001011",
  37343=>"010110000",
  37344=>"110110110",
  37345=>"100100000",
  37346=>"111111010",
  37347=>"010000111",
  37348=>"110011111",
  37349=>"010011011",
  37350=>"010101010",
  37351=>"000010101",
  37352=>"111111110",
  37353=>"001111001",
  37354=>"010000100",
  37355=>"101110101",
  37356=>"111000111",
  37357=>"000000000",
  37358=>"100001100",
  37359=>"100000100",
  37360=>"100110100",
  37361=>"101001011",
  37362=>"101110011",
  37363=>"001100111",
  37364=>"001000011",
  37365=>"110111000",
  37366=>"010101110",
  37367=>"011010001",
  37368=>"100100000",
  37369=>"111011100",
  37370=>"101111101",
  37371=>"111100000",
  37372=>"101001000",
  37373=>"101111110",
  37374=>"101001010",
  37375=>"100010101",
  37376=>"001111111",
  37377=>"100001011",
  37378=>"111101011",
  37379=>"011001011",
  37380=>"010100010",
  37381=>"010101000",
  37382=>"110011011",
  37383=>"101000100",
  37384=>"110011000",
  37385=>"010110101",
  37386=>"010101110",
  37387=>"110000001",
  37388=>"111011100",
  37389=>"111001111",
  37390=>"000001101",
  37391=>"010001111",
  37392=>"001001101",
  37393=>"000010100",
  37394=>"101100000",
  37395=>"010111101",
  37396=>"011100011",
  37397=>"010110001",
  37398=>"011111100",
  37399=>"011110111",
  37400=>"101100001",
  37401=>"000111100",
  37402=>"001100000",
  37403=>"000100101",
  37404=>"000001100",
  37405=>"001101001",
  37406=>"100100001",
  37407=>"011001010",
  37408=>"001111000",
  37409=>"111011011",
  37410=>"011000101",
  37411=>"100010101",
  37412=>"100110110",
  37413=>"011101101",
  37414=>"001010110",
  37415=>"100101100",
  37416=>"111011110",
  37417=>"010011000",
  37418=>"100001010",
  37419=>"110011011",
  37420=>"111110001",
  37421=>"111010011",
  37422=>"011010101",
  37423=>"000001111",
  37424=>"101110000",
  37425=>"111011110",
  37426=>"100111101",
  37427=>"111011001",
  37428=>"011100110",
  37429=>"110111000",
  37430=>"101010000",
  37431=>"100010011",
  37432=>"100111111",
  37433=>"001111001",
  37434=>"110110000",
  37435=>"110101000",
  37436=>"000100000",
  37437=>"011100101",
  37438=>"010101000",
  37439=>"100010101",
  37440=>"000001000",
  37441=>"101101101",
  37442=>"111100111",
  37443=>"011110001",
  37444=>"101001100",
  37445=>"011001001",
  37446=>"011000000",
  37447=>"000101100",
  37448=>"010110111",
  37449=>"101111001",
  37450=>"110110110",
  37451=>"110000001",
  37452=>"101011100",
  37453=>"101011001",
  37454=>"111000100",
  37455=>"011001100",
  37456=>"110000110",
  37457=>"001011000",
  37458=>"010111001",
  37459=>"110011010",
  37460=>"101111011",
  37461=>"011001010",
  37462=>"101000000",
  37463=>"001111100",
  37464=>"110011000",
  37465=>"100010001",
  37466=>"011001011",
  37467=>"000110100",
  37468=>"100100110",
  37469=>"011100000",
  37470=>"000011101",
  37471=>"101110011",
  37472=>"011001110",
  37473=>"010011011",
  37474=>"011100000",
  37475=>"111101001",
  37476=>"011011001",
  37477=>"011100111",
  37478=>"100101110",
  37479=>"000000100",
  37480=>"110100010",
  37481=>"110010110",
  37482=>"000110100",
  37483=>"111110000",
  37484=>"110001001",
  37485=>"100100100",
  37486=>"110010100",
  37487=>"010001111",
  37488=>"110000101",
  37489=>"111111100",
  37490=>"010000111",
  37491=>"110000110",
  37492=>"011011000",
  37493=>"100000000",
  37494=>"011001011",
  37495=>"100010110",
  37496=>"110010101",
  37497=>"101010110",
  37498=>"000011010",
  37499=>"111111010",
  37500=>"000011111",
  37501=>"010101011",
  37502=>"110101100",
  37503=>"011110110",
  37504=>"010101010",
  37505=>"101111100",
  37506=>"111101111",
  37507=>"001000000",
  37508=>"000000000",
  37509=>"110000110",
  37510=>"011110111",
  37511=>"111110100",
  37512=>"000010111",
  37513=>"110011010",
  37514=>"000101111",
  37515=>"011011111",
  37516=>"001000010",
  37517=>"011000100",
  37518=>"110001010",
  37519=>"001100110",
  37520=>"001111101",
  37521=>"110011110",
  37522=>"111110111",
  37523=>"100011010",
  37524=>"100100111",
  37525=>"100110111",
  37526=>"001110000",
  37527=>"101110000",
  37528=>"001010010",
  37529=>"111110110",
  37530=>"110100110",
  37531=>"101010101",
  37532=>"000100110",
  37533=>"100010010",
  37534=>"101000000",
  37535=>"000111100",
  37536=>"111010010",
  37537=>"101000101",
  37538=>"001000101",
  37539=>"011011010",
  37540=>"110101101",
  37541=>"011101110",
  37542=>"101111101",
  37543=>"111001001",
  37544=>"110000010",
  37545=>"011010100",
  37546=>"001101000",
  37547=>"010010000",
  37548=>"000000011",
  37549=>"100000100",
  37550=>"010010111",
  37551=>"001000110",
  37552=>"101100101",
  37553=>"100001111",
  37554=>"100001011",
  37555=>"111110101",
  37556=>"100100110",
  37557=>"100000111",
  37558=>"001001001",
  37559=>"100000011",
  37560=>"110001010",
  37561=>"101011000",
  37562=>"011100110",
  37563=>"000111111",
  37564=>"111110000",
  37565=>"010001000",
  37566=>"001001100",
  37567=>"110001111",
  37568=>"101101111",
  37569=>"101101010",
  37570=>"001010101",
  37571=>"011001110",
  37572=>"010010001",
  37573=>"100011101",
  37574=>"111000101",
  37575=>"001001010",
  37576=>"110010101",
  37577=>"000001010",
  37578=>"101010001",
  37579=>"001001111",
  37580=>"001111000",
  37581=>"110000110",
  37582=>"001010111",
  37583=>"010011110",
  37584=>"010111100",
  37585=>"001100101",
  37586=>"100010010",
  37587=>"011000010",
  37588=>"010000100",
  37589=>"111011101",
  37590=>"011110100",
  37591=>"000000101",
  37592=>"100110000",
  37593=>"000000111",
  37594=>"101001010",
  37595=>"100001100",
  37596=>"101101111",
  37597=>"100000001",
  37598=>"010101101",
  37599=>"111100110",
  37600=>"001000110",
  37601=>"101000110",
  37602=>"010100101",
  37603=>"110011101",
  37604=>"011001010",
  37605=>"010101000",
  37606=>"100000100",
  37607=>"110111001",
  37608=>"000011010",
  37609=>"011001011",
  37610=>"100000110",
  37611=>"101011011",
  37612=>"010011000",
  37613=>"010010001",
  37614=>"001011100",
  37615=>"110001111",
  37616=>"110010001",
  37617=>"101011111",
  37618=>"111111001",
  37619=>"110110011",
  37620=>"001010001",
  37621=>"111110010",
  37622=>"110110101",
  37623=>"111101101",
  37624=>"101101111",
  37625=>"000001010",
  37626=>"101000111",
  37627=>"000001001",
  37628=>"110011110",
  37629=>"001110100",
  37630=>"011000001",
  37631=>"110111011",
  37632=>"011010110",
  37633=>"110000000",
  37634=>"111111101",
  37635=>"101000000",
  37636=>"000001101",
  37637=>"100000011",
  37638=>"111011010",
  37639=>"001101111",
  37640=>"000011110",
  37641=>"110111011",
  37642=>"010000001",
  37643=>"000011100",
  37644=>"110110011",
  37645=>"010110100",
  37646=>"011101000",
  37647=>"100011010",
  37648=>"111011001",
  37649=>"101101101",
  37650=>"000111000",
  37651=>"100011011",
  37652=>"101111100",
  37653=>"010001111",
  37654=>"010001111",
  37655=>"111011111",
  37656=>"000101111",
  37657=>"011110000",
  37658=>"000100010",
  37659=>"111000011",
  37660=>"011000000",
  37661=>"111101010",
  37662=>"001000110",
  37663=>"100111010",
  37664=>"101110111",
  37665=>"110011101",
  37666=>"011011010",
  37667=>"011011000",
  37668=>"111001100",
  37669=>"101000100",
  37670=>"111011000",
  37671=>"101101101",
  37672=>"110100111",
  37673=>"110001001",
  37674=>"110001101",
  37675=>"100010001",
  37676=>"110011111",
  37677=>"010011110",
  37678=>"000001000",
  37679=>"000010001",
  37680=>"011100011",
  37681=>"100000110",
  37682=>"001011111",
  37683=>"101001100",
  37684=>"101100001",
  37685=>"110101100",
  37686=>"110000010",
  37687=>"000000110",
  37688=>"001111011",
  37689=>"001001001",
  37690=>"011011001",
  37691=>"111110101",
  37692=>"010101111",
  37693=>"010010111",
  37694=>"101011011",
  37695=>"000000001",
  37696=>"011000110",
  37697=>"100110100",
  37698=>"101100001",
  37699=>"001010110",
  37700=>"000000010",
  37701=>"110100011",
  37702=>"110100001",
  37703=>"001100100",
  37704=>"010101110",
  37705=>"001100100",
  37706=>"000110001",
  37707=>"100111011",
  37708=>"011000000",
  37709=>"101001001",
  37710=>"111000001",
  37711=>"110111010",
  37712=>"001101010",
  37713=>"101011000",
  37714=>"000100010",
  37715=>"001111111",
  37716=>"100001101",
  37717=>"000000001",
  37718=>"001110001",
  37719=>"001110010",
  37720=>"010000011",
  37721=>"110101010",
  37722=>"001001000",
  37723=>"001100011",
  37724=>"000000010",
  37725=>"101111000",
  37726=>"001111000",
  37727=>"001110010",
  37728=>"000001000",
  37729=>"010011001",
  37730=>"110101001",
  37731=>"101000110",
  37732=>"011101010",
  37733=>"001101111",
  37734=>"100100001",
  37735=>"011010001",
  37736=>"111010000",
  37737=>"100101101",
  37738=>"011110000",
  37739=>"001111110",
  37740=>"011110000",
  37741=>"101000011",
  37742=>"111100011",
  37743=>"011111101",
  37744=>"111000100",
  37745=>"001101101",
  37746=>"111110101",
  37747=>"100001000",
  37748=>"000001001",
  37749=>"000101101",
  37750=>"010000011",
  37751=>"100101010",
  37752=>"011000010",
  37753=>"100010011",
  37754=>"101011011",
  37755=>"101100101",
  37756=>"100001100",
  37757=>"110101001",
  37758=>"111111111",
  37759=>"100000100",
  37760=>"011110010",
  37761=>"111001110",
  37762=>"001000011",
  37763=>"001001101",
  37764=>"110100111",
  37765=>"111111111",
  37766=>"011111110",
  37767=>"001001000",
  37768=>"101110011",
  37769=>"111111000",
  37770=>"111100100",
  37771=>"011010000",
  37772=>"111100000",
  37773=>"011111111",
  37774=>"110001110",
  37775=>"011011100",
  37776=>"000011100",
  37777=>"000000001",
  37778=>"001101001",
  37779=>"001000101",
  37780=>"001100001",
  37781=>"111010000",
  37782=>"011011010",
  37783=>"000111100",
  37784=>"010100100",
  37785=>"011000010",
  37786=>"010011111",
  37787=>"011000101",
  37788=>"010101010",
  37789=>"110001101",
  37790=>"010100110",
  37791=>"010110001",
  37792=>"000001001",
  37793=>"000110001",
  37794=>"100111001",
  37795=>"101001110",
  37796=>"001001010",
  37797=>"100111110",
  37798=>"010100010",
  37799=>"110000101",
  37800=>"010101110",
  37801=>"101100011",
  37802=>"111110010",
  37803=>"111001111",
  37804=>"000001110",
  37805=>"000110001",
  37806=>"101010110",
  37807=>"100101000",
  37808=>"000001100",
  37809=>"110101101",
  37810=>"001011000",
  37811=>"001110011",
  37812=>"100111111",
  37813=>"110000101",
  37814=>"110111100",
  37815=>"011110001",
  37816=>"001001001",
  37817=>"000011110",
  37818=>"011010000",
  37819=>"001111110",
  37820=>"010000011",
  37821=>"111010001",
  37822=>"101000000",
  37823=>"000001000",
  37824=>"110111010",
  37825=>"001011100",
  37826=>"101101110",
  37827=>"001111010",
  37828=>"110100001",
  37829=>"101000111",
  37830=>"111101110",
  37831=>"000100101",
  37832=>"100110110",
  37833=>"011100000",
  37834=>"010100010",
  37835=>"010101000",
  37836=>"000101110",
  37837=>"001100101",
  37838=>"010111110",
  37839=>"011101111",
  37840=>"111111001",
  37841=>"011110010",
  37842=>"000110010",
  37843=>"010101101",
  37844=>"000000010",
  37845=>"111010010",
  37846=>"010111011",
  37847=>"110000100",
  37848=>"001000000",
  37849=>"111000010",
  37850=>"101100111",
  37851=>"001010110",
  37852=>"010010110",
  37853=>"000010010",
  37854=>"111010000",
  37855=>"100100001",
  37856=>"101101111",
  37857=>"010011001",
  37858=>"011110110",
  37859=>"010100110",
  37860=>"010100100",
  37861=>"010001111",
  37862=>"110100111",
  37863=>"000110001",
  37864=>"001000111",
  37865=>"000010100",
  37866=>"101000011",
  37867=>"110100000",
  37868=>"100011110",
  37869=>"001100011",
  37870=>"001000010",
  37871=>"111011010",
  37872=>"000000001",
  37873=>"000000101",
  37874=>"101111100",
  37875=>"101110001",
  37876=>"101011110",
  37877=>"001000101",
  37878=>"111100001",
  37879=>"101010101",
  37880=>"101011110",
  37881=>"110101110",
  37882=>"100111101",
  37883=>"110110111",
  37884=>"000001100",
  37885=>"011110110",
  37886=>"100001011",
  37887=>"100011000",
  37888=>"110101110",
  37889=>"101100100",
  37890=>"100011010",
  37891=>"001010011",
  37892=>"000111110",
  37893=>"111001010",
  37894=>"110011111",
  37895=>"000100000",
  37896=>"000001100",
  37897=>"111010001",
  37898=>"011100000",
  37899=>"111110110",
  37900=>"001001001",
  37901=>"101111111",
  37902=>"110101010",
  37903=>"011100110",
  37904=>"101110111",
  37905=>"110100100",
  37906=>"110111100",
  37907=>"111001011",
  37908=>"000000101",
  37909=>"111100101",
  37910=>"110110000",
  37911=>"000000111",
  37912=>"001101010",
  37913=>"110100001",
  37914=>"011000110",
  37915=>"000100110",
  37916=>"111010101",
  37917=>"100111101",
  37918=>"111011010",
  37919=>"100001100",
  37920=>"000001011",
  37921=>"111100001",
  37922=>"011001010",
  37923=>"010011100",
  37924=>"100011110",
  37925=>"011001100",
  37926=>"110100010",
  37927=>"100110000",
  37928=>"001101001",
  37929=>"001010100",
  37930=>"101110010",
  37931=>"010010000",
  37932=>"101111101",
  37933=>"011010010",
  37934=>"011011101",
  37935=>"111010100",
  37936=>"110000011",
  37937=>"111100111",
  37938=>"110011110",
  37939=>"010001011",
  37940=>"010000100",
  37941=>"101111110",
  37942=>"110000000",
  37943=>"000111010",
  37944=>"000100100",
  37945=>"111011111",
  37946=>"000000001",
  37947=>"011000000",
  37948=>"110111110",
  37949=>"001110010",
  37950=>"011100011",
  37951=>"111001100",
  37952=>"011001001",
  37953=>"100000100",
  37954=>"011110111",
  37955=>"001011001",
  37956=>"010100101",
  37957=>"001111011",
  37958=>"100011001",
  37959=>"000011000",
  37960=>"100011010",
  37961=>"001010100",
  37962=>"110001011",
  37963=>"000011100",
  37964=>"000100010",
  37965=>"111101010",
  37966=>"011111001",
  37967=>"111011000",
  37968=>"110011001",
  37969=>"010011011",
  37970=>"101010100",
  37971=>"101101110",
  37972=>"001001000",
  37973=>"000000000",
  37974=>"100001110",
  37975=>"011111111",
  37976=>"000111011",
  37977=>"010111111",
  37978=>"111101010",
  37979=>"001011000",
  37980=>"000110001",
  37981=>"011010000",
  37982=>"010011000",
  37983=>"100001001",
  37984=>"110000110",
  37985=>"111010000",
  37986=>"100001010",
  37987=>"011001001",
  37988=>"000100011",
  37989=>"010111011",
  37990=>"000010111",
  37991=>"010100111",
  37992=>"110100001",
  37993=>"110011011",
  37994=>"010010101",
  37995=>"100100101",
  37996=>"000111110",
  37997=>"000011000",
  37998=>"111010000",
  37999=>"100001000",
  38000=>"011000000",
  38001=>"010101110",
  38002=>"000111010",
  38003=>"001100011",
  38004=>"011011110",
  38005=>"001011111",
  38006=>"110101010",
  38007=>"101010100",
  38008=>"110111101",
  38009=>"000110010",
  38010=>"100100101",
  38011=>"001111101",
  38012=>"111000010",
  38013=>"010100100",
  38014=>"111111100",
  38015=>"001011101",
  38016=>"000010001",
  38017=>"101001111",
  38018=>"110101101",
  38019=>"001000100",
  38020=>"011100100",
  38021=>"110110110",
  38022=>"001011101",
  38023=>"000001100",
  38024=>"000110101",
  38025=>"100000010",
  38026=>"010011011",
  38027=>"010010100",
  38028=>"111111110",
  38029=>"000001110",
  38030=>"001001011",
  38031=>"001101000",
  38032=>"110001000",
  38033=>"111111100",
  38034=>"101010111",
  38035=>"011111011",
  38036=>"100101101",
  38037=>"011100111",
  38038=>"100110011",
  38039=>"011010100",
  38040=>"110001010",
  38041=>"011010100",
  38042=>"111101110",
  38043=>"111111100",
  38044=>"100011010",
  38045=>"010000011",
  38046=>"001111110",
  38047=>"010101110",
  38048=>"010001110",
  38049=>"011011101",
  38050=>"010011100",
  38051=>"001110100",
  38052=>"111101010",
  38053=>"100011101",
  38054=>"000011000",
  38055=>"010100000",
  38056=>"001000111",
  38057=>"100111101",
  38058=>"000010110",
  38059=>"100011101",
  38060=>"111101011",
  38061=>"011110111",
  38062=>"100011111",
  38063=>"011010101",
  38064=>"110001011",
  38065=>"000100001",
  38066=>"001100010",
  38067=>"100000110",
  38068=>"011010010",
  38069=>"000011000",
  38070=>"111100011",
  38071=>"000011111",
  38072=>"100010101",
  38073=>"000011000",
  38074=>"001001000",
  38075=>"000100001",
  38076=>"101110111",
  38077=>"110100000",
  38078=>"011110100",
  38079=>"001011100",
  38080=>"100111110",
  38081=>"101110000",
  38082=>"000101111",
  38083=>"010111101",
  38084=>"100111000",
  38085=>"110100010",
  38086=>"111100101",
  38087=>"100010110",
  38088=>"100001100",
  38089=>"011000011",
  38090=>"101001101",
  38091=>"101000000",
  38092=>"101100111",
  38093=>"010100100",
  38094=>"001010110",
  38095=>"110010111",
  38096=>"110010010",
  38097=>"100110100",
  38098=>"111111010",
  38099=>"110101011",
  38100=>"000011111",
  38101=>"001011111",
  38102=>"010110101",
  38103=>"100010101",
  38104=>"110110100",
  38105=>"001111000",
  38106=>"101011000",
  38107=>"010010000",
  38108=>"100010111",
  38109=>"000101011",
  38110=>"000011111",
  38111=>"001010001",
  38112=>"101111000",
  38113=>"100100111",
  38114=>"110000100",
  38115=>"110100010",
  38116=>"010011000",
  38117=>"110000110",
  38118=>"000110010",
  38119=>"100100111",
  38120=>"000111011",
  38121=>"000100000",
  38122=>"001111100",
  38123=>"101011011",
  38124=>"100011000",
  38125=>"010100110",
  38126=>"010101011",
  38127=>"110101000",
  38128=>"111110011",
  38129=>"100111101",
  38130=>"101000010",
  38131=>"001010010",
  38132=>"011111101",
  38133=>"001011010",
  38134=>"100010011",
  38135=>"010100001",
  38136=>"010100010",
  38137=>"111110111",
  38138=>"100110101",
  38139=>"101111100",
  38140=>"111001011",
  38141=>"001101000",
  38142=>"010001100",
  38143=>"101110101",
  38144=>"101000100",
  38145=>"001111010",
  38146=>"101000111",
  38147=>"101011100",
  38148=>"010100010",
  38149=>"011110010",
  38150=>"011010110",
  38151=>"110111001",
  38152=>"101101001",
  38153=>"001011011",
  38154=>"111101101",
  38155=>"000010001",
  38156=>"000100001",
  38157=>"101110100",
  38158=>"010100000",
  38159=>"100011100",
  38160=>"100001000",
  38161=>"011101101",
  38162=>"001011110",
  38163=>"000001011",
  38164=>"110011101",
  38165=>"000100011",
  38166=>"001100100",
  38167=>"111110110",
  38168=>"010000011",
  38169=>"111100010",
  38170=>"111101101",
  38171=>"110100010",
  38172=>"110000000",
  38173=>"000011010",
  38174=>"000100001",
  38175=>"100110000",
  38176=>"010010011",
  38177=>"000001101",
  38178=>"101000001",
  38179=>"000001000",
  38180=>"011101110",
  38181=>"011100110",
  38182=>"110100010",
  38183=>"101011011",
  38184=>"010100001",
  38185=>"011111111",
  38186=>"010111100",
  38187=>"100110000",
  38188=>"000010101",
  38189=>"101011100",
  38190=>"000010000",
  38191=>"010101110",
  38192=>"011001101",
  38193=>"000010010",
  38194=>"001010101",
  38195=>"000000000",
  38196=>"010111100",
  38197=>"100010100",
  38198=>"110000111",
  38199=>"111101111",
  38200=>"011111111",
  38201=>"011000101",
  38202=>"000100110",
  38203=>"011000111",
  38204=>"111101011",
  38205=>"101001111",
  38206=>"100110100",
  38207=>"101111111",
  38208=>"010100111",
  38209=>"011000101",
  38210=>"100100100",
  38211=>"111010011",
  38212=>"001110011",
  38213=>"000000111",
  38214=>"110100001",
  38215=>"100001010",
  38216=>"100010101",
  38217=>"110000110",
  38218=>"101001101",
  38219=>"001111011",
  38220=>"111000111",
  38221=>"110001010",
  38222=>"010000101",
  38223=>"101101001",
  38224=>"101000101",
  38225=>"011011111",
  38226=>"010010101",
  38227=>"001011011",
  38228=>"000010101",
  38229=>"011010001",
  38230=>"110000000",
  38231=>"000111010",
  38232=>"011001111",
  38233=>"001111001",
  38234=>"000100100",
  38235=>"110001100",
  38236=>"111001011",
  38237=>"100001010",
  38238=>"111000000",
  38239=>"001011001",
  38240=>"001001010",
  38241=>"000011100",
  38242=>"001011001",
  38243=>"110110000",
  38244=>"111010001",
  38245=>"100100011",
  38246=>"011111111",
  38247=>"011110110",
  38248=>"111111111",
  38249=>"001001001",
  38250=>"100111101",
  38251=>"000010010",
  38252=>"101100010",
  38253=>"011111111",
  38254=>"101001111",
  38255=>"011010101",
  38256=>"110000111",
  38257=>"110000111",
  38258=>"110011110",
  38259=>"111110001",
  38260=>"011010111",
  38261=>"011100110",
  38262=>"001101010",
  38263=>"110001110",
  38264=>"100111101",
  38265=>"100111111",
  38266=>"100101010",
  38267=>"101001000",
  38268=>"101000101",
  38269=>"001110010",
  38270=>"001010010",
  38271=>"000111100",
  38272=>"011001000",
  38273=>"000100110",
  38274=>"100110001",
  38275=>"010001010",
  38276=>"100011110",
  38277=>"101011010",
  38278=>"101001011",
  38279=>"011110100",
  38280=>"001110010",
  38281=>"011000110",
  38282=>"010001011",
  38283=>"011100110",
  38284=>"101000111",
  38285=>"100010001",
  38286=>"000000100",
  38287=>"111111011",
  38288=>"110111101",
  38289=>"000110001",
  38290=>"010101011",
  38291=>"100110001",
  38292=>"001100100",
  38293=>"000110100",
  38294=>"110010100",
  38295=>"100110111",
  38296=>"111100010",
  38297=>"011101010",
  38298=>"100101011",
  38299=>"100001011",
  38300=>"101110110",
  38301=>"011010100",
  38302=>"111000000",
  38303=>"110100001",
  38304=>"011100100",
  38305=>"111111111",
  38306=>"111000011",
  38307=>"011011001",
  38308=>"101111110",
  38309=>"111010111",
  38310=>"111011111",
  38311=>"001001001",
  38312=>"011111010",
  38313=>"001100000",
  38314=>"100000110",
  38315=>"110010001",
  38316=>"001000000",
  38317=>"111111010",
  38318=>"010110000",
  38319=>"000001111",
  38320=>"001111010",
  38321=>"010110111",
  38322=>"100110011",
  38323=>"011111001",
  38324=>"010011100",
  38325=>"111110100",
  38326=>"010001011",
  38327=>"000100111",
  38328=>"111011000",
  38329=>"011001001",
  38330=>"000011000",
  38331=>"111011110",
  38332=>"010101010",
  38333=>"110101100",
  38334=>"010100101",
  38335=>"011010001",
  38336=>"010010100",
  38337=>"001011000",
  38338=>"010110011",
  38339=>"101101110",
  38340=>"100000001",
  38341=>"111011111",
  38342=>"100001110",
  38343=>"001001000",
  38344=>"100000110",
  38345=>"111110000",
  38346=>"111101001",
  38347=>"010001100",
  38348=>"100111110",
  38349=>"101000110",
  38350=>"111110000",
  38351=>"101001001",
  38352=>"110010110",
  38353=>"011110000",
  38354=>"101001011",
  38355=>"110011011",
  38356=>"111010110",
  38357=>"110011100",
  38358=>"101101111",
  38359=>"110000010",
  38360=>"111101110",
  38361=>"100010001",
  38362=>"110100010",
  38363=>"010100111",
  38364=>"010110110",
  38365=>"010010001",
  38366=>"001111001",
  38367=>"101011100",
  38368=>"010010111",
  38369=>"000111111",
  38370=>"010011110",
  38371=>"111010001",
  38372=>"001001001",
  38373=>"010000000",
  38374=>"100110111",
  38375=>"100100001",
  38376=>"111001001",
  38377=>"000000100",
  38378=>"110100101",
  38379=>"000010101",
  38380=>"101100001",
  38381=>"011110000",
  38382=>"000001111",
  38383=>"011110000",
  38384=>"101010010",
  38385=>"111101011",
  38386=>"000101110",
  38387=>"101001001",
  38388=>"000000100",
  38389=>"000101111",
  38390=>"011101000",
  38391=>"000101000",
  38392=>"010100110",
  38393=>"011100010",
  38394=>"011011110",
  38395=>"110100001",
  38396=>"010100010",
  38397=>"001111100",
  38398=>"010111000",
  38399=>"001110000",
  38400=>"010101010",
  38401=>"100010011",
  38402=>"010010110",
  38403=>"001101011",
  38404=>"001010110",
  38405=>"001100110",
  38406=>"010100011",
  38407=>"101100010",
  38408=>"110110001",
  38409=>"000000110",
  38410=>"110111001",
  38411=>"111100011",
  38412=>"000011101",
  38413=>"111111000",
  38414=>"100100101",
  38415=>"101101000",
  38416=>"111101010",
  38417=>"011010001",
  38418=>"001011110",
  38419=>"111010101",
  38420=>"010110100",
  38421=>"001111111",
  38422=>"010010111",
  38423=>"010001101",
  38424=>"001011100",
  38425=>"100000111",
  38426=>"111011101",
  38427=>"110000101",
  38428=>"100011111",
  38429=>"100100010",
  38430=>"100110110",
  38431=>"111101110",
  38432=>"010110000",
  38433=>"110101010",
  38434=>"000111000",
  38435=>"101001000",
  38436=>"111000000",
  38437=>"100110010",
  38438=>"011011001",
  38439=>"101001100",
  38440=>"100000000",
  38441=>"100011111",
  38442=>"011010010",
  38443=>"101100111",
  38444=>"111010011",
  38445=>"001111110",
  38446=>"011101000",
  38447=>"001111110",
  38448=>"000001101",
  38449=>"001001010",
  38450=>"011001111",
  38451=>"111011001",
  38452=>"010000010",
  38453=>"110011001",
  38454=>"001111111",
  38455=>"001011001",
  38456=>"001100100",
  38457=>"110110101",
  38458=>"011100101",
  38459=>"011000010",
  38460=>"111111111",
  38461=>"000000100",
  38462=>"101111101",
  38463=>"100000000",
  38464=>"110001101",
  38465=>"000111010",
  38466=>"100000101",
  38467=>"000110100",
  38468=>"100000110",
  38469=>"001100010",
  38470=>"010011100",
  38471=>"101101010",
  38472=>"111000111",
  38473=>"110110001",
  38474=>"110011101",
  38475=>"110110110",
  38476=>"011101000",
  38477=>"010000010",
  38478=>"111101000",
  38479=>"011010001",
  38480=>"100000011",
  38481=>"100010000",
  38482=>"100000010",
  38483=>"110111011",
  38484=>"010000100",
  38485=>"111010010",
  38486=>"000010111",
  38487=>"011000000",
  38488=>"111111010",
  38489=>"010110011",
  38490=>"001000000",
  38491=>"001000111",
  38492=>"011100100",
  38493=>"101110010",
  38494=>"101000110",
  38495=>"011001110",
  38496=>"000000011",
  38497=>"001101000",
  38498=>"011010110",
  38499=>"010111101",
  38500=>"001001101",
  38501=>"100011001",
  38502=>"010100110",
  38503=>"000111010",
  38504=>"010001000",
  38505=>"011100001",
  38506=>"101111100",
  38507=>"110101010",
  38508=>"001101101",
  38509=>"001111010",
  38510=>"111001001",
  38511=>"001111000",
  38512=>"110011001",
  38513=>"111000100",
  38514=>"010011101",
  38515=>"100101110",
  38516=>"011010110",
  38517=>"101000001",
  38518=>"000110010",
  38519=>"101010100",
  38520=>"101001101",
  38521=>"010010010",
  38522=>"011110111",
  38523=>"000100111",
  38524=>"001011111",
  38525=>"101111100",
  38526=>"100100000",
  38527=>"111000110",
  38528=>"110101001",
  38529=>"110011010",
  38530=>"110100101",
  38531=>"001110011",
  38532=>"011010100",
  38533=>"001000001",
  38534=>"100010100",
  38535=>"101011110",
  38536=>"010011010",
  38537=>"000000111",
  38538=>"000000111",
  38539=>"001010101",
  38540=>"101111011",
  38541=>"100111100",
  38542=>"111110001",
  38543=>"101110110",
  38544=>"001110001",
  38545=>"100001111",
  38546=>"000000111",
  38547=>"000010101",
  38548=>"010110010",
  38549=>"000110110",
  38550=>"010110111",
  38551=>"000001000",
  38552=>"110111100",
  38553=>"000111100",
  38554=>"000000000",
  38555=>"011100001",
  38556=>"000000101",
  38557=>"100100101",
  38558=>"110111010",
  38559=>"110000011",
  38560=>"000010010",
  38561=>"111101111",
  38562=>"101111010",
  38563=>"000000110",
  38564=>"101110000",
  38565=>"000011100",
  38566=>"100010001",
  38567=>"110100100",
  38568=>"110000100",
  38569=>"000111110",
  38570=>"010100001",
  38571=>"101101011",
  38572=>"100110000",
  38573=>"101011100",
  38574=>"001110100",
  38575=>"111000111",
  38576=>"100011100",
  38577=>"110101111",
  38578=>"010000010",
  38579=>"000100100",
  38580=>"000010110",
  38581=>"110111011",
  38582=>"001001110",
  38583=>"011001110",
  38584=>"111100100",
  38585=>"101100010",
  38586=>"001011101",
  38587=>"111100001",
  38588=>"101101110",
  38589=>"101000111",
  38590=>"110101010",
  38591=>"101000000",
  38592=>"101011110",
  38593=>"011010000",
  38594=>"100010111",
  38595=>"111111111",
  38596=>"111111000",
  38597=>"000100100",
  38598=>"000100111",
  38599=>"111001011",
  38600=>"101011010",
  38601=>"100011011",
  38602=>"011000000",
  38603=>"110001101",
  38604=>"110111111",
  38605=>"001111110",
  38606=>"000010101",
  38607=>"000100001",
  38608=>"011111010",
  38609=>"000000110",
  38610=>"111011010",
  38611=>"110011000",
  38612=>"111010101",
  38613=>"011110001",
  38614=>"010100110",
  38615=>"011110100",
  38616=>"010100011",
  38617=>"001000111",
  38618=>"110010111",
  38619=>"101001001",
  38620=>"000011111",
  38621=>"101000000",
  38622=>"110010010",
  38623=>"000011000",
  38624=>"001011110",
  38625=>"000111101",
  38626=>"010001001",
  38627=>"111111110",
  38628=>"111100110",
  38629=>"100010110",
  38630=>"100000001",
  38631=>"010100010",
  38632=>"001110010",
  38633=>"110110001",
  38634=>"101010100",
  38635=>"100100010",
  38636=>"101111100",
  38637=>"010001110",
  38638=>"000111111",
  38639=>"001001000",
  38640=>"101001110",
  38641=>"001011001",
  38642=>"010100111",
  38643=>"111111110",
  38644=>"001000111",
  38645=>"100001000",
  38646=>"111101000",
  38647=>"000011100",
  38648=>"101111111",
  38649=>"100101010",
  38650=>"001101101",
  38651=>"001000000",
  38652=>"100111100",
  38653=>"110000111",
  38654=>"110001111",
  38655=>"011110111",
  38656=>"100101101",
  38657=>"101000000",
  38658=>"001110100",
  38659=>"110001100",
  38660=>"110111001",
  38661=>"011111010",
  38662=>"110010101",
  38663=>"111101011",
  38664=>"001011001",
  38665=>"110011010",
  38666=>"111100101",
  38667=>"001101100",
  38668=>"011110001",
  38669=>"111000100",
  38670=>"011100001",
  38671=>"010100000",
  38672=>"100101000",
  38673=>"110111111",
  38674=>"101001011",
  38675=>"100110100",
  38676=>"010000110",
  38677=>"000010000",
  38678=>"110101111",
  38679=>"010001111",
  38680=>"001000000",
  38681=>"100011110",
  38682=>"010011100",
  38683=>"011010111",
  38684=>"000011001",
  38685=>"000110101",
  38686=>"101011111",
  38687=>"110010010",
  38688=>"101011101",
  38689=>"111001001",
  38690=>"000101110",
  38691=>"000111010",
  38692=>"101011100",
  38693=>"100000100",
  38694=>"100000100",
  38695=>"001000110",
  38696=>"110100000",
  38697=>"110110100",
  38698=>"010010001",
  38699=>"100101110",
  38700=>"101100110",
  38701=>"000000111",
  38702=>"000110010",
  38703=>"010001111",
  38704=>"001011100",
  38705=>"110010100",
  38706=>"010111001",
  38707=>"100111011",
  38708=>"101001001",
  38709=>"100001001",
  38710=>"101101010",
  38711=>"100111001",
  38712=>"000100101",
  38713=>"001000100",
  38714=>"100001010",
  38715=>"000101011",
  38716=>"110001001",
  38717=>"011100011",
  38718=>"010101000",
  38719=>"000111001",
  38720=>"100011010",
  38721=>"010100110",
  38722=>"010011010",
  38723=>"010111001",
  38724=>"100010010",
  38725=>"101110010",
  38726=>"101001101",
  38727=>"000001011",
  38728=>"000011110",
  38729=>"000111010",
  38730=>"001010101",
  38731=>"011100000",
  38732=>"011101011",
  38733=>"001110110",
  38734=>"100110000",
  38735=>"010010010",
  38736=>"111101010",
  38737=>"000001110",
  38738=>"000110000",
  38739=>"111001101",
  38740=>"001011001",
  38741=>"110001111",
  38742=>"100110100",
  38743=>"010011100",
  38744=>"110011110",
  38745=>"101011011",
  38746=>"001111111",
  38747=>"111000011",
  38748=>"000010001",
  38749=>"011110111",
  38750=>"001100101",
  38751=>"100010000",
  38752=>"101100010",
  38753=>"111010111",
  38754=>"011010100",
  38755=>"010110101",
  38756=>"010101000",
  38757=>"110110011",
  38758=>"101111000",
  38759=>"001101011",
  38760=>"000100110",
  38761=>"100101001",
  38762=>"000010101",
  38763=>"010101000",
  38764=>"110110000",
  38765=>"001001100",
  38766=>"011111100",
  38767=>"010100100",
  38768=>"001011001",
  38769=>"101000001",
  38770=>"000010001",
  38771=>"011010000",
  38772=>"101101000",
  38773=>"011011010",
  38774=>"110100111",
  38775=>"110000101",
  38776=>"010111110",
  38777=>"000111010",
  38778=>"010111011",
  38779=>"101110100",
  38780=>"010100100",
  38781=>"101001000",
  38782=>"001111101",
  38783=>"000110111",
  38784=>"111001011",
  38785=>"111100011",
  38786=>"011111100",
  38787=>"101000100",
  38788=>"010101111",
  38789=>"111100011",
  38790=>"111000000",
  38791=>"001000001",
  38792=>"110110010",
  38793=>"111011011",
  38794=>"110111101",
  38795=>"100010001",
  38796=>"010101100",
  38797=>"011111001",
  38798=>"110110110",
  38799=>"101101101",
  38800=>"111010010",
  38801=>"100100111",
  38802=>"110010111",
  38803=>"001100110",
  38804=>"001001111",
  38805=>"111001111",
  38806=>"000011110",
  38807=>"010001000",
  38808=>"111110001",
  38809=>"010101100",
  38810=>"101101111",
  38811=>"110100101",
  38812=>"111111001",
  38813=>"000110100",
  38814=>"101100101",
  38815=>"111010000",
  38816=>"011111101",
  38817=>"100010001",
  38818=>"011010000",
  38819=>"111110111",
  38820=>"000100000",
  38821=>"100010000",
  38822=>"111100011",
  38823=>"000001100",
  38824=>"000001101",
  38825=>"001010101",
  38826=>"100111010",
  38827=>"001010110",
  38828=>"001000011",
  38829=>"110011100",
  38830=>"011110111",
  38831=>"000111000",
  38832=>"000011000",
  38833=>"111101110",
  38834=>"100001001",
  38835=>"011110100",
  38836=>"110101110",
  38837=>"001100111",
  38838=>"110110000",
  38839=>"100111011",
  38840=>"011011010",
  38841=>"001001010",
  38842=>"101010111",
  38843=>"011100001",
  38844=>"000011000",
  38845=>"001001011",
  38846=>"000010100",
  38847=>"110101011",
  38848=>"001000111",
  38849=>"100101010",
  38850=>"101111100",
  38851=>"111011110",
  38852=>"111101000",
  38853=>"100010111",
  38854=>"110101001",
  38855=>"010110011",
  38856=>"111100100",
  38857=>"001010001",
  38858=>"010100010",
  38859=>"011100001",
  38860=>"010000000",
  38861=>"110000110",
  38862=>"111101111",
  38863=>"101011101",
  38864=>"100101011",
  38865=>"011001111",
  38866=>"001001000",
  38867=>"110100100",
  38868=>"101100001",
  38869=>"000100011",
  38870=>"100000011",
  38871=>"010000101",
  38872=>"000111001",
  38873=>"111011111",
  38874=>"111010011",
  38875=>"111110011",
  38876=>"011100001",
  38877=>"010100110",
  38878=>"000101001",
  38879=>"111111010",
  38880=>"010010011",
  38881=>"101001000",
  38882=>"010011101",
  38883=>"001001100",
  38884=>"100010101",
  38885=>"001111110",
  38886=>"101111111",
  38887=>"110100010",
  38888=>"110011110",
  38889=>"011110011",
  38890=>"011000101",
  38891=>"100011001",
  38892=>"000001001",
  38893=>"011111101",
  38894=>"110001111",
  38895=>"101101110",
  38896=>"111010010",
  38897=>"110101110",
  38898=>"110010001",
  38899=>"000000000",
  38900=>"010101100",
  38901=>"100010101",
  38902=>"010111000",
  38903=>"101111101",
  38904=>"000100101",
  38905=>"010000010",
  38906=>"000010010",
  38907=>"110100010",
  38908=>"001001011",
  38909=>"101001011",
  38910=>"100100000",
  38911=>"100000101",
  38912=>"100100000",
  38913=>"011000000",
  38914=>"110100100",
  38915=>"101010111",
  38916=>"111100110",
  38917=>"000110010",
  38918=>"111001000",
  38919=>"011111100",
  38920=>"001011100",
  38921=>"100111001",
  38922=>"100110011",
  38923=>"110110001",
  38924=>"111000101",
  38925=>"011010001",
  38926=>"011010011",
  38927=>"110111111",
  38928=>"100100000",
  38929=>"101111010",
  38930=>"111101110",
  38931=>"111001000",
  38932=>"010010000",
  38933=>"111100001",
  38934=>"011010011",
  38935=>"000001010",
  38936=>"111111101",
  38937=>"001011110",
  38938=>"101100100",
  38939=>"111010111",
  38940=>"010010010",
  38941=>"110110000",
  38942=>"101101100",
  38943=>"000001000",
  38944=>"011100111",
  38945=>"000101111",
  38946=>"101110101",
  38947=>"101010101",
  38948=>"101100110",
  38949=>"001100101",
  38950=>"101010001",
  38951=>"110010111",
  38952=>"100011111",
  38953=>"001011001",
  38954=>"001011001",
  38955=>"100001100",
  38956=>"001001101",
  38957=>"101010010",
  38958=>"000111111",
  38959=>"001101010",
  38960=>"010111100",
  38961=>"000000101",
  38962=>"011101110",
  38963=>"100100000",
  38964=>"110010000",
  38965=>"010010010",
  38966=>"000100011",
  38967=>"100111111",
  38968=>"001000010",
  38969=>"100011110",
  38970=>"000010011",
  38971=>"001111101",
  38972=>"010100000",
  38973=>"000001111",
  38974=>"110010010",
  38975=>"000110101",
  38976=>"010110011",
  38977=>"010101110",
  38978=>"000000101",
  38979=>"100000000",
  38980=>"111011001",
  38981=>"000101111",
  38982=>"101101110",
  38983=>"101111001",
  38984=>"110010111",
  38985=>"100111011",
  38986=>"011101101",
  38987=>"001111110",
  38988=>"001000011",
  38989=>"011100111",
  38990=>"001110101",
  38991=>"101110110",
  38992=>"101101101",
  38993=>"111110101",
  38994=>"010000001",
  38995=>"001011111",
  38996=>"000101010",
  38997=>"101011001",
  38998=>"101100000",
  38999=>"001001001",
  39000=>"010110011",
  39001=>"010001010",
  39002=>"101100101",
  39003=>"100010001",
  39004=>"011001011",
  39005=>"100111111",
  39006=>"100010000",
  39007=>"001000101",
  39008=>"011011100",
  39009=>"100101100",
  39010=>"011000001",
  39011=>"010000101",
  39012=>"010100100",
  39013=>"001000001",
  39014=>"100010110",
  39015=>"111001000",
  39016=>"100010001",
  39017=>"110100111",
  39018=>"101111100",
  39019=>"111000111",
  39020=>"000110101",
  39021=>"000110100",
  39022=>"111000101",
  39023=>"111101111",
  39024=>"111011011",
  39025=>"100000101",
  39026=>"101110011",
  39027=>"000110000",
  39028=>"011111011",
  39029=>"110010100",
  39030=>"001010110",
  39031=>"010011111",
  39032=>"010100011",
  39033=>"010111111",
  39034=>"100110011",
  39035=>"011111010",
  39036=>"010001010",
  39037=>"110001010",
  39038=>"011110011",
  39039=>"100100100",
  39040=>"001110000",
  39041=>"110000110",
  39042=>"011010111",
  39043=>"100100001",
  39044=>"110011000",
  39045=>"000010010",
  39046=>"001001011",
  39047=>"011110011",
  39048=>"101000101",
  39049=>"101010100",
  39050=>"100001101",
  39051=>"000010001",
  39052=>"010010111",
  39053=>"010110111",
  39054=>"111010110",
  39055=>"100110100",
  39056=>"000010011",
  39057=>"111000110",
  39058=>"101100001",
  39059=>"100000010",
  39060=>"011110001",
  39061=>"000001001",
  39062=>"001001101",
  39063=>"001011010",
  39064=>"010000011",
  39065=>"001011101",
  39066=>"100111011",
  39067=>"010000010",
  39068=>"101001111",
  39069=>"110000110",
  39070=>"001111000",
  39071=>"011000100",
  39072=>"101110111",
  39073=>"110001111",
  39074=>"101100101",
  39075=>"001011000",
  39076=>"001101000",
  39077=>"011110111",
  39078=>"011011100",
  39079=>"111001011",
  39080=>"101101111",
  39081=>"000001001",
  39082=>"100111101",
  39083=>"101001011",
  39084=>"011110000",
  39085=>"100101011",
  39086=>"100111111",
  39087=>"001011100",
  39088=>"000100011",
  39089=>"010110011",
  39090=>"000001101",
  39091=>"001001101",
  39092=>"011101010",
  39093=>"000010110",
  39094=>"001011000",
  39095=>"001101101",
  39096=>"001110101",
  39097=>"101100001",
  39098=>"010010011",
  39099=>"010011000",
  39100=>"101001011",
  39101=>"010010110",
  39102=>"100111111",
  39103=>"000110110",
  39104=>"000101011",
  39105=>"101101111",
  39106=>"000001010",
  39107=>"011011011",
  39108=>"010101111",
  39109=>"001101001",
  39110=>"001110110",
  39111=>"010110110",
  39112=>"000111111",
  39113=>"000000001",
  39114=>"110100000",
  39115=>"010000000",
  39116=>"001010111",
  39117=>"101111110",
  39118=>"110011000",
  39119=>"101111100",
  39120=>"010010010",
  39121=>"111011001",
  39122=>"100100010",
  39123=>"111110101",
  39124=>"000001000",
  39125=>"010111001",
  39126=>"011111000",
  39127=>"100100010",
  39128=>"101110001",
  39129=>"101110000",
  39130=>"011111010",
  39131=>"111011110",
  39132=>"111011110",
  39133=>"000000010",
  39134=>"101101001",
  39135=>"000100101",
  39136=>"110111101",
  39137=>"111111000",
  39138=>"000111101",
  39139=>"111101011",
  39140=>"100111010",
  39141=>"101011100",
  39142=>"101111110",
  39143=>"010110000",
  39144=>"110011001",
  39145=>"110000010",
  39146=>"001000001",
  39147=>"001101100",
  39148=>"010010110",
  39149=>"100100001",
  39150=>"001011111",
  39151=>"110010000",
  39152=>"110000100",
  39153=>"011101101",
  39154=>"001010010",
  39155=>"000000000",
  39156=>"101000101",
  39157=>"100110010",
  39158=>"010011011",
  39159=>"001001110",
  39160=>"111010100",
  39161=>"000110110",
  39162=>"100011110",
  39163=>"111000101",
  39164=>"000101100",
  39165=>"000111010",
  39166=>"110110111",
  39167=>"001101010",
  39168=>"110100011",
  39169=>"011111000",
  39170=>"001100000",
  39171=>"101001001",
  39172=>"101011010",
  39173=>"011111110",
  39174=>"110111111",
  39175=>"101110001",
  39176=>"101000110",
  39177=>"111001111",
  39178=>"001001111",
  39179=>"011000110",
  39180=>"010011010",
  39181=>"000111011",
  39182=>"000010111",
  39183=>"001001010",
  39184=>"100001000",
  39185=>"011110010",
  39186=>"111110111",
  39187=>"010101010",
  39188=>"010111010",
  39189=>"111100110",
  39190=>"101100010",
  39191=>"100000010",
  39192=>"111011000",
  39193=>"010100000",
  39194=>"100001001",
  39195=>"010000011",
  39196=>"000010110",
  39197=>"000111011",
  39198=>"000111010",
  39199=>"001110111",
  39200=>"111011100",
  39201=>"010011111",
  39202=>"111111100",
  39203=>"100000010",
  39204=>"001110000",
  39205=>"101111010",
  39206=>"101101011",
  39207=>"100001111",
  39208=>"000101110",
  39209=>"000100011",
  39210=>"100010100",
  39211=>"110100010",
  39212=>"110000010",
  39213=>"101011001",
  39214=>"001101001",
  39215=>"000110001",
  39216=>"001111110",
  39217=>"100011001",
  39218=>"111110010",
  39219=>"010000100",
  39220=>"000100011",
  39221=>"010101001",
  39222=>"110100101",
  39223=>"011000010",
  39224=>"100101000",
  39225=>"110111011",
  39226=>"100110101",
  39227=>"010111011",
  39228=>"101101101",
  39229=>"100101100",
  39230=>"111011111",
  39231=>"010100111",
  39232=>"010111000",
  39233=>"100001110",
  39234=>"101101100",
  39235=>"010100001",
  39236=>"100110000",
  39237=>"101001110",
  39238=>"110101011",
  39239=>"010010010",
  39240=>"010111010",
  39241=>"000000110",
  39242=>"001001001",
  39243=>"110111001",
  39244=>"110001011",
  39245=>"010001010",
  39246=>"111010101",
  39247=>"100001101",
  39248=>"010110011",
  39249=>"000100101",
  39250=>"100111111",
  39251=>"100101000",
  39252=>"110101111",
  39253=>"001110111",
  39254=>"111111100",
  39255=>"000101010",
  39256=>"000100110",
  39257=>"101100001",
  39258=>"000011000",
  39259=>"000011000",
  39260=>"101100100",
  39261=>"001010001",
  39262=>"010010000",
  39263=>"011000000",
  39264=>"000000000",
  39265=>"011011001",
  39266=>"011010010",
  39267=>"001110110",
  39268=>"111010101",
  39269=>"101100101",
  39270=>"100111110",
  39271=>"100111101",
  39272=>"001010110",
  39273=>"010111110",
  39274=>"001010110",
  39275=>"000000111",
  39276=>"100001001",
  39277=>"010011001",
  39278=>"110100101",
  39279=>"100011000",
  39280=>"001011000",
  39281=>"001001011",
  39282=>"101000111",
  39283=>"101111100",
  39284=>"000101011",
  39285=>"001110100",
  39286=>"100100100",
  39287=>"110101110",
  39288=>"110110010",
  39289=>"011110110",
  39290=>"011011111",
  39291=>"001100101",
  39292=>"010100010",
  39293=>"000100000",
  39294=>"111110000",
  39295=>"101000101",
  39296=>"000011101",
  39297=>"010110111",
  39298=>"110110101",
  39299=>"001101010",
  39300=>"111111111",
  39301=>"110111111",
  39302=>"000100001",
  39303=>"101111101",
  39304=>"000000011",
  39305=>"011010001",
  39306=>"111010101",
  39307=>"000010010",
  39308=>"101101111",
  39309=>"111000001",
  39310=>"100001000",
  39311=>"010111101",
  39312=>"010010000",
  39313=>"110000011",
  39314=>"000110111",
  39315=>"001011110",
  39316=>"100000110",
  39317=>"100000011",
  39318=>"101111000",
  39319=>"110010101",
  39320=>"111111111",
  39321=>"001010100",
  39322=>"100110101",
  39323=>"111010101",
  39324=>"000011111",
  39325=>"011011001",
  39326=>"111001101",
  39327=>"111110010",
  39328=>"100101101",
  39329=>"101010100",
  39330=>"111011100",
  39331=>"001000000",
  39332=>"110001000",
  39333=>"101010010",
  39334=>"000001001",
  39335=>"011100010",
  39336=>"101011101",
  39337=>"001001101",
  39338=>"001000100",
  39339=>"111101101",
  39340=>"011010100",
  39341=>"010011100",
  39342=>"011111101",
  39343=>"100100101",
  39344=>"100111011",
  39345=>"100101100",
  39346=>"001010000",
  39347=>"001000011",
  39348=>"000010001",
  39349=>"000000110",
  39350=>"111110100",
  39351=>"010010001",
  39352=>"110101011",
  39353=>"010110110",
  39354=>"001011101",
  39355=>"111100001",
  39356=>"011000010",
  39357=>"110110100",
  39358=>"011010101",
  39359=>"000101101",
  39360=>"001010000",
  39361=>"101000100",
  39362=>"101101010",
  39363=>"101101010",
  39364=>"111010110",
  39365=>"010101000",
  39366=>"100000110",
  39367=>"011101100",
  39368=>"001000111",
  39369=>"000100100",
  39370=>"010100101",
  39371=>"000001011",
  39372=>"101111101",
  39373=>"000110100",
  39374=>"100110101",
  39375=>"000000100",
  39376=>"100100101",
  39377=>"110111111",
  39378=>"100001110",
  39379=>"000000101",
  39380=>"011011010",
  39381=>"111110010",
  39382=>"000001110",
  39383=>"000110011",
  39384=>"100010001",
  39385=>"011101011",
  39386=>"010111011",
  39387=>"011010101",
  39388=>"000101010",
  39389=>"000110101",
  39390=>"010110101",
  39391=>"111110110",
  39392=>"000010101",
  39393=>"010001101",
  39394=>"111111101",
  39395=>"100010111",
  39396=>"101111101",
  39397=>"101101111",
  39398=>"010011100",
  39399=>"111110000",
  39400=>"111101101",
  39401=>"111101010",
  39402=>"010110100",
  39403=>"011001101",
  39404=>"010010111",
  39405=>"001111011",
  39406=>"010111010",
  39407=>"110110100",
  39408=>"101010100",
  39409=>"101000010",
  39410=>"001000010",
  39411=>"100000000",
  39412=>"100111100",
  39413=>"010100111",
  39414=>"100100010",
  39415=>"000010010",
  39416=>"101101011",
  39417=>"010110000",
  39418=>"101001111",
  39419=>"111110110",
  39420=>"111100101",
  39421=>"101101101",
  39422=>"101111010",
  39423=>"000011000",
  39424=>"111100100",
  39425=>"101111010",
  39426=>"111010011",
  39427=>"000111001",
  39428=>"111111001",
  39429=>"010111010",
  39430=>"110010110",
  39431=>"010110101",
  39432=>"010011001",
  39433=>"110101110",
  39434=>"010010101",
  39435=>"001000010",
  39436=>"001011110",
  39437=>"000111010",
  39438=>"001101000",
  39439=>"010011001",
  39440=>"010100101",
  39441=>"101010000",
  39442=>"111011100",
  39443=>"011101010",
  39444=>"010111101",
  39445=>"101001111",
  39446=>"111111100",
  39447=>"110110011",
  39448=>"111000110",
  39449=>"011110110",
  39450=>"001101111",
  39451=>"010111110",
  39452=>"011001011",
  39453=>"011100100",
  39454=>"000000101",
  39455=>"000000000",
  39456=>"001010010",
  39457=>"011011000",
  39458=>"000000000",
  39459=>"001000111",
  39460=>"110011001",
  39461=>"011001001",
  39462=>"100001000",
  39463=>"010110101",
  39464=>"000101111",
  39465=>"111110001",
  39466=>"011000110",
  39467=>"100000101",
  39468=>"000101110",
  39469=>"011010000",
  39470=>"001100111",
  39471=>"010111111",
  39472=>"110010000",
  39473=>"100010100",
  39474=>"000101011",
  39475=>"111000111",
  39476=>"000110111",
  39477=>"101011111",
  39478=>"111001010",
  39479=>"010010111",
  39480=>"100000111",
  39481=>"101110101",
  39482=>"001011001",
  39483=>"011010010",
  39484=>"111100111",
  39485=>"000101111",
  39486=>"000100011",
  39487=>"110000001",
  39488=>"011011010",
  39489=>"010100011",
  39490=>"001100000",
  39491=>"100110011",
  39492=>"000100100",
  39493=>"011001111",
  39494=>"000000111",
  39495=>"000111100",
  39496=>"101100100",
  39497=>"000011001",
  39498=>"101001111",
  39499=>"111111001",
  39500=>"000010110",
  39501=>"100000110",
  39502=>"110010110",
  39503=>"001000000",
  39504=>"101111011",
  39505=>"001010110",
  39506=>"101001001",
  39507=>"010011001",
  39508=>"110101001",
  39509=>"000000010",
  39510=>"111000000",
  39511=>"001110100",
  39512=>"111001010",
  39513=>"001011100",
  39514=>"000001001",
  39515=>"000111000",
  39516=>"111000000",
  39517=>"100100001",
  39518=>"000010010",
  39519=>"001100101",
  39520=>"111000000",
  39521=>"011001000",
  39522=>"010100011",
  39523=>"101000001",
  39524=>"011101101",
  39525=>"000100000",
  39526=>"111010010",
  39527=>"000000000",
  39528=>"000100000",
  39529=>"011101110",
  39530=>"111010110",
  39531=>"101111010",
  39532=>"111100010",
  39533=>"100001111",
  39534=>"010011100",
  39535=>"010000110",
  39536=>"010010101",
  39537=>"001100010",
  39538=>"110011001",
  39539=>"000001000",
  39540=>"111111001",
  39541=>"000001001",
  39542=>"110000100",
  39543=>"101011100",
  39544=>"110000101",
  39545=>"110111111",
  39546=>"000001000",
  39547=>"000000111",
  39548=>"110000010",
  39549=>"010001110",
  39550=>"101100101",
  39551=>"001001101",
  39552=>"011101101",
  39553=>"101011100",
  39554=>"001011101",
  39555=>"011000001",
  39556=>"101001000",
  39557=>"101101000",
  39558=>"000010000",
  39559=>"101010010",
  39560=>"010000101",
  39561=>"001110110",
  39562=>"010110010",
  39563=>"010010100",
  39564=>"000010101",
  39565=>"001000010",
  39566=>"111001011",
  39567=>"000110100",
  39568=>"111111000",
  39569=>"100010000",
  39570=>"110111100",
  39571=>"110110010",
  39572=>"010110100",
  39573=>"000111100",
  39574=>"010010100",
  39575=>"111011011",
  39576=>"111011101",
  39577=>"010101101",
  39578=>"000001001",
  39579=>"110011011",
  39580=>"011101111",
  39581=>"111100110",
  39582=>"111111110",
  39583=>"100001000",
  39584=>"011111111",
  39585=>"110101010",
  39586=>"000000000",
  39587=>"010010010",
  39588=>"101111110",
  39589=>"101100100",
  39590=>"000000100",
  39591=>"101101101",
  39592=>"101111001",
  39593=>"000000010",
  39594=>"100100100",
  39595=>"100001100",
  39596=>"010011000",
  39597=>"101100100",
  39598=>"001011101",
  39599=>"011101111",
  39600=>"001000001",
  39601=>"011100011",
  39602=>"001111110",
  39603=>"101110001",
  39604=>"000011001",
  39605=>"010111110",
  39606=>"111111111",
  39607=>"100000111",
  39608=>"010010000",
  39609=>"101011100",
  39610=>"110010101",
  39611=>"110101100",
  39612=>"101111111",
  39613=>"111111001",
  39614=>"001101100",
  39615=>"101000101",
  39616=>"101011010",
  39617=>"010000110",
  39618=>"111110011",
  39619=>"111000010",
  39620=>"010101111",
  39621=>"111111010",
  39622=>"011100111",
  39623=>"010000010",
  39624=>"000101100",
  39625=>"011001001",
  39626=>"001100100",
  39627=>"010011000",
  39628=>"100010001",
  39629=>"101100000",
  39630=>"011101110",
  39631=>"111101010",
  39632=>"010000001",
  39633=>"000010011",
  39634=>"000101101",
  39635=>"000001000",
  39636=>"001111011",
  39637=>"000001100",
  39638=>"000101001",
  39639=>"011000101",
  39640=>"000011111",
  39641=>"011001010",
  39642=>"101101101",
  39643=>"000000101",
  39644=>"100000100",
  39645=>"100010100",
  39646=>"011000100",
  39647=>"000000000",
  39648=>"101110110",
  39649=>"011001011",
  39650=>"111100110",
  39651=>"100010010",
  39652=>"110011010",
  39653=>"101110010",
  39654=>"000100100",
  39655=>"011011111",
  39656=>"000010010",
  39657=>"101010001",
  39658=>"000001011",
  39659=>"001100110",
  39660=>"000000100",
  39661=>"000110111",
  39662=>"010001110",
  39663=>"011110111",
  39664=>"011010110",
  39665=>"100010011",
  39666=>"110111000",
  39667=>"101001010",
  39668=>"000001110",
  39669=>"010101010",
  39670=>"101001010",
  39671=>"111010100",
  39672=>"001101001",
  39673=>"110011010",
  39674=>"111010111",
  39675=>"101011100",
  39676=>"001001110",
  39677=>"011111010",
  39678=>"110011011",
  39679=>"110111010",
  39680=>"001010001",
  39681=>"111010111",
  39682=>"000000001",
  39683=>"011000010",
  39684=>"111110001",
  39685=>"010000101",
  39686=>"010110101",
  39687=>"000010101",
  39688=>"010101000",
  39689=>"111000011",
  39690=>"001010110",
  39691=>"111110111",
  39692=>"101010101",
  39693=>"010110001",
  39694=>"111111010",
  39695=>"110010000",
  39696=>"000001001",
  39697=>"100000000",
  39698=>"110000000",
  39699=>"111001101",
  39700=>"110101111",
  39701=>"110111010",
  39702=>"110010110",
  39703=>"000001010",
  39704=>"001001001",
  39705=>"010011011",
  39706=>"001100010",
  39707=>"000000100",
  39708=>"111101100",
  39709=>"000001101",
  39710=>"111111110",
  39711=>"011001111",
  39712=>"001100101",
  39713=>"101000100",
  39714=>"010000011",
  39715=>"101011011",
  39716=>"101010100",
  39717=>"101001000",
  39718=>"001100100",
  39719=>"101011011",
  39720=>"010100010",
  39721=>"010001011",
  39722=>"000111111",
  39723=>"010010010",
  39724=>"110010100",
  39725=>"010001101",
  39726=>"001101010",
  39727=>"000101101",
  39728=>"000101100",
  39729=>"010010100",
  39730=>"000100000",
  39731=>"011000000",
  39732=>"011001000",
  39733=>"100011000",
  39734=>"011110101",
  39735=>"011111101",
  39736=>"010110111",
  39737=>"100100001",
  39738=>"001100000",
  39739=>"010110011",
  39740=>"001001000",
  39741=>"000111111",
  39742=>"100101001",
  39743=>"000010010",
  39744=>"101010101",
  39745=>"111111100",
  39746=>"011100001",
  39747=>"101101010",
  39748=>"011001111",
  39749=>"110011110",
  39750=>"101100101",
  39751=>"100111111",
  39752=>"010011010",
  39753=>"000000101",
  39754=>"010111010",
  39755=>"100001001",
  39756=>"111000010",
  39757=>"000000000",
  39758=>"000100100",
  39759=>"100000000",
  39760=>"111100111",
  39761=>"000100001",
  39762=>"000011100",
  39763=>"000010000",
  39764=>"100011010",
  39765=>"001010001",
  39766=>"000101110",
  39767=>"010000100",
  39768=>"110000111",
  39769=>"000111001",
  39770=>"100000011",
  39771=>"100011011",
  39772=>"111001110",
  39773=>"000000100",
  39774=>"010111000",
  39775=>"101100111",
  39776=>"010001101",
  39777=>"110100100",
  39778=>"011111001",
  39779=>"011111001",
  39780=>"011111001",
  39781=>"111110100",
  39782=>"100110110",
  39783=>"010110110",
  39784=>"000011000",
  39785=>"001101111",
  39786=>"100001001",
  39787=>"011100101",
  39788=>"010000110",
  39789=>"001001001",
  39790=>"000000100",
  39791=>"110101101",
  39792=>"001110011",
  39793=>"000001001",
  39794=>"101101111",
  39795=>"110100111",
  39796=>"001101010",
  39797=>"101111101",
  39798=>"011111111",
  39799=>"000000101",
  39800=>"101111010",
  39801=>"110111001",
  39802=>"101001101",
  39803=>"001110110",
  39804=>"101111111",
  39805=>"111110110",
  39806=>"101000100",
  39807=>"011101101",
  39808=>"100010101",
  39809=>"001101000",
  39810=>"000100001",
  39811=>"111010111",
  39812=>"110100001",
  39813=>"000100000",
  39814=>"100100111",
  39815=>"100001100",
  39816=>"110001111",
  39817=>"001001010",
  39818=>"001100011",
  39819=>"111000000",
  39820=>"001011100",
  39821=>"010011010",
  39822=>"100011100",
  39823=>"000111100",
  39824=>"111100000",
  39825=>"100010010",
  39826=>"100101100",
  39827=>"011111110",
  39828=>"111001001",
  39829=>"100101111",
  39830=>"111101111",
  39831=>"000001010",
  39832=>"011100001",
  39833=>"101001101",
  39834=>"001011111",
  39835=>"110110011",
  39836=>"010000101",
  39837=>"100100001",
  39838=>"000111000",
  39839=>"000010010",
  39840=>"011010011",
  39841=>"100100101",
  39842=>"000010011",
  39843=>"000000110",
  39844=>"000100111",
  39845=>"011100000",
  39846=>"110100111",
  39847=>"111110100",
  39848=>"110010010",
  39849=>"010011000",
  39850=>"111100110",
  39851=>"110010110",
  39852=>"101001101",
  39853=>"111011111",
  39854=>"001010101",
  39855=>"100110101",
  39856=>"100010011",
  39857=>"111111101",
  39858=>"111101101",
  39859=>"111010111",
  39860=>"101110110",
  39861=>"010110111",
  39862=>"101101110",
  39863=>"101001111",
  39864=>"000010101",
  39865=>"110001011",
  39866=>"000111001",
  39867=>"011000001",
  39868=>"001000011",
  39869=>"111101011",
  39870=>"101101110",
  39871=>"000111101",
  39872=>"100101010",
  39873=>"001000001",
  39874=>"111100011",
  39875=>"000101101",
  39876=>"111101100",
  39877=>"100100100",
  39878=>"010010000",
  39879=>"100000000",
  39880=>"011010010",
  39881=>"001110111",
  39882=>"011001001",
  39883=>"101101101",
  39884=>"110000110",
  39885=>"010000100",
  39886=>"001000001",
  39887=>"111010110",
  39888=>"010001000",
  39889=>"110010010",
  39890=>"110110100",
  39891=>"111111111",
  39892=>"101001110",
  39893=>"111011100",
  39894=>"110111100",
  39895=>"010010000",
  39896=>"010010110",
  39897=>"011010110",
  39898=>"000000001",
  39899=>"111011100",
  39900=>"000110011",
  39901=>"100111100",
  39902=>"011011000",
  39903=>"100011100",
  39904=>"110101100",
  39905=>"101101010",
  39906=>"010101110",
  39907=>"011001101",
  39908=>"000101110",
  39909=>"001101000",
  39910=>"001100011",
  39911=>"001111101",
  39912=>"101110101",
  39913=>"000011000",
  39914=>"011001000",
  39915=>"101010101",
  39916=>"011010000",
  39917=>"001011101",
  39918=>"110101101",
  39919=>"110001001",
  39920=>"101111101",
  39921=>"101110111",
  39922=>"001011001",
  39923=>"101101011",
  39924=>"001100000",
  39925=>"001101101",
  39926=>"011110010",
  39927=>"000001011",
  39928=>"100100010",
  39929=>"011000001",
  39930=>"001101110",
  39931=>"000010011",
  39932=>"101111101",
  39933=>"001010001",
  39934=>"101101101",
  39935=>"010110010",
  39936=>"000011011",
  39937=>"010110011",
  39938=>"110111011",
  39939=>"110110011",
  39940=>"011101101",
  39941=>"011110110",
  39942=>"000011100",
  39943=>"111111001",
  39944=>"001100000",
  39945=>"110000010",
  39946=>"001010000",
  39947=>"110011010",
  39948=>"100101100",
  39949=>"011000100",
  39950=>"010010000",
  39951=>"001000010",
  39952=>"010110100",
  39953=>"011001100",
  39954=>"110000110",
  39955=>"011001100",
  39956=>"001001001",
  39957=>"110110111",
  39958=>"010110000",
  39959=>"011111001",
  39960=>"100011010",
  39961=>"100000001",
  39962=>"011111000",
  39963=>"011011000",
  39964=>"001101101",
  39965=>"111101110",
  39966=>"001011110",
  39967=>"101100110",
  39968=>"001000110",
  39969=>"000101110",
  39970=>"010100010",
  39971=>"011000101",
  39972=>"000001100",
  39973=>"110000010",
  39974=>"110001011",
  39975=>"100010101",
  39976=>"110101011",
  39977=>"101111001",
  39978=>"000101000",
  39979=>"010000001",
  39980=>"010010110",
  39981=>"000001011",
  39982=>"001001010",
  39983=>"101010010",
  39984=>"011001001",
  39985=>"011110111",
  39986=>"101111010",
  39987=>"110101101",
  39988=>"110111010",
  39989=>"101011111",
  39990=>"100110100",
  39991=>"100010100",
  39992=>"111111011",
  39993=>"110000110",
  39994=>"011101010",
  39995=>"001001100",
  39996=>"100101101",
  39997=>"011000110",
  39998=>"100000111",
  39999=>"000000011",
  40000=>"011011111",
  40001=>"001001000",
  40002=>"101011000",
  40003=>"100111111",
  40004=>"000000110",
  40005=>"001100110",
  40006=>"000110101",
  40007=>"100101100",
  40008=>"001110101",
  40009=>"100100110",
  40010=>"001011000",
  40011=>"000000000",
  40012=>"101001001",
  40013=>"111000100",
  40014=>"101101011",
  40015=>"101101011",
  40016=>"100111011",
  40017=>"010100000",
  40018=>"100111011",
  40019=>"110100111",
  40020=>"111101110",
  40021=>"101100101",
  40022=>"100011011",
  40023=>"101111001",
  40024=>"101011110",
  40025=>"000111000",
  40026=>"001101110",
  40027=>"111011111",
  40028=>"110011011",
  40029=>"001100001",
  40030=>"110001010",
  40031=>"010110011",
  40032=>"001001000",
  40033=>"000100001",
  40034=>"100000001",
  40035=>"010000001",
  40036=>"111100010",
  40037=>"011110011",
  40038=>"011110001",
  40039=>"100101010",
  40040=>"101001111",
  40041=>"001101011",
  40042=>"101110100",
  40043=>"100100100",
  40044=>"110010110",
  40045=>"000000000",
  40046=>"000001011",
  40047=>"001111011",
  40048=>"101011011",
  40049=>"111001001",
  40050=>"000101101",
  40051=>"000111011",
  40052=>"001001101",
  40053=>"010011111",
  40054=>"001010101",
  40055=>"101111011",
  40056=>"000000110",
  40057=>"001010011",
  40058=>"011001110",
  40059=>"010011100",
  40060=>"110111100",
  40061=>"100111000",
  40062=>"001001100",
  40063=>"011000100",
  40064=>"011111110",
  40065=>"101101110",
  40066=>"000100010",
  40067=>"111101110",
  40068=>"011001100",
  40069=>"011101001",
  40070=>"000100110",
  40071=>"011111101",
  40072=>"111101101",
  40073=>"100111010",
  40074=>"001011001",
  40075=>"001010111",
  40076=>"100111111",
  40077=>"110000010",
  40078=>"100000000",
  40079=>"101110111",
  40080=>"000000000",
  40081=>"100110011",
  40082=>"111000001",
  40083=>"001011011",
  40084=>"100110100",
  40085=>"011110111",
  40086=>"110100000",
  40087=>"101100111",
  40088=>"010010111",
  40089=>"000100110",
  40090=>"010011010",
  40091=>"010110000",
  40092=>"101000000",
  40093=>"100011111",
  40094=>"111100000",
  40095=>"001011111",
  40096=>"001010001",
  40097=>"000010110",
  40098=>"010100000",
  40099=>"001101111",
  40100=>"101010110",
  40101=>"000100010",
  40102=>"101110000",
  40103=>"001011001",
  40104=>"010100100",
  40105=>"001001011",
  40106=>"000110000",
  40107=>"101000001",
  40108=>"000001111",
  40109=>"000111001",
  40110=>"101101110",
  40111=>"010100001",
  40112=>"010100001",
  40113=>"100011110",
  40114=>"101101000",
  40115=>"100000100",
  40116=>"110101100",
  40117=>"001010010",
  40118=>"011010101",
  40119=>"111010101",
  40120=>"001110101",
  40121=>"111000101",
  40122=>"001011011",
  40123=>"110011000",
  40124=>"010001100",
  40125=>"001001011",
  40126=>"011110111",
  40127=>"010001100",
  40128=>"000111010",
  40129=>"110110011",
  40130=>"110100110",
  40131=>"001001110",
  40132=>"111111001",
  40133=>"010000110",
  40134=>"111001110",
  40135=>"101011110",
  40136=>"110010100",
  40137=>"110111101",
  40138=>"101111111",
  40139=>"110100010",
  40140=>"000110110",
  40141=>"100001001",
  40142=>"101111001",
  40143=>"111111101",
  40144=>"001010100",
  40145=>"100000101",
  40146=>"100111110",
  40147=>"001101010",
  40148=>"111101100",
  40149=>"010011011",
  40150=>"110001110",
  40151=>"001111101",
  40152=>"101101100",
  40153=>"111001001",
  40154=>"001011011",
  40155=>"111111110",
  40156=>"001100000",
  40157=>"011101111",
  40158=>"000000000",
  40159=>"011000111",
  40160=>"101001001",
  40161=>"110001110",
  40162=>"011110100",
  40163=>"010110101",
  40164=>"000000111",
  40165=>"000100001",
  40166=>"110011001",
  40167=>"111001001",
  40168=>"010000000",
  40169=>"110101101",
  40170=>"011001111",
  40171=>"100110001",
  40172=>"111110111",
  40173=>"100111000",
  40174=>"001111100",
  40175=>"011101011",
  40176=>"111110100",
  40177=>"110110110",
  40178=>"111010101",
  40179=>"111000000",
  40180=>"011110011",
  40181=>"111100101",
  40182=>"101111010",
  40183=>"101110000",
  40184=>"001010111",
  40185=>"001101110",
  40186=>"010000111",
  40187=>"001010111",
  40188=>"010110011",
  40189=>"100011001",
  40190=>"001101100",
  40191=>"100010000",
  40192=>"001100000",
  40193=>"010110111",
  40194=>"010101110",
  40195=>"101111110",
  40196=>"100010011",
  40197=>"101111101",
  40198=>"010010000",
  40199=>"000001101",
  40200=>"110100101",
  40201=>"011101011",
  40202=>"000110001",
  40203=>"001100111",
  40204=>"011111100",
  40205=>"111001110",
  40206=>"101011101",
  40207=>"000100101",
  40208=>"010010000",
  40209=>"100001100",
  40210=>"000000101",
  40211=>"100100000",
  40212=>"000001111",
  40213=>"000000001",
  40214=>"110010001",
  40215=>"101010000",
  40216=>"011010010",
  40217=>"001001010",
  40218=>"001010110",
  40219=>"100001111",
  40220=>"011100001",
  40221=>"001111000",
  40222=>"100101100",
  40223=>"111001001",
  40224=>"001001110",
  40225=>"000110000",
  40226=>"000111001",
  40227=>"001110001",
  40228=>"011101111",
  40229=>"001111001",
  40230=>"010010110",
  40231=>"011000100",
  40232=>"101000001",
  40233=>"010110110",
  40234=>"011101001",
  40235=>"001011000",
  40236=>"111110110",
  40237=>"000011101",
  40238=>"110011000",
  40239=>"001100001",
  40240=>"100110110",
  40241=>"111100110",
  40242=>"001111001",
  40243=>"000101010",
  40244=>"010100001",
  40245=>"101111000",
  40246=>"110101011",
  40247=>"111100101",
  40248=>"001100011",
  40249=>"100001011",
  40250=>"001011100",
  40251=>"000111101",
  40252=>"101101101",
  40253=>"011101101",
  40254=>"110011111",
  40255=>"000100111",
  40256=>"001011011",
  40257=>"101111000",
  40258=>"110100111",
  40259=>"011111110",
  40260=>"010110010",
  40261=>"010110110",
  40262=>"000111010",
  40263=>"001101101",
  40264=>"010010000",
  40265=>"101000001",
  40266=>"100010101",
  40267=>"111110000",
  40268=>"001111000",
  40269=>"010011111",
  40270=>"110111001",
  40271=>"001110001",
  40272=>"010000001",
  40273=>"111111110",
  40274=>"011001011",
  40275=>"001001001",
  40276=>"101101010",
  40277=>"111001001",
  40278=>"111011110",
  40279=>"100001011",
  40280=>"110010010",
  40281=>"111111111",
  40282=>"011001111",
  40283=>"111111010",
  40284=>"010011101",
  40285=>"010000011",
  40286=>"110100011",
  40287=>"111101000",
  40288=>"100010111",
  40289=>"000010001",
  40290=>"111101001",
  40291=>"100100001",
  40292=>"101001101",
  40293=>"000011100",
  40294=>"110111101",
  40295=>"100110001",
  40296=>"000001010",
  40297=>"011001100",
  40298=>"110111111",
  40299=>"011000101",
  40300=>"000111100",
  40301=>"110100110",
  40302=>"111100000",
  40303=>"011010011",
  40304=>"011101010",
  40305=>"010011100",
  40306=>"111100100",
  40307=>"110111000",
  40308=>"000010011",
  40309=>"010001001",
  40310=>"011010100",
  40311=>"011110101",
  40312=>"011001011",
  40313=>"111100111",
  40314=>"010001101",
  40315=>"111101101",
  40316=>"000100110",
  40317=>"101101010",
  40318=>"110010000",
  40319=>"110111111",
  40320=>"001000011",
  40321=>"101110001",
  40322=>"000101011",
  40323=>"010010100",
  40324=>"000100000",
  40325=>"100111100",
  40326=>"100011011",
  40327=>"101010010",
  40328=>"111101010",
  40329=>"010000001",
  40330=>"011111111",
  40331=>"000011010",
  40332=>"100001100",
  40333=>"111110010",
  40334=>"011110100",
  40335=>"101000000",
  40336=>"011110010",
  40337=>"111101111",
  40338=>"111010010",
  40339=>"001011011",
  40340=>"110100101",
  40341=>"011010010",
  40342=>"001001110",
  40343=>"101111011",
  40344=>"001011111",
  40345=>"010000001",
  40346=>"110100110",
  40347=>"001101111",
  40348=>"001111010",
  40349=>"011010011",
  40350=>"110110110",
  40351=>"111010001",
  40352=>"101011110",
  40353=>"101000101",
  40354=>"010001110",
  40355=>"011110000",
  40356=>"110010101",
  40357=>"111011110",
  40358=>"001011111",
  40359=>"001001001",
  40360=>"111010001",
  40361=>"011000000",
  40362=>"111100000",
  40363=>"010110111",
  40364=>"000100010",
  40365=>"100100101",
  40366=>"111100011",
  40367=>"101010011",
  40368=>"010011011",
  40369=>"110101000",
  40370=>"000010000",
  40371=>"011001001",
  40372=>"000101100",
  40373=>"100011001",
  40374=>"011101100",
  40375=>"100001101",
  40376=>"100101001",
  40377=>"100000010",
  40378=>"010001001",
  40379=>"000001000",
  40380=>"001000110",
  40381=>"010111001",
  40382=>"101010000",
  40383=>"000011111",
  40384=>"110100010",
  40385=>"110111000",
  40386=>"100010011",
  40387=>"010100010",
  40388=>"010010000",
  40389=>"111011011",
  40390=>"111010110",
  40391=>"111100000",
  40392=>"001110101",
  40393=>"010000110",
  40394=>"110000100",
  40395=>"111101011",
  40396=>"001010111",
  40397=>"001100001",
  40398=>"001110011",
  40399=>"010100110",
  40400=>"111100000",
  40401=>"001110101",
  40402=>"010110000",
  40403=>"011101100",
  40404=>"110011110",
  40405=>"101110100",
  40406=>"001010011",
  40407=>"110001001",
  40408=>"101011010",
  40409=>"101100011",
  40410=>"101001001",
  40411=>"010010110",
  40412=>"001110011",
  40413=>"000011100",
  40414=>"101110111",
  40415=>"000000000",
  40416=>"000110000",
  40417=>"101111010",
  40418=>"111010111",
  40419=>"111001101",
  40420=>"101001101",
  40421=>"111000100",
  40422=>"011111000",
  40423=>"001101100",
  40424=>"100111010",
  40425=>"010110010",
  40426=>"010100001",
  40427=>"010111100",
  40428=>"110100000",
  40429=>"001011101",
  40430=>"011011000",
  40431=>"111010110",
  40432=>"110000111",
  40433=>"000011111",
  40434=>"010010010",
  40435=>"001101101",
  40436=>"101100110",
  40437=>"110111100",
  40438=>"100101101",
  40439=>"010010011",
  40440=>"011101100",
  40441=>"111011000",
  40442=>"000010011",
  40443=>"110001011",
  40444=>"100001001",
  40445=>"110101000",
  40446=>"001101001",
  40447=>"111111100",
  40448=>"001010110",
  40449=>"011000010",
  40450=>"001111010",
  40451=>"011011100",
  40452=>"100110111",
  40453=>"110010010",
  40454=>"111000111",
  40455=>"001101110",
  40456=>"001001100",
  40457=>"010000010",
  40458=>"101000110",
  40459=>"011100111",
  40460=>"000001110",
  40461=>"011010010",
  40462=>"111100100",
  40463=>"011110111",
  40464=>"100000111",
  40465=>"101010111",
  40466=>"101001100",
  40467=>"000110111",
  40468=>"111111000",
  40469=>"111010011",
  40470=>"111011011",
  40471=>"101101011",
  40472=>"000110010",
  40473=>"100011001",
  40474=>"100101010",
  40475=>"000100011",
  40476=>"101111101",
  40477=>"101100110",
  40478=>"100111101",
  40479=>"101100110",
  40480=>"010011101",
  40481=>"100011111",
  40482=>"001010000",
  40483=>"100110011",
  40484=>"110010110",
  40485=>"110011100",
  40486=>"011011010",
  40487=>"110001000",
  40488=>"100111111",
  40489=>"110111011",
  40490=>"010011100",
  40491=>"000100110",
  40492=>"111100100",
  40493=>"000110100",
  40494=>"101110000",
  40495=>"100110101",
  40496=>"101000001",
  40497=>"111011110",
  40498=>"101101001",
  40499=>"010110010",
  40500=>"110100100",
  40501=>"000010010",
  40502=>"111000110",
  40503=>"101110011",
  40504=>"100101010",
  40505=>"010111110",
  40506=>"011001111",
  40507=>"111011110",
  40508=>"011101101",
  40509=>"110110101",
  40510=>"100101010",
  40511=>"111101111",
  40512=>"111001101",
  40513=>"111101011",
  40514=>"110110010",
  40515=>"000101110",
  40516=>"100000001",
  40517=>"000100111",
  40518=>"101000000",
  40519=>"111010010",
  40520=>"111110000",
  40521=>"000101011",
  40522=>"010011010",
  40523=>"001001101",
  40524=>"010011101",
  40525=>"000100001",
  40526=>"010000000",
  40527=>"000100011",
  40528=>"101100000",
  40529=>"000000110",
  40530=>"011001110",
  40531=>"001010011",
  40532=>"011100010",
  40533=>"000000100",
  40534=>"100010000",
  40535=>"011101110",
  40536=>"101000000",
  40537=>"111100100",
  40538=>"001110000",
  40539=>"100110010",
  40540=>"101011001",
  40541=>"100110100",
  40542=>"010000100",
  40543=>"010100101",
  40544=>"000111111",
  40545=>"011011000",
  40546=>"010000000",
  40547=>"111110010",
  40548=>"010111101",
  40549=>"011011100",
  40550=>"110011101",
  40551=>"011000101",
  40552=>"110011011",
  40553=>"000011010",
  40554=>"011000111",
  40555=>"011011001",
  40556=>"100110111",
  40557=>"100010010",
  40558=>"011011010",
  40559=>"110111111",
  40560=>"100011100",
  40561=>"000011001",
  40562=>"010010001",
  40563=>"010100110",
  40564=>"100111001",
  40565=>"111010010",
  40566=>"101010101",
  40567=>"101011111",
  40568=>"010111001",
  40569=>"010101000",
  40570=>"111111111",
  40571=>"101101111",
  40572=>"101011000",
  40573=>"000011111",
  40574=>"100101111",
  40575=>"001001001",
  40576=>"111100100",
  40577=>"100001000",
  40578=>"000011101",
  40579=>"101011001",
  40580=>"000011011",
  40581=>"101001000",
  40582=>"100100101",
  40583=>"110100110",
  40584=>"011010011",
  40585=>"100100010",
  40586=>"001011000",
  40587=>"101101111",
  40588=>"000101101",
  40589=>"101101001",
  40590=>"000010011",
  40591=>"011111000",
  40592=>"100010100",
  40593=>"110110000",
  40594=>"001011000",
  40595=>"111001011",
  40596=>"000011011",
  40597=>"010000001",
  40598=>"100001001",
  40599=>"110101100",
  40600=>"001100011",
  40601=>"111000011",
  40602=>"101001001",
  40603=>"111100100",
  40604=>"110111101",
  40605=>"101011100",
  40606=>"110000010",
  40607=>"010111101",
  40608=>"011010110",
  40609=>"110101001",
  40610=>"011110101",
  40611=>"110000011",
  40612=>"001001001",
  40613=>"111111100",
  40614=>"101111101",
  40615=>"001001010",
  40616=>"100000101",
  40617=>"110110100",
  40618=>"000000110",
  40619=>"110100110",
  40620=>"010011010",
  40621=>"101101111",
  40622=>"111100111",
  40623=>"110001001",
  40624=>"010100011",
  40625=>"111111001",
  40626=>"111011011",
  40627=>"011100100",
  40628=>"000000111",
  40629=>"001011100",
  40630=>"010110100",
  40631=>"101001111",
  40632=>"100101101",
  40633=>"000000101",
  40634=>"101110001",
  40635=>"100000110",
  40636=>"101100001",
  40637=>"010000000",
  40638=>"001101101",
  40639=>"010000001",
  40640=>"110001010",
  40641=>"011100011",
  40642=>"111111110",
  40643=>"000011010",
  40644=>"001011101",
  40645=>"001000100",
  40646=>"100110111",
  40647=>"101100111",
  40648=>"000110110",
  40649=>"011110101",
  40650=>"101101000",
  40651=>"001010011",
  40652=>"101000111",
  40653=>"000100011",
  40654=>"001010100",
  40655=>"011010100",
  40656=>"000000010",
  40657=>"100000101",
  40658=>"000111111",
  40659=>"101000001",
  40660=>"110010010",
  40661=>"011000111",
  40662=>"000101000",
  40663=>"111000100",
  40664=>"000111000",
  40665=>"110110111",
  40666=>"001101011",
  40667=>"101101101",
  40668=>"101001000",
  40669=>"110101011",
  40670=>"110011101",
  40671=>"110111111",
  40672=>"011001111",
  40673=>"001111000",
  40674=>"110010100",
  40675=>"111111100",
  40676=>"000010100",
  40677=>"110100011",
  40678=>"000010010",
  40679=>"011010010",
  40680=>"110111100",
  40681=>"111100000",
  40682=>"110001001",
  40683=>"010100000",
  40684=>"110110110",
  40685=>"111011011",
  40686=>"111010111",
  40687=>"011010100",
  40688=>"101001100",
  40689=>"100111001",
  40690=>"010100100",
  40691=>"011011111",
  40692=>"111100000",
  40693=>"100100100",
  40694=>"010001000",
  40695=>"000110111",
  40696=>"011011110",
  40697=>"101011111",
  40698=>"000101101",
  40699=>"100000100",
  40700=>"111010011",
  40701=>"111111100",
  40702=>"010000000",
  40703=>"100100110",
  40704=>"010011000",
  40705=>"111000001",
  40706=>"000110011",
  40707=>"110111110",
  40708=>"110010110",
  40709=>"001000100",
  40710=>"100001000",
  40711=>"010010110",
  40712=>"101110001",
  40713=>"001010101",
  40714=>"011001100",
  40715=>"110011101",
  40716=>"001101111",
  40717=>"000100110",
  40718=>"011111110",
  40719=>"001010110",
  40720=>"100100001",
  40721=>"011001110",
  40722=>"101111110",
  40723=>"111110001",
  40724=>"001011001",
  40725=>"101011001",
  40726=>"010100101",
  40727=>"000111100",
  40728=>"111001101",
  40729=>"110001100",
  40730=>"110101111",
  40731=>"110101000",
  40732=>"101110010",
  40733=>"010110101",
  40734=>"101110110",
  40735=>"101111010",
  40736=>"100001110",
  40737=>"010101001",
  40738=>"001001111",
  40739=>"000100100",
  40740=>"110110001",
  40741=>"100001111",
  40742=>"011000001",
  40743=>"011100000",
  40744=>"101001110",
  40745=>"111100111",
  40746=>"111000001",
  40747=>"000110001",
  40748=>"010011010",
  40749=>"000100001",
  40750=>"101101101",
  40751=>"001110000",
  40752=>"001110000",
  40753=>"010110001",
  40754=>"101011100",
  40755=>"010011100",
  40756=>"101011010",
  40757=>"110001011",
  40758=>"100111011",
  40759=>"111011111",
  40760=>"000010101",
  40761=>"110001010",
  40762=>"100011111",
  40763=>"110111100",
  40764=>"100001000",
  40765=>"111111011",
  40766=>"011110000",
  40767=>"100001001",
  40768=>"000000011",
  40769=>"011101111",
  40770=>"100010100",
  40771=>"011011100",
  40772=>"001111111",
  40773=>"100001111",
  40774=>"001110000",
  40775=>"010111011",
  40776=>"110111100",
  40777=>"111000011",
  40778=>"001111111",
  40779=>"111111011",
  40780=>"100010100",
  40781=>"001110101",
  40782=>"111010100",
  40783=>"001001001",
  40784=>"000100001",
  40785=>"111111110",
  40786=>"011011100",
  40787=>"101010001",
  40788=>"111101110",
  40789=>"010111001",
  40790=>"001010100",
  40791=>"010110000",
  40792=>"011011100",
  40793=>"000011010",
  40794=>"111111000",
  40795=>"000110101",
  40796=>"111000111",
  40797=>"001111010",
  40798=>"110000000",
  40799=>"110000011",
  40800=>"101101011",
  40801=>"100110010",
  40802=>"101101110",
  40803=>"001010110",
  40804=>"100000101",
  40805=>"001111001",
  40806=>"000000011",
  40807=>"010111101",
  40808=>"101100110",
  40809=>"000001111",
  40810=>"011101111",
  40811=>"010010110",
  40812=>"000011110",
  40813=>"001001101",
  40814=>"001000110",
  40815=>"001100100",
  40816=>"100111100",
  40817=>"000000111",
  40818=>"100111101",
  40819=>"100011000",
  40820=>"111001001",
  40821=>"100011110",
  40822=>"000001000",
  40823=>"001101001",
  40824=>"110100010",
  40825=>"011011111",
  40826=>"101101111",
  40827=>"010001100",
  40828=>"010001000",
  40829=>"010000011",
  40830=>"110000011",
  40831=>"011110011",
  40832=>"100011001",
  40833=>"101000111",
  40834=>"011100111",
  40835=>"100011101",
  40836=>"011101010",
  40837=>"100001100",
  40838=>"000110000",
  40839=>"010110001",
  40840=>"111111001",
  40841=>"101001010",
  40842=>"001101010",
  40843=>"000001101",
  40844=>"101101001",
  40845=>"111101100",
  40846=>"001111101",
  40847=>"101000000",
  40848=>"101100101",
  40849=>"111100111",
  40850=>"111100100",
  40851=>"011000001",
  40852=>"111001011",
  40853=>"001100000",
  40854=>"101101011",
  40855=>"110000010",
  40856=>"010011110",
  40857=>"111001110",
  40858=>"001000011",
  40859=>"000100001",
  40860=>"000111101",
  40861=>"011001101",
  40862=>"011001000",
  40863=>"101111011",
  40864=>"101111111",
  40865=>"110111110",
  40866=>"110000110",
  40867=>"001010100",
  40868=>"010001000",
  40869=>"110110010",
  40870=>"000010011",
  40871=>"110111011",
  40872=>"111010101",
  40873=>"111011001",
  40874=>"110111111",
  40875=>"110010111",
  40876=>"010010101",
  40877=>"110101111",
  40878=>"110000001",
  40879=>"001001110",
  40880=>"010110100",
  40881=>"100011100",
  40882=>"100011000",
  40883=>"110110001",
  40884=>"000011101",
  40885=>"111110000",
  40886=>"100110011",
  40887=>"011101011",
  40888=>"111101001",
  40889=>"001110111",
  40890=>"110111011",
  40891=>"000101110",
  40892=>"110001010",
  40893=>"010110000",
  40894=>"100010110",
  40895=>"100010000",
  40896=>"101000000",
  40897=>"000001010",
  40898=>"010101011",
  40899=>"011110011",
  40900=>"101101101",
  40901=>"110100001",
  40902=>"000110100",
  40903=>"001111000",
  40904=>"001000101",
  40905=>"100011110",
  40906=>"000011111",
  40907=>"111101101",
  40908=>"101110101",
  40909=>"111110000",
  40910=>"111111110",
  40911=>"101001111",
  40912=>"010000111",
  40913=>"000101011",
  40914=>"100100100",
  40915=>"100000100",
  40916=>"000000110",
  40917=>"000000010",
  40918=>"111001011",
  40919=>"101011110",
  40920=>"100001011",
  40921=>"101011000",
  40922=>"101100100",
  40923=>"001101010",
  40924=>"100100100",
  40925=>"010001011",
  40926=>"110101100",
  40927=>"000100010",
  40928=>"001100100",
  40929=>"000000000",
  40930=>"010001101",
  40931=>"101110000",
  40932=>"101010111",
  40933=>"111011111",
  40934=>"011100001",
  40935=>"111011110",
  40936=>"011100101",
  40937=>"001000101",
  40938=>"011001000",
  40939=>"011011110",
  40940=>"000110011",
  40941=>"111000001",
  40942=>"110011111",
  40943=>"110001011",
  40944=>"000100100",
  40945=>"001100010",
  40946=>"000100000",
  40947=>"100011101",
  40948=>"000001101",
  40949=>"001110000",
  40950=>"000100110",
  40951=>"101000110",
  40952=>"011001111",
  40953=>"110101011",
  40954=>"111010000",
  40955=>"010011100",
  40956=>"111111100",
  40957=>"011001110",
  40958=>"011100100",
  40959=>"000000011",
  40960=>"010000011",
  40961=>"011111001",
  40962=>"010100111",
  40963=>"101110010",
  40964=>"000001110",
  40965=>"000000010",
  40966=>"110011100",
  40967=>"000111111",
  40968=>"111101000",
  40969=>"000000111",
  40970=>"010011010",
  40971=>"010001001",
  40972=>"001010101",
  40973=>"101110110",
  40974=>"001001000",
  40975=>"000111111",
  40976=>"010110100",
  40977=>"100100111",
  40978=>"000101100",
  40979=>"101000101",
  40980=>"110000001",
  40981=>"110000110",
  40982=>"111011100",
  40983=>"111111111",
  40984=>"111111110",
  40985=>"110010011",
  40986=>"010001101",
  40987=>"000100000",
  40988=>"001010001",
  40989=>"001010011",
  40990=>"110110100",
  40991=>"110011111",
  40992=>"001000100",
  40993=>"111010000",
  40994=>"101100000",
  40995=>"100110010",
  40996=>"101111110",
  40997=>"001010010",
  40998=>"011110111",
  40999=>"010011100",
  41000=>"000001011",
  41001=>"110100110",
  41002=>"101100100",
  41003=>"100110001",
  41004=>"001111001",
  41005=>"101111000",
  41006=>"001010110",
  41007=>"110111011",
  41008=>"111101111",
  41009=>"000000011",
  41010=>"000001001",
  41011=>"010110100",
  41012=>"111111100",
  41013=>"001010000",
  41014=>"001011100",
  41015=>"100100110",
  41016=>"101110100",
  41017=>"100011010",
  41018=>"001011011",
  41019=>"111111001",
  41020=>"111110101",
  41021=>"011011101",
  41022=>"101011000",
  41023=>"111101111",
  41024=>"010101101",
  41025=>"000000110",
  41026=>"110010011",
  41027=>"100100101",
  41028=>"011010000",
  41029=>"100110011",
  41030=>"000111100",
  41031=>"101110011",
  41032=>"110000000",
  41033=>"000010111",
  41034=>"010110001",
  41035=>"100100101",
  41036=>"011010011",
  41037=>"010110011",
  41038=>"000111111",
  41039=>"101000000",
  41040=>"000100101",
  41041=>"000110110",
  41042=>"100011001",
  41043=>"111100100",
  41044=>"110011001",
  41045=>"100111000",
  41046=>"111000011",
  41047=>"010000000",
  41048=>"111101111",
  41049=>"011000000",
  41050=>"110111100",
  41051=>"000001110",
  41052=>"111001100",
  41053=>"100010000",
  41054=>"000011111",
  41055=>"111101000",
  41056=>"001001100",
  41057=>"111110011",
  41058=>"100110111",
  41059=>"011100010",
  41060=>"100011010",
  41061=>"101101111",
  41062=>"110000010",
  41063=>"011111010",
  41064=>"101101101",
  41065=>"111010010",
  41066=>"101101010",
  41067=>"110110001",
  41068=>"011101000",
  41069=>"110100111",
  41070=>"101101011",
  41071=>"010111101",
  41072=>"100011000",
  41073=>"110000000",
  41074=>"101000000",
  41075=>"100110110",
  41076=>"001010000",
  41077=>"100011011",
  41078=>"100000110",
  41079=>"100110110",
  41080=>"100110001",
  41081=>"101110000",
  41082=>"100101101",
  41083=>"010010000",
  41084=>"100010011",
  41085=>"011000111",
  41086=>"011100111",
  41087=>"111100110",
  41088=>"101100111",
  41089=>"000100000",
  41090=>"110100000",
  41091=>"100100111",
  41092=>"000111011",
  41093=>"111011011",
  41094=>"000101000",
  41095=>"000001010",
  41096=>"111111011",
  41097=>"110110100",
  41098=>"010100000",
  41099=>"111001011",
  41100=>"100111111",
  41101=>"000010110",
  41102=>"011001011",
  41103=>"011110100",
  41104=>"101000110",
  41105=>"101001111",
  41106=>"111000010",
  41107=>"110111101",
  41108=>"100000101",
  41109=>"100110000",
  41110=>"011000000",
  41111=>"111011111",
  41112=>"000100100",
  41113=>"011000111",
  41114=>"011100101",
  41115=>"011010010",
  41116=>"111011111",
  41117=>"001111110",
  41118=>"100110010",
  41119=>"101100111",
  41120=>"001000001",
  41121=>"011111101",
  41122=>"010101001",
  41123=>"100111101",
  41124=>"111110011",
  41125=>"000110001",
  41126=>"011011111",
  41127=>"101010110",
  41128=>"011000100",
  41129=>"011010110",
  41130=>"101011010",
  41131=>"110011011",
  41132=>"001111111",
  41133=>"111100110",
  41134=>"000011011",
  41135=>"010001011",
  41136=>"011000011",
  41137=>"001011010",
  41138=>"000100000",
  41139=>"000111000",
  41140=>"100111000",
  41141=>"100010011",
  41142=>"111111010",
  41143=>"001011000",
  41144=>"100000001",
  41145=>"001100011",
  41146=>"000100000",
  41147=>"011110011",
  41148=>"011001101",
  41149=>"011001011",
  41150=>"100000100",
  41151=>"001100001",
  41152=>"010111110",
  41153=>"000010000",
  41154=>"100111100",
  41155=>"011000001",
  41156=>"011001000",
  41157=>"101111110",
  41158=>"000111111",
  41159=>"110101001",
  41160=>"111000001",
  41161=>"001110011",
  41162=>"001000010",
  41163=>"000001010",
  41164=>"010000111",
  41165=>"001001101",
  41166=>"011100110",
  41167=>"101101001",
  41168=>"011010111",
  41169=>"100110000",
  41170=>"101001010",
  41171=>"010101110",
  41172=>"101110011",
  41173=>"000101001",
  41174=>"001000101",
  41175=>"001000010",
  41176=>"111001110",
  41177=>"000101010",
  41178=>"111010010",
  41179=>"100111100",
  41180=>"110010011",
  41181=>"100111100",
  41182=>"100010001",
  41183=>"001010010",
  41184=>"000011110",
  41185=>"010111110",
  41186=>"111111000",
  41187=>"100000110",
  41188=>"000111110",
  41189=>"000001001",
  41190=>"101001111",
  41191=>"000010000",
  41192=>"001010000",
  41193=>"110011000",
  41194=>"111010000",
  41195=>"100111111",
  41196=>"011100001",
  41197=>"111001010",
  41198=>"100111010",
  41199=>"010010000",
  41200=>"111110010",
  41201=>"010110101",
  41202=>"000110010",
  41203=>"001110010",
  41204=>"011111100",
  41205=>"110100000",
  41206=>"001011001",
  41207=>"111111001",
  41208=>"010111110",
  41209=>"010001001",
  41210=>"000110100",
  41211=>"010000011",
  41212=>"011100101",
  41213=>"111111111",
  41214=>"001011000",
  41215=>"111011100",
  41216=>"000100110",
  41217=>"000111010",
  41218=>"000011000",
  41219=>"110001101",
  41220=>"111110001",
  41221=>"011010010",
  41222=>"011101100",
  41223=>"010011111",
  41224=>"000101011",
  41225=>"111111010",
  41226=>"110110010",
  41227=>"001101000",
  41228=>"010101110",
  41229=>"010000100",
  41230=>"110100000",
  41231=>"111110111",
  41232=>"101100011",
  41233=>"000111110",
  41234=>"001111111",
  41235=>"111111001",
  41236=>"100111011",
  41237=>"111101011",
  41238=>"011100011",
  41239=>"100111000",
  41240=>"011101111",
  41241=>"001001100",
  41242=>"001011001",
  41243=>"110001100",
  41244=>"010010101",
  41245=>"001001001",
  41246=>"010110010",
  41247=>"111010001",
  41248=>"010000110",
  41249=>"101101010",
  41250=>"111000100",
  41251=>"100110110",
  41252=>"011111010",
  41253=>"110100010",
  41254=>"111010001",
  41255=>"111111000",
  41256=>"011100011",
  41257=>"000000000",
  41258=>"110100001",
  41259=>"110101011",
  41260=>"111100011",
  41261=>"100010100",
  41262=>"001010011",
  41263=>"100110101",
  41264=>"000110001",
  41265=>"001101101",
  41266=>"111100100",
  41267=>"111011011",
  41268=>"011001110",
  41269=>"001100100",
  41270=>"100100000",
  41271=>"110100110",
  41272=>"100101011",
  41273=>"000100010",
  41274=>"111010101",
  41275=>"110111011",
  41276=>"001000000",
  41277=>"111011110",
  41278=>"001011001",
  41279=>"101000011",
  41280=>"011011110",
  41281=>"011100101",
  41282=>"000001010",
  41283=>"011011110",
  41284=>"010000000",
  41285=>"010001111",
  41286=>"011000101",
  41287=>"011111101",
  41288=>"111001101",
  41289=>"000000110",
  41290=>"011100010",
  41291=>"011100100",
  41292=>"111011110",
  41293=>"111110111",
  41294=>"000001100",
  41295=>"111101101",
  41296=>"011010001",
  41297=>"100000001",
  41298=>"011011101",
  41299=>"010001100",
  41300=>"101001000",
  41301=>"110111111",
  41302=>"011111001",
  41303=>"100011001",
  41304=>"110111111",
  41305=>"100001101",
  41306=>"110110111",
  41307=>"110110100",
  41308=>"111101000",
  41309=>"000011010",
  41310=>"001011101",
  41311=>"000011010",
  41312=>"011001000",
  41313=>"001010011",
  41314=>"100000110",
  41315=>"011111000",
  41316=>"110001010",
  41317=>"010001111",
  41318=>"011100010",
  41319=>"010010110",
  41320=>"010101000",
  41321=>"100001011",
  41322=>"010010100",
  41323=>"100010010",
  41324=>"011000000",
  41325=>"011100001",
  41326=>"100111000",
  41327=>"000111110",
  41328=>"101000101",
  41329=>"010100011",
  41330=>"111100111",
  41331=>"010111000",
  41332=>"001101110",
  41333=>"101001111",
  41334=>"001000000",
  41335=>"010010000",
  41336=>"001010111",
  41337=>"000110101",
  41338=>"010010011",
  41339=>"011001011",
  41340=>"100100000",
  41341=>"110111100",
  41342=>"000000111",
  41343=>"110000000",
  41344=>"001000110",
  41345=>"100011111",
  41346=>"000010111",
  41347=>"111101111",
  41348=>"000101111",
  41349=>"101101110",
  41350=>"000000010",
  41351=>"001000111",
  41352=>"010100110",
  41353=>"001010110",
  41354=>"110001001",
  41355=>"010001001",
  41356=>"000101110",
  41357=>"110101100",
  41358=>"101110110",
  41359=>"110101010",
  41360=>"011000101",
  41361=>"101111001",
  41362=>"100000010",
  41363=>"001001010",
  41364=>"000001100",
  41365=>"001000100",
  41366=>"110000101",
  41367=>"110111100",
  41368=>"110110111",
  41369=>"000010110",
  41370=>"000101011",
  41371=>"010001010",
  41372=>"110010000",
  41373=>"110111011",
  41374=>"011010010",
  41375=>"010111101",
  41376=>"111100100",
  41377=>"101011100",
  41378=>"001011010",
  41379=>"010110000",
  41380=>"111001111",
  41381=>"011110111",
  41382=>"100110101",
  41383=>"110110010",
  41384=>"000011100",
  41385=>"010101100",
  41386=>"000011010",
  41387=>"001110000",
  41388=>"110010110",
  41389=>"000000110",
  41390=>"100001000",
  41391=>"100100110",
  41392=>"111010001",
  41393=>"100010010",
  41394=>"010000111",
  41395=>"001000000",
  41396=>"011011111",
  41397=>"100101110",
  41398=>"011010001",
  41399=>"010101000",
  41400=>"111000000",
  41401=>"010001011",
  41402=>"111001011",
  41403=>"011000011",
  41404=>"011101110",
  41405=>"011100010",
  41406=>"111001100",
  41407=>"011001011",
  41408=>"100010100",
  41409=>"011011001",
  41410=>"000011010",
  41411=>"111100000",
  41412=>"000000111",
  41413=>"000011000",
  41414=>"001000011",
  41415=>"111011111",
  41416=>"011101010",
  41417=>"010000010",
  41418=>"111000000",
  41419=>"000001010",
  41420=>"101101110",
  41421=>"111001111",
  41422=>"000110100",
  41423=>"101000010",
  41424=>"001001101",
  41425=>"000011111",
  41426=>"001110010",
  41427=>"101100100",
  41428=>"001011111",
  41429=>"000100110",
  41430=>"101110110",
  41431=>"110001100",
  41432=>"011100100",
  41433=>"011010000",
  41434=>"001010110",
  41435=>"001111001",
  41436=>"010101111",
  41437=>"111101110",
  41438=>"010101100",
  41439=>"000010100",
  41440=>"001101000",
  41441=>"011101101",
  41442=>"011101110",
  41443=>"111000011",
  41444=>"110001010",
  41445=>"110001010",
  41446=>"100000101",
  41447=>"001000000",
  41448=>"010000000",
  41449=>"011010110",
  41450=>"010011110",
  41451=>"101000110",
  41452=>"101101110",
  41453=>"101110010",
  41454=>"010000110",
  41455=>"011101000",
  41456=>"000111011",
  41457=>"101100100",
  41458=>"100110111",
  41459=>"000110100",
  41460=>"100000000",
  41461=>"011110101",
  41462=>"100010101",
  41463=>"101011001",
  41464=>"001111100",
  41465=>"111100011",
  41466=>"110111111",
  41467=>"100000000",
  41468=>"111111110",
  41469=>"100111001",
  41470=>"010110101",
  41471=>"010100101",
  41472=>"011001000",
  41473=>"001101001",
  41474=>"100101111",
  41475=>"010001110",
  41476=>"101001010",
  41477=>"100100101",
  41478=>"010001000",
  41479=>"010110011",
  41480=>"111111011",
  41481=>"001111111",
  41482=>"110001010",
  41483=>"000000110",
  41484=>"111101010",
  41485=>"011001010",
  41486=>"000110110",
  41487=>"010010010",
  41488=>"101001010",
  41489=>"010000010",
  41490=>"010000100",
  41491=>"100101111",
  41492=>"110110100",
  41493=>"010010000",
  41494=>"001001000",
  41495=>"001010101",
  41496=>"100110100",
  41497=>"001100010",
  41498=>"100100101",
  41499=>"110011000",
  41500=>"111110100",
  41501=>"110000001",
  41502=>"111101111",
  41503=>"101111011",
  41504=>"001101100",
  41505=>"011101011",
  41506=>"000001100",
  41507=>"011101100",
  41508=>"010001010",
  41509=>"101101000",
  41510=>"011000000",
  41511=>"001011001",
  41512=>"000001000",
  41513=>"100000011",
  41514=>"111110001",
  41515=>"101001110",
  41516=>"010111010",
  41517=>"001101111",
  41518=>"111100011",
  41519=>"110000010",
  41520=>"011000000",
  41521=>"001111110",
  41522=>"110101011",
  41523=>"001101011",
  41524=>"010100110",
  41525=>"010110001",
  41526=>"000010001",
  41527=>"100110010",
  41528=>"010001110",
  41529=>"001110001",
  41530=>"100001100",
  41531=>"001001111",
  41532=>"110011110",
  41533=>"101111101",
  41534=>"000110101",
  41535=>"011001111",
  41536=>"000001010",
  41537=>"000011011",
  41538=>"100111101",
  41539=>"010001111",
  41540=>"101000010",
  41541=>"010111110",
  41542=>"101010111",
  41543=>"000000000",
  41544=>"000010111",
  41545=>"010011100",
  41546=>"010001011",
  41547=>"000010010",
  41548=>"001000111",
  41549=>"110011010",
  41550=>"001000000",
  41551=>"011111000",
  41552=>"111000000",
  41553=>"011110011",
  41554=>"110110101",
  41555=>"000111010",
  41556=>"101111100",
  41557=>"110000000",
  41558=>"100110110",
  41559=>"111111101",
  41560=>"011101110",
  41561=>"000010100",
  41562=>"001111110",
  41563=>"000100110",
  41564=>"010000110",
  41565=>"111111101",
  41566=>"010100100",
  41567=>"000110100",
  41568=>"001110100",
  41569=>"010100110",
  41570=>"110010011",
  41571=>"110100111",
  41572=>"000010100",
  41573=>"100100000",
  41574=>"101000010",
  41575=>"010011010",
  41576=>"111101011",
  41577=>"000011001",
  41578=>"001100011",
  41579=>"011000000",
  41580=>"000100111",
  41581=>"011100100",
  41582=>"101010001",
  41583=>"111111100",
  41584=>"101111011",
  41585=>"001110011",
  41586=>"110111001",
  41587=>"000010000",
  41588=>"000111111",
  41589=>"010110001",
  41590=>"001111001",
  41591=>"000001001",
  41592=>"100001000",
  41593=>"000011010",
  41594=>"110101010",
  41595=>"010101110",
  41596=>"101000111",
  41597=>"111110010",
  41598=>"111010001",
  41599=>"001111110",
  41600=>"010001001",
  41601=>"000100001",
  41602=>"111001001",
  41603=>"101001000",
  41604=>"000101001",
  41605=>"010001000",
  41606=>"101111011",
  41607=>"001011111",
  41608=>"000000011",
  41609=>"011101001",
  41610=>"000100111",
  41611=>"001110110",
  41612=>"101011010",
  41613=>"010110011",
  41614=>"110111100",
  41615=>"000100110",
  41616=>"001001111",
  41617=>"010111001",
  41618=>"011010110",
  41619=>"000110001",
  41620=>"000101100",
  41621=>"100001011",
  41622=>"111110011",
  41623=>"101000110",
  41624=>"001000001",
  41625=>"010000000",
  41626=>"101101001",
  41627=>"001100110",
  41628=>"000001100",
  41629=>"101010111",
  41630=>"110101000",
  41631=>"011101010",
  41632=>"111011010",
  41633=>"110011011",
  41634=>"111101101",
  41635=>"101110001",
  41636=>"101011011",
  41637=>"110111011",
  41638=>"101111101",
  41639=>"010010111",
  41640=>"011001010",
  41641=>"000010100",
  41642=>"101000011",
  41643=>"001010001",
  41644=>"111111011",
  41645=>"011100111",
  41646=>"110101011",
  41647=>"111000101",
  41648=>"001100111",
  41649=>"101100110",
  41650=>"100010101",
  41651=>"010011111",
  41652=>"000101101",
  41653=>"101011011",
  41654=>"011110110",
  41655=>"110011110",
  41656=>"101101100",
  41657=>"000010001",
  41658=>"101010000",
  41659=>"011010010",
  41660=>"110001110",
  41661=>"011001001",
  41662=>"000100110",
  41663=>"111001110",
  41664=>"001111000",
  41665=>"101111110",
  41666=>"001010001",
  41667=>"110100010",
  41668=>"000111001",
  41669=>"110010000",
  41670=>"110001110",
  41671=>"001010001",
  41672=>"101111100",
  41673=>"110111101",
  41674=>"111101100",
  41675=>"111111101",
  41676=>"001001110",
  41677=>"111101011",
  41678=>"101001110",
  41679=>"111011010",
  41680=>"011101011",
  41681=>"111001010",
  41682=>"101011000",
  41683=>"000001000",
  41684=>"100100001",
  41685=>"010010010",
  41686=>"111000011",
  41687=>"011111111",
  41688=>"000111100",
  41689=>"101111011",
  41690=>"000110000",
  41691=>"011010010",
  41692=>"000000010",
  41693=>"100010110",
  41694=>"100111111",
  41695=>"100100010",
  41696=>"100110000",
  41697=>"110110101",
  41698=>"101111010",
  41699=>"010110111",
  41700=>"110001011",
  41701=>"011111011",
  41702=>"010011100",
  41703=>"100100101",
  41704=>"100110110",
  41705=>"011010110",
  41706=>"011010111",
  41707=>"001110110",
  41708=>"111010111",
  41709=>"001010100",
  41710=>"011101001",
  41711=>"111001100",
  41712=>"001000111",
  41713=>"011011111",
  41714=>"110011110",
  41715=>"110110010",
  41716=>"111111101",
  41717=>"101001111",
  41718=>"100110111",
  41719=>"101001101",
  41720=>"011101111",
  41721=>"111001100",
  41722=>"111100100",
  41723=>"010111110",
  41724=>"000011100",
  41725=>"110010010",
  41726=>"001010110",
  41727=>"101111001",
  41728=>"101110010",
  41729=>"001100100",
  41730=>"000010110",
  41731=>"011101000",
  41732=>"110100111",
  41733=>"010110110",
  41734=>"001000101",
  41735=>"010100100",
  41736=>"000100101",
  41737=>"011010101",
  41738=>"000000011",
  41739=>"010100111",
  41740=>"011001101",
  41741=>"000110111",
  41742=>"101010011",
  41743=>"101111111",
  41744=>"010011010",
  41745=>"111001111",
  41746=>"000110001",
  41747=>"001110010",
  41748=>"111000111",
  41749=>"000000000",
  41750=>"010110001",
  41751=>"101101111",
  41752=>"001001110",
  41753=>"000111111",
  41754=>"011100001",
  41755=>"010010100",
  41756=>"001011111",
  41757=>"110010010",
  41758=>"000000001",
  41759=>"111100011",
  41760=>"010101101",
  41761=>"010000111",
  41762=>"101111111",
  41763=>"100011100",
  41764=>"101000001",
  41765=>"010111100",
  41766=>"010000111",
  41767=>"110000111",
  41768=>"001101000",
  41769=>"001000111",
  41770=>"111110011",
  41771=>"111111011",
  41772=>"001101000",
  41773=>"110111111",
  41774=>"001111001",
  41775=>"110110101",
  41776=>"111100000",
  41777=>"010110011",
  41778=>"100001100",
  41779=>"101111110",
  41780=>"110010010",
  41781=>"001011100",
  41782=>"111000001",
  41783=>"111110010",
  41784=>"011000011",
  41785=>"101000011",
  41786=>"010101000",
  41787=>"000011010",
  41788=>"010011111",
  41789=>"111001011",
  41790=>"000010001",
  41791=>"011101100",
  41792=>"000100110",
  41793=>"011000001",
  41794=>"111001010",
  41795=>"100100001",
  41796=>"011001001",
  41797=>"001011101",
  41798=>"000000010",
  41799=>"011001101",
  41800=>"111100110",
  41801=>"100011111",
  41802=>"011001111",
  41803=>"000011110",
  41804=>"011000010",
  41805=>"001100101",
  41806=>"010101000",
  41807=>"000000010",
  41808=>"011001010",
  41809=>"110011000",
  41810=>"001000111",
  41811=>"010000000",
  41812=>"000010101",
  41813=>"110011100",
  41814=>"000100110",
  41815=>"101010000",
  41816=>"010010110",
  41817=>"011110100",
  41818=>"100000000",
  41819=>"000110101",
  41820=>"011000010",
  41821=>"010011101",
  41822=>"000000110",
  41823=>"000100110",
  41824=>"100001001",
  41825=>"011001100",
  41826=>"101100000",
  41827=>"011010010",
  41828=>"000010100",
  41829=>"111000001",
  41830=>"101111110",
  41831=>"010110100",
  41832=>"000011010",
  41833=>"101010011",
  41834=>"111010000",
  41835=>"110100010",
  41836=>"000110101",
  41837=>"111101001",
  41838=>"110100111",
  41839=>"011001001",
  41840=>"010010101",
  41841=>"100010111",
  41842=>"000010110",
  41843=>"000000001",
  41844=>"000010001",
  41845=>"111111100",
  41846=>"111010111",
  41847=>"110000110",
  41848=>"100100000",
  41849=>"101111101",
  41850=>"110011010",
  41851=>"101101110",
  41852=>"010111001",
  41853=>"011100001",
  41854=>"011000010",
  41855=>"001001100",
  41856=>"010110010",
  41857=>"011101001",
  41858=>"001100110",
  41859=>"000001011",
  41860=>"010111111",
  41861=>"000001110",
  41862=>"001011100",
  41863=>"101011000",
  41864=>"010110001",
  41865=>"100000111",
  41866=>"100100101",
  41867=>"110100010",
  41868=>"000100000",
  41869=>"100001110",
  41870=>"111101001",
  41871=>"011011010",
  41872=>"110001000",
  41873=>"100000101",
  41874=>"110010101",
  41875=>"111100000",
  41876=>"011001010",
  41877=>"100011100",
  41878=>"000010111",
  41879=>"111110111",
  41880=>"100011000",
  41881=>"010111111",
  41882=>"110010111",
  41883=>"010110001",
  41884=>"000111001",
  41885=>"101000000",
  41886=>"101001001",
  41887=>"111110011",
  41888=>"000110100",
  41889=>"111101100",
  41890=>"110011001",
  41891=>"011001001",
  41892=>"110111011",
  41893=>"100100000",
  41894=>"110100010",
  41895=>"010100101",
  41896=>"100111111",
  41897=>"110110010",
  41898=>"011101110",
  41899=>"111001111",
  41900=>"001110100",
  41901=>"010011000",
  41902=>"000100111",
  41903=>"001100000",
  41904=>"000001111",
  41905=>"110000111",
  41906=>"001001110",
  41907=>"110001101",
  41908=>"000111100",
  41909=>"011100100",
  41910=>"001111101",
  41911=>"010010010",
  41912=>"001011011",
  41913=>"000000010",
  41914=>"110100101",
  41915=>"011110011",
  41916=>"111111100",
  41917=>"000010010",
  41918=>"000000100",
  41919=>"010101000",
  41920=>"101000011",
  41921=>"011111110",
  41922=>"010011010",
  41923=>"001101100",
  41924=>"101100000",
  41925=>"011111111",
  41926=>"101001111",
  41927=>"111100000",
  41928=>"101101110",
  41929=>"100000100",
  41930=>"011000111",
  41931=>"101011110",
  41932=>"100010001",
  41933=>"110001111",
  41934=>"100100000",
  41935=>"111100001",
  41936=>"001111000",
  41937=>"010011001",
  41938=>"101101100",
  41939=>"110010000",
  41940=>"010000000",
  41941=>"011010011",
  41942=>"001010100",
  41943=>"010100000",
  41944=>"010010010",
  41945=>"010100110",
  41946=>"001101111",
  41947=>"111011111",
  41948=>"000110110",
  41949=>"001000110",
  41950=>"001001111",
  41951=>"100001001",
  41952=>"000000000",
  41953=>"100111110",
  41954=>"011001010",
  41955=>"111011001",
  41956=>"000100110",
  41957=>"001011011",
  41958=>"101010101",
  41959=>"110011000",
  41960=>"111110000",
  41961=>"010010010",
  41962=>"001110111",
  41963=>"000111101",
  41964=>"110011011",
  41965=>"000011100",
  41966=>"010000011",
  41967=>"011101101",
  41968=>"011011100",
  41969=>"001100100",
  41970=>"100101111",
  41971=>"001100110",
  41972=>"100010101",
  41973=>"110010101",
  41974=>"000010001",
  41975=>"000111111",
  41976=>"100000110",
  41977=>"011010011",
  41978=>"100100010",
  41979=>"011110000",
  41980=>"000101011",
  41981=>"001001100",
  41982=>"101111100",
  41983=>"100100111",
  41984=>"101001110",
  41985=>"000011010",
  41986=>"101100000",
  41987=>"101111010",
  41988=>"000000000",
  41989=>"011100000",
  41990=>"011111000",
  41991=>"001101100",
  41992=>"000100011",
  41993=>"001101100",
  41994=>"000010011",
  41995=>"111011110",
  41996=>"100110111",
  41997=>"101011101",
  41998=>"100101000",
  41999=>"110000010",
  42000=>"101101111",
  42001=>"000001100",
  42002=>"111000010",
  42003=>"100110001",
  42004=>"001111001",
  42005=>"010010110",
  42006=>"000010011",
  42007=>"110100011",
  42008=>"010110101",
  42009=>"000001101",
  42010=>"110110100",
  42011=>"010011011",
  42012=>"011001110",
  42013=>"111001001",
  42014=>"100100011",
  42015=>"011110101",
  42016=>"011100011",
  42017=>"011111010",
  42018=>"011110100",
  42019=>"000110010",
  42020=>"100010001",
  42021=>"110011101",
  42022=>"000001100",
  42023=>"110000111",
  42024=>"111111110",
  42025=>"100011000",
  42026=>"010111111",
  42027=>"110111011",
  42028=>"110111001",
  42029=>"011010000",
  42030=>"111100101",
  42031=>"101101000",
  42032=>"011110011",
  42033=>"000100111",
  42034=>"111010000",
  42035=>"100001111",
  42036=>"100100000",
  42037=>"010010001",
  42038=>"011010000",
  42039=>"011111110",
  42040=>"000110011",
  42041=>"110010010",
  42042=>"000111100",
  42043=>"000110111",
  42044=>"000000111",
  42045=>"111000000",
  42046=>"111000001",
  42047=>"111101101",
  42048=>"011111100",
  42049=>"000000001",
  42050=>"011110000",
  42051=>"101101001",
  42052=>"110010100",
  42053=>"111010010",
  42054=>"010110101",
  42055=>"001011011",
  42056=>"101001100",
  42057=>"011001100",
  42058=>"011101101",
  42059=>"011011111",
  42060=>"000000010",
  42061=>"000100101",
  42062=>"010101000",
  42063=>"011100011",
  42064=>"000001100",
  42065=>"110111111",
  42066=>"101001000",
  42067=>"010011100",
  42068=>"000111101",
  42069=>"010011010",
  42070=>"010001101",
  42071=>"010000011",
  42072=>"010101000",
  42073=>"111110000",
  42074=>"000110100",
  42075=>"010001001",
  42076=>"000100011",
  42077=>"100101010",
  42078=>"011100001",
  42079=>"001001011",
  42080=>"001001110",
  42081=>"011101111",
  42082=>"100001100",
  42083=>"111101111",
  42084=>"111111011",
  42085=>"000000111",
  42086=>"001000001",
  42087=>"011100110",
  42088=>"001110100",
  42089=>"011010000",
  42090=>"110110111",
  42091=>"000001001",
  42092=>"001100110",
  42093=>"101100010",
  42094=>"110010101",
  42095=>"100111011",
  42096=>"101110111",
  42097=>"001011110",
  42098=>"111100010",
  42099=>"011010111",
  42100=>"000001110",
  42101=>"000101100",
  42102=>"101101110",
  42103=>"010011101",
  42104=>"001100001",
  42105=>"011010011",
  42106=>"101000010",
  42107=>"000100101",
  42108=>"101100110",
  42109=>"110000011",
  42110=>"000000101",
  42111=>"000101111",
  42112=>"000011000",
  42113=>"000010011",
  42114=>"010010010",
  42115=>"111101011",
  42116=>"011001100",
  42117=>"010100101",
  42118=>"111011111",
  42119=>"110110000",
  42120=>"011010110",
  42121=>"111001011",
  42122=>"100001111",
  42123=>"111101001",
  42124=>"111000010",
  42125=>"100001011",
  42126=>"001101010",
  42127=>"100001110",
  42128=>"000001011",
  42129=>"110111000",
  42130=>"000101111",
  42131=>"101010011",
  42132=>"000111111",
  42133=>"000100111",
  42134=>"010010110",
  42135=>"110010010",
  42136=>"000100111",
  42137=>"010100100",
  42138=>"010100101",
  42139=>"111001000",
  42140=>"000101011",
  42141=>"110010001",
  42142=>"011011100",
  42143=>"000111111",
  42144=>"101111110",
  42145=>"111001001",
  42146=>"101010100",
  42147=>"011010001",
  42148=>"110010101",
  42149=>"010110111",
  42150=>"101111100",
  42151=>"100110011",
  42152=>"011010010",
  42153=>"111000011",
  42154=>"110110100",
  42155=>"101110100",
  42156=>"000001111",
  42157=>"100100111",
  42158=>"011010001",
  42159=>"101000110",
  42160=>"001000100",
  42161=>"000100101",
  42162=>"110100011",
  42163=>"100000101",
  42164=>"100000101",
  42165=>"000101011",
  42166=>"001000000",
  42167=>"101100111",
  42168=>"000110001",
  42169=>"010000010",
  42170=>"001110110",
  42171=>"110111110",
  42172=>"011100001",
  42173=>"111001001",
  42174=>"010111111",
  42175=>"001111001",
  42176=>"110111000",
  42177=>"100010101",
  42178=>"111101100",
  42179=>"011100000",
  42180=>"101000111",
  42181=>"100011110",
  42182=>"000110111",
  42183=>"011110100",
  42184=>"111001110",
  42185=>"100111001",
  42186=>"111001111",
  42187=>"101110111",
  42188=>"010110101",
  42189=>"100010110",
  42190=>"000000100",
  42191=>"011101010",
  42192=>"000101111",
  42193=>"001100101",
  42194=>"001000001",
  42195=>"100011101",
  42196=>"100001111",
  42197=>"000000011",
  42198=>"001101001",
  42199=>"100110001",
  42200=>"001000001",
  42201=>"110011111",
  42202=>"110110111",
  42203=>"001000100",
  42204=>"111010110",
  42205=>"110001011",
  42206=>"001011010",
  42207=>"011011000",
  42208=>"001000110",
  42209=>"100111011",
  42210=>"100111111",
  42211=>"011001011",
  42212=>"000010000",
  42213=>"000110111",
  42214=>"101111010",
  42215=>"101010011",
  42216=>"000000010",
  42217=>"111100110",
  42218=>"111011111",
  42219=>"000001001",
  42220=>"011010011",
  42221=>"011011110",
  42222=>"111110010",
  42223=>"111100110",
  42224=>"010001110",
  42225=>"101110110",
  42226=>"111111010",
  42227=>"111111110",
  42228=>"111101111",
  42229=>"111011010",
  42230=>"110001101",
  42231=>"101110100",
  42232=>"000001101",
  42233=>"000100101",
  42234=>"100010100",
  42235=>"001111110",
  42236=>"011011101",
  42237=>"111010011",
  42238=>"110110100",
  42239=>"101111000",
  42240=>"110100110",
  42241=>"100101101",
  42242=>"010011010",
  42243=>"010101100",
  42244=>"110001111",
  42245=>"001011111",
  42246=>"011001110",
  42247=>"110001010",
  42248=>"000001000",
  42249=>"001101001",
  42250=>"001010111",
  42251=>"101110100",
  42252=>"001001001",
  42253=>"110010010",
  42254=>"100110000",
  42255=>"010111001",
  42256=>"001110001",
  42257=>"001100110",
  42258=>"111100010",
  42259=>"110010110",
  42260=>"010001110",
  42261=>"111001011",
  42262=>"111110100",
  42263=>"000000100",
  42264=>"100101110",
  42265=>"001100010",
  42266=>"110000101",
  42267=>"101100000",
  42268=>"011010011",
  42269=>"100100010",
  42270=>"011111110",
  42271=>"110110000",
  42272=>"100011000",
  42273=>"111111001",
  42274=>"100111001",
  42275=>"111001111",
  42276=>"110101111",
  42277=>"010010011",
  42278=>"000100000",
  42279=>"111010100",
  42280=>"010100011",
  42281=>"011011011",
  42282=>"100100010",
  42283=>"101011010",
  42284=>"111100000",
  42285=>"001000100",
  42286=>"001000111",
  42287=>"101101010",
  42288=>"000111011",
  42289=>"011010011",
  42290=>"000001101",
  42291=>"011011011",
  42292=>"110010000",
  42293=>"101100001",
  42294=>"101000100",
  42295=>"101010100",
  42296=>"000001001",
  42297=>"000100110",
  42298=>"010100010",
  42299=>"110111000",
  42300=>"100101001",
  42301=>"110101110",
  42302=>"010001100",
  42303=>"101100000",
  42304=>"000010110",
  42305=>"000110110",
  42306=>"100111110",
  42307=>"110101001",
  42308=>"000001011",
  42309=>"111100000",
  42310=>"101000001",
  42311=>"111010000",
  42312=>"000011100",
  42313=>"100000111",
  42314=>"000001110",
  42315=>"000011111",
  42316=>"111110011",
  42317=>"100010111",
  42318=>"110010101",
  42319=>"011100000",
  42320=>"101110000",
  42321=>"010011011",
  42322=>"100000001",
  42323=>"001001001",
  42324=>"001100100",
  42325=>"010001110",
  42326=>"001110101",
  42327=>"111111001",
  42328=>"111010111",
  42329=>"101011011",
  42330=>"001110111",
  42331=>"101111000",
  42332=>"100001111",
  42333=>"110101000",
  42334=>"100000000",
  42335=>"010101011",
  42336=>"011100001",
  42337=>"111010001",
  42338=>"011111010",
  42339=>"000001101",
  42340=>"011101010",
  42341=>"010010100",
  42342=>"111110010",
  42343=>"011010001",
  42344=>"110000101",
  42345=>"000000000",
  42346=>"001101010",
  42347=>"111011001",
  42348=>"110001101",
  42349=>"011011000",
  42350=>"101100110",
  42351=>"010110000",
  42352=>"001000000",
  42353=>"001010111",
  42354=>"100101001",
  42355=>"101001111",
  42356=>"010000101",
  42357=>"001111110",
  42358=>"000001010",
  42359=>"101101101",
  42360=>"010001101",
  42361=>"110110011",
  42362=>"100110010",
  42363=>"000010010",
  42364=>"000100111",
  42365=>"001011001",
  42366=>"111000001",
  42367=>"011110110",
  42368=>"110111001",
  42369=>"011111011",
  42370=>"011001000",
  42371=>"001101110",
  42372=>"000100110",
  42373=>"111001011",
  42374=>"110011001",
  42375=>"110110010",
  42376=>"000000011",
  42377=>"010001011",
  42378=>"100000010",
  42379=>"110000000",
  42380=>"101001001",
  42381=>"110101111",
  42382=>"100000111",
  42383=>"100011001",
  42384=>"110101110",
  42385=>"001000011",
  42386=>"100001110",
  42387=>"101100111",
  42388=>"110101110",
  42389=>"001100110",
  42390=>"101100110",
  42391=>"110001101",
  42392=>"100101001",
  42393=>"001100000",
  42394=>"100011000",
  42395=>"011100010",
  42396=>"001101000",
  42397=>"001101111",
  42398=>"100000001",
  42399=>"001101100",
  42400=>"110101100",
  42401=>"010000111",
  42402=>"001000001",
  42403=>"000000000",
  42404=>"101011110",
  42405=>"100100100",
  42406=>"101110111",
  42407=>"110010110",
  42408=>"111111100",
  42409=>"110011000",
  42410=>"000101100",
  42411=>"100101100",
  42412=>"010110001",
  42413=>"100011001",
  42414=>"111011110",
  42415=>"100110001",
  42416=>"000000101",
  42417=>"010111111",
  42418=>"001101011",
  42419=>"001100111",
  42420=>"110111101",
  42421=>"110001111",
  42422=>"101011000",
  42423=>"110000100",
  42424=>"110001111",
  42425=>"111001011",
  42426=>"110100110",
  42427=>"001001110",
  42428=>"000000000",
  42429=>"100001110",
  42430=>"011001001",
  42431=>"101011110",
  42432=>"111011001",
  42433=>"011001001",
  42434=>"100100011",
  42435=>"011011101",
  42436=>"000011000",
  42437=>"111100111",
  42438=>"010010101",
  42439=>"111100110",
  42440=>"001010011",
  42441=>"000110000",
  42442=>"100001010",
  42443=>"001101111",
  42444=>"000101001",
  42445=>"110110101",
  42446=>"100011010",
  42447=>"101101000",
  42448=>"001111011",
  42449=>"011011011",
  42450=>"011010001",
  42451=>"010111011",
  42452=>"011100101",
  42453=>"110110101",
  42454=>"110011111",
  42455=>"100001000",
  42456=>"000111100",
  42457=>"101000100",
  42458=>"101010101",
  42459=>"100100001",
  42460=>"110011011",
  42461=>"110100011",
  42462=>"010001001",
  42463=>"101101011",
  42464=>"010100000",
  42465=>"011001000",
  42466=>"110100100",
  42467=>"101101100",
  42468=>"000110110",
  42469=>"101011010",
  42470=>"100001010",
  42471=>"101001100",
  42472=>"010110110",
  42473=>"011110011",
  42474=>"110010111",
  42475=>"110011000",
  42476=>"101100101",
  42477=>"001111001",
  42478=>"111000110",
  42479=>"000101010",
  42480=>"110110010",
  42481=>"000110001",
  42482=>"111111001",
  42483=>"111100010",
  42484=>"001011101",
  42485=>"101010001",
  42486=>"110101101",
  42487=>"101010111",
  42488=>"100001100",
  42489=>"011001001",
  42490=>"110010010",
  42491=>"111110001",
  42492=>"000001000",
  42493=>"100100110",
  42494=>"101111110",
  42495=>"111111111",
  42496=>"100001110",
  42497=>"001000100",
  42498=>"111101110",
  42499=>"111100000",
  42500=>"111010100",
  42501=>"110101000",
  42502=>"011010110",
  42503=>"011011111",
  42504=>"100000101",
  42505=>"010111101",
  42506=>"000101100",
  42507=>"011010001",
  42508=>"111001101",
  42509=>"101000000",
  42510=>"101001000",
  42511=>"101010001",
  42512=>"111001110",
  42513=>"010111100",
  42514=>"000110000",
  42515=>"100010011",
  42516=>"110011011",
  42517=>"001001111",
  42518=>"011001111",
  42519=>"101000010",
  42520=>"101101010",
  42521=>"101001000",
  42522=>"000111110",
  42523=>"101001110",
  42524=>"000100111",
  42525=>"000000111",
  42526=>"100001010",
  42527=>"101100111",
  42528=>"101111101",
  42529=>"111100101",
  42530=>"001001001",
  42531=>"001000100",
  42532=>"011011000",
  42533=>"000011101",
  42534=>"001010001",
  42535=>"111101000",
  42536=>"000010101",
  42537=>"110001000",
  42538=>"110000100",
  42539=>"011101111",
  42540=>"011100000",
  42541=>"001101010",
  42542=>"000010001",
  42543=>"000110010",
  42544=>"110000000",
  42545=>"100101000",
  42546=>"110001110",
  42547=>"000010110",
  42548=>"000011110",
  42549=>"000110110",
  42550=>"000101010",
  42551=>"001111000",
  42552=>"110101011",
  42553=>"101110011",
  42554=>"100011000",
  42555=>"011001101",
  42556=>"010100000",
  42557=>"110000011",
  42558=>"101101011",
  42559=>"100000100",
  42560=>"111100101",
  42561=>"000100111",
  42562=>"010001010",
  42563=>"011110111",
  42564=>"101000101",
  42565=>"010011010",
  42566=>"001010001",
  42567=>"000110001",
  42568=>"001000100",
  42569=>"011001011",
  42570=>"111001111",
  42571=>"100110110",
  42572=>"011111001",
  42573=>"011001111",
  42574=>"101000011",
  42575=>"111010001",
  42576=>"110111011",
  42577=>"101101110",
  42578=>"000001110",
  42579=>"001000010",
  42580=>"101101101",
  42581=>"011101100",
  42582=>"000100000",
  42583=>"110111001",
  42584=>"001000100",
  42585=>"001100100",
  42586=>"111001110",
  42587=>"101111000",
  42588=>"000010101",
  42589=>"011110100",
  42590=>"011111100",
  42591=>"011101000",
  42592=>"001001001",
  42593=>"011010110",
  42594=>"010001010",
  42595=>"110000001",
  42596=>"011101010",
  42597=>"110110000",
  42598=>"000001010",
  42599=>"100100011",
  42600=>"000000100",
  42601=>"101101101",
  42602=>"110100001",
  42603=>"100111101",
  42604=>"111010111",
  42605=>"011101000",
  42606=>"111000110",
  42607=>"000000000",
  42608=>"001100111",
  42609=>"101010000",
  42610=>"110001110",
  42611=>"011001000",
  42612=>"000110110",
  42613=>"000100101",
  42614=>"101100110",
  42615=>"000010010",
  42616=>"100000001",
  42617=>"100110001",
  42618=>"000011111",
  42619=>"100001000",
  42620=>"111111100",
  42621=>"001111010",
  42622=>"100001110",
  42623=>"111010100",
  42624=>"011100001",
  42625=>"101000001",
  42626=>"100010011",
  42627=>"100010101",
  42628=>"011011011",
  42629=>"100100000",
  42630=>"011011111",
  42631=>"110101001",
  42632=>"011101011",
  42633=>"000001010",
  42634=>"100111011",
  42635=>"000001101",
  42636=>"111000101",
  42637=>"110110000",
  42638=>"011000001",
  42639=>"000011101",
  42640=>"010110100",
  42641=>"011010011",
  42642=>"101000111",
  42643=>"101101000",
  42644=>"101100011",
  42645=>"000111101",
  42646=>"110110100",
  42647=>"000000011",
  42648=>"011011110",
  42649=>"010010100",
  42650=>"011000110",
  42651=>"001011111",
  42652=>"000100001",
  42653=>"110100010",
  42654=>"010101100",
  42655=>"001001110",
  42656=>"101111011",
  42657=>"010001111",
  42658=>"010101001",
  42659=>"001011110",
  42660=>"011111101",
  42661=>"000011001",
  42662=>"010010100",
  42663=>"001101101",
  42664=>"110001000",
  42665=>"011101001",
  42666=>"011101100",
  42667=>"000010111",
  42668=>"010110000",
  42669=>"010100011",
  42670=>"001011000",
  42671=>"101011000",
  42672=>"010011101",
  42673=>"010101101",
  42674=>"111000111",
  42675=>"010101001",
  42676=>"000000110",
  42677=>"111101010",
  42678=>"100011101",
  42679=>"010100010",
  42680=>"000111000",
  42681=>"101001011",
  42682=>"010011110",
  42683=>"011000001",
  42684=>"110111000",
  42685=>"011110010",
  42686=>"111101111",
  42687=>"100110100",
  42688=>"110011010",
  42689=>"111111000",
  42690=>"000000110",
  42691=>"111110111",
  42692=>"011101000",
  42693=>"001011001",
  42694=>"101000100",
  42695=>"111101000",
  42696=>"110001001",
  42697=>"110110011",
  42698=>"101111110",
  42699=>"110111001",
  42700=>"111110101",
  42701=>"000100100",
  42702=>"001001001",
  42703=>"001111100",
  42704=>"100001111",
  42705=>"000100011",
  42706=>"000010011",
  42707=>"001011100",
  42708=>"001000011",
  42709=>"000111011",
  42710=>"110110000",
  42711=>"000001001",
  42712=>"001010111",
  42713=>"111101010",
  42714=>"001001011",
  42715=>"100010001",
  42716=>"001101111",
  42717=>"000010001",
  42718=>"101101001",
  42719=>"001000101",
  42720=>"000100000",
  42721=>"110111001",
  42722=>"010111110",
  42723=>"001101101",
  42724=>"110110101",
  42725=>"000001000",
  42726=>"100111000",
  42727=>"101011100",
  42728=>"001011010",
  42729=>"010101010",
  42730=>"100010100",
  42731=>"001111000",
  42732=>"001100001",
  42733=>"000000000",
  42734=>"010001111",
  42735=>"000011011",
  42736=>"010110100",
  42737=>"000010110",
  42738=>"010011111",
  42739=>"000010000",
  42740=>"100101010",
  42741=>"000100000",
  42742=>"001000101",
  42743=>"110010111",
  42744=>"110001001",
  42745=>"110100001",
  42746=>"111011011",
  42747=>"000001000",
  42748=>"100111101",
  42749=>"000110101",
  42750=>"000011111",
  42751=>"101110110",
  42752=>"101011111",
  42753=>"001000111",
  42754=>"010000000",
  42755=>"011010101",
  42756=>"100010001",
  42757=>"111000001",
  42758=>"101110111",
  42759=>"010001010",
  42760=>"100100100",
  42761=>"000101111",
  42762=>"001101100",
  42763=>"001000000",
  42764=>"011000110",
  42765=>"001011011",
  42766=>"111111100",
  42767=>"011111101",
  42768=>"101101111",
  42769=>"101011001",
  42770=>"100101000",
  42771=>"101001000",
  42772=>"100000010",
  42773=>"011101100",
  42774=>"110111101",
  42775=>"000101011",
  42776=>"000001110",
  42777=>"010000101",
  42778=>"000000100",
  42779=>"011111001",
  42780=>"101011000",
  42781=>"111101010",
  42782=>"111100110",
  42783=>"001011010",
  42784=>"000101100",
  42785=>"100001101",
  42786=>"001011001",
  42787=>"111010111",
  42788=>"101110011",
  42789=>"100100101",
  42790=>"100101111",
  42791=>"100011110",
  42792=>"011111111",
  42793=>"011000000",
  42794=>"101100000",
  42795=>"110101101",
  42796=>"101100101",
  42797=>"100001000",
  42798=>"101101110",
  42799=>"110010100",
  42800=>"001100000",
  42801=>"011011101",
  42802=>"101111010",
  42803=>"011011111",
  42804=>"110011001",
  42805=>"010000001",
  42806=>"101001000",
  42807=>"010010001",
  42808=>"000111011",
  42809=>"001000010",
  42810=>"111010000",
  42811=>"000000001",
  42812=>"000110001",
  42813=>"000011111",
  42814=>"001000111",
  42815=>"010001011",
  42816=>"001101011",
  42817=>"000110100",
  42818=>"001001111",
  42819=>"001010110",
  42820=>"011000100",
  42821=>"010000101",
  42822=>"010000000",
  42823=>"010000100",
  42824=>"000000100",
  42825=>"101111101",
  42826=>"011101000",
  42827=>"101011110",
  42828=>"000001011",
  42829=>"101010010",
  42830=>"011101110",
  42831=>"100101011",
  42832=>"110110011",
  42833=>"100000110",
  42834=>"101000111",
  42835=>"010010001",
  42836=>"001000101",
  42837=>"101000110",
  42838=>"100110100",
  42839=>"001110010",
  42840=>"010011001",
  42841=>"011110001",
  42842=>"000000101",
  42843=>"100010110",
  42844=>"010000001",
  42845=>"000100111",
  42846=>"011010011",
  42847=>"001101110",
  42848=>"010010011",
  42849=>"010000100",
  42850=>"001000010",
  42851=>"110110010",
  42852=>"010011010",
  42853=>"010101101",
  42854=>"001100001",
  42855=>"011110110",
  42856=>"100100010",
  42857=>"011010101",
  42858=>"100100010",
  42859=>"110000010",
  42860=>"010111110",
  42861=>"001100100",
  42862=>"100101101",
  42863=>"011111111",
  42864=>"000110100",
  42865=>"000111011",
  42866=>"010111101",
  42867=>"001000001",
  42868=>"000011011",
  42869=>"001000001",
  42870=>"110010111",
  42871=>"100110011",
  42872=>"001001111",
  42873=>"100110111",
  42874=>"001101110",
  42875=>"000000111",
  42876=>"000100011",
  42877=>"111001001",
  42878=>"101111110",
  42879=>"111110100",
  42880=>"001010110",
  42881=>"100001110",
  42882=>"100001011",
  42883=>"010100111",
  42884=>"101111000",
  42885=>"001101100",
  42886=>"001011011",
  42887=>"100010010",
  42888=>"100100000",
  42889=>"111100110",
  42890=>"111001010",
  42891=>"100010101",
  42892=>"111101000",
  42893=>"011001000",
  42894=>"110011010",
  42895=>"111010100",
  42896=>"100000001",
  42897=>"010001100",
  42898=>"110110111",
  42899=>"111100011",
  42900=>"000001010",
  42901=>"001111111",
  42902=>"100101100",
  42903=>"111001101",
  42904=>"010000100",
  42905=>"101100010",
  42906=>"010011010",
  42907=>"100110001",
  42908=>"010101001",
  42909=>"111110001",
  42910=>"001011110",
  42911=>"011000111",
  42912=>"000001111",
  42913=>"011100010",
  42914=>"011101000",
  42915=>"101100111",
  42916=>"110110111",
  42917=>"000111011",
  42918=>"010010011",
  42919=>"001100011",
  42920=>"100010000",
  42921=>"011011111",
  42922=>"100101101",
  42923=>"100101100",
  42924=>"000110011",
  42925=>"101000100",
  42926=>"110111011",
  42927=>"111010110",
  42928=>"101101110",
  42929=>"110110011",
  42930=>"001001101",
  42931=>"011110110",
  42932=>"001011011",
  42933=>"001001111",
  42934=>"000010101",
  42935=>"000000000",
  42936=>"011000100",
  42937=>"101100101",
  42938=>"100110111",
  42939=>"001011011",
  42940=>"000100011",
  42941=>"000000001",
  42942=>"111010111",
  42943=>"100001111",
  42944=>"001000111",
  42945=>"001010110",
  42946=>"110000110",
  42947=>"001010101",
  42948=>"100011010",
  42949=>"110111101",
  42950=>"111111100",
  42951=>"110001110",
  42952=>"000101110",
  42953=>"000010100",
  42954=>"100001100",
  42955=>"000110011",
  42956=>"110111111",
  42957=>"110101101",
  42958=>"010111010",
  42959=>"001100001",
  42960=>"011010011",
  42961=>"000100011",
  42962=>"100100100",
  42963=>"011001100",
  42964=>"100000100",
  42965=>"001001000",
  42966=>"101000100",
  42967=>"011110101",
  42968=>"000010110",
  42969=>"001101001",
  42970=>"111101001",
  42971=>"111101111",
  42972=>"101011101",
  42973=>"100011000",
  42974=>"010100101",
  42975=>"110011101",
  42976=>"010111110",
  42977=>"101100100",
  42978=>"110111111",
  42979=>"011001010",
  42980=>"101100110",
  42981=>"100100111",
  42982=>"111111011",
  42983=>"100110100",
  42984=>"010000101",
  42985=>"010011001",
  42986=>"100010010",
  42987=>"010011000",
  42988=>"100011011",
  42989=>"010111001",
  42990=>"101101011",
  42991=>"110101110",
  42992=>"111101010",
  42993=>"000110101",
  42994=>"000000000",
  42995=>"100100110",
  42996=>"110010110",
  42997=>"001010101",
  42998=>"110000001",
  42999=>"001010010",
  43000=>"110000100",
  43001=>"011111110",
  43002=>"010001100",
  43003=>"100011001",
  43004=>"110110011",
  43005=>"010110010",
  43006=>"001101101",
  43007=>"100111111",
  43008=>"101010100",
  43009=>"000111111",
  43010=>"110100110",
  43011=>"000000111",
  43012=>"001000110",
  43013=>"011101001",
  43014=>"110101111",
  43015=>"011010000",
  43016=>"010011010",
  43017=>"110001100",
  43018=>"101101000",
  43019=>"010111101",
  43020=>"111101110",
  43021=>"110111001",
  43022=>"000011101",
  43023=>"101010001",
  43024=>"111100111",
  43025=>"101100110",
  43026=>"111001011",
  43027=>"101001111",
  43028=>"011101110",
  43029=>"010011101",
  43030=>"100111101",
  43031=>"011110110",
  43032=>"000001111",
  43033=>"001111011",
  43034=>"101111001",
  43035=>"100111000",
  43036=>"011100000",
  43037=>"000101100",
  43038=>"001110011",
  43039=>"100000110",
  43040=>"011010010",
  43041=>"000011010",
  43042=>"010010010",
  43043=>"110011100",
  43044=>"110011010",
  43045=>"110001000",
  43046=>"110001000",
  43047=>"000111110",
  43048=>"000100110",
  43049=>"100010011",
  43050=>"101010100",
  43051=>"010100010",
  43052=>"011011110",
  43053=>"001100101",
  43054=>"111100100",
  43055=>"000100110",
  43056=>"010110010",
  43057=>"000110011",
  43058=>"101100111",
  43059=>"010000001",
  43060=>"110111000",
  43061=>"111110100",
  43062=>"100000110",
  43063=>"100101001",
  43064=>"001100110",
  43065=>"101001110",
  43066=>"011001101",
  43067=>"001110110",
  43068=>"100011111",
  43069=>"111011011",
  43070=>"100100000",
  43071=>"111101110",
  43072=>"011101010",
  43073=>"101000011",
  43074=>"100100000",
  43075=>"111101110",
  43076=>"001001101",
  43077=>"001011100",
  43078=>"010011000",
  43079=>"111100100",
  43080=>"101101011",
  43081=>"011011011",
  43082=>"011011011",
  43083=>"101111000",
  43084=>"010110111",
  43085=>"100110111",
  43086=>"001111101",
  43087=>"110111010",
  43088=>"010001100",
  43089=>"101111011",
  43090=>"100110110",
  43091=>"011000101",
  43092=>"011110101",
  43093=>"000000010",
  43094=>"000110010",
  43095=>"101101100",
  43096=>"100001001",
  43097=>"111101110",
  43098=>"101010000",
  43099=>"111100110",
  43100=>"001001011",
  43101=>"010001000",
  43102=>"001100111",
  43103=>"010100001",
  43104=>"111010001",
  43105=>"110010011",
  43106=>"000011000",
  43107=>"111101111",
  43108=>"101100100",
  43109=>"111100111",
  43110=>"100110001",
  43111=>"110101101",
  43112=>"010011101",
  43113=>"010000000",
  43114=>"101000011",
  43115=>"011110110",
  43116=>"010011000",
  43117=>"110110000",
  43118=>"010011101",
  43119=>"001000100",
  43120=>"110101001",
  43121=>"101010110",
  43122=>"111001101",
  43123=>"100101100",
  43124=>"100101100",
  43125=>"111111111",
  43126=>"100011111",
  43127=>"000001010",
  43128=>"010100011",
  43129=>"011101101",
  43130=>"001101111",
  43131=>"011111011",
  43132=>"111110011",
  43133=>"000110001",
  43134=>"100010110",
  43135=>"010111000",
  43136=>"100111000",
  43137=>"011000110",
  43138=>"010001110",
  43139=>"000101110",
  43140=>"111000000",
  43141=>"100110110",
  43142=>"100000000",
  43143=>"100011000",
  43144=>"010100000",
  43145=>"000010001",
  43146=>"101000011",
  43147=>"111010101",
  43148=>"110111000",
  43149=>"011100100",
  43150=>"110011111",
  43151=>"101000101",
  43152=>"001111101",
  43153=>"110011000",
  43154=>"011101010",
  43155=>"011011001",
  43156=>"000010001",
  43157=>"011000110",
  43158=>"101001111",
  43159=>"101100000",
  43160=>"000000001",
  43161=>"001101100",
  43162=>"101100101",
  43163=>"100110000",
  43164=>"101011001",
  43165=>"011000011",
  43166=>"110011010",
  43167=>"110110000",
  43168=>"000100110",
  43169=>"001011010",
  43170=>"100100000",
  43171=>"111011110",
  43172=>"110110101",
  43173=>"101010011",
  43174=>"111001011",
  43175=>"000000001",
  43176=>"000010010",
  43177=>"011111100",
  43178=>"101100001",
  43179=>"110000011",
  43180=>"111110111",
  43181=>"101100110",
  43182=>"001101110",
  43183=>"101111011",
  43184=>"010010000",
  43185=>"010010011",
  43186=>"011110100",
  43187=>"010101100",
  43188=>"111001011",
  43189=>"001011011",
  43190=>"001001001",
  43191=>"010011000",
  43192=>"101010110",
  43193=>"101001010",
  43194=>"110100110",
  43195=>"010111000",
  43196=>"101110001",
  43197=>"111101011",
  43198=>"010000011",
  43199=>"110100110",
  43200=>"100010010",
  43201=>"101101011",
  43202=>"101111110",
  43203=>"101001101",
  43204=>"111011111",
  43205=>"011001001",
  43206=>"110111110",
  43207=>"101011000",
  43208=>"111111000",
  43209=>"010100001",
  43210=>"000010000",
  43211=>"001100110",
  43212=>"001100111",
  43213=>"101101111",
  43214=>"100100010",
  43215=>"001101001",
  43216=>"101101110",
  43217=>"111001000",
  43218=>"101010111",
  43219=>"001011111",
  43220=>"101111101",
  43221=>"111110100",
  43222=>"101001000",
  43223=>"101100000",
  43224=>"010100000",
  43225=>"010111010",
  43226=>"011110110",
  43227=>"111111000",
  43228=>"010000001",
  43229=>"010110000",
  43230=>"100011110",
  43231=>"111101111",
  43232=>"010111001",
  43233=>"011001101",
  43234=>"100010001",
  43235=>"011011011",
  43236=>"110111110",
  43237=>"001101111",
  43238=>"011011011",
  43239=>"011001011",
  43240=>"010011100",
  43241=>"101101000",
  43242=>"000101110",
  43243=>"010100101",
  43244=>"100101101",
  43245=>"101111110",
  43246=>"101010100",
  43247=>"101110010",
  43248=>"111101011",
  43249=>"111011100",
  43250=>"011100100",
  43251=>"100001100",
  43252=>"101101000",
  43253=>"100010111",
  43254=>"101101111",
  43255=>"101100010",
  43256=>"011011001",
  43257=>"110111000",
  43258=>"101100100",
  43259=>"110111101",
  43260=>"101101010",
  43261=>"101100111",
  43262=>"001100110",
  43263=>"111111101",
  43264=>"101001001",
  43265=>"001100000",
  43266=>"111110011",
  43267=>"100100000",
  43268=>"001110110",
  43269=>"001110000",
  43270=>"100000100",
  43271=>"011110110",
  43272=>"110110001",
  43273=>"100101000",
  43274=>"011100100",
  43275=>"111010001",
  43276=>"101111011",
  43277=>"010000010",
  43278=>"111100111",
  43279=>"101110010",
  43280=>"010111100",
  43281=>"100011111",
  43282=>"101001001",
  43283=>"100101111",
  43284=>"101000010",
  43285=>"101100010",
  43286=>"010101001",
  43287=>"100101000",
  43288=>"111101101",
  43289=>"101101000",
  43290=>"100001110",
  43291=>"101110000",
  43292=>"110000000",
  43293=>"100110111",
  43294=>"011000111",
  43295=>"000101000",
  43296=>"000000110",
  43297=>"001111010",
  43298=>"010100011",
  43299=>"101000000",
  43300=>"010001000",
  43301=>"110110110",
  43302=>"010111111",
  43303=>"011100011",
  43304=>"100001011",
  43305=>"000111111",
  43306=>"000111100",
  43307=>"011100000",
  43308=>"111010011",
  43309=>"110100111",
  43310=>"111101100",
  43311=>"100010110",
  43312=>"001001101",
  43313=>"110100000",
  43314=>"100000000",
  43315=>"000100011",
  43316=>"011011000",
  43317=>"111011011",
  43318=>"101011001",
  43319=>"001001101",
  43320=>"010011110",
  43321=>"111001100",
  43322=>"000110100",
  43323=>"100000010",
  43324=>"010111011",
  43325=>"110011111",
  43326=>"000000111",
  43327=>"000001010",
  43328=>"100111001",
  43329=>"000000011",
  43330=>"011111110",
  43331=>"100000000",
  43332=>"011010001",
  43333=>"010010101",
  43334=>"001100100",
  43335=>"011011001",
  43336=>"010001000",
  43337=>"001000000",
  43338=>"100001111",
  43339=>"011111000",
  43340=>"101001000",
  43341=>"011111110",
  43342=>"100111011",
  43343=>"111111100",
  43344=>"100110101",
  43345=>"101000001",
  43346=>"011110111",
  43347=>"100110011",
  43348=>"000000100",
  43349=>"100111100",
  43350=>"000000111",
  43351=>"001100100",
  43352=>"000101100",
  43353=>"000110110",
  43354=>"010011111",
  43355=>"000010100",
  43356=>"010100100",
  43357=>"000111010",
  43358=>"011010110",
  43359=>"000110111",
  43360=>"010111110",
  43361=>"001101110",
  43362=>"001001111",
  43363=>"000001111",
  43364=>"001001001",
  43365=>"100000000",
  43366=>"010100111",
  43367=>"000111010",
  43368=>"011111111",
  43369=>"101001011",
  43370=>"000000000",
  43371=>"111111001",
  43372=>"101101100",
  43373=>"001100000",
  43374=>"111011011",
  43375=>"111111001",
  43376=>"100101100",
  43377=>"110010010",
  43378=>"111110101",
  43379=>"000000101",
  43380=>"110110100",
  43381=>"101001111",
  43382=>"111110101",
  43383=>"011100110",
  43384=>"110111111",
  43385=>"001000110",
  43386=>"010110011",
  43387=>"110111000",
  43388=>"000110010",
  43389=>"100111101",
  43390=>"001101111",
  43391=>"100000011",
  43392=>"100010111",
  43393=>"011010100",
  43394=>"000010001",
  43395=>"111110010",
  43396=>"001010010",
  43397=>"000000000",
  43398=>"110101000",
  43399=>"001010101",
  43400=>"001000111",
  43401=>"100101010",
  43402=>"100101101",
  43403=>"000111110",
  43404=>"001000000",
  43405=>"000110110",
  43406=>"111010111",
  43407=>"100101111",
  43408=>"110100010",
  43409=>"010101011",
  43410=>"110100001",
  43411=>"001001001",
  43412=>"001100101",
  43413=>"000100011",
  43414=>"111010000",
  43415=>"101100000",
  43416=>"111000100",
  43417=>"101010100",
  43418=>"101001000",
  43419=>"010100010",
  43420=>"001001001",
  43421=>"100011101",
  43422=>"100101000",
  43423=>"001110011",
  43424=>"000010000",
  43425=>"110110001",
  43426=>"011100101",
  43427=>"101001110",
  43428=>"111110101",
  43429=>"011101111",
  43430=>"111011011",
  43431=>"110000101",
  43432=>"110111010",
  43433=>"101011100",
  43434=>"101001101",
  43435=>"010011011",
  43436=>"001011101",
  43437=>"010011001",
  43438=>"010001001",
  43439=>"001001100",
  43440=>"000000011",
  43441=>"110010000",
  43442=>"000011111",
  43443=>"000000111",
  43444=>"100111011",
  43445=>"000111110",
  43446=>"000010011",
  43447=>"110010110",
  43448=>"111101110",
  43449=>"100100010",
  43450=>"010011010",
  43451=>"010001000",
  43452=>"000110110",
  43453=>"010100101",
  43454=>"011110101",
  43455=>"010100001",
  43456=>"001100010",
  43457=>"001110100",
  43458=>"101111110",
  43459=>"000000101",
  43460=>"001011101",
  43461=>"010110010",
  43462=>"111011010",
  43463=>"110110010",
  43464=>"110000111",
  43465=>"110111111",
  43466=>"101100001",
  43467=>"011001101",
  43468=>"010100100",
  43469=>"111100000",
  43470=>"101000001",
  43471=>"110111000",
  43472=>"000000111",
  43473=>"001011001",
  43474=>"011000010",
  43475=>"011100111",
  43476=>"100011011",
  43477=>"001000000",
  43478=>"111111001",
  43479=>"101011101",
  43480=>"001001100",
  43481=>"010010000",
  43482=>"111111111",
  43483=>"000110111",
  43484=>"011010101",
  43485=>"000000101",
  43486=>"111100110",
  43487=>"000101111",
  43488=>"111100000",
  43489=>"001111001",
  43490=>"001101111",
  43491=>"101001001",
  43492=>"000100101",
  43493=>"010100001",
  43494=>"100011001",
  43495=>"001100110",
  43496=>"011010011",
  43497=>"111011100",
  43498=>"111110000",
  43499=>"100101001",
  43500=>"011011101",
  43501=>"101010101",
  43502=>"010001100",
  43503=>"110001101",
  43504=>"001011001",
  43505=>"110111100",
  43506=>"111000010",
  43507=>"001110101",
  43508=>"101111101",
  43509=>"110101100",
  43510=>"110011110",
  43511=>"110101111",
  43512=>"110001001",
  43513=>"010101101",
  43514=>"000110000",
  43515=>"110001010",
  43516=>"000011000",
  43517=>"001000110",
  43518=>"111011000",
  43519=>"011110101",
  43520=>"101111010",
  43521=>"000110111",
  43522=>"001011001",
  43523=>"011100111",
  43524=>"101101101",
  43525=>"101101110",
  43526=>"111000110",
  43527=>"010000111",
  43528=>"111010111",
  43529=>"100010100",
  43530=>"011101101",
  43531=>"010100000",
  43532=>"100000011",
  43533=>"101111001",
  43534=>"100001001",
  43535=>"111111010",
  43536=>"001010101",
  43537=>"110110101",
  43538=>"100111000",
  43539=>"101011110",
  43540=>"010110000",
  43541=>"001011001",
  43542=>"000000001",
  43543=>"101000101",
  43544=>"101011000",
  43545=>"101100011",
  43546=>"110111000",
  43547=>"011011101",
  43548=>"001100110",
  43549=>"101111000",
  43550=>"100110000",
  43551=>"010000101",
  43552=>"111011011",
  43553=>"110001111",
  43554=>"111011010",
  43555=>"000101000",
  43556=>"011000010",
  43557=>"100000100",
  43558=>"011110111",
  43559=>"000001100",
  43560=>"100100101",
  43561=>"001011011",
  43562=>"110000000",
  43563=>"011110101",
  43564=>"010111100",
  43565=>"000111111",
  43566=>"101101010",
  43567=>"011100100",
  43568=>"000110011",
  43569=>"111111000",
  43570=>"011110101",
  43571=>"101011011",
  43572=>"110111000",
  43573=>"110111110",
  43574=>"001101101",
  43575=>"100010000",
  43576=>"000000101",
  43577=>"001101001",
  43578=>"001111011",
  43579=>"101100110",
  43580=>"101110000",
  43581=>"111011000",
  43582=>"100000010",
  43583=>"000100100",
  43584=>"101001111",
  43585=>"011110101",
  43586=>"011101000",
  43587=>"110011011",
  43588=>"111011100",
  43589=>"000011001",
  43590=>"001001000",
  43591=>"001011111",
  43592=>"010011010",
  43593=>"111101101",
  43594=>"010110010",
  43595=>"101101001",
  43596=>"101101001",
  43597=>"010001011",
  43598=>"010010001",
  43599=>"000101100",
  43600=>"011111011",
  43601=>"110001000",
  43602=>"010101011",
  43603=>"101000100",
  43604=>"000101110",
  43605=>"111001101",
  43606=>"000111111",
  43607=>"000010110",
  43608=>"100101110",
  43609=>"000000001",
  43610=>"111100100",
  43611=>"011110110",
  43612=>"100010000",
  43613=>"000000010",
  43614=>"111100111",
  43615=>"111011011",
  43616=>"011001000",
  43617=>"001111001",
  43618=>"101111011",
  43619=>"010100000",
  43620=>"011000000",
  43621=>"011001100",
  43622=>"110011001",
  43623=>"010110101",
  43624=>"101100111",
  43625=>"010011101",
  43626=>"101100110",
  43627=>"110001101",
  43628=>"010101011",
  43629=>"001110110",
  43630=>"110101010",
  43631=>"101001101",
  43632=>"101011001",
  43633=>"011101000",
  43634=>"011000011",
  43635=>"111110001",
  43636=>"001011001",
  43637=>"011110110",
  43638=>"001110110",
  43639=>"111101001",
  43640=>"111100001",
  43641=>"001101101",
  43642=>"011111001",
  43643=>"001001001",
  43644=>"101110100",
  43645=>"100110001",
  43646=>"010111101",
  43647=>"010010010",
  43648=>"001111011",
  43649=>"011010011",
  43650=>"000001011",
  43651=>"010000100",
  43652=>"100000011",
  43653=>"011010010",
  43654=>"010100110",
  43655=>"011101110",
  43656=>"111111001",
  43657=>"100100111",
  43658=>"110010101",
  43659=>"110101001",
  43660=>"111000011",
  43661=>"100001000",
  43662=>"011000011",
  43663=>"011000001",
  43664=>"111111111",
  43665=>"110011011",
  43666=>"001101110",
  43667=>"011101010",
  43668=>"011011011",
  43669=>"000100101",
  43670=>"001001101",
  43671=>"001010000",
  43672=>"101010000",
  43673=>"011111110",
  43674=>"000111101",
  43675=>"001100000",
  43676=>"101000001",
  43677=>"010010010",
  43678=>"110011000",
  43679=>"111011011",
  43680=>"101001010",
  43681=>"110101011",
  43682=>"000010101",
  43683=>"001111100",
  43684=>"111011001",
  43685=>"000000110",
  43686=>"100101001",
  43687=>"011001000",
  43688=>"110101010",
  43689=>"001100011",
  43690=>"000100100",
  43691=>"101011110",
  43692=>"101110000",
  43693=>"110010111",
  43694=>"100011001",
  43695=>"000101010",
  43696=>"101011000",
  43697=>"111110110",
  43698=>"001101110",
  43699=>"011010000",
  43700=>"010100011",
  43701=>"111111011",
  43702=>"000000101",
  43703=>"000010001",
  43704=>"111000111",
  43705=>"010001000",
  43706=>"100001100",
  43707=>"111110011",
  43708=>"000100110",
  43709=>"001011101",
  43710=>"011111000",
  43711=>"101010111",
  43712=>"101001110",
  43713=>"000101000",
  43714=>"001000011",
  43715=>"100100000",
  43716=>"111011000",
  43717=>"010101111",
  43718=>"101000110",
  43719=>"110010111",
  43720=>"100011000",
  43721=>"110110101",
  43722=>"100000000",
  43723=>"101100100",
  43724=>"011101110",
  43725=>"111011110",
  43726=>"110101011",
  43727=>"100011001",
  43728=>"111011011",
  43729=>"000100111",
  43730=>"111001000",
  43731=>"000001001",
  43732=>"000000110",
  43733=>"010000011",
  43734=>"000001111",
  43735=>"101010111",
  43736=>"001011011",
  43737=>"110111100",
  43738=>"000000110",
  43739=>"111011011",
  43740=>"100010111",
  43741=>"110100000",
  43742=>"000001101",
  43743=>"100111101",
  43744=>"100110000",
  43745=>"110110000",
  43746=>"000101011",
  43747=>"101000011",
  43748=>"100011101",
  43749=>"010110000",
  43750=>"000101101",
  43751=>"101101001",
  43752=>"010100011",
  43753=>"110011101",
  43754=>"000001110",
  43755=>"110100011",
  43756=>"000111000",
  43757=>"100101111",
  43758=>"110100110",
  43759=>"011001101",
  43760=>"001101011",
  43761=>"011011000",
  43762=>"101001111",
  43763=>"001010000",
  43764=>"110101000",
  43765=>"110100111",
  43766=>"101000011",
  43767=>"001110100",
  43768=>"000000001",
  43769=>"111100111",
  43770=>"001111011",
  43771=>"101110000",
  43772=>"101001010",
  43773=>"000001100",
  43774=>"111000010",
  43775=>"000111101",
  43776=>"111110000",
  43777=>"101010000",
  43778=>"000110110",
  43779=>"110011111",
  43780=>"011011011",
  43781=>"001110001",
  43782=>"101111001",
  43783=>"001101100",
  43784=>"100010010",
  43785=>"000010110",
  43786=>"110100011",
  43787=>"011100100",
  43788=>"100110100",
  43789=>"011011101",
  43790=>"101000000",
  43791=>"101010001",
  43792=>"111111100",
  43793=>"011001011",
  43794=>"011111010",
  43795=>"001001000",
  43796=>"111010101",
  43797=>"010000101",
  43798=>"111000100",
  43799=>"000101001",
  43800=>"101101101",
  43801=>"001001111",
  43802=>"100001000",
  43803=>"010000010",
  43804=>"010000001",
  43805=>"111111010",
  43806=>"000000011",
  43807=>"010110101",
  43808=>"001101101",
  43809=>"100100001",
  43810=>"110100111",
  43811=>"010100111",
  43812=>"111001100",
  43813=>"010110010",
  43814=>"010000010",
  43815=>"010101011",
  43816=>"000011000",
  43817=>"110111001",
  43818=>"011011011",
  43819=>"011010001",
  43820=>"110001001",
  43821=>"101101010",
  43822=>"111101001",
  43823=>"001001010",
  43824=>"100100111",
  43825=>"000000110",
  43826=>"100110110",
  43827=>"010011010",
  43828=>"100001011",
  43829=>"111000111",
  43830=>"000000100",
  43831=>"100100011",
  43832=>"100001001",
  43833=>"010101011",
  43834=>"101000110",
  43835=>"110111111",
  43836=>"110111010",
  43837=>"000011001",
  43838=>"110001000",
  43839=>"111001111",
  43840=>"110000100",
  43841=>"101001010",
  43842=>"000000011",
  43843=>"100110100",
  43844=>"000001111",
  43845=>"001001110",
  43846=>"011010100",
  43847=>"100111010",
  43848=>"101110001",
  43849=>"011000001",
  43850=>"010110011",
  43851=>"010001001",
  43852=>"001001010",
  43853=>"110101110",
  43854=>"110001100",
  43855=>"100001010",
  43856=>"100101010",
  43857=>"100000010",
  43858=>"011111011",
  43859=>"010011001",
  43860=>"011110011",
  43861=>"111100110",
  43862=>"011101011",
  43863=>"010110011",
  43864=>"100010000",
  43865=>"110101010",
  43866=>"001101010",
  43867=>"000100010",
  43868=>"011101111",
  43869=>"100100100",
  43870=>"011010011",
  43871=>"111000111",
  43872=>"010100010",
  43873=>"101001111",
  43874=>"110011101",
  43875=>"011111111",
  43876=>"010000011",
  43877=>"010111111",
  43878=>"011011000",
  43879=>"100011000",
  43880=>"111010001",
  43881=>"011110101",
  43882=>"000010011",
  43883=>"001010001",
  43884=>"101000100",
  43885=>"001001011",
  43886=>"000101000",
  43887=>"111101110",
  43888=>"001001001",
  43889=>"111110011",
  43890=>"001011001",
  43891=>"110011100",
  43892=>"000000000",
  43893=>"101110111",
  43894=>"100000000",
  43895=>"100111101",
  43896=>"101010010",
  43897=>"011110011",
  43898=>"001000100",
  43899=>"110011111",
  43900=>"010001111",
  43901=>"000001001",
  43902=>"100111011",
  43903=>"010100010",
  43904=>"010010001",
  43905=>"010010010",
  43906=>"010111000",
  43907=>"011110000",
  43908=>"111011110",
  43909=>"101101101",
  43910=>"000111010",
  43911=>"110000111",
  43912=>"101101100",
  43913=>"000100010",
  43914=>"101000001",
  43915=>"000001010",
  43916=>"011011110",
  43917=>"110000101",
  43918=>"010001100",
  43919=>"101110110",
  43920=>"001001000",
  43921=>"001001101",
  43922=>"000001000",
  43923=>"100111101",
  43924=>"110110101",
  43925=>"000010001",
  43926=>"011110011",
  43927=>"100101001",
  43928=>"011110100",
  43929=>"001011111",
  43930=>"011010011",
  43931=>"011000000",
  43932=>"010101101",
  43933=>"000100100",
  43934=>"111001100",
  43935=>"001110001",
  43936=>"001111010",
  43937=>"011000000",
  43938=>"111001110",
  43939=>"000101010",
  43940=>"010001101",
  43941=>"011111010",
  43942=>"000110000",
  43943=>"010000011",
  43944=>"001111100",
  43945=>"101110010",
  43946=>"100100010",
  43947=>"001100101",
  43948=>"011000011",
  43949=>"001011110",
  43950=>"010100001",
  43951=>"110001000",
  43952=>"011001011",
  43953=>"011010001",
  43954=>"011001111",
  43955=>"100101110",
  43956=>"111000100",
  43957=>"101101110",
  43958=>"011001110",
  43959=>"110100100",
  43960=>"000101110",
  43961=>"000010001",
  43962=>"111000010",
  43963=>"001011101",
  43964=>"101111100",
  43965=>"100000000",
  43966=>"010001110",
  43967=>"000011010",
  43968=>"011110000",
  43969=>"011100001",
  43970=>"100001011",
  43971=>"000110000",
  43972=>"010100110",
  43973=>"001011101",
  43974=>"001111000",
  43975=>"111100000",
  43976=>"000110010",
  43977=>"100101110",
  43978=>"001010101",
  43979=>"000111100",
  43980=>"001111111",
  43981=>"110111000",
  43982=>"001000111",
  43983=>"011011001",
  43984=>"101110100",
  43985=>"001101111",
  43986=>"111110000",
  43987=>"001000101",
  43988=>"011000101",
  43989=>"111010100",
  43990=>"000111111",
  43991=>"111010001",
  43992=>"110000111",
  43993=>"101011000",
  43994=>"111101010",
  43995=>"110100101",
  43996=>"010110110",
  43997=>"000010010",
  43998=>"110011001",
  43999=>"100110101",
  44000=>"011000110",
  44001=>"111010011",
  44002=>"001001010",
  44003=>"011011011",
  44004=>"001001000",
  44005=>"010000100",
  44006=>"010111001",
  44007=>"110011100",
  44008=>"110100100",
  44009=>"011000100",
  44010=>"100011111",
  44011=>"011101001",
  44012=>"001101110",
  44013=>"110100010",
  44014=>"101111101",
  44015=>"000110110",
  44016=>"100111101",
  44017=>"011011001",
  44018=>"001110111",
  44019=>"011001001",
  44020=>"010101000",
  44021=>"000101110",
  44022=>"111111001",
  44023=>"000010111",
  44024=>"010001001",
  44025=>"101010011",
  44026=>"101010010",
  44027=>"000011010",
  44028=>"001001001",
  44029=>"000011000",
  44030=>"110111110",
  44031=>"000100010",
  44032=>"010001101",
  44033=>"000011101",
  44034=>"101011001",
  44035=>"011110001",
  44036=>"010001000",
  44037=>"001101010",
  44038=>"011010111",
  44039=>"010100010",
  44040=>"111000001",
  44041=>"100011011",
  44042=>"111010101",
  44043=>"101001101",
  44044=>"011010110",
  44045=>"000001111",
  44046=>"001101101",
  44047=>"110001000",
  44048=>"110000111",
  44049=>"100011011",
  44050=>"001111100",
  44051=>"110010010",
  44052=>"101010101",
  44053=>"011010111",
  44054=>"110101000",
  44055=>"010001001",
  44056=>"001000101",
  44057=>"100100000",
  44058=>"111010111",
  44059=>"001110111",
  44060=>"111010101",
  44061=>"101000111",
  44062=>"001101101",
  44063=>"111010001",
  44064=>"010111101",
  44065=>"111101000",
  44066=>"111111011",
  44067=>"001101101",
  44068=>"101101011",
  44069=>"010100111",
  44070=>"111011010",
  44071=>"110101010",
  44072=>"110111000",
  44073=>"001110000",
  44074=>"000001111",
  44075=>"000010011",
  44076=>"010011111",
  44077=>"001100111",
  44078=>"010000000",
  44079=>"000110111",
  44080=>"111011000",
  44081=>"100001111",
  44082=>"100111100",
  44083=>"101110110",
  44084=>"000011000",
  44085=>"011011001",
  44086=>"111101111",
  44087=>"000001101",
  44088=>"011000000",
  44089=>"000111010",
  44090=>"011110000",
  44091=>"111101111",
  44092=>"111010000",
  44093=>"011011001",
  44094=>"011011000",
  44095=>"111111011",
  44096=>"000000010",
  44097=>"010110101",
  44098=>"000011000",
  44099=>"010110001",
  44100=>"010010111",
  44101=>"001010001",
  44102=>"011111010",
  44103=>"110001111",
  44104=>"100111010",
  44105=>"010000110",
  44106=>"011011110",
  44107=>"011101010",
  44108=>"100110000",
  44109=>"100100011",
  44110=>"000011100",
  44111=>"100111110",
  44112=>"100110001",
  44113=>"011110111",
  44114=>"100000110",
  44115=>"000000100",
  44116=>"001101111",
  44117=>"011011010",
  44118=>"111010000",
  44119=>"110000100",
  44120=>"000101000",
  44121=>"111001101",
  44122=>"011001001",
  44123=>"001000011",
  44124=>"101000111",
  44125=>"100010111",
  44126=>"000001100",
  44127=>"010111110",
  44128=>"010101011",
  44129=>"000111110",
  44130=>"010111100",
  44131=>"110111011",
  44132=>"100001100",
  44133=>"100101111",
  44134=>"111001001",
  44135=>"100101111",
  44136=>"100110100",
  44137=>"111100111",
  44138=>"001100010",
  44139=>"111100110",
  44140=>"111010100",
  44141=>"001110001",
  44142=>"100011000",
  44143=>"011011000",
  44144=>"010101110",
  44145=>"001111111",
  44146=>"111101111",
  44147=>"011101001",
  44148=>"010000010",
  44149=>"110010100",
  44150=>"110011111",
  44151=>"110101110",
  44152=>"011101110",
  44153=>"111000000",
  44154=>"001011011",
  44155=>"000010100",
  44156=>"001100011",
  44157=>"101100110",
  44158=>"010011101",
  44159=>"100011000",
  44160=>"011101110",
  44161=>"101111011",
  44162=>"001001000",
  44163=>"101110111",
  44164=>"100100101",
  44165=>"111110110",
  44166=>"000101000",
  44167=>"110111001",
  44168=>"101111010",
  44169=>"000010111",
  44170=>"001101011",
  44171=>"000000011",
  44172=>"111001111",
  44173=>"100100110",
  44174=>"100010001",
  44175=>"101101001",
  44176=>"110011111",
  44177=>"101011111",
  44178=>"001010100",
  44179=>"001001100",
  44180=>"100000000",
  44181=>"000100000",
  44182=>"100111101",
  44183=>"010000010",
  44184=>"011100010",
  44185=>"101110011",
  44186=>"101010011",
  44187=>"101010110",
  44188=>"100110110",
  44189=>"111100010",
  44190=>"001100011",
  44191=>"001101011",
  44192=>"000011000",
  44193=>"111110001",
  44194=>"111111111",
  44195=>"010011010",
  44196=>"011000000",
  44197=>"011000101",
  44198=>"110001101",
  44199=>"011101111",
  44200=>"111001110",
  44201=>"010011100",
  44202=>"110100000",
  44203=>"111011011",
  44204=>"001010011",
  44205=>"000011100",
  44206=>"010001000",
  44207=>"111110011",
  44208=>"101101110",
  44209=>"011010100",
  44210=>"001100100",
  44211=>"110101011",
  44212=>"101000111",
  44213=>"000010001",
  44214=>"101000011",
  44215=>"111110110",
  44216=>"100100111",
  44217=>"110000011",
  44218=>"000010011",
  44219=>"111101110",
  44220=>"011001001",
  44221=>"101011100",
  44222=>"100010110",
  44223=>"010010010",
  44224=>"001111010",
  44225=>"101001001",
  44226=>"111101111",
  44227=>"010000001",
  44228=>"101000000",
  44229=>"011111001",
  44230=>"100000110",
  44231=>"000001101",
  44232=>"010010011",
  44233=>"111111100",
  44234=>"110010010",
  44235=>"011101011",
  44236=>"000101110",
  44237=>"100000010",
  44238=>"111111111",
  44239=>"110000000",
  44240=>"110000010",
  44241=>"101010010",
  44242=>"111011111",
  44243=>"111111010",
  44244=>"100110001",
  44245=>"111100001",
  44246=>"111111010",
  44247=>"110000000",
  44248=>"011000110",
  44249=>"101001010",
  44250=>"111011111",
  44251=>"110001111",
  44252=>"001001001",
  44253=>"111111100",
  44254=>"011001110",
  44255=>"101000110",
  44256=>"111010100",
  44257=>"010001000",
  44258=>"000000011",
  44259=>"111101001",
  44260=>"100101010",
  44261=>"001101110",
  44262=>"010100011",
  44263=>"000010110",
  44264=>"101100110",
  44265=>"011011111",
  44266=>"010110010",
  44267=>"100100100",
  44268=>"110000111",
  44269=>"101011101",
  44270=>"000001100",
  44271=>"111110011",
  44272=>"010001111",
  44273=>"000101101",
  44274=>"001001111",
  44275=>"011000001",
  44276=>"100110001",
  44277=>"100000000",
  44278=>"001110011",
  44279=>"110110000",
  44280=>"000001010",
  44281=>"101101100",
  44282=>"011111100",
  44283=>"001001000",
  44284=>"111011100",
  44285=>"011110110",
  44286=>"011000111",
  44287=>"111110111",
  44288=>"110100100",
  44289=>"011011001",
  44290=>"100000100",
  44291=>"011001000",
  44292=>"110111101",
  44293=>"001000100",
  44294=>"000001000",
  44295=>"011011011",
  44296=>"001100110",
  44297=>"110110001",
  44298=>"010011111",
  44299=>"100001100",
  44300=>"011010010",
  44301=>"110010011",
  44302=>"011110101",
  44303=>"001100101",
  44304=>"110101010",
  44305=>"010011100",
  44306=>"011101000",
  44307=>"110101000",
  44308=>"101000010",
  44309=>"001110001",
  44310=>"010000001",
  44311=>"011100001",
  44312=>"110011011",
  44313=>"101001110",
  44314=>"011101011",
  44315=>"000001011",
  44316=>"010001010",
  44317=>"100010001",
  44318=>"101111110",
  44319=>"001000110",
  44320=>"100010000",
  44321=>"100101011",
  44322=>"010001011",
  44323=>"001101111",
  44324=>"000001011",
  44325=>"010101111",
  44326=>"110110011",
  44327=>"001101101",
  44328=>"010100100",
  44329=>"000001111",
  44330=>"010010111",
  44331=>"110000110",
  44332=>"111110110",
  44333=>"111001100",
  44334=>"000011000",
  44335=>"111101100",
  44336=>"010010000",
  44337=>"101001110",
  44338=>"101111111",
  44339=>"000101110",
  44340=>"011011111",
  44341=>"101011101",
  44342=>"010101011",
  44343=>"010010001",
  44344=>"001010110",
  44345=>"111111011",
  44346=>"111111001",
  44347=>"011111001",
  44348=>"001100000",
  44349=>"011000100",
  44350=>"101000010",
  44351=>"010101100",
  44352=>"001001000",
  44353=>"100101101",
  44354=>"010010011",
  44355=>"001000001",
  44356=>"110111011",
  44357=>"100101000",
  44358=>"011111100",
  44359=>"100100001",
  44360=>"111111001",
  44361=>"100010110",
  44362=>"110011111",
  44363=>"111101000",
  44364=>"111100000",
  44365=>"000001110",
  44366=>"101110111",
  44367=>"100111110",
  44368=>"101001110",
  44369=>"001111111",
  44370=>"110100000",
  44371=>"111110011",
  44372=>"011011011",
  44373=>"101101001",
  44374=>"100111110",
  44375=>"010001110",
  44376=>"010010001",
  44377=>"111111111",
  44378=>"111110110",
  44379=>"001111100",
  44380=>"001000111",
  44381=>"111110100",
  44382=>"000111011",
  44383=>"001010000",
  44384=>"111110000",
  44385=>"101110010",
  44386=>"000000110",
  44387=>"010010000",
  44388=>"100011010",
  44389=>"010100001",
  44390=>"111011100",
  44391=>"010001100",
  44392=>"000111110",
  44393=>"010011101",
  44394=>"010111001",
  44395=>"110101101",
  44396=>"110000000",
  44397=>"000101111",
  44398=>"000000010",
  44399=>"011111111",
  44400=>"010011011",
  44401=>"011001011",
  44402=>"100000111",
  44403=>"111010100",
  44404=>"110111110",
  44405=>"001011101",
  44406=>"101101011",
  44407=>"111110101",
  44408=>"111100110",
  44409=>"000000011",
  44410=>"101011010",
  44411=>"011000001",
  44412=>"010111101",
  44413=>"001010000",
  44414=>"111010101",
  44415=>"000111001",
  44416=>"110100100",
  44417=>"101010100",
  44418=>"010011011",
  44419=>"010000000",
  44420=>"001101001",
  44421=>"111101111",
  44422=>"001101010",
  44423=>"111011111",
  44424=>"110100101",
  44425=>"010100111",
  44426=>"001111010",
  44427=>"111101100",
  44428=>"010010100",
  44429=>"100000011",
  44430=>"111010111",
  44431=>"111111100",
  44432=>"110000010",
  44433=>"010011111",
  44434=>"010100101",
  44435=>"010111110",
  44436=>"101011010",
  44437=>"001110011",
  44438=>"011000010",
  44439=>"011011011",
  44440=>"100001001",
  44441=>"000000010",
  44442=>"110101000",
  44443=>"010110111",
  44444=>"110101010",
  44445=>"000000001",
  44446=>"000010010",
  44447=>"110110000",
  44448=>"101101101",
  44449=>"001010010",
  44450=>"101110101",
  44451=>"010001000",
  44452=>"111011000",
  44453=>"000100001",
  44454=>"110101110",
  44455=>"010101001",
  44456=>"001111100",
  44457=>"110111101",
  44458=>"101101111",
  44459=>"100001101",
  44460=>"110101100",
  44461=>"111101001",
  44462=>"111101000",
  44463=>"000100111",
  44464=>"111111101",
  44465=>"000100101",
  44466=>"010110001",
  44467=>"000110111",
  44468=>"100001111",
  44469=>"000111100",
  44470=>"001001001",
  44471=>"100101101",
  44472=>"001000111",
  44473=>"010101110",
  44474=>"001010011",
  44475=>"001110000",
  44476=>"110010100",
  44477=>"010100000",
  44478=>"111011001",
  44479=>"000111101",
  44480=>"000111100",
  44481=>"100101011",
  44482=>"110001010",
  44483=>"011111100",
  44484=>"100000000",
  44485=>"010101010",
  44486=>"100101010",
  44487=>"111010110",
  44488=>"111000101",
  44489=>"101111110",
  44490=>"001001011",
  44491=>"000110100",
  44492=>"010001011",
  44493=>"010000000",
  44494=>"101011001",
  44495=>"011111001",
  44496=>"100010110",
  44497=>"010011010",
  44498=>"100010110",
  44499=>"101100011",
  44500=>"011111100",
  44501=>"100010000",
  44502=>"100001100",
  44503=>"001101110",
  44504=>"110000000",
  44505=>"111110111",
  44506=>"111111110",
  44507=>"001000101",
  44508=>"111000111",
  44509=>"111011110",
  44510=>"001110100",
  44511=>"111110010",
  44512=>"100010011",
  44513=>"110000010",
  44514=>"110101011",
  44515=>"110111001",
  44516=>"001100000",
  44517=>"100110101",
  44518=>"110000011",
  44519=>"000101001",
  44520=>"000111111",
  44521=>"010111001",
  44522=>"101001000",
  44523=>"100110011",
  44524=>"111111111",
  44525=>"101000011",
  44526=>"001000011",
  44527=>"101100011",
  44528=>"110101010",
  44529=>"101001001",
  44530=>"101011111",
  44531=>"011110000",
  44532=>"000000010",
  44533=>"000100110",
  44534=>"101100000",
  44535=>"110001010",
  44536=>"111111011",
  44537=>"010101100",
  44538=>"011001111",
  44539=>"101111010",
  44540=>"100101011",
  44541=>"000011101",
  44542=>"010100101",
  44543=>"111110111",
  44544=>"010011100",
  44545=>"100110000",
  44546=>"001010111",
  44547=>"110101011",
  44548=>"101011110",
  44549=>"011100010",
  44550=>"100011011",
  44551=>"011111001",
  44552=>"010100110",
  44553=>"001111111",
  44554=>"000000111",
  44555=>"001100000",
  44556=>"001111010",
  44557=>"001110010",
  44558=>"000111010",
  44559=>"011101010",
  44560=>"011000010",
  44561=>"111000110",
  44562=>"000001010",
  44563=>"111101111",
  44564=>"011001001",
  44565=>"111101001",
  44566=>"101001101",
  44567=>"001010001",
  44568=>"100110111",
  44569=>"011111101",
  44570=>"010001010",
  44571=>"110010110",
  44572=>"010000010",
  44573=>"110110010",
  44574=>"110111011",
  44575=>"110010000",
  44576=>"110001001",
  44577=>"100010011",
  44578=>"011101001",
  44579=>"110110010",
  44580=>"101010111",
  44581=>"001000111",
  44582=>"001111000",
  44583=>"010001111",
  44584=>"100110111",
  44585=>"111001000",
  44586=>"011100000",
  44587=>"100001101",
  44588=>"000100111",
  44589=>"000001010",
  44590=>"001110100",
  44591=>"100001100",
  44592=>"111101110",
  44593=>"110100100",
  44594=>"100111101",
  44595=>"110111000",
  44596=>"001111011",
  44597=>"100110111",
  44598=>"010000001",
  44599=>"111101101",
  44600=>"001010001",
  44601=>"001000111",
  44602=>"111110011",
  44603=>"100111100",
  44604=>"111101000",
  44605=>"001100110",
  44606=>"111001111",
  44607=>"101100010",
  44608=>"001100000",
  44609=>"101101101",
  44610=>"000010011",
  44611=>"011111010",
  44612=>"101101101",
  44613=>"010100010",
  44614=>"010000111",
  44615=>"001010110",
  44616=>"000110011",
  44617=>"010110010",
  44618=>"010000011",
  44619=>"000011111",
  44620=>"110100110",
  44621=>"101001011",
  44622=>"110001000",
  44623=>"101001111",
  44624=>"011011010",
  44625=>"100111110",
  44626=>"101111100",
  44627=>"101101100",
  44628=>"000100111",
  44629=>"101111101",
  44630=>"010010000",
  44631=>"101010001",
  44632=>"000011010",
  44633=>"001100111",
  44634=>"100000001",
  44635=>"011110010",
  44636=>"101000001",
  44637=>"101101111",
  44638=>"101110110",
  44639=>"111110111",
  44640=>"000110001",
  44641=>"100101011",
  44642=>"000101000",
  44643=>"100000100",
  44644=>"001100010",
  44645=>"110011101",
  44646=>"010000010",
  44647=>"000111111",
  44648=>"111011010",
  44649=>"100000110",
  44650=>"110001000",
  44651=>"111101110",
  44652=>"000110000",
  44653=>"101000001",
  44654=>"001101101",
  44655=>"000110110",
  44656=>"001011011",
  44657=>"111111001",
  44658=>"010000000",
  44659=>"101101110",
  44660=>"010011000",
  44661=>"110010000",
  44662=>"111010110",
  44663=>"100001010",
  44664=>"111001111",
  44665=>"101001001",
  44666=>"011000010",
  44667=>"011111000",
  44668=>"111001010",
  44669=>"100010001",
  44670=>"011110100",
  44671=>"010011000",
  44672=>"001001110",
  44673=>"100001101",
  44674=>"010001110",
  44675=>"010110100",
  44676=>"001101010",
  44677=>"100000010",
  44678=>"001011010",
  44679=>"011000010",
  44680=>"111010001",
  44681=>"001101111",
  44682=>"101111011",
  44683=>"010010010",
  44684=>"100001110",
  44685=>"100110001",
  44686=>"001100010",
  44687=>"100100110",
  44688=>"100000010",
  44689=>"010001110",
  44690=>"000110101",
  44691=>"100001000",
  44692=>"100111010",
  44693=>"110110001",
  44694=>"010010110",
  44695=>"101111111",
  44696=>"111110110",
  44697=>"000000010",
  44698=>"100010110",
  44699=>"101101010",
  44700=>"111101001",
  44701=>"101110101",
  44702=>"010000000",
  44703=>"110011101",
  44704=>"001000010",
  44705=>"010010101",
  44706=>"110101111",
  44707=>"111100100",
  44708=>"110010010",
  44709=>"001100001",
  44710=>"110010001",
  44711=>"000111010",
  44712=>"001101001",
  44713=>"001101100",
  44714=>"000110110",
  44715=>"011001111",
  44716=>"110101011",
  44717=>"101111001",
  44718=>"100000100",
  44719=>"000000100",
  44720=>"001100011",
  44721=>"000100101",
  44722=>"011110101",
  44723=>"101100111",
  44724=>"110001111",
  44725=>"100010000",
  44726=>"111001000",
  44727=>"110100010",
  44728=>"001001110",
  44729=>"110100001",
  44730=>"111001001",
  44731=>"101001001",
  44732=>"100010100",
  44733=>"101111011",
  44734=>"101100001",
  44735=>"000100111",
  44736=>"000000010",
  44737=>"100111010",
  44738=>"110001111",
  44739=>"100100111",
  44740=>"010000110",
  44741=>"001001001",
  44742=>"111100110",
  44743=>"001100110",
  44744=>"111011001",
  44745=>"100100101",
  44746=>"100001000",
  44747=>"010110001",
  44748=>"001100011",
  44749=>"001101010",
  44750=>"010111011",
  44751=>"011100100",
  44752=>"010111001",
  44753=>"011000001",
  44754=>"000000001",
  44755=>"011001010",
  44756=>"101101010",
  44757=>"010011101",
  44758=>"001101011",
  44759=>"101001010",
  44760=>"011000101",
  44761=>"110110001",
  44762=>"111011111",
  44763=>"100100111",
  44764=>"001000000",
  44765=>"001010010",
  44766=>"111011110",
  44767=>"101001111",
  44768=>"111111110",
  44769=>"000000101",
  44770=>"100100001",
  44771=>"011010111",
  44772=>"001100000",
  44773=>"011101001",
  44774=>"110011110",
  44775=>"101111111",
  44776=>"110010111",
  44777=>"101111110",
  44778=>"001100011",
  44779=>"001000000",
  44780=>"010110101",
  44781=>"011000011",
  44782=>"000001111",
  44783=>"011110110",
  44784=>"000011101",
  44785=>"001101011",
  44786=>"110010001",
  44787=>"111110110",
  44788=>"110110011",
  44789=>"111100000",
  44790=>"001000110",
  44791=>"011111100",
  44792=>"000001110",
  44793=>"001001001",
  44794=>"001011000",
  44795=>"001111010",
  44796=>"110010100",
  44797=>"111100010",
  44798=>"001011010",
  44799=>"010010011",
  44800=>"100000011",
  44801=>"101000101",
  44802=>"101000111",
  44803=>"101000001",
  44804=>"011101110",
  44805=>"100000111",
  44806=>"101110000",
  44807=>"101101001",
  44808=>"010001010",
  44809=>"011010110",
  44810=>"011111011",
  44811=>"001101110",
  44812=>"100101101",
  44813=>"100011101",
  44814=>"011010001",
  44815=>"100101100",
  44816=>"100101000",
  44817=>"011100110",
  44818=>"101000101",
  44819=>"100000000",
  44820=>"101001101",
  44821=>"110011100",
  44822=>"011111100",
  44823=>"100001101",
  44824=>"001111010",
  44825=>"010010111",
  44826=>"101000011",
  44827=>"100110010",
  44828=>"111011000",
  44829=>"010010011",
  44830=>"000001010",
  44831=>"000001001",
  44832=>"001111111",
  44833=>"110101001",
  44834=>"011101111",
  44835=>"111000000",
  44836=>"100100011",
  44837=>"101100110",
  44838=>"000000110",
  44839=>"011111001",
  44840=>"111001101",
  44841=>"100001010",
  44842=>"111010100",
  44843=>"111100000",
  44844=>"001100011",
  44845=>"011100000",
  44846=>"000110010",
  44847=>"111011111",
  44848=>"100101010",
  44849=>"110101001",
  44850=>"110000101",
  44851=>"010011101",
  44852=>"011101000",
  44853=>"110110110",
  44854=>"100110000",
  44855=>"100111000",
  44856=>"001000110",
  44857=>"111010100",
  44858=>"000000111",
  44859=>"110101001",
  44860=>"001000100",
  44861=>"000001010",
  44862=>"111101001",
  44863=>"111110110",
  44864=>"001010101",
  44865=>"011000000",
  44866=>"010101100",
  44867=>"110011011",
  44868=>"001110001",
  44869=>"010101110",
  44870=>"100000001",
  44871=>"011111001",
  44872=>"100000010",
  44873=>"101000010",
  44874=>"111011100",
  44875=>"110101100",
  44876=>"111001101",
  44877=>"110010101",
  44878=>"100010111",
  44879=>"011010011",
  44880=>"110100110",
  44881=>"000010100",
  44882=>"111000101",
  44883=>"010101010",
  44884=>"011001101",
  44885=>"011001001",
  44886=>"100001100",
  44887=>"001001011",
  44888=>"011111100",
  44889=>"101000000",
  44890=>"000001000",
  44891=>"000111101",
  44892=>"101110110",
  44893=>"000101010",
  44894=>"100001001",
  44895=>"111100001",
  44896=>"111100110",
  44897=>"001000100",
  44898=>"000000111",
  44899=>"101110100",
  44900=>"000000010",
  44901=>"010101111",
  44902=>"000101100",
  44903=>"100000010",
  44904=>"100011000",
  44905=>"100101100",
  44906=>"011111110",
  44907=>"101011010",
  44908=>"001001000",
  44909=>"100111000",
  44910=>"010010010",
  44911=>"011100000",
  44912=>"111100001",
  44913=>"111011000",
  44914=>"001101011",
  44915=>"000001110",
  44916=>"110010011",
  44917=>"000000111",
  44918=>"111111011",
  44919=>"101100000",
  44920=>"010000000",
  44921=>"100000001",
  44922=>"100111111",
  44923=>"001000111",
  44924=>"100100100",
  44925=>"111111101",
  44926=>"010110101",
  44927=>"010001001",
  44928=>"000101010",
  44929=>"000000001",
  44930=>"100001010",
  44931=>"010100100",
  44932=>"011010101",
  44933=>"111111100",
  44934=>"100111000",
  44935=>"010101111",
  44936=>"011100000",
  44937=>"000101111",
  44938=>"111101110",
  44939=>"110011110",
  44940=>"100001011",
  44941=>"101111111",
  44942=>"111101000",
  44943=>"101111000",
  44944=>"111111111",
  44945=>"101000000",
  44946=>"001111000",
  44947=>"111110110",
  44948=>"101110001",
  44949=>"100001010",
  44950=>"100110100",
  44951=>"111111000",
  44952=>"101010001",
  44953=>"111001000",
  44954=>"011010000",
  44955=>"111111111",
  44956=>"000110011",
  44957=>"100010111",
  44958=>"000010001",
  44959=>"011110110",
  44960=>"011010111",
  44961=>"000000000",
  44962=>"001001101",
  44963=>"101110111",
  44964=>"011111011",
  44965=>"101111010",
  44966=>"011101000",
  44967=>"000001111",
  44968=>"101101010",
  44969=>"111000010",
  44970=>"101111001",
  44971=>"001100010",
  44972=>"011011011",
  44973=>"111000010",
  44974=>"101111111",
  44975=>"100000011",
  44976=>"101100000",
  44977=>"110100001",
  44978=>"110011111",
  44979=>"101010010",
  44980=>"001111010",
  44981=>"111001010",
  44982=>"000100110",
  44983=>"111101001",
  44984=>"000101001",
  44985=>"110111011",
  44986=>"000110011",
  44987=>"000101111",
  44988=>"101111010",
  44989=>"111100010",
  44990=>"011011000",
  44991=>"000001010",
  44992=>"101100111",
  44993=>"100111011",
  44994=>"111110000",
  44995=>"100110010",
  44996=>"100110101",
  44997=>"111000010",
  44998=>"010001000",
  44999=>"011100101",
  45000=>"110000000",
  45001=>"000101101",
  45002=>"000100111",
  45003=>"111110111",
  45004=>"100000010",
  45005=>"000011100",
  45006=>"110011000",
  45007=>"100110010",
  45008=>"100101000",
  45009=>"001001010",
  45010=>"010000110",
  45011=>"000010100",
  45012=>"110111111",
  45013=>"010001111",
  45014=>"100001010",
  45015=>"010001000",
  45016=>"111001101",
  45017=>"000001101",
  45018=>"010110111",
  45019=>"001101011",
  45020=>"001011001",
  45021=>"000111001",
  45022=>"000101100",
  45023=>"001010001",
  45024=>"110111000",
  45025=>"100100001",
  45026=>"011001110",
  45027=>"110111101",
  45028=>"111101101",
  45029=>"011010011",
  45030=>"111000100",
  45031=>"111000001",
  45032=>"100001110",
  45033=>"011010011",
  45034=>"101101000",
  45035=>"000010011",
  45036=>"110101100",
  45037=>"010001010",
  45038=>"101011111",
  45039=>"011010100",
  45040=>"001111111",
  45041=>"110011000",
  45042=>"011101010",
  45043=>"101101111",
  45044=>"010101111",
  45045=>"011011000",
  45046=>"010101001",
  45047=>"011101101",
  45048=>"110110101",
  45049=>"000010100",
  45050=>"000011011",
  45051=>"101100000",
  45052=>"000110001",
  45053=>"010101011",
  45054=>"000011000",
  45055=>"110011111",
  45056=>"111101001",
  45057=>"101011111",
  45058=>"010010001",
  45059=>"110010111",
  45060=>"111011111",
  45061=>"100010111",
  45062=>"001001101",
  45063=>"010111100",
  45064=>"100111110",
  45065=>"100100110",
  45066=>"000100000",
  45067=>"001111100",
  45068=>"010111101",
  45069=>"110000011",
  45070=>"100000110",
  45071=>"110101011",
  45072=>"101101110",
  45073=>"001000100",
  45074=>"000011011",
  45075=>"011110101",
  45076=>"000000100",
  45077=>"111011010",
  45078=>"100101101",
  45079=>"010011100",
  45080=>"010000101",
  45081=>"111010110",
  45082=>"101010011",
  45083=>"101100001",
  45084=>"000001000",
  45085=>"011101000",
  45086=>"011000101",
  45087=>"000101110",
  45088=>"010100111",
  45089=>"100110111",
  45090=>"011100001",
  45091=>"000010111",
  45092=>"010011100",
  45093=>"100100000",
  45094=>"010010111",
  45095=>"010010101",
  45096=>"000100101",
  45097=>"110000010",
  45098=>"111010101",
  45099=>"011001000",
  45100=>"111111001",
  45101=>"001000011",
  45102=>"011011011",
  45103=>"001011111",
  45104=>"011000100",
  45105=>"100011100",
  45106=>"011001000",
  45107=>"001101001",
  45108=>"110100101",
  45109=>"011000001",
  45110=>"111011010",
  45111=>"000110010",
  45112=>"100001110",
  45113=>"000001111",
  45114=>"100101001",
  45115=>"000010101",
  45116=>"010101110",
  45117=>"101100010",
  45118=>"111101101",
  45119=>"011001110",
  45120=>"111100110",
  45121=>"001010001",
  45122=>"111001010",
  45123=>"101101100",
  45124=>"111111111",
  45125=>"000110100",
  45126=>"001000000",
  45127=>"010000001",
  45128=>"110111001",
  45129=>"000111111",
  45130=>"100001100",
  45131=>"111110000",
  45132=>"001101010",
  45133=>"001001000",
  45134=>"000101000",
  45135=>"001111111",
  45136=>"111010101",
  45137=>"111011001",
  45138=>"100001000",
  45139=>"111110010",
  45140=>"010111110",
  45141=>"000100000",
  45142=>"100001011",
  45143=>"100100101",
  45144=>"101001111",
  45145=>"110011010",
  45146=>"011100010",
  45147=>"101101101",
  45148=>"001011000",
  45149=>"000001000",
  45150=>"000110110",
  45151=>"010101001",
  45152=>"000100110",
  45153=>"110110000",
  45154=>"110110010",
  45155=>"000011101",
  45156=>"110111101",
  45157=>"000100111",
  45158=>"100011000",
  45159=>"111000001",
  45160=>"010001010",
  45161=>"001001001",
  45162=>"011101000",
  45163=>"110110001",
  45164=>"100111101",
  45165=>"000011010",
  45166=>"011110010",
  45167=>"111111011",
  45168=>"100111101",
  45169=>"111110100",
  45170=>"111000111",
  45171=>"000110111",
  45172=>"000011011",
  45173=>"000101001",
  45174=>"011011010",
  45175=>"011001101",
  45176=>"000001001",
  45177=>"000110010",
  45178=>"011101110",
  45179=>"000010011",
  45180=>"001001001",
  45181=>"111110010",
  45182=>"100010111",
  45183=>"000001101",
  45184=>"111100110",
  45185=>"001100101",
  45186=>"111001100",
  45187=>"001100011",
  45188=>"111001011",
  45189=>"111010110",
  45190=>"111010110",
  45191=>"010111011",
  45192=>"111000001",
  45193=>"001000000",
  45194=>"001010100",
  45195=>"010110000",
  45196=>"101100001",
  45197=>"111110000",
  45198=>"101011000",
  45199=>"011111010",
  45200=>"001110101",
  45201=>"110100110",
  45202=>"000110000",
  45203=>"000111001",
  45204=>"111000111",
  45205=>"000011111",
  45206=>"011001100",
  45207=>"001100110",
  45208=>"001010111",
  45209=>"000110000",
  45210=>"000101001",
  45211=>"101100111",
  45212=>"100010001",
  45213=>"010100011",
  45214=>"000100011",
  45215=>"000001110",
  45216=>"101011111",
  45217=>"011011111",
  45218=>"111100001",
  45219=>"111000101",
  45220=>"010000010",
  45221=>"000011111",
  45222=>"010000011",
  45223=>"111001101",
  45224=>"010101000",
  45225=>"100101110",
  45226=>"111011101",
  45227=>"101011101",
  45228=>"001111100",
  45229=>"100110100",
  45230=>"100111000",
  45231=>"110101111",
  45232=>"000100110",
  45233=>"000001010",
  45234=>"001001111",
  45235=>"001010010",
  45236=>"000101111",
  45237=>"001011100",
  45238=>"111100010",
  45239=>"000101010",
  45240=>"101010011",
  45241=>"011001110",
  45242=>"001000100",
  45243=>"100101011",
  45244=>"010010100",
  45245=>"101000100",
  45246=>"001011101",
  45247=>"100110010",
  45248=>"000110010",
  45249=>"011111000",
  45250=>"110111100",
  45251=>"001010001",
  45252=>"010100001",
  45253=>"000001101",
  45254=>"010100101",
  45255=>"100011100",
  45256=>"110111100",
  45257=>"100010110",
  45258=>"000011011",
  45259=>"001000010",
  45260=>"011001011",
  45261=>"111111101",
  45262=>"010110001",
  45263=>"010100000",
  45264=>"010010001",
  45265=>"010101101",
  45266=>"010100000",
  45267=>"111000001",
  45268=>"110110110",
  45269=>"101110111",
  45270=>"101111011",
  45271=>"001011110",
  45272=>"101100001",
  45273=>"111011011",
  45274=>"110001001",
  45275=>"001110100",
  45276=>"110101110",
  45277=>"011011101",
  45278=>"000111110",
  45279=>"100100011",
  45280=>"101011110",
  45281=>"111001010",
  45282=>"100110010",
  45283=>"110011110",
  45284=>"110101000",
  45285=>"111000010",
  45286=>"010101011",
  45287=>"101111111",
  45288=>"010111000",
  45289=>"111111100",
  45290=>"101100011",
  45291=>"110010100",
  45292=>"100111110",
  45293=>"101101011",
  45294=>"000001110",
  45295=>"010010000",
  45296=>"010101001",
  45297=>"111110000",
  45298=>"000101000",
  45299=>"100001000",
  45300=>"000001100",
  45301=>"001110111",
  45302=>"100001101",
  45303=>"010111111",
  45304=>"111101011",
  45305=>"001100010",
  45306=>"100110100",
  45307=>"000110100",
  45308=>"011010010",
  45309=>"011010101",
  45310=>"000000001",
  45311=>"011101010",
  45312=>"111001111",
  45313=>"001011010",
  45314=>"101110100",
  45315=>"011111000",
  45316=>"000111010",
  45317=>"100111000",
  45318=>"101001010",
  45319=>"100011000",
  45320=>"110000000",
  45321=>"100011101",
  45322=>"000101100",
  45323=>"111101110",
  45324=>"011000100",
  45325=>"100010100",
  45326=>"000001010",
  45327=>"101000101",
  45328=>"000011110",
  45329=>"000000000",
  45330=>"111101110",
  45331=>"001101110",
  45332=>"010010110",
  45333=>"100011010",
  45334=>"001000101",
  45335=>"000101111",
  45336=>"000001011",
  45337=>"010011011",
  45338=>"010100010",
  45339=>"100011100",
  45340=>"100000100",
  45341=>"001001011",
  45342=>"011110011",
  45343=>"111000111",
  45344=>"001011100",
  45345=>"001010111",
  45346=>"111010011",
  45347=>"011110110",
  45348=>"110001010",
  45349=>"001001001",
  45350=>"010010010",
  45351=>"110001000",
  45352=>"001111101",
  45353=>"000010101",
  45354=>"101000101",
  45355=>"011100000",
  45356=>"010001010",
  45357=>"000001000",
  45358=>"110100111",
  45359=>"101111010",
  45360=>"100101011",
  45361=>"101100111",
  45362=>"100001010",
  45363=>"110111001",
  45364=>"111111010",
  45365=>"011010010",
  45366=>"000110001",
  45367=>"110111110",
  45368=>"000000000",
  45369=>"000110111",
  45370=>"010111100",
  45371=>"000011011",
  45372=>"000011110",
  45373=>"110100100",
  45374=>"110100011",
  45375=>"011100111",
  45376=>"100001010",
  45377=>"110100000",
  45378=>"000011000",
  45379=>"000111101",
  45380=>"111110100",
  45381=>"010011100",
  45382=>"000000100",
  45383=>"000011100",
  45384=>"101000110",
  45385=>"000011010",
  45386=>"010110111",
  45387=>"010100111",
  45388=>"101010110",
  45389=>"111011011",
  45390=>"001000011",
  45391=>"101100001",
  45392=>"101000010",
  45393=>"000111011",
  45394=>"101100111",
  45395=>"100110001",
  45396=>"101101000",
  45397=>"100011011",
  45398=>"000011010",
  45399=>"101010111",
  45400=>"110000100",
  45401=>"100011111",
  45402=>"110100110",
  45403=>"111111110",
  45404=>"110101110",
  45405=>"011001000",
  45406=>"111000001",
  45407=>"110000111",
  45408=>"001000011",
  45409=>"111111110",
  45410=>"011110111",
  45411=>"110000011",
  45412=>"000100011",
  45413=>"001101000",
  45414=>"000011110",
  45415=>"011001001",
  45416=>"011000011",
  45417=>"111010010",
  45418=>"001101000",
  45419=>"110100010",
  45420=>"010000101",
  45421=>"010001111",
  45422=>"001010110",
  45423=>"011101101",
  45424=>"000101001",
  45425=>"111101001",
  45426=>"000100010",
  45427=>"111111111",
  45428=>"100111001",
  45429=>"000110001",
  45430=>"000000011",
  45431=>"101001111",
  45432=>"011101110",
  45433=>"000001111",
  45434=>"101010110",
  45435=>"001111101",
  45436=>"001011010",
  45437=>"000000110",
  45438=>"001001000",
  45439=>"010011100",
  45440=>"000011001",
  45441=>"000001100",
  45442=>"010100000",
  45443=>"100011111",
  45444=>"001001010",
  45445=>"111001001",
  45446=>"110100110",
  45447=>"101111100",
  45448=>"100101101",
  45449=>"011100011",
  45450=>"011001011",
  45451=>"011011110",
  45452=>"100000100",
  45453=>"001000110",
  45454=>"110011111",
  45455=>"101101011",
  45456=>"110110001",
  45457=>"101001100",
  45458=>"111011000",
  45459=>"100011101",
  45460=>"100110000",
  45461=>"011100110",
  45462=>"010111000",
  45463=>"011101100",
  45464=>"011100001",
  45465=>"101000110",
  45466=>"010111010",
  45467=>"001110011",
  45468=>"001101101",
  45469=>"010001011",
  45470=>"101010101",
  45471=>"001101101",
  45472=>"110011000",
  45473=>"010011110",
  45474=>"101110000",
  45475=>"010101001",
  45476=>"010000110",
  45477=>"001000011",
  45478=>"100111010",
  45479=>"101000111",
  45480=>"000011011",
  45481=>"101111100",
  45482=>"110001000",
  45483=>"000010001",
  45484=>"100010100",
  45485=>"000101000",
  45486=>"000101000",
  45487=>"010011111",
  45488=>"100100001",
  45489=>"001111110",
  45490=>"111101000",
  45491=>"011111111",
  45492=>"001110101",
  45493=>"110010100",
  45494=>"111111000",
  45495=>"101101100",
  45496=>"100100001",
  45497=>"000000011",
  45498=>"101011111",
  45499=>"101000101",
  45500=>"001111000",
  45501=>"001000101",
  45502=>"101001000",
  45503=>"110110111",
  45504=>"111000000",
  45505=>"100010010",
  45506=>"001001001",
  45507=>"100110000",
  45508=>"111101011",
  45509=>"010010101",
  45510=>"010100000",
  45511=>"000001000",
  45512=>"001100000",
  45513=>"101100010",
  45514=>"111101100",
  45515=>"111101110",
  45516=>"010111000",
  45517=>"101110001",
  45518=>"000000011",
  45519=>"001011100",
  45520=>"000111011",
  45521=>"101101111",
  45522=>"000101110",
  45523=>"000111001",
  45524=>"100001000",
  45525=>"100000111",
  45526=>"001110001",
  45527=>"100001100",
  45528=>"110000001",
  45529=>"111101011",
  45530=>"000011001",
  45531=>"000001100",
  45532=>"000010000",
  45533=>"010110010",
  45534=>"100001011",
  45535=>"011000101",
  45536=>"100011111",
  45537=>"010001111",
  45538=>"101010110",
  45539=>"100110001",
  45540=>"010110001",
  45541=>"110100001",
  45542=>"000100010",
  45543=>"000000011",
  45544=>"111111101",
  45545=>"000111011",
  45546=>"111100000",
  45547=>"010010111",
  45548=>"000111110",
  45549=>"011111101",
  45550=>"100010110",
  45551=>"100100001",
  45552=>"111010011",
  45553=>"101111101",
  45554=>"111110110",
  45555=>"011010110",
  45556=>"111001101",
  45557=>"111011000",
  45558=>"000110100",
  45559=>"010010001",
  45560=>"111011001",
  45561=>"110011110",
  45562=>"011010100",
  45563=>"100000011",
  45564=>"000110110",
  45565=>"011111000",
  45566=>"110111111",
  45567=>"100100111",
  45568=>"011000010",
  45569=>"100110011",
  45570=>"100001011",
  45571=>"110110010",
  45572=>"000010110",
  45573=>"100111101",
  45574=>"001010000",
  45575=>"000110000",
  45576=>"111111011",
  45577=>"011000101",
  45578=>"010011111",
  45579=>"111101100",
  45580=>"000110100",
  45581=>"101101110",
  45582=>"001101010",
  45583=>"100011011",
  45584=>"001111000",
  45585=>"010010010",
  45586=>"010011110",
  45587=>"111101011",
  45588=>"000100110",
  45589=>"110001111",
  45590=>"001100100",
  45591=>"100010110",
  45592=>"101111110",
  45593=>"100111111",
  45594=>"001111100",
  45595=>"001111011",
  45596=>"011110100",
  45597=>"101100000",
  45598=>"100001111",
  45599=>"100101010",
  45600=>"001101110",
  45601=>"100100100",
  45602=>"000010101",
  45603=>"010100000",
  45604=>"110000010",
  45605=>"111001111",
  45606=>"001101001",
  45607=>"000101100",
  45608=>"010101011",
  45609=>"100000000",
  45610=>"100111011",
  45611=>"111010011",
  45612=>"010111001",
  45613=>"101100110",
  45614=>"101000001",
  45615=>"110011101",
  45616=>"011010101",
  45617=>"100010111",
  45618=>"000100101",
  45619=>"110001001",
  45620=>"111010011",
  45621=>"111100001",
  45622=>"001101001",
  45623=>"011101011",
  45624=>"010010001",
  45625=>"111010110",
  45626=>"001010001",
  45627=>"000110000",
  45628=>"111000001",
  45629=>"101111101",
  45630=>"100101001",
  45631=>"010001111",
  45632=>"010001000",
  45633=>"011110001",
  45634=>"000001011",
  45635=>"010000001",
  45636=>"111010110",
  45637=>"110101100",
  45638=>"010010110",
  45639=>"100011000",
  45640=>"011011111",
  45641=>"111100000",
  45642=>"011011001",
  45643=>"101011011",
  45644=>"110101001",
  45645=>"000010111",
  45646=>"111011100",
  45647=>"000000010",
  45648=>"100101101",
  45649=>"101010010",
  45650=>"000100000",
  45651=>"000111001",
  45652=>"110110001",
  45653=>"100010000",
  45654=>"000011100",
  45655=>"011011010",
  45656=>"111100001",
  45657=>"110111000",
  45658=>"011101010",
  45659=>"100011111",
  45660=>"101110101",
  45661=>"010000110",
  45662=>"001001011",
  45663=>"001111000",
  45664=>"001010011",
  45665=>"010111111",
  45666=>"100110000",
  45667=>"101001100",
  45668=>"010101010",
  45669=>"101000111",
  45670=>"101110110",
  45671=>"011011010",
  45672=>"010111000",
  45673=>"010010010",
  45674=>"000101111",
  45675=>"001110100",
  45676=>"100010001",
  45677=>"001111100",
  45678=>"011000111",
  45679=>"010010100",
  45680=>"100100110",
  45681=>"000110111",
  45682=>"110111100",
  45683=>"011010111",
  45684=>"000010110",
  45685=>"000101001",
  45686=>"001111111",
  45687=>"011110100",
  45688=>"011000001",
  45689=>"001100111",
  45690=>"001000100",
  45691=>"110100110",
  45692=>"101011111",
  45693=>"101010110",
  45694=>"100000001",
  45695=>"111111101",
  45696=>"001001100",
  45697=>"110011011",
  45698=>"100110011",
  45699=>"000101101",
  45700=>"100010011",
  45701=>"101101111",
  45702=>"101101110",
  45703=>"100110110",
  45704=>"100110001",
  45705=>"110111101",
  45706=>"010111101",
  45707=>"001011010",
  45708=>"010000111",
  45709=>"000011000",
  45710=>"101101111",
  45711=>"010011110",
  45712=>"111000001",
  45713=>"010110000",
  45714=>"001011100",
  45715=>"000100111",
  45716=>"110101111",
  45717=>"100000111",
  45718=>"100110010",
  45719=>"001101110",
  45720=>"111011011",
  45721=>"110101110",
  45722=>"010000011",
  45723=>"011000111",
  45724=>"000101001",
  45725=>"011011101",
  45726=>"001100000",
  45727=>"001001010",
  45728=>"010010100",
  45729=>"100001110",
  45730=>"001000010",
  45731=>"001011111",
  45732=>"110001111",
  45733=>"110111100",
  45734=>"010010000",
  45735=>"011011010",
  45736=>"001110010",
  45737=>"110010000",
  45738=>"100100111",
  45739=>"101100100",
  45740=>"000101001",
  45741=>"110111110",
  45742=>"100100011",
  45743=>"011000011",
  45744=>"000100001",
  45745=>"010010110",
  45746=>"010001010",
  45747=>"001001000",
  45748=>"000000000",
  45749=>"011000101",
  45750=>"100110011",
  45751=>"000111000",
  45752=>"000100010",
  45753=>"111000001",
  45754=>"111111010",
  45755=>"111101010",
  45756=>"110010011",
  45757=>"001000100",
  45758=>"101010010",
  45759=>"000110101",
  45760=>"001100000",
  45761=>"111001000",
  45762=>"111101011",
  45763=>"010110001",
  45764=>"000101000",
  45765=>"001111111",
  45766=>"110001010",
  45767=>"100001001",
  45768=>"110111110",
  45769=>"000110000",
  45770=>"100001111",
  45771=>"101000001",
  45772=>"011101101",
  45773=>"100001011",
  45774=>"100010010",
  45775=>"111110000",
  45776=>"100011110",
  45777=>"101101111",
  45778=>"000111110",
  45779=>"011101001",
  45780=>"011011101",
  45781=>"111011111",
  45782=>"110000011",
  45783=>"001101010",
  45784=>"011011111",
  45785=>"011000111",
  45786=>"110011010",
  45787=>"101000010",
  45788=>"111011101",
  45789=>"010101010",
  45790=>"110110101",
  45791=>"000001011",
  45792=>"000011110",
  45793=>"111000000",
  45794=>"100000011",
  45795=>"000111010",
  45796=>"101010111",
  45797=>"100110001",
  45798=>"100011101",
  45799=>"010000001",
  45800=>"001001000",
  45801=>"100011101",
  45802=>"110011001",
  45803=>"010010001",
  45804=>"100000110",
  45805=>"011000100",
  45806=>"001011011",
  45807=>"101100000",
  45808=>"110001111",
  45809=>"000101000",
  45810=>"011000010",
  45811=>"111011011",
  45812=>"100110111",
  45813=>"010100101",
  45814=>"001100011",
  45815=>"011011111",
  45816=>"010011100",
  45817=>"110001000",
  45818=>"000001111",
  45819=>"100001001",
  45820=>"000111000",
  45821=>"101101010",
  45822=>"100101011",
  45823=>"001111100",
  45824=>"101010110",
  45825=>"110110011",
  45826=>"100101000",
  45827=>"100001101",
  45828=>"101011111",
  45829=>"010100001",
  45830=>"001101001",
  45831=>"000100111",
  45832=>"010011010",
  45833=>"111000100",
  45834=>"111111111",
  45835=>"000000010",
  45836=>"001111000",
  45837=>"000110001",
  45838=>"100100111",
  45839=>"110000000",
  45840=>"111110000",
  45841=>"100100110",
  45842=>"111011011",
  45843=>"001110010",
  45844=>"101110101",
  45845=>"100010000",
  45846=>"100010001",
  45847=>"001110010",
  45848=>"000101011",
  45849=>"001000101",
  45850=>"100111101",
  45851=>"011110011",
  45852=>"011011101",
  45853=>"111111101",
  45854=>"110001101",
  45855=>"101011011",
  45856=>"011101000",
  45857=>"000011100",
  45858=>"000010110",
  45859=>"001000000",
  45860=>"111101011",
  45861=>"110001010",
  45862=>"100111100",
  45863=>"101100101",
  45864=>"001111110",
  45865=>"001000001",
  45866=>"111100110",
  45867=>"101011000",
  45868=>"101000111",
  45869=>"001101101",
  45870=>"011101101",
  45871=>"110010111",
  45872=>"000100101",
  45873=>"001100010",
  45874=>"011110011",
  45875=>"010011000",
  45876=>"101001000",
  45877=>"001101100",
  45878=>"111110010",
  45879=>"111001111",
  45880=>"111100101",
  45881=>"011110101",
  45882=>"101100000",
  45883=>"001111111",
  45884=>"011111010",
  45885=>"000100000",
  45886=>"111101101",
  45887=>"000000110",
  45888=>"101111001",
  45889=>"001110011",
  45890=>"000011111",
  45891=>"110101110",
  45892=>"000001101",
  45893=>"111100001",
  45894=>"110110010",
  45895=>"111001110",
  45896=>"101000011",
  45897=>"000100110",
  45898=>"010010000",
  45899=>"010100010",
  45900=>"110000101",
  45901=>"010000111",
  45902=>"000111100",
  45903=>"001011100",
  45904=>"011111100",
  45905=>"101100101",
  45906=>"100101110",
  45907=>"000110000",
  45908=>"011011110",
  45909=>"011101000",
  45910=>"000000110",
  45911=>"100000100",
  45912=>"100001101",
  45913=>"100000100",
  45914=>"010010011",
  45915=>"100101110",
  45916=>"100001001",
  45917=>"010111000",
  45918=>"001000000",
  45919=>"101100000",
  45920=>"011111111",
  45921=>"111001001",
  45922=>"000100010",
  45923=>"101000000",
  45924=>"101010110",
  45925=>"011000000",
  45926=>"000100011",
  45927=>"111101010",
  45928=>"111010011",
  45929=>"001100001",
  45930=>"001100101",
  45931=>"010111001",
  45932=>"001011010",
  45933=>"110101000",
  45934=>"110011100",
  45935=>"110101010",
  45936=>"010101010",
  45937=>"010001011",
  45938=>"110010100",
  45939=>"010101110",
  45940=>"100110011",
  45941=>"010110101",
  45942=>"000011001",
  45943=>"001111110",
  45944=>"111011110",
  45945=>"011010001",
  45946=>"010100111",
  45947=>"001001011",
  45948=>"000100001",
  45949=>"011010010",
  45950=>"000001011",
  45951=>"100000111",
  45952=>"100111000",
  45953=>"111011000",
  45954=>"000111111",
  45955=>"001111100",
  45956=>"111100110",
  45957=>"101001111",
  45958=>"110101000",
  45959=>"100010011",
  45960=>"101001110",
  45961=>"100110100",
  45962=>"100000101",
  45963=>"010000010",
  45964=>"100001011",
  45965=>"000001001",
  45966=>"101110001",
  45967=>"000101000",
  45968=>"111010100",
  45969=>"011010000",
  45970=>"110110011",
  45971=>"101111100",
  45972=>"000101100",
  45973=>"011001011",
  45974=>"001011011",
  45975=>"110100101",
  45976=>"101100111",
  45977=>"011101100",
  45978=>"100011110",
  45979=>"100111011",
  45980=>"001110110",
  45981=>"100111011",
  45982=>"010001110",
  45983=>"001110001",
  45984=>"110110010",
  45985=>"001010011",
  45986=>"100000010",
  45987=>"000000100",
  45988=>"010100101",
  45989=>"110010111",
  45990=>"010110010",
  45991=>"111111110",
  45992=>"010111010",
  45993=>"101111011",
  45994=>"110111111",
  45995=>"000001100",
  45996=>"001110010",
  45997=>"011100100",
  45998=>"111000011",
  45999=>"101010110",
  46000=>"001101110",
  46001=>"010000110",
  46002=>"001110010",
  46003=>"100100111",
  46004=>"011110101",
  46005=>"100001010",
  46006=>"111000101",
  46007=>"101010100",
  46008=>"001001001",
  46009=>"001010011",
  46010=>"101110011",
  46011=>"111001111",
  46012=>"110111000",
  46013=>"111001001",
  46014=>"010000100",
  46015=>"010000000",
  46016=>"110011100",
  46017=>"101010010",
  46018=>"101101011",
  46019=>"110010100",
  46020=>"010000000",
  46021=>"000111010",
  46022=>"101110000",
  46023=>"100110101",
  46024=>"000110100",
  46025=>"110110000",
  46026=>"010101111",
  46027=>"010000010",
  46028=>"110110101",
  46029=>"011001000",
  46030=>"000101111",
  46031=>"001010101",
  46032=>"000001000",
  46033=>"011001110",
  46034=>"001011001",
  46035=>"101000001",
  46036=>"111001111",
  46037=>"100010100",
  46038=>"100000011",
  46039=>"111010000",
  46040=>"110110010",
  46041=>"110110001",
  46042=>"001000000",
  46043=>"000000011",
  46044=>"001010110",
  46045=>"110111111",
  46046=>"110000001",
  46047=>"001010001",
  46048=>"100100011",
  46049=>"100101001",
  46050=>"110010000",
  46051=>"111011101",
  46052=>"011110100",
  46053=>"000000011",
  46054=>"100011101",
  46055=>"100000011",
  46056=>"000111010",
  46057=>"000110110",
  46058=>"111001111",
  46059=>"110001001",
  46060=>"101001000",
  46061=>"000111010",
  46062=>"101110001",
  46063=>"011100010",
  46064=>"110010000",
  46065=>"101111001",
  46066=>"110110111",
  46067=>"110011111",
  46068=>"001011000",
  46069=>"101001110",
  46070=>"100000001",
  46071=>"010100010",
  46072=>"001001001",
  46073=>"111000110",
  46074=>"001011111",
  46075=>"000001010",
  46076=>"110110000",
  46077=>"110100111",
  46078=>"000010000",
  46079=>"001001101",
  46080=>"110000000",
  46081=>"010001000",
  46082=>"111011000",
  46083=>"010101010",
  46084=>"010010110",
  46085=>"001100101",
  46086=>"000101100",
  46087=>"111010100",
  46088=>"010101011",
  46089=>"001011000",
  46090=>"000011000",
  46091=>"111110101",
  46092=>"110011100",
  46093=>"111011101",
  46094=>"001110001",
  46095=>"100111111",
  46096=>"111110111",
  46097=>"000010111",
  46098=>"100100000",
  46099=>"100011010",
  46100=>"111110111",
  46101=>"100100000",
  46102=>"101100110",
  46103=>"100111100",
  46104=>"100101110",
  46105=>"011111011",
  46106=>"000110111",
  46107=>"010111001",
  46108=>"100000111",
  46109=>"010110000",
  46110=>"011001100",
  46111=>"001101101",
  46112=>"000001000",
  46113=>"101111111",
  46114=>"001100010",
  46115=>"011101001",
  46116=>"101000010",
  46117=>"010000011",
  46118=>"001000110",
  46119=>"000010000",
  46120=>"100001001",
  46121=>"011011101",
  46122=>"111001111",
  46123=>"100110110",
  46124=>"101110011",
  46125=>"101101000",
  46126=>"000011010",
  46127=>"110100011",
  46128=>"110111001",
  46129=>"010111100",
  46130=>"001110000",
  46131=>"010001110",
  46132=>"100001111",
  46133=>"101010111",
  46134=>"001110011",
  46135=>"111001111",
  46136=>"000000000",
  46137=>"001000001",
  46138=>"111101011",
  46139=>"000101011",
  46140=>"111110110",
  46141=>"101000001",
  46142=>"010010010",
  46143=>"101110100",
  46144=>"100011000",
  46145=>"100010111",
  46146=>"001011101",
  46147=>"100110001",
  46148=>"110000011",
  46149=>"101111011",
  46150=>"010100110",
  46151=>"000111011",
  46152=>"010101010",
  46153=>"111000000",
  46154=>"110100110",
  46155=>"101011110",
  46156=>"011000011",
  46157=>"001011111",
  46158=>"001111001",
  46159=>"010000111",
  46160=>"111101101",
  46161=>"000000110",
  46162=>"010100000",
  46163=>"000011110",
  46164=>"101111101",
  46165=>"111101001",
  46166=>"001000000",
  46167=>"101011111",
  46168=>"110000011",
  46169=>"101011010",
  46170=>"011011011",
  46171=>"000001000",
  46172=>"101000001",
  46173=>"111000010",
  46174=>"010101001",
  46175=>"010001000",
  46176=>"001001111",
  46177=>"010000000",
  46178=>"100000110",
  46179=>"010101100",
  46180=>"010110000",
  46181=>"100100111",
  46182=>"001000101",
  46183=>"110001001",
  46184=>"001010110",
  46185=>"111111101",
  46186=>"001001001",
  46187=>"010010100",
  46188=>"010111010",
  46189=>"101011011",
  46190=>"101111111",
  46191=>"111110000",
  46192=>"111100111",
  46193=>"011001001",
  46194=>"101010100",
  46195=>"010111000",
  46196=>"000000110",
  46197=>"111001101",
  46198=>"010000110",
  46199=>"110100001",
  46200=>"010111111",
  46201=>"001111101",
  46202=>"110110100",
  46203=>"010000001",
  46204=>"110111110",
  46205=>"100110001",
  46206=>"000011110",
  46207=>"101100110",
  46208=>"011111111",
  46209=>"101101111",
  46210=>"111011111",
  46211=>"111110101",
  46212=>"111011101",
  46213=>"100001100",
  46214=>"010111000",
  46215=>"011001111",
  46216=>"011000110",
  46217=>"110110011",
  46218=>"101011010",
  46219=>"100010010",
  46220=>"011100001",
  46221=>"001101111",
  46222=>"110011101",
  46223=>"101110010",
  46224=>"010101100",
  46225=>"011111000",
  46226=>"011111111",
  46227=>"110010100",
  46228=>"101011110",
  46229=>"110000100",
  46230=>"110100011",
  46231=>"110001110",
  46232=>"011101010",
  46233=>"000101000",
  46234=>"000010101",
  46235=>"010101100",
  46236=>"001100110",
  46237=>"100011011",
  46238=>"001011000",
  46239=>"000011000",
  46240=>"100100001",
  46241=>"011100101",
  46242=>"000010100",
  46243=>"100001011",
  46244=>"010011011",
  46245=>"010011111",
  46246=>"001001110",
  46247=>"111001101",
  46248=>"001010110",
  46249=>"001000111",
  46250=>"110001011",
  46251=>"100011000",
  46252=>"010000001",
  46253=>"011110010",
  46254=>"110111001",
  46255=>"000010110",
  46256=>"010000101",
  46257=>"001101110",
  46258=>"001101011",
  46259=>"111111001",
  46260=>"010001001",
  46261=>"101010110",
  46262=>"110001101",
  46263=>"011101111",
  46264=>"000000100",
  46265=>"111010010",
  46266=>"111010100",
  46267=>"111100111",
  46268=>"001101011",
  46269=>"000111001",
  46270=>"010001010",
  46271=>"011101010",
  46272=>"001100010",
  46273=>"000110101",
  46274=>"100100100",
  46275=>"110110110",
  46276=>"010010011",
  46277=>"110001100",
  46278=>"110000000",
  46279=>"011111101",
  46280=>"100001000",
  46281=>"110010111",
  46282=>"110001111",
  46283=>"111010101",
  46284=>"001001011",
  46285=>"100000111",
  46286=>"001010010",
  46287=>"100001010",
  46288=>"010101010",
  46289=>"100001011",
  46290=>"111100011",
  46291=>"001101100",
  46292=>"000000010",
  46293=>"001101000",
  46294=>"110111011",
  46295=>"001010001",
  46296=>"110011101",
  46297=>"101010010",
  46298=>"001000110",
  46299=>"001100001",
  46300=>"100110010",
  46301=>"001001000",
  46302=>"111011101",
  46303=>"011101111",
  46304=>"000100011",
  46305=>"010000011",
  46306=>"010111111",
  46307=>"000111111",
  46308=>"100100110",
  46309=>"011000001",
  46310=>"110011100",
  46311=>"010110001",
  46312=>"101100001",
  46313=>"111000101",
  46314=>"001111000",
  46315=>"011001110",
  46316=>"000110100",
  46317=>"111000011",
  46318=>"000011101",
  46319=>"111111001",
  46320=>"101111100",
  46321=>"111111000",
  46322=>"101110010",
  46323=>"101111011",
  46324=>"001011100",
  46325=>"000000110",
  46326=>"110010100",
  46327=>"111001001",
  46328=>"100110011",
  46329=>"100100100",
  46330=>"100100000",
  46331=>"001101100",
  46332=>"010101011",
  46333=>"110001101",
  46334=>"010101010",
  46335=>"010111111",
  46336=>"111010100",
  46337=>"011111101",
  46338=>"111111011",
  46339=>"110101011",
  46340=>"001100100",
  46341=>"101110010",
  46342=>"111110100",
  46343=>"111010111",
  46344=>"011001011",
  46345=>"101100110",
  46346=>"110011101",
  46347=>"100000000",
  46348=>"010000100",
  46349=>"010001111",
  46350=>"101001011",
  46351=>"111110001",
  46352=>"111010001",
  46353=>"010000011",
  46354=>"010100000",
  46355=>"000100001",
  46356=>"110011000",
  46357=>"111001100",
  46358=>"110011000",
  46359=>"011000010",
  46360=>"001110000",
  46361=>"101110010",
  46362=>"101001110",
  46363=>"001100000",
  46364=>"110100010",
  46365=>"110010111",
  46366=>"001111010",
  46367=>"100110010",
  46368=>"011101111",
  46369=>"000000000",
  46370=>"100011000",
  46371=>"101010001",
  46372=>"111010100",
  46373=>"001101000",
  46374=>"111100010",
  46375=>"001010100",
  46376=>"100001111",
  46377=>"110001011",
  46378=>"101110100",
  46379=>"110011111",
  46380=>"011001011",
  46381=>"011001000",
  46382=>"111001001",
  46383=>"101100011",
  46384=>"010001100",
  46385=>"110011000",
  46386=>"001111000",
  46387=>"001111101",
  46388=>"110110011",
  46389=>"101100011",
  46390=>"011000001",
  46391=>"011011010",
  46392=>"010010010",
  46393=>"000010100",
  46394=>"010000000",
  46395=>"001101101",
  46396=>"011001111",
  46397=>"101011101",
  46398=>"100001011",
  46399=>"110111000",
  46400=>"111000001",
  46401=>"101110100",
  46402=>"100100011",
  46403=>"011011000",
  46404=>"001111101",
  46405=>"001101110",
  46406=>"101101000",
  46407=>"001110000",
  46408=>"011111100",
  46409=>"100100110",
  46410=>"111110001",
  46411=>"000111111",
  46412=>"111100101",
  46413=>"110000101",
  46414=>"100111010",
  46415=>"101010001",
  46416=>"101011110",
  46417=>"110111000",
  46418=>"010000010",
  46419=>"001011100",
  46420=>"111110100",
  46421=>"111100101",
  46422=>"011101001",
  46423=>"010011010",
  46424=>"111111111",
  46425=>"000110111",
  46426=>"001000110",
  46427=>"011100001",
  46428=>"011110111",
  46429=>"111101001",
  46430=>"100000100",
  46431=>"011010000",
  46432=>"000101011",
  46433=>"100010111",
  46434=>"011111010",
  46435=>"001010000",
  46436=>"110100011",
  46437=>"111010000",
  46438=>"101000000",
  46439=>"000100100",
  46440=>"100110001",
  46441=>"010011001",
  46442=>"101110111",
  46443=>"111000110",
  46444=>"101110001",
  46445=>"111111011",
  46446=>"100010001",
  46447=>"111111010",
  46448=>"011100010",
  46449=>"101011001",
  46450=>"111101011",
  46451=>"000110011",
  46452=>"100000000",
  46453=>"111110110",
  46454=>"110010000",
  46455=>"001101010",
  46456=>"111001101",
  46457=>"100000010",
  46458=>"100001110",
  46459=>"110111111",
  46460=>"101011010",
  46461=>"101001001",
  46462=>"000111110",
  46463=>"001100111",
  46464=>"011110101",
  46465=>"011100000",
  46466=>"101010011",
  46467=>"000010001",
  46468=>"011100101",
  46469=>"101101101",
  46470=>"010101111",
  46471=>"111001001",
  46472=>"011111110",
  46473=>"111010101",
  46474=>"110110100",
  46475=>"111000111",
  46476=>"100100101",
  46477=>"101010101",
  46478=>"111001100",
  46479=>"001110110",
  46480=>"101001110",
  46481=>"010100111",
  46482=>"110110010",
  46483=>"000101011",
  46484=>"000011101",
  46485=>"001011001",
  46486=>"001110000",
  46487=>"111100111",
  46488=>"000011110",
  46489=>"111101011",
  46490=>"100000110",
  46491=>"001010101",
  46492=>"001100010",
  46493=>"000000000",
  46494=>"001110010",
  46495=>"100010101",
  46496=>"011101011",
  46497=>"010000101",
  46498=>"001000111",
  46499=>"011111010",
  46500=>"101111010",
  46501=>"000001011",
  46502=>"000000001",
  46503=>"100001011",
  46504=>"110101010",
  46505=>"110100100",
  46506=>"000100000",
  46507=>"110100101",
  46508=>"000000011",
  46509=>"110110011",
  46510=>"100011110",
  46511=>"010101000",
  46512=>"010111101",
  46513=>"100010100",
  46514=>"001000101",
  46515=>"011110111",
  46516=>"010100000",
  46517=>"100101111",
  46518=>"010100111",
  46519=>"101110110",
  46520=>"011001100",
  46521=>"000001111",
  46522=>"101000011",
  46523=>"111101110",
  46524=>"110001011",
  46525=>"000000110",
  46526=>"000110110",
  46527=>"001001101",
  46528=>"110010011",
  46529=>"110110010",
  46530=>"000001011",
  46531=>"001100111",
  46532=>"000010110",
  46533=>"011111111",
  46534=>"110100101",
  46535=>"110100111",
  46536=>"011001111",
  46537=>"101000000",
  46538=>"111011011",
  46539=>"010010110",
  46540=>"000000101",
  46541=>"010110101",
  46542=>"001010111",
  46543=>"011111110",
  46544=>"011110001",
  46545=>"010011100",
  46546=>"011000010",
  46547=>"000100001",
  46548=>"110111001",
  46549=>"101101101",
  46550=>"000010001",
  46551=>"010001100",
  46552=>"101001000",
  46553=>"110000000",
  46554=>"000000011",
  46555=>"010100001",
  46556=>"011101001",
  46557=>"100111010",
  46558=>"000101000",
  46559=>"111000111",
  46560=>"111100000",
  46561=>"101000000",
  46562=>"100011101",
  46563=>"001010001",
  46564=>"110111111",
  46565=>"110011010",
  46566=>"011001110",
  46567=>"111001100",
  46568=>"001101101",
  46569=>"110010110",
  46570=>"001001100",
  46571=>"010011001",
  46572=>"100001111",
  46573=>"111001101",
  46574=>"101101011",
  46575=>"111101000",
  46576=>"100011110",
  46577=>"111001010",
  46578=>"000101100",
  46579=>"000010100",
  46580=>"110111110",
  46581=>"001000100",
  46582=>"110100000",
  46583=>"000101100",
  46584=>"110100110",
  46585=>"100000010",
  46586=>"111010100",
  46587=>"110111100",
  46588=>"111010111",
  46589=>"000001000",
  46590=>"000110101",
  46591=>"110110111",
  46592=>"110011001",
  46593=>"001101001",
  46594=>"101011110",
  46595=>"110000111",
  46596=>"001110101",
  46597=>"001010100",
  46598=>"100011000",
  46599=>"011001010",
  46600=>"100111010",
  46601=>"011111010",
  46602=>"101010110",
  46603=>"100110010",
  46604=>"101001100",
  46605=>"001101000",
  46606=>"100111010",
  46607=>"000101000",
  46608=>"110001011",
  46609=>"100010110",
  46610=>"000010000",
  46611=>"111010011",
  46612=>"011111010",
  46613=>"010101101",
  46614=>"011110010",
  46615=>"101001100",
  46616=>"000011100",
  46617=>"110011010",
  46618=>"101110100",
  46619=>"010011100",
  46620=>"011100110",
  46621=>"011100000",
  46622=>"111000011",
  46623=>"001000111",
  46624=>"000111010",
  46625=>"101100101",
  46626=>"101110100",
  46627=>"101011001",
  46628=>"000011101",
  46629=>"000000101",
  46630=>"110000101",
  46631=>"100110100",
  46632=>"111001100",
  46633=>"110111111",
  46634=>"010001001",
  46635=>"101110010",
  46636=>"011001000",
  46637=>"111100001",
  46638=>"001110011",
  46639=>"110010110",
  46640=>"000000110",
  46641=>"100101111",
  46642=>"110111011",
  46643=>"111111001",
  46644=>"111001000",
  46645=>"110110100",
  46646=>"110001000",
  46647=>"111100000",
  46648=>"010000101",
  46649=>"000110100",
  46650=>"001100100",
  46651=>"011111001",
  46652=>"000000110",
  46653=>"001110010",
  46654=>"010111100",
  46655=>"011101111",
  46656=>"001000111",
  46657=>"100000101",
  46658=>"010110010",
  46659=>"011001100",
  46660=>"110110011",
  46661=>"001011101",
  46662=>"110100110",
  46663=>"000101100",
  46664=>"001110001",
  46665=>"110010110",
  46666=>"001000001",
  46667=>"101000111",
  46668=>"000111110",
  46669=>"000000001",
  46670=>"100000000",
  46671=>"100000110",
  46672=>"010111100",
  46673=>"000110101",
  46674=>"011111101",
  46675=>"011000010",
  46676=>"011010010",
  46677=>"010011001",
  46678=>"010011100",
  46679=>"011111101",
  46680=>"110100010",
  46681=>"000100000",
  46682=>"000011011",
  46683=>"110100100",
  46684=>"011010111",
  46685=>"110000000",
  46686=>"000000011",
  46687=>"110111101",
  46688=>"111011011",
  46689=>"101110110",
  46690=>"000010101",
  46691=>"110000111",
  46692=>"111000101",
  46693=>"001101010",
  46694=>"001010001",
  46695=>"011000100",
  46696=>"001101000",
  46697=>"100001000",
  46698=>"111001100",
  46699=>"001110000",
  46700=>"101100111",
  46701=>"000101110",
  46702=>"010111000",
  46703=>"000111110",
  46704=>"110000000",
  46705=>"000001101",
  46706=>"111111111",
  46707=>"100100011",
  46708=>"011000011",
  46709=>"010101111",
  46710=>"011010100",
  46711=>"011101100",
  46712=>"011011010",
  46713=>"100111011",
  46714=>"110111010",
  46715=>"011110111",
  46716=>"001000010",
  46717=>"000111111",
  46718=>"001010100",
  46719=>"000000110",
  46720=>"000000001",
  46721=>"000111011",
  46722=>"110100100",
  46723=>"010110111",
  46724=>"101100011",
  46725=>"001001101",
  46726=>"110001111",
  46727=>"100000001",
  46728=>"010011000",
  46729=>"010100110",
  46730=>"101010101",
  46731=>"000111011",
  46732=>"001001001",
  46733=>"111111110",
  46734=>"001001001",
  46735=>"001111111",
  46736=>"100110110",
  46737=>"100111111",
  46738=>"111010111",
  46739=>"011001111",
  46740=>"110001101",
  46741=>"011001001",
  46742=>"011000111",
  46743=>"000011011",
  46744=>"010011001",
  46745=>"100110011",
  46746=>"110011000",
  46747=>"010001001",
  46748=>"011011000",
  46749=>"100011110",
  46750=>"001011111",
  46751=>"100101000",
  46752=>"010001100",
  46753=>"000001011",
  46754=>"111001010",
  46755=>"000000011",
  46756=>"110100001",
  46757=>"101101000",
  46758=>"110000110",
  46759=>"110011101",
  46760=>"001000110",
  46761=>"111111010",
  46762=>"001101100",
  46763=>"101000000",
  46764=>"000110111",
  46765=>"111000000",
  46766=>"000110111",
  46767=>"111111110",
  46768=>"000110101",
  46769=>"010101010",
  46770=>"001100010",
  46771=>"011110110",
  46772=>"111010011",
  46773=>"111100000",
  46774=>"111011001",
  46775=>"010110000",
  46776=>"101101010",
  46777=>"010001010",
  46778=>"110100110",
  46779=>"000001011",
  46780=>"111010001",
  46781=>"110111010",
  46782=>"010110110",
  46783=>"110111011",
  46784=>"100011011",
  46785=>"001001110",
  46786=>"110010101",
  46787=>"001011011",
  46788=>"101101111",
  46789=>"001011100",
  46790=>"001010111",
  46791=>"101001000",
  46792=>"111101111",
  46793=>"010110111",
  46794=>"111001011",
  46795=>"111100000",
  46796=>"010101110",
  46797=>"101010110",
  46798=>"001010110",
  46799=>"000011111",
  46800=>"001000011",
  46801=>"101111011",
  46802=>"110111100",
  46803=>"111011000",
  46804=>"011011100",
  46805=>"111101001",
  46806=>"011111001",
  46807=>"010001001",
  46808=>"000001000",
  46809=>"010110101",
  46810=>"010111011",
  46811=>"010100011",
  46812=>"110001001",
  46813=>"010001000",
  46814=>"000101000",
  46815=>"101001001",
  46816=>"000110010",
  46817=>"101000001",
  46818=>"001100110",
  46819=>"011010011",
  46820=>"111110010",
  46821=>"100001000",
  46822=>"010101111",
  46823=>"001010010",
  46824=>"000100001",
  46825=>"111011010",
  46826=>"011000110",
  46827=>"010101111",
  46828=>"010011010",
  46829=>"110001100",
  46830=>"001111101",
  46831=>"000101110",
  46832=>"011111111",
  46833=>"110110101",
  46834=>"011100111",
  46835=>"110101001",
  46836=>"010001001",
  46837=>"110010010",
  46838=>"001110101",
  46839=>"111110111",
  46840=>"100010100",
  46841=>"101010001",
  46842=>"000101111",
  46843=>"001001001",
  46844=>"101100011",
  46845=>"010010011",
  46846=>"011111001",
  46847=>"110101011",
  46848=>"001110100",
  46849=>"000001110",
  46850=>"001001011",
  46851=>"111101010",
  46852=>"010000001",
  46853=>"001110110",
  46854=>"111001001",
  46855=>"101101010",
  46856=>"101001001",
  46857=>"100111101",
  46858=>"111000011",
  46859=>"110111100",
  46860=>"001101011",
  46861=>"111000111",
  46862=>"000100011",
  46863=>"101010110",
  46864=>"000001000",
  46865=>"101001110",
  46866=>"111110111",
  46867=>"100001001",
  46868=>"011000110",
  46869=>"100100111",
  46870=>"101110111",
  46871=>"001000010",
  46872=>"111111011",
  46873=>"011001000",
  46874=>"101011011",
  46875=>"101110010",
  46876=>"000011110",
  46877=>"101011110",
  46878=>"010011100",
  46879=>"111101100",
  46880=>"100011110",
  46881=>"000100101",
  46882=>"000010010",
  46883=>"011101000",
  46884=>"100000011",
  46885=>"100111000",
  46886=>"111111011",
  46887=>"010010111",
  46888=>"111100101",
  46889=>"011100111",
  46890=>"000100010",
  46891=>"101000101",
  46892=>"100111101",
  46893=>"001101000",
  46894=>"010001010",
  46895=>"000100010",
  46896=>"000011100",
  46897=>"110000011",
  46898=>"010111111",
  46899=>"011011100",
  46900=>"011110000",
  46901=>"011110000",
  46902=>"111101111",
  46903=>"111001101",
  46904=>"000010110",
  46905=>"010000110",
  46906=>"111000100",
  46907=>"001100001",
  46908=>"101100100",
  46909=>"001110010",
  46910=>"111011101",
  46911=>"010110010",
  46912=>"001111000",
  46913=>"000110101",
  46914=>"000101010",
  46915=>"001111001",
  46916=>"000011111",
  46917=>"001001001",
  46918=>"111011001",
  46919=>"110111101",
  46920=>"011110011",
  46921=>"001000100",
  46922=>"111010100",
  46923=>"100110101",
  46924=>"011100100",
  46925=>"011010110",
  46926=>"010010100",
  46927=>"111100111",
  46928=>"111000110",
  46929=>"010001110",
  46930=>"000000100",
  46931=>"100111000",
  46932=>"110111000",
  46933=>"111011100",
  46934=>"011011001",
  46935=>"001110110",
  46936=>"010111111",
  46937=>"011110000",
  46938=>"110010000",
  46939=>"011001000",
  46940=>"100011000",
  46941=>"101001111",
  46942=>"111000000",
  46943=>"000101011",
  46944=>"111000110",
  46945=>"000001101",
  46946=>"101001100",
  46947=>"101010100",
  46948=>"110011011",
  46949=>"100100010",
  46950=>"010001011",
  46951=>"001101100",
  46952=>"011111111",
  46953=>"011100011",
  46954=>"110111011",
  46955=>"000011010",
  46956=>"001011111",
  46957=>"011110000",
  46958=>"000101110",
  46959=>"111000101",
  46960=>"000100101",
  46961=>"011110111",
  46962=>"011100011",
  46963=>"000010111",
  46964=>"111010011",
  46965=>"000000011",
  46966=>"110001000",
  46967=>"001011101",
  46968=>"000001011",
  46969=>"011000011",
  46970=>"100000100",
  46971=>"110101011",
  46972=>"100110010",
  46973=>"101111110",
  46974=>"010001100",
  46975=>"000001010",
  46976=>"000100010",
  46977=>"011011100",
  46978=>"010100000",
  46979=>"100011000",
  46980=>"100101111",
  46981=>"011000001",
  46982=>"111010110",
  46983=>"010000010",
  46984=>"000001110",
  46985=>"110110111",
  46986=>"101011000",
  46987=>"111100101",
  46988=>"110110011",
  46989=>"000100101",
  46990=>"000011011",
  46991=>"001101000",
  46992=>"000110101",
  46993=>"001010001",
  46994=>"111101000",
  46995=>"100001010",
  46996=>"111110001",
  46997=>"101000110",
  46998=>"100101001",
  46999=>"110110000",
  47000=>"110001010",
  47001=>"001101000",
  47002=>"100001111",
  47003=>"000000110",
  47004=>"110001000",
  47005=>"000011100",
  47006=>"101001100",
  47007=>"100010000",
  47008=>"000011001",
  47009=>"000010110",
  47010=>"111010111",
  47011=>"111000000",
  47012=>"011001001",
  47013=>"001000001",
  47014=>"010100111",
  47015=>"001111111",
  47016=>"100010010",
  47017=>"111101100",
  47018=>"111101101",
  47019=>"001011101",
  47020=>"011111101",
  47021=>"000100001",
  47022=>"010100110",
  47023=>"010110001",
  47024=>"101000100",
  47025=>"000010011",
  47026=>"100101001",
  47027=>"010110111",
  47028=>"111010101",
  47029=>"010100011",
  47030=>"010111111",
  47031=>"110111011",
  47032=>"011010011",
  47033=>"110010000",
  47034=>"011111100",
  47035=>"110001100",
  47036=>"111101111",
  47037=>"100011101",
  47038=>"101011011",
  47039=>"010101110",
  47040=>"011010011",
  47041=>"010100110",
  47042=>"010001111",
  47043=>"011111000",
  47044=>"101001000",
  47045=>"111001011",
  47046=>"001001110",
  47047=>"000001010",
  47048=>"000000010",
  47049=>"111111110",
  47050=>"010110101",
  47051=>"011111110",
  47052=>"110010101",
  47053=>"101000111",
  47054=>"110001110",
  47055=>"110101111",
  47056=>"111101000",
  47057=>"011101100",
  47058=>"001010111",
  47059=>"100111100",
  47060=>"111100111",
  47061=>"110110011",
  47062=>"000010110",
  47063=>"000010011",
  47064=>"110000010",
  47065=>"101000111",
  47066=>"010001011",
  47067=>"000011110",
  47068=>"101011000",
  47069=>"101111100",
  47070=>"100010111",
  47071=>"101101001",
  47072=>"010110001",
  47073=>"001010001",
  47074=>"000011111",
  47075=>"000110101",
  47076=>"110010010",
  47077=>"000111111",
  47078=>"110011111",
  47079=>"110001001",
  47080=>"100001100",
  47081=>"010101001",
  47082=>"011001011",
  47083=>"000101001",
  47084=>"111001000",
  47085=>"010100000",
  47086=>"101100100",
  47087=>"000110110",
  47088=>"001100010",
  47089=>"000101010",
  47090=>"111000111",
  47091=>"101011101",
  47092=>"111111110",
  47093=>"010111110",
  47094=>"000000101",
  47095=>"010001100",
  47096=>"101101101",
  47097=>"101001000",
  47098=>"110100101",
  47099=>"100010101",
  47100=>"100110010",
  47101=>"011011000",
  47102=>"010000110",
  47103=>"011011100",
  47104=>"100000000",
  47105=>"011001100",
  47106=>"001010111",
  47107=>"011100110",
  47108=>"100101000",
  47109=>"000101001",
  47110=>"101110100",
  47111=>"100001111",
  47112=>"100100010",
  47113=>"001101100",
  47114=>"110011011",
  47115=>"000110001",
  47116=>"111111010",
  47117=>"100011100",
  47118=>"010011000",
  47119=>"000111000",
  47120=>"011000011",
  47121=>"001101010",
  47122=>"011101111",
  47123=>"001101110",
  47124=>"100101100",
  47125=>"001011001",
  47126=>"110001101",
  47127=>"011011110",
  47128=>"000100111",
  47129=>"001001011",
  47130=>"101101100",
  47131=>"011101000",
  47132=>"001011011",
  47133=>"100100101",
  47134=>"111100000",
  47135=>"011000000",
  47136=>"100100011",
  47137=>"100001000",
  47138=>"101000101",
  47139=>"001100100",
  47140=>"010011010",
  47141=>"010110010",
  47142=>"000111001",
  47143=>"110100101",
  47144=>"000001010",
  47145=>"101101000",
  47146=>"110100100",
  47147=>"010001111",
  47148=>"001111100",
  47149=>"111010000",
  47150=>"000000111",
  47151=>"000010001",
  47152=>"000100001",
  47153=>"001111100",
  47154=>"001100110",
  47155=>"111111000",
  47156=>"000101111",
  47157=>"110111001",
  47158=>"100100010",
  47159=>"010001110",
  47160=>"000001111",
  47161=>"010101001",
  47162=>"110100110",
  47163=>"000111001",
  47164=>"111011010",
  47165=>"000010110",
  47166=>"011100011",
  47167=>"100111101",
  47168=>"011001101",
  47169=>"101000000",
  47170=>"000101010",
  47171=>"110100010",
  47172=>"101001000",
  47173=>"010011111",
  47174=>"011010100",
  47175=>"111011100",
  47176=>"001110110",
  47177=>"011110000",
  47178=>"111010010",
  47179=>"000011000",
  47180=>"010000010",
  47181=>"100000110",
  47182=>"011010101",
  47183=>"001011000",
  47184=>"000110001",
  47185=>"000000010",
  47186=>"010111101",
  47187=>"100100100",
  47188=>"001110011",
  47189=>"101100010",
  47190=>"100010111",
  47191=>"101110111",
  47192=>"111111000",
  47193=>"000001101",
  47194=>"000011011",
  47195=>"010100010",
  47196=>"001000010",
  47197=>"000010000",
  47198=>"001001001",
  47199=>"001101110",
  47200=>"000100100",
  47201=>"111111110",
  47202=>"000001100",
  47203=>"101000110",
  47204=>"011101001",
  47205=>"110101101",
  47206=>"100010100",
  47207=>"001000101",
  47208=>"100010100",
  47209=>"000001010",
  47210=>"111111111",
  47211=>"110100110",
  47212=>"111110000",
  47213=>"100011110",
  47214=>"010111010",
  47215=>"000001101",
  47216=>"100001000",
  47217=>"011011011",
  47218=>"110110001",
  47219=>"011010000",
  47220=>"110011110",
  47221=>"100011001",
  47222=>"111011111",
  47223=>"111010011",
  47224=>"111011100",
  47225=>"111100010",
  47226=>"010000101",
  47227=>"000111001",
  47228=>"111010101",
  47229=>"010101100",
  47230=>"110110111",
  47231=>"111111110",
  47232=>"011110110",
  47233=>"000000110",
  47234=>"101101110",
  47235=>"000101001",
  47236=>"010101111",
  47237=>"100100101",
  47238=>"011100101",
  47239=>"001110001",
  47240=>"100011010",
  47241=>"100110000",
  47242=>"100111011",
  47243=>"000110010",
  47244=>"100001010",
  47245=>"010111101",
  47246=>"101101100",
  47247=>"010011011",
  47248=>"110000011",
  47249=>"011010101",
  47250=>"010111001",
  47251=>"110010110",
  47252=>"010001100",
  47253=>"110001101",
  47254=>"101011110",
  47255=>"111001001",
  47256=>"101111100",
  47257=>"101101111",
  47258=>"000010110",
  47259=>"000111111",
  47260=>"100000011",
  47261=>"011000010",
  47262=>"110110111",
  47263=>"000100000",
  47264=>"010001101",
  47265=>"010000001",
  47266=>"111110111",
  47267=>"011101001",
  47268=>"010111000",
  47269=>"111010110",
  47270=>"111101001",
  47271=>"111111110",
  47272=>"000110010",
  47273=>"111110111",
  47274=>"100011110",
  47275=>"000010001",
  47276=>"111110011",
  47277=>"001010010",
  47278=>"011101110",
  47279=>"011001110",
  47280=>"001010000",
  47281=>"010011100",
  47282=>"101100111",
  47283=>"101111100",
  47284=>"000000111",
  47285=>"111010010",
  47286=>"111100000",
  47287=>"100100111",
  47288=>"001111001",
  47289=>"101101111",
  47290=>"000000001",
  47291=>"111111101",
  47292=>"110101000",
  47293=>"100100110",
  47294=>"001010001",
  47295=>"000011010",
  47296=>"011010011",
  47297=>"011111101",
  47298=>"111100101",
  47299=>"110100110",
  47300=>"111110110",
  47301=>"100101010",
  47302=>"111010100",
  47303=>"111001111",
  47304=>"111100000",
  47305=>"100111011",
  47306=>"110111110",
  47307=>"101000100",
  47308=>"001001111",
  47309=>"111000011",
  47310=>"111110010",
  47311=>"010000111",
  47312=>"101010101",
  47313=>"110101110",
  47314=>"111110001",
  47315=>"110100010",
  47316=>"101000101",
  47317=>"110101010",
  47318=>"111010001",
  47319=>"010001011",
  47320=>"100011001",
  47321=>"010110100",
  47322=>"010110101",
  47323=>"000000000",
  47324=>"111111000",
  47325=>"101000111",
  47326=>"010001000",
  47327=>"000001111",
  47328=>"000010101",
  47329=>"100100110",
  47330=>"000000010",
  47331=>"101100110",
  47332=>"101001111",
  47333=>"110001000",
  47334=>"000000011",
  47335=>"000101111",
  47336=>"001111010",
  47337=>"000101111",
  47338=>"110001111",
  47339=>"000000011",
  47340=>"101001010",
  47341=>"001110001",
  47342=>"100101101",
  47343=>"101101100",
  47344=>"011101111",
  47345=>"001101111",
  47346=>"101101000",
  47347=>"010010110",
  47348=>"100010010",
  47349=>"001100111",
  47350=>"101101110",
  47351=>"101000000",
  47352=>"010100011",
  47353=>"100011001",
  47354=>"000001101",
  47355=>"100001101",
  47356=>"011110010",
  47357=>"100100110",
  47358=>"101001000",
  47359=>"010010011",
  47360=>"011001110",
  47361=>"010110011",
  47362=>"000011101",
  47363=>"011110001",
  47364=>"011101110",
  47365=>"000101110",
  47366=>"000111001",
  47367=>"111111001",
  47368=>"101000011",
  47369=>"000111011",
  47370=>"011100110",
  47371=>"000000100",
  47372=>"000101111",
  47373=>"100000100",
  47374=>"010001101",
  47375=>"000101100",
  47376=>"101010000",
  47377=>"110101101",
  47378=>"101101010",
  47379=>"110000110",
  47380=>"101011011",
  47381=>"110110000",
  47382=>"000100101",
  47383=>"010001111",
  47384=>"110000010",
  47385=>"001100111",
  47386=>"110000001",
  47387=>"100010110",
  47388=>"110010001",
  47389=>"101100111",
  47390=>"011010011",
  47391=>"000001011",
  47392=>"000000001",
  47393=>"000111110",
  47394=>"000111101",
  47395=>"111011000",
  47396=>"101010011",
  47397=>"101001010",
  47398=>"111100001",
  47399=>"011001100",
  47400=>"101001000",
  47401=>"111011111",
  47402=>"111010101",
  47403=>"111000110",
  47404=>"111111111",
  47405=>"000110110",
  47406=>"010111010",
  47407=>"000101011",
  47408=>"000011101",
  47409=>"110110100",
  47410=>"111100101",
  47411=>"110010111",
  47412=>"110001011",
  47413=>"000101100",
  47414=>"000111101",
  47415=>"001011000",
  47416=>"001101111",
  47417=>"110110000",
  47418=>"101001111",
  47419=>"101100001",
  47420=>"001010110",
  47421=>"111111110",
  47422=>"011010000",
  47423=>"110000100",
  47424=>"011000100",
  47425=>"000101100",
  47426=>"111001111",
  47427=>"100100111",
  47428=>"100101111",
  47429=>"110011111",
  47430=>"100010111",
  47431=>"100101001",
  47432=>"001011001",
  47433=>"100111100",
  47434=>"011110000",
  47435=>"010000000",
  47436=>"100000110",
  47437=>"110011001",
  47438=>"001000100",
  47439=>"111000110",
  47440=>"100011000",
  47441=>"101101010",
  47442=>"001100001",
  47443=>"110110010",
  47444=>"010110001",
  47445=>"000100100",
  47446=>"011100000",
  47447=>"101111111",
  47448=>"101101000",
  47449=>"100000100",
  47450=>"000111110",
  47451=>"001100000",
  47452=>"101111000",
  47453=>"000101001",
  47454=>"111011010",
  47455=>"010100100",
  47456=>"110100001",
  47457=>"100001101",
  47458=>"110110011",
  47459=>"001001111",
  47460=>"011010001",
  47461=>"111111011",
  47462=>"010101111",
  47463=>"010100100",
  47464=>"000000000",
  47465=>"001000000",
  47466=>"000000000",
  47467=>"101001110",
  47468=>"010111010",
  47469=>"100010101",
  47470=>"001101000",
  47471=>"001000100",
  47472=>"011110110",
  47473=>"010111111",
  47474=>"010001010",
  47475=>"100001110",
  47476=>"101101001",
  47477=>"010001010",
  47478=>"111111111",
  47479=>"111111111",
  47480=>"111100101",
  47481=>"111101111",
  47482=>"010010101",
  47483=>"010100010",
  47484=>"111011001",
  47485=>"110101010",
  47486=>"101000100",
  47487=>"100001001",
  47488=>"110010100",
  47489=>"000010111",
  47490=>"101000011",
  47491=>"110101000",
  47492=>"000011100",
  47493=>"010011101",
  47494=>"001100110",
  47495=>"111111000",
  47496=>"101000010",
  47497=>"100100000",
  47498=>"100110110",
  47499=>"100010101",
  47500=>"100101010",
  47501=>"001111111",
  47502=>"001011001",
  47503=>"101100000",
  47504=>"100010001",
  47505=>"100001011",
  47506=>"001100011",
  47507=>"011110011",
  47508=>"110001110",
  47509=>"110000110",
  47510=>"101100000",
  47511=>"101110000",
  47512=>"100000000",
  47513=>"101100010",
  47514=>"100111110",
  47515=>"010101000",
  47516=>"001011011",
  47517=>"111111111",
  47518=>"111000001",
  47519=>"100101011",
  47520=>"110001100",
  47521=>"111110101",
  47522=>"100110101",
  47523=>"000000001",
  47524=>"110011110",
  47525=>"000110110",
  47526=>"011000001",
  47527=>"111000010",
  47528=>"001000100",
  47529=>"010010101",
  47530=>"100000001",
  47531=>"111111000",
  47532=>"101001101",
  47533=>"011111010",
  47534=>"100111100",
  47535=>"111001011",
  47536=>"000101100",
  47537=>"101111100",
  47538=>"111100111",
  47539=>"111110110",
  47540=>"111001010",
  47541=>"100101010",
  47542=>"101000100",
  47543=>"100110100",
  47544=>"001110010",
  47545=>"001001111",
  47546=>"000100111",
  47547=>"000011011",
  47548=>"000101010",
  47549=>"111101110",
  47550=>"011110100",
  47551=>"000010101",
  47552=>"001001010",
  47553=>"001011001",
  47554=>"111110111",
  47555=>"010011001",
  47556=>"000001000",
  47557=>"110000011",
  47558=>"010000001",
  47559=>"011100000",
  47560=>"101001111",
  47561=>"100101011",
  47562=>"000101110",
  47563=>"111010101",
  47564=>"011110100",
  47565=>"100110010",
  47566=>"100000000",
  47567=>"100110001",
  47568=>"101001001",
  47569=>"000101101",
  47570=>"110100011",
  47571=>"000111111",
  47572=>"011000100",
  47573=>"011010110",
  47574=>"010010011",
  47575=>"101111010",
  47576=>"000111001",
  47577=>"110011011",
  47578=>"000001110",
  47579=>"101100111",
  47580=>"100000100",
  47581=>"100000111",
  47582=>"010001001",
  47583=>"001010100",
  47584=>"111101111",
  47585=>"001100010",
  47586=>"101111101",
  47587=>"111000001",
  47588=>"010100010",
  47589=>"111011110",
  47590=>"110000000",
  47591=>"110010011",
  47592=>"100000100",
  47593=>"101010101",
  47594=>"001110000",
  47595=>"010101001",
  47596=>"111110101",
  47597=>"011101101",
  47598=>"010010001",
  47599=>"010100100",
  47600=>"100111001",
  47601=>"000001011",
  47602=>"100100001",
  47603=>"010011100",
  47604=>"011011010",
  47605=>"001111110",
  47606=>"110010100",
  47607=>"111100010",
  47608=>"001001111",
  47609=>"110101010",
  47610=>"001000101",
  47611=>"111111101",
  47612=>"100110110",
  47613=>"011110001",
  47614=>"011110010",
  47615=>"010111000",
  47616=>"111000010",
  47617=>"001110110",
  47618=>"001001001",
  47619=>"111100111",
  47620=>"001110011",
  47621=>"100000011",
  47622=>"110111111",
  47623=>"010111111",
  47624=>"110111010",
  47625=>"101111100",
  47626=>"111010010",
  47627=>"101001010",
  47628=>"000011100",
  47629=>"110101100",
  47630=>"000100010",
  47631=>"100000101",
  47632=>"000111110",
  47633=>"110101110",
  47634=>"101001111",
  47635=>"100101111",
  47636=>"011000101",
  47637=>"110111111",
  47638=>"000000001",
  47639=>"001110000",
  47640=>"110111001",
  47641=>"100011001",
  47642=>"100111110",
  47643=>"100110000",
  47644=>"000100011",
  47645=>"000011010",
  47646=>"110010010",
  47647=>"011110011",
  47648=>"010000010",
  47649=>"111011100",
  47650=>"101000000",
  47651=>"111011001",
  47652=>"100000010",
  47653=>"000100000",
  47654=>"000111101",
  47655=>"001010010",
  47656=>"001101111",
  47657=>"000111111",
  47658=>"101100001",
  47659=>"010101010",
  47660=>"010000011",
  47661=>"011101000",
  47662=>"101111111",
  47663=>"111011011",
  47664=>"000000111",
  47665=>"001100111",
  47666=>"100100111",
  47667=>"000011101",
  47668=>"111001110",
  47669=>"111111000",
  47670=>"011011100",
  47671=>"000000100",
  47672=>"101101100",
  47673=>"000000010",
  47674=>"100011010",
  47675=>"011001000",
  47676=>"000100000",
  47677=>"000000000",
  47678=>"011001011",
  47679=>"100000001",
  47680=>"101100010",
  47681=>"101011101",
  47682=>"101011100",
  47683=>"100100111",
  47684=>"000011100",
  47685=>"000000110",
  47686=>"000010001",
  47687=>"111000010",
  47688=>"100010011",
  47689=>"101011111",
  47690=>"100000111",
  47691=>"010010010",
  47692=>"100111000",
  47693=>"111101101",
  47694=>"011111110",
  47695=>"001101011",
  47696=>"100001110",
  47697=>"010011000",
  47698=>"100100011",
  47699=>"010000011",
  47700=>"001010000",
  47701=>"001000110",
  47702=>"001101000",
  47703=>"010001111",
  47704=>"010001111",
  47705=>"001010010",
  47706=>"001101010",
  47707=>"001101011",
  47708=>"100011010",
  47709=>"111101010",
  47710=>"101111110",
  47711=>"110100011",
  47712=>"101001101",
  47713=>"110110010",
  47714=>"001101000",
  47715=>"000000001",
  47716=>"000111010",
  47717=>"100101000",
  47718=>"000001010",
  47719=>"101101111",
  47720=>"000101010",
  47721=>"110111000",
  47722=>"010000110",
  47723=>"100110000",
  47724=>"000000001",
  47725=>"010011011",
  47726=>"110100001",
  47727=>"110111110",
  47728=>"101101110",
  47729=>"000011011",
  47730=>"111110011",
  47731=>"010011101",
  47732=>"100010010",
  47733=>"100000010",
  47734=>"101001100",
  47735=>"011100101",
  47736=>"001011101",
  47737=>"001001001",
  47738=>"010111011",
  47739=>"010010111",
  47740=>"110101001",
  47741=>"110111001",
  47742=>"010000011",
  47743=>"001000010",
  47744=>"001100110",
  47745=>"101100011",
  47746=>"001110000",
  47747=>"110110000",
  47748=>"110010101",
  47749=>"000001000",
  47750=>"111000111",
  47751=>"101011111",
  47752=>"001110001",
  47753=>"110101011",
  47754=>"111011011",
  47755=>"001100100",
  47756=>"000001000",
  47757=>"110101111",
  47758=>"110101000",
  47759=>"100001011",
  47760=>"010110011",
  47761=>"000100111",
  47762=>"101100000",
  47763=>"001010000",
  47764=>"111110000",
  47765=>"000010111",
  47766=>"101010010",
  47767=>"001000010",
  47768=>"000000010",
  47769=>"100011001",
  47770=>"000100011",
  47771=>"101111010",
  47772=>"100010100",
  47773=>"111111000",
  47774=>"110110010",
  47775=>"010100110",
  47776=>"000111011",
  47777=>"110000010",
  47778=>"111100011",
  47779=>"000111111",
  47780=>"111010110",
  47781=>"011011110",
  47782=>"101110010",
  47783=>"101100011",
  47784=>"011111110",
  47785=>"000001001",
  47786=>"000100011",
  47787=>"011000011",
  47788=>"101110001",
  47789=>"011101010",
  47790=>"111111100",
  47791=>"101100100",
  47792=>"111110000",
  47793=>"011001010",
  47794=>"100011111",
  47795=>"001010101",
  47796=>"110100101",
  47797=>"010110110",
  47798=>"111110100",
  47799=>"111110111",
  47800=>"000110000",
  47801=>"101110110",
  47802=>"100101010",
  47803=>"110010010",
  47804=>"001011011",
  47805=>"110101101",
  47806=>"111011001",
  47807=>"110100000",
  47808=>"111001111",
  47809=>"010000111",
  47810=>"010111001",
  47811=>"010110110",
  47812=>"000001000",
  47813=>"111011010",
  47814=>"001010111",
  47815=>"010111010",
  47816=>"001011001",
  47817=>"100010110",
  47818=>"001111011",
  47819=>"011011101",
  47820=>"101000011",
  47821=>"111111011",
  47822=>"100000110",
  47823=>"100011100",
  47824=>"011011111",
  47825=>"010011110",
  47826=>"110101011",
  47827=>"011010011",
  47828=>"100010000",
  47829=>"100101000",
  47830=>"011110011",
  47831=>"101000111",
  47832=>"100101001",
  47833=>"010011110",
  47834=>"010000100",
  47835=>"100111100",
  47836=>"001101011",
  47837=>"001001111",
  47838=>"110110101",
  47839=>"100011100",
  47840=>"111011001",
  47841=>"000100001",
  47842=>"000010011",
  47843=>"110101101",
  47844=>"001100101",
  47845=>"001101111",
  47846=>"011110000",
  47847=>"001100000",
  47848=>"100001010",
  47849=>"010111110",
  47850=>"011110111",
  47851=>"101010100",
  47852=>"101001000",
  47853=>"100111101",
  47854=>"110011111",
  47855=>"110100101",
  47856=>"010110111",
  47857=>"001010011",
  47858=>"111110100",
  47859=>"011010011",
  47860=>"101011101",
  47861=>"000010111",
  47862=>"101000110",
  47863=>"110100001",
  47864=>"011010010",
  47865=>"111110111",
  47866=>"000110101",
  47867=>"100111110",
  47868=>"100101100",
  47869=>"111010101",
  47870=>"000101011",
  47871=>"100001000",
  47872=>"100100111",
  47873=>"011111011",
  47874=>"110011011",
  47875=>"001100011",
  47876=>"010110011",
  47877=>"010001000",
  47878=>"001101101",
  47879=>"000100100",
  47880=>"101011000",
  47881=>"000100001",
  47882=>"000100100",
  47883=>"000000000",
  47884=>"010101000",
  47885=>"111110111",
  47886=>"101011011",
  47887=>"110000101",
  47888=>"001101001",
  47889=>"000000101",
  47890=>"110110110",
  47891=>"001100000",
  47892=>"010111011",
  47893=>"111011111",
  47894=>"110011101",
  47895=>"110011111",
  47896=>"001101100",
  47897=>"001101010",
  47898=>"100000000",
  47899=>"011101001",
  47900=>"101101101",
  47901=>"000101100",
  47902=>"110010001",
  47903=>"100001000",
  47904=>"111000100",
  47905=>"111110111",
  47906=>"001101101",
  47907=>"000100000",
  47908=>"101011100",
  47909=>"110000011",
  47910=>"101111111",
  47911=>"101111110",
  47912=>"000000100",
  47913=>"101010101",
  47914=>"010001100",
  47915=>"000101010",
  47916=>"010111111",
  47917=>"110101110",
  47918=>"101111001",
  47919=>"010110100",
  47920=>"110001011",
  47921=>"010101001",
  47922=>"110111000",
  47923=>"011000110",
  47924=>"010001110",
  47925=>"110111101",
  47926=>"101111000",
  47927=>"111001011",
  47928=>"011000101",
  47929=>"110001000",
  47930=>"111001001",
  47931=>"111100111",
  47932=>"111101000",
  47933=>"110011010",
  47934=>"010010110",
  47935=>"011100001",
  47936=>"000000111",
  47937=>"011001111",
  47938=>"010111010",
  47939=>"010101001",
  47940=>"010111000",
  47941=>"111100010",
  47942=>"101101001",
  47943=>"101100000",
  47944=>"101000101",
  47945=>"000001101",
  47946=>"000101111",
  47947=>"010110110",
  47948=>"111011100",
  47949=>"000011011",
  47950=>"101000110",
  47951=>"000101001",
  47952=>"010000001",
  47953=>"101001111",
  47954=>"100100000",
  47955=>"001000101",
  47956=>"011000000",
  47957=>"001010111",
  47958=>"010110010",
  47959=>"010110101",
  47960=>"111110100",
  47961=>"110111001",
  47962=>"111110110",
  47963=>"001010000",
  47964=>"110111001",
  47965=>"010101101",
  47966=>"100000111",
  47967=>"100110011",
  47968=>"110011000",
  47969=>"001001000",
  47970=>"011001000",
  47971=>"100101011",
  47972=>"010111001",
  47973=>"001000001",
  47974=>"000101100",
  47975=>"110011101",
  47976=>"001101111",
  47977=>"011010101",
  47978=>"000110100",
  47979=>"010100101",
  47980=>"110011000",
  47981=>"111110101",
  47982=>"011001001",
  47983=>"111000100",
  47984=>"010010000",
  47985=>"011111111",
  47986=>"001011100",
  47987=>"111101001",
  47988=>"001000100",
  47989=>"010010010",
  47990=>"110011101",
  47991=>"100101110",
  47992=>"010010110",
  47993=>"111110101",
  47994=>"111100101",
  47995=>"111010000",
  47996=>"011001001",
  47997=>"001011101",
  47998=>"011111000",
  47999=>"100101111",
  48000=>"111001001",
  48001=>"100101111",
  48002=>"101111010",
  48003=>"011101011",
  48004=>"111100000",
  48005=>"011111111",
  48006=>"100100111",
  48007=>"110010001",
  48008=>"011111011",
  48009=>"010000000",
  48010=>"000111010",
  48011=>"101010000",
  48012=>"000111010",
  48013=>"111001100",
  48014=>"000100101",
  48015=>"011010110",
  48016=>"001100111",
  48017=>"110011001",
  48018=>"010000110",
  48019=>"001000011",
  48020=>"001001000",
  48021=>"000010111",
  48022=>"010001101",
  48023=>"001001010",
  48024=>"011100000",
  48025=>"111111100",
  48026=>"110001001",
  48027=>"110000110",
  48028=>"000000000",
  48029=>"001010101",
  48030=>"000001101",
  48031=>"111011110",
  48032=>"010110100",
  48033=>"111101011",
  48034=>"110000011",
  48035=>"100000100",
  48036=>"100111110",
  48037=>"010011000",
  48038=>"111001110",
  48039=>"111100111",
  48040=>"111001000",
  48041=>"101000100",
  48042=>"010110001",
  48043=>"011010010",
  48044=>"000110110",
  48045=>"110000111",
  48046=>"000110011",
  48047=>"111111001",
  48048=>"001010100",
  48049=>"100100101",
  48050=>"001011010",
  48051=>"100000011",
  48052=>"010100001",
  48053=>"011000010",
  48054=>"111111110",
  48055=>"100101100",
  48056=>"100110001",
  48057=>"000001010",
  48058=>"100010001",
  48059=>"111010101",
  48060=>"101000110",
  48061=>"101010101",
  48062=>"001001010",
  48063=>"010000000",
  48064=>"110100110",
  48065=>"110100101",
  48066=>"001101101",
  48067=>"010001000",
  48068=>"001101111",
  48069=>"001110100",
  48070=>"110000001",
  48071=>"110100110",
  48072=>"010101100",
  48073=>"111000111",
  48074=>"010111100",
  48075=>"010000100",
  48076=>"110110111",
  48077=>"001110101",
  48078=>"100110000",
  48079=>"011000101",
  48080=>"111110001",
  48081=>"000011010",
  48082=>"110010101",
  48083=>"000000100",
  48084=>"000101001",
  48085=>"010010101",
  48086=>"110101000",
  48087=>"101100001",
  48088=>"010100011",
  48089=>"001101110",
  48090=>"011011111",
  48091=>"011110111",
  48092=>"101110101",
  48093=>"010110101",
  48094=>"010111111",
  48095=>"010011100",
  48096=>"000110101",
  48097=>"000111001",
  48098=>"101100001",
  48099=>"100100010",
  48100=>"000011010",
  48101=>"011111001",
  48102=>"110000000",
  48103=>"100111011",
  48104=>"101001100",
  48105=>"001011001",
  48106=>"111100100",
  48107=>"100000100",
  48108=>"111101101",
  48109=>"001100110",
  48110=>"100001001",
  48111=>"110110110",
  48112=>"100010010",
  48113=>"101101001",
  48114=>"000011100",
  48115=>"101110000",
  48116=>"111110111",
  48117=>"011100111",
  48118=>"010000010",
  48119=>"011000001",
  48120=>"010111000",
  48121=>"111110101",
  48122=>"000010001",
  48123=>"001000001",
  48124=>"111000000",
  48125=>"110101101",
  48126=>"100100101",
  48127=>"101010101",
  48128=>"011001111",
  48129=>"110011010",
  48130=>"111100111",
  48131=>"010011101",
  48132=>"001010100",
  48133=>"010011010",
  48134=>"000111111",
  48135=>"110000100",
  48136=>"010010000",
  48137=>"001010001",
  48138=>"000110100",
  48139=>"000001111",
  48140=>"010000001",
  48141=>"110011111",
  48142=>"111011000",
  48143=>"011010000",
  48144=>"101100100",
  48145=>"000111111",
  48146=>"010000100",
  48147=>"000101110",
  48148=>"011000011",
  48149=>"000011100",
  48150=>"100111000",
  48151=>"011000000",
  48152=>"000111001",
  48153=>"000000111",
  48154=>"000010010",
  48155=>"101001101",
  48156=>"100100110",
  48157=>"000001000",
  48158=>"110000100",
  48159=>"101111100",
  48160=>"001001100",
  48161=>"010001111",
  48162=>"100000110",
  48163=>"111010100",
  48164=>"011111000",
  48165=>"111000110",
  48166=>"010110011",
  48167=>"011101110",
  48168=>"001110001",
  48169=>"011010100",
  48170=>"111000011",
  48171=>"111011101",
  48172=>"001101001",
  48173=>"110011101",
  48174=>"011010010",
  48175=>"111011000",
  48176=>"101010010",
  48177=>"011100110",
  48178=>"010111111",
  48179=>"100110000",
  48180=>"010110010",
  48181=>"000001010",
  48182=>"010010000",
  48183=>"010101101",
  48184=>"100010000",
  48185=>"001111111",
  48186=>"000001101",
  48187=>"101111100",
  48188=>"010011011",
  48189=>"111011000",
  48190=>"001001011",
  48191=>"101011111",
  48192=>"100011001",
  48193=>"100011010",
  48194=>"010001010",
  48195=>"100100111",
  48196=>"110010111",
  48197=>"000110011",
  48198=>"110010100",
  48199=>"010101100",
  48200=>"001110011",
  48201=>"011100010",
  48202=>"110010000",
  48203=>"000000000",
  48204=>"001110011",
  48205=>"010011111",
  48206=>"100001011",
  48207=>"111110011",
  48208=>"101001010",
  48209=>"001111110",
  48210=>"011100101",
  48211=>"101111010",
  48212=>"101101100",
  48213=>"010100111",
  48214=>"011101111",
  48215=>"001101100",
  48216=>"110100110",
  48217=>"110011111",
  48218=>"101010100",
  48219=>"010100100",
  48220=>"000001111",
  48221=>"100100111",
  48222=>"110100001",
  48223=>"011101100",
  48224=>"111011000",
  48225=>"111010111",
  48226=>"110101001",
  48227=>"001000100",
  48228=>"000100001",
  48229=>"100010000",
  48230=>"001010010",
  48231=>"100101011",
  48232=>"000010000",
  48233=>"000111101",
  48234=>"111100000",
  48235=>"100101110",
  48236=>"011000110",
  48237=>"110001100",
  48238=>"100000100",
  48239=>"001100100",
  48240=>"101110111",
  48241=>"101100000",
  48242=>"101101101",
  48243=>"110000011",
  48244=>"000101110",
  48245=>"111001111",
  48246=>"001100101",
  48247=>"011110111",
  48248=>"000011110",
  48249=>"000010000",
  48250=>"001000100",
  48251=>"101111111",
  48252=>"001100111",
  48253=>"111111110",
  48254=>"000100001",
  48255=>"000001110",
  48256=>"001101110",
  48257=>"101111011",
  48258=>"000000111",
  48259=>"011110110",
  48260=>"011000100",
  48261=>"101110101",
  48262=>"001010000",
  48263=>"101110110",
  48264=>"111111101",
  48265=>"101111111",
  48266=>"001010100",
  48267=>"010110001",
  48268=>"000011110",
  48269=>"100000001",
  48270=>"001101000",
  48271=>"001011011",
  48272=>"110101010",
  48273=>"011100101",
  48274=>"101110110",
  48275=>"001000101",
  48276=>"001100001",
  48277=>"101010011",
  48278=>"001110000",
  48279=>"110100001",
  48280=>"001001000",
  48281=>"010000010",
  48282=>"100001010",
  48283=>"010111100",
  48284=>"101010100",
  48285=>"100101000",
  48286=>"000000101",
  48287=>"101110001",
  48288=>"011010000",
  48289=>"110011001",
  48290=>"110000100",
  48291=>"010100101",
  48292=>"110100111",
  48293=>"111001110",
  48294=>"101110000",
  48295=>"110111000",
  48296=>"010100111",
  48297=>"100111110",
  48298=>"101110110",
  48299=>"010010111",
  48300=>"111001001",
  48301=>"010100100",
  48302=>"011110000",
  48303=>"001110010",
  48304=>"101000011",
  48305=>"101011111",
  48306=>"001110111",
  48307=>"111111011",
  48308=>"000100100",
  48309=>"001110100",
  48310=>"011111001",
  48311=>"101011101",
  48312=>"100000001",
  48313=>"000001011",
  48314=>"001001100",
  48315=>"111011000",
  48316=>"101111101",
  48317=>"111101111",
  48318=>"100010100",
  48319=>"110000101",
  48320=>"010100100",
  48321=>"011000111",
  48322=>"111100011",
  48323=>"001000101",
  48324=>"111000010",
  48325=>"011110110",
  48326=>"111101110",
  48327=>"000110101",
  48328=>"001000101",
  48329=>"011010001",
  48330=>"111100011",
  48331=>"011101110",
  48332=>"110101011",
  48333=>"011101101",
  48334=>"111110011",
  48335=>"111100011",
  48336=>"100010011",
  48337=>"000101111",
  48338=>"101011000",
  48339=>"000000011",
  48340=>"000001000",
  48341=>"100010110",
  48342=>"111100001",
  48343=>"001010101",
  48344=>"000100100",
  48345=>"101000001",
  48346=>"001000100",
  48347=>"100000010",
  48348=>"100101001",
  48349=>"101010111",
  48350=>"100000011",
  48351=>"101011000",
  48352=>"111110111",
  48353=>"111000111",
  48354=>"010001100",
  48355=>"110101010",
  48356=>"011010101",
  48357=>"000001100",
  48358=>"110000011",
  48359=>"011101101",
  48360=>"000111011",
  48361=>"101001000",
  48362=>"100010110",
  48363=>"101000001",
  48364=>"101001000",
  48365=>"011100101",
  48366=>"001011011",
  48367=>"101000110",
  48368=>"100011100",
  48369=>"101101011",
  48370=>"110100110",
  48371=>"001011010",
  48372=>"111101001",
  48373=>"000000101",
  48374=>"101100100",
  48375=>"000100001",
  48376=>"111010001",
  48377=>"011101100",
  48378=>"001011000",
  48379=>"101100000",
  48380=>"111010111",
  48381=>"110110011",
  48382=>"100111011",
  48383=>"001010111",
  48384=>"010001010",
  48385=>"101010101",
  48386=>"000110110",
  48387=>"010101101",
  48388=>"001111100",
  48389=>"011010111",
  48390=>"111111111",
  48391=>"111001011",
  48392=>"001111000",
  48393=>"000011000",
  48394=>"100011111",
  48395=>"100001010",
  48396=>"001111110",
  48397=>"111011110",
  48398=>"000000110",
  48399=>"100000111",
  48400=>"011111010",
  48401=>"001110101",
  48402=>"100010010",
  48403=>"111100111",
  48404=>"000001010",
  48405=>"101101111",
  48406=>"000010100",
  48407=>"000100001",
  48408=>"111111000",
  48409=>"000011110",
  48410=>"111011110",
  48411=>"110111000",
  48412=>"001011100",
  48413=>"110110001",
  48414=>"011110100",
  48415=>"100001001",
  48416=>"001111111",
  48417=>"111100110",
  48418=>"111101000",
  48419=>"011001011",
  48420=>"101001110",
  48421=>"100001101",
  48422=>"100111010",
  48423=>"011111110",
  48424=>"111011000",
  48425=>"100110110",
  48426=>"101111100",
  48427=>"100111101",
  48428=>"001000010",
  48429=>"011011100",
  48430=>"001111101",
  48431=>"111000010",
  48432=>"000001110",
  48433=>"101111001",
  48434=>"010101100",
  48435=>"101010001",
  48436=>"110011110",
  48437=>"100000000",
  48438=>"001000001",
  48439=>"001111110",
  48440=>"010100011",
  48441=>"000100010",
  48442=>"011011001",
  48443=>"101000101",
  48444=>"111111101",
  48445=>"001110110",
  48446=>"111010111",
  48447=>"101100111",
  48448=>"010010101",
  48449=>"001110011",
  48450=>"001000111",
  48451=>"010010001",
  48452=>"010000100",
  48453=>"001000101",
  48454=>"000001001",
  48455=>"001011000",
  48456=>"110101101",
  48457=>"101001010",
  48458=>"011100001",
  48459=>"100010010",
  48460=>"101011010",
  48461=>"100000010",
  48462=>"000001000",
  48463=>"000010001",
  48464=>"101101001",
  48465=>"001011011",
  48466=>"111011001",
  48467=>"000001001",
  48468=>"000001101",
  48469=>"011010110",
  48470=>"111010100",
  48471=>"100010011",
  48472=>"100111011",
  48473=>"110101000",
  48474=>"001100001",
  48475=>"110011000",
  48476=>"011100111",
  48477=>"100001011",
  48478=>"010000110",
  48479=>"001000010",
  48480=>"010111011",
  48481=>"011001110",
  48482=>"110000111",
  48483=>"001100101",
  48484=>"101110011",
  48485=>"101011010",
  48486=>"011110010",
  48487=>"111111011",
  48488=>"111111111",
  48489=>"100110000",
  48490=>"110111011",
  48491=>"000100001",
  48492=>"101010111",
  48493=>"000010001",
  48494=>"111101110",
  48495=>"011011011",
  48496=>"000010010",
  48497=>"111001111",
  48498=>"010010111",
  48499=>"111000100",
  48500=>"011000101",
  48501=>"011100000",
  48502=>"100110000",
  48503=>"110111001",
  48504=>"001001001",
  48505=>"110001001",
  48506=>"011001111",
  48507=>"101010010",
  48508=>"001101000",
  48509=>"100101000",
  48510=>"000010011",
  48511=>"001101001",
  48512=>"001000110",
  48513=>"001010101",
  48514=>"101111101",
  48515=>"011010000",
  48516=>"010101010",
  48517=>"001001100",
  48518=>"010110111",
  48519=>"110011001",
  48520=>"110001101",
  48521=>"111000100",
  48522=>"111111111",
  48523=>"100000111",
  48524=>"001000100",
  48525=>"101000110",
  48526=>"101010100",
  48527=>"110001101",
  48528=>"011011011",
  48529=>"010111001",
  48530=>"101101001",
  48531=>"010010000",
  48532=>"000011000",
  48533=>"011111000",
  48534=>"110111110",
  48535=>"111100100",
  48536=>"111010001",
  48537=>"010011000",
  48538=>"100000100",
  48539=>"001011100",
  48540=>"011111000",
  48541=>"110011000",
  48542=>"000100110",
  48543=>"000001001",
  48544=>"101100000",
  48545=>"010101111",
  48546=>"100000011",
  48547=>"010111101",
  48548=>"010011111",
  48549=>"000101001",
  48550=>"001001101",
  48551=>"010011001",
  48552=>"000001111",
  48553=>"001011100",
  48554=>"011001001",
  48555=>"010110110",
  48556=>"110110001",
  48557=>"001111111",
  48558=>"000000000",
  48559=>"001001000",
  48560=>"101110111",
  48561=>"001010010",
  48562=>"000001010",
  48563=>"000001011",
  48564=>"100001010",
  48565=>"010100011",
  48566=>"100111011",
  48567=>"100001110",
  48568=>"011101010",
  48569=>"000100011",
  48570=>"101010110",
  48571=>"101110000",
  48572=>"000010010",
  48573=>"111001011",
  48574=>"010010111",
  48575=>"110001101",
  48576=>"010101010",
  48577=>"011110110",
  48578=>"001001011",
  48579=>"011101111",
  48580=>"000100011",
  48581=>"000001000",
  48582=>"100001011",
  48583=>"001100010",
  48584=>"110010001",
  48585=>"000000100",
  48586=>"010011111",
  48587=>"101010101",
  48588=>"100101111",
  48589=>"000110111",
  48590=>"111011111",
  48591=>"110100111",
  48592=>"011010011",
  48593=>"000010111",
  48594=>"111000001",
  48595=>"101110010",
  48596=>"011001101",
  48597=>"101010001",
  48598=>"010010110",
  48599=>"001001100",
  48600=>"100010000",
  48601=>"001010010",
  48602=>"101101100",
  48603=>"101101001",
  48604=>"100110011",
  48605=>"100111010",
  48606=>"001001111",
  48607=>"110001001",
  48608=>"111101010",
  48609=>"000000110",
  48610=>"110100011",
  48611=>"110101000",
  48612=>"110011000",
  48613=>"101010110",
  48614=>"010111000",
  48615=>"000011001",
  48616=>"111101111",
  48617=>"100011111",
  48618=>"011110000",
  48619=>"010101100",
  48620=>"101000101",
  48621=>"101000010",
  48622=>"010000111",
  48623=>"010001011",
  48624=>"110101011",
  48625=>"101111011",
  48626=>"000110000",
  48627=>"100001010",
  48628=>"000110011",
  48629=>"110001100",
  48630=>"100011111",
  48631=>"000101100",
  48632=>"001101010",
  48633=>"110100110",
  48634=>"000011100",
  48635=>"111110101",
  48636=>"100100110",
  48637=>"010100101",
  48638=>"000001100",
  48639=>"101010110",
  48640=>"101011001",
  48641=>"110000111",
  48642=>"000110000",
  48643=>"011010011",
  48644=>"000111010",
  48645=>"000011001",
  48646=>"110110101",
  48647=>"101111110",
  48648=>"110101010",
  48649=>"001001010",
  48650=>"110011111",
  48651=>"001100111",
  48652=>"000100000",
  48653=>"110000100",
  48654=>"000111000",
  48655=>"001110011",
  48656=>"110011010",
  48657=>"100111000",
  48658=>"001001011",
  48659=>"010101101",
  48660=>"110011001",
  48661=>"010010110",
  48662=>"100100101",
  48663=>"101011101",
  48664=>"111001010",
  48665=>"110001001",
  48666=>"001001101",
  48667=>"101010001",
  48668=>"011000011",
  48669=>"101010010",
  48670=>"011011001",
  48671=>"101100001",
  48672=>"001011000",
  48673=>"010001110",
  48674=>"110011010",
  48675=>"100011100",
  48676=>"011111101",
  48677=>"100110001",
  48678=>"001111110",
  48679=>"000111001",
  48680=>"101010000",
  48681=>"110011100",
  48682=>"001100000",
  48683=>"101101000",
  48684=>"011101111",
  48685=>"011001011",
  48686=>"111110000",
  48687=>"111001011",
  48688=>"111010100",
  48689=>"100000011",
  48690=>"000100100",
  48691=>"000001100",
  48692=>"001000010",
  48693=>"110100100",
  48694=>"111000010",
  48695=>"111011100",
  48696=>"101111001",
  48697=>"011111111",
  48698=>"101001101",
  48699=>"101111110",
  48700=>"011101010",
  48701=>"100100000",
  48702=>"101001001",
  48703=>"100010101",
  48704=>"111110000",
  48705=>"111111100",
  48706=>"000001101",
  48707=>"001010111",
  48708=>"100000111",
  48709=>"100100110",
  48710=>"111000100",
  48711=>"011010000",
  48712=>"011110111",
  48713=>"011000001",
  48714=>"001010000",
  48715=>"111100100",
  48716=>"110010000",
  48717=>"101110111",
  48718=>"001010101",
  48719=>"011011111",
  48720=>"101010011",
  48721=>"001001010",
  48722=>"100100111",
  48723=>"111011000",
  48724=>"001011100",
  48725=>"001100101",
  48726=>"010100011",
  48727=>"001001011",
  48728=>"001011110",
  48729=>"110010111",
  48730=>"101000010",
  48731=>"010010011",
  48732=>"011101100",
  48733=>"000010001",
  48734=>"001101101",
  48735=>"100100010",
  48736=>"111000111",
  48737=>"010101110",
  48738=>"010110001",
  48739=>"001101110",
  48740=>"111100111",
  48741=>"011010111",
  48742=>"001000100",
  48743=>"110101011",
  48744=>"111000000",
  48745=>"000100101",
  48746=>"101011011",
  48747=>"111011000",
  48748=>"010110111",
  48749=>"101100011",
  48750=>"111101111",
  48751=>"011101011",
  48752=>"010011101",
  48753=>"011000100",
  48754=>"010101111",
  48755=>"011100101",
  48756=>"000011111",
  48757=>"100001000",
  48758=>"010011110",
  48759=>"001010001",
  48760=>"100101100",
  48761=>"110101101",
  48762=>"100011101",
  48763=>"000000110",
  48764=>"011001001",
  48765=>"000101000",
  48766=>"000101000",
  48767=>"100101100",
  48768=>"111111110",
  48769=>"110111110",
  48770=>"001011000",
  48771=>"011110000",
  48772=>"001011111",
  48773=>"000000011",
  48774=>"000000100",
  48775=>"001011011",
  48776=>"111010100",
  48777=>"100100011",
  48778=>"111110101",
  48779=>"011110110",
  48780=>"111011000",
  48781=>"011101101",
  48782=>"111011010",
  48783=>"100111010",
  48784=>"110001000",
  48785=>"110111011",
  48786=>"100011101",
  48787=>"010010110",
  48788=>"111110101",
  48789=>"101100011",
  48790=>"100001100",
  48791=>"101001011",
  48792=>"111110101",
  48793=>"000001011",
  48794=>"010111101",
  48795=>"001010011",
  48796=>"000011100",
  48797=>"010001111",
  48798=>"000010111",
  48799=>"010001100",
  48800=>"010100000",
  48801=>"011100011",
  48802=>"010010100",
  48803=>"011100011",
  48804=>"001101010",
  48805=>"101011011",
  48806=>"111111011",
  48807=>"111001111",
  48808=>"101111111",
  48809=>"010001101",
  48810=>"011100000",
  48811=>"101101000",
  48812=>"011101000",
  48813=>"001000110",
  48814=>"101000000",
  48815=>"000100111",
  48816=>"101001100",
  48817=>"110110001",
  48818=>"001010101",
  48819=>"000010011",
  48820=>"001100110",
  48821=>"010011100",
  48822=>"001100011",
  48823=>"101010000",
  48824=>"101101001",
  48825=>"010101101",
  48826=>"101100010",
  48827=>"010101100",
  48828=>"001110000",
  48829=>"000011011",
  48830=>"001000000",
  48831=>"111000100",
  48832=>"001111001",
  48833=>"100100011",
  48834=>"111011111",
  48835=>"011111011",
  48836=>"111010110",
  48837=>"111111010",
  48838=>"010101111",
  48839=>"010101110",
  48840=>"101001010",
  48841=>"100000000",
  48842=>"111101101",
  48843=>"010111110",
  48844=>"011110001",
  48845=>"101101111",
  48846=>"101111010",
  48847=>"100010011",
  48848=>"011000010",
  48849=>"100011110",
  48850=>"111000011",
  48851=>"111111001",
  48852=>"100010100",
  48853=>"011111110",
  48854=>"101100010",
  48855=>"000000000",
  48856=>"001100000",
  48857=>"010010001",
  48858=>"000111111",
  48859=>"100010001",
  48860=>"110110111",
  48861=>"001101000",
  48862=>"111111101",
  48863=>"001010011",
  48864=>"011111110",
  48865=>"001010110",
  48866=>"100000110",
  48867=>"111010010",
  48868=>"101011101",
  48869=>"010000011",
  48870=>"100000001",
  48871=>"011110110",
  48872=>"000110011",
  48873=>"101110100",
  48874=>"000011101",
  48875=>"111011011",
  48876=>"110000111",
  48877=>"110010011",
  48878=>"010011110",
  48879=>"000111100",
  48880=>"001101001",
  48881=>"011011010",
  48882=>"100010111",
  48883=>"010010010",
  48884=>"111100100",
  48885=>"010001011",
  48886=>"010010011",
  48887=>"101100010",
  48888=>"101001010",
  48889=>"111000110",
  48890=>"000100010",
  48891=>"111001100",
  48892=>"111111000",
  48893=>"100000000",
  48894=>"100001110",
  48895=>"001100100",
  48896=>"100001001",
  48897=>"111000010",
  48898=>"001110111",
  48899=>"101000001",
  48900=>"111101100",
  48901=>"011000110",
  48902=>"101000001",
  48903=>"111110001",
  48904=>"011011111",
  48905=>"111101111",
  48906=>"010111100",
  48907=>"010110110",
  48908=>"011011110",
  48909=>"111111110",
  48910=>"000000101",
  48911=>"011010000",
  48912=>"111110001",
  48913=>"010101111",
  48914=>"010111111",
  48915=>"111111110",
  48916=>"100100111",
  48917=>"010011111",
  48918=>"100010011",
  48919=>"100001101",
  48920=>"010100011",
  48921=>"000100010",
  48922=>"010011110",
  48923=>"110010111",
  48924=>"110011100",
  48925=>"101000010",
  48926=>"010010101",
  48927=>"010100011",
  48928=>"000001100",
  48929=>"011010010",
  48930=>"000100010",
  48931=>"111010010",
  48932=>"011110001",
  48933=>"001101101",
  48934=>"111111000",
  48935=>"000110101",
  48936=>"101111000",
  48937=>"010111000",
  48938=>"011100011",
  48939=>"011000101",
  48940=>"111101111",
  48941=>"111011101",
  48942=>"101110110",
  48943=>"111000001",
  48944=>"110001011",
  48945=>"100011101",
  48946=>"001110001",
  48947=>"101011101",
  48948=>"000001111",
  48949=>"111010111",
  48950=>"100111010",
  48951=>"101110010",
  48952=>"111110111",
  48953=>"111101100",
  48954=>"000110010",
  48955=>"100101100",
  48956=>"110011100",
  48957=>"000010000",
  48958=>"101110011",
  48959=>"101000010",
  48960=>"011000001",
  48961=>"111001100",
  48962=>"001000100",
  48963=>"011011001",
  48964=>"011000101",
  48965=>"001100010",
  48966=>"011101110",
  48967=>"000111110",
  48968=>"000110011",
  48969=>"100100000",
  48970=>"111010011",
  48971=>"001010101",
  48972=>"011101000",
  48973=>"110111011",
  48974=>"000000110",
  48975=>"010101000",
  48976=>"000000010",
  48977=>"111000011",
  48978=>"010011000",
  48979=>"011110010",
  48980=>"100110101",
  48981=>"010101001",
  48982=>"011000010",
  48983=>"110110110",
  48984=>"111011101",
  48985=>"111111101",
  48986=>"000000111",
  48987=>"101000110",
  48988=>"011000001",
  48989=>"110001100",
  48990=>"011110111",
  48991=>"100110011",
  48992=>"100110100",
  48993=>"010010011",
  48994=>"101100000",
  48995=>"110110001",
  48996=>"011001101",
  48997=>"100100011",
  48998=>"101101110",
  48999=>"100100111",
  49000=>"001100010",
  49001=>"110001011",
  49002=>"101101001",
  49003=>"000100001",
  49004=>"010111111",
  49005=>"001111010",
  49006=>"101111100",
  49007=>"001101100",
  49008=>"100000000",
  49009=>"011010000",
  49010=>"101001111",
  49011=>"111111010",
  49012=>"000001000",
  49013=>"101101110",
  49014=>"000000101",
  49015=>"000000110",
  49016=>"011110111",
  49017=>"101110011",
  49018=>"001111100",
  49019=>"011101100",
  49020=>"000001101",
  49021=>"100001110",
  49022=>"110100100",
  49023=>"111110011",
  49024=>"011101000",
  49025=>"101001111",
  49026=>"000111010",
  49027=>"001100000",
  49028=>"001000100",
  49029=>"111100000",
  49030=>"010100111",
  49031=>"101010010",
  49032=>"010000010",
  49033=>"100011001",
  49034=>"011010111",
  49035=>"100011011",
  49036=>"100001000",
  49037=>"100111010",
  49038=>"000001010",
  49039=>"100111101",
  49040=>"001000101",
  49041=>"111100001",
  49042=>"100011001",
  49043=>"101010000",
  49044=>"110101000",
  49045=>"110110010",
  49046=>"100000010",
  49047=>"000011100",
  49048=>"111110000",
  49049=>"000100010",
  49050=>"110110100",
  49051=>"100010110",
  49052=>"010001011",
  49053=>"110011110",
  49054=>"101101010",
  49055=>"010010001",
  49056=>"000110100",
  49057=>"111000001",
  49058=>"111010010",
  49059=>"101000100",
  49060=>"001010101",
  49061=>"000111001",
  49062=>"011010101",
  49063=>"011101001",
  49064=>"101110110",
  49065=>"110001000",
  49066=>"000011111",
  49067=>"100001010",
  49068=>"001001111",
  49069=>"111011111",
  49070=>"001000100",
  49071=>"010100110",
  49072=>"010010110",
  49073=>"110100011",
  49074=>"100001100",
  49075=>"110001011",
  49076=>"111010011",
  49077=>"100011000",
  49078=>"010010101",
  49079=>"111000100",
  49080=>"011001001",
  49081=>"001001010",
  49082=>"000110010",
  49083=>"111110010",
  49084=>"101000100",
  49085=>"000000000",
  49086=>"000100111",
  49087=>"001110000",
  49088=>"011101011",
  49089=>"111100000",
  49090=>"111110011",
  49091=>"110001111",
  49092=>"011011011",
  49093=>"011101111",
  49094=>"100110110",
  49095=>"010000001",
  49096=>"110000001",
  49097=>"011111001",
  49098=>"001110001",
  49099=>"010001010",
  49100=>"111011110",
  49101=>"010000100",
  49102=>"001110100",
  49103=>"111001110",
  49104=>"000010101",
  49105=>"000111000",
  49106=>"101110111",
  49107=>"000101000",
  49108=>"011111010",
  49109=>"101111001",
  49110=>"101110111",
  49111=>"011000110",
  49112=>"011111001",
  49113=>"010111111",
  49114=>"100100100",
  49115=>"100101111",
  49116=>"100001011",
  49117=>"100001110",
  49118=>"100011010",
  49119=>"000110100",
  49120=>"110001110",
  49121=>"001110101",
  49122=>"101101111",
  49123=>"001010100",
  49124=>"000110000",
  49125=>"100011101",
  49126=>"100100010",
  49127=>"110000011",
  49128=>"101101010",
  49129=>"111001011",
  49130=>"100011010",
  49131=>"100111101",
  49132=>"111010101",
  49133=>"100101000",
  49134=>"011001010",
  49135=>"100100000",
  49136=>"000010111",
  49137=>"011101011",
  49138=>"011010100",
  49139=>"001011011",
  49140=>"110100000",
  49141=>"000100110",
  49142=>"011110000",
  49143=>"000100011",
  49144=>"101000101",
  49145=>"011011001",
  49146=>"011110010",
  49147=>"001111001",
  49148=>"110101111",
  49149=>"010000110",
  49150=>"010000001",
  49151=>"100100110",
  49152=>"100110110",
  49153=>"111011011",
  49154=>"011110011",
  49155=>"010101110",
  49156=>"111111111",
  49157=>"011000111",
  49158=>"010001010",
  49159=>"011101100",
  49160=>"001001001",
  49161=>"100110010",
  49162=>"000010001",
  49163=>"100100000",
  49164=>"001000111",
  49165=>"100001100",
  49166=>"101000011",
  49167=>"111010100",
  49168=>"011111001",
  49169=>"010001011",
  49170=>"101000101",
  49171=>"101001100",
  49172=>"111111100",
  49173=>"010000101",
  49174=>"101101100",
  49175=>"001100011",
  49176=>"110111000",
  49177=>"011010111",
  49178=>"100000001",
  49179=>"110001011",
  49180=>"011101001",
  49181=>"100100101",
  49182=>"000001001",
  49183=>"110111010",
  49184=>"000101011",
  49185=>"110101101",
  49186=>"101001100",
  49187=>"010100010",
  49188=>"100111110",
  49189=>"011000010",
  49190=>"101010000",
  49191=>"110001000",
  49192=>"010101001",
  49193=>"001110000",
  49194=>"110100000",
  49195=>"010100011",
  49196=>"111111001",
  49197=>"010010111",
  49198=>"010101001",
  49199=>"101010100",
  49200=>"111110100",
  49201=>"001101011",
  49202=>"100100010",
  49203=>"110101001",
  49204=>"111101000",
  49205=>"101101111",
  49206=>"000010110",
  49207=>"001011101",
  49208=>"101101101",
  49209=>"111011111",
  49210=>"000001101",
  49211=>"011111000",
  49212=>"100010001",
  49213=>"111000100",
  49214=>"101001010",
  49215=>"100101110",
  49216=>"010110110",
  49217=>"001001111",
  49218=>"011000100",
  49219=>"101000001",
  49220=>"011110101",
  49221=>"000010001",
  49222=>"001011110",
  49223=>"000011101",
  49224=>"001100011",
  49225=>"011100001",
  49226=>"100101100",
  49227=>"101001010",
  49228=>"010000010",
  49229=>"000111000",
  49230=>"000011001",
  49231=>"000110110",
  49232=>"010001101",
  49233=>"000000111",
  49234=>"000010100",
  49235=>"101001100",
  49236=>"100000010",
  49237=>"110101101",
  49238=>"110110110",
  49239=>"101111100",
  49240=>"111100110",
  49241=>"001001000",
  49242=>"010111001",
  49243=>"101111101",
  49244=>"001101000",
  49245=>"001011001",
  49246=>"000100100",
  49247=>"010010111",
  49248=>"100111110",
  49249=>"010101011",
  49250=>"010011111",
  49251=>"011000101",
  49252=>"000000110",
  49253=>"011000011",
  49254=>"010000111",
  49255=>"000001101",
  49256=>"111001000",
  49257=>"111011110",
  49258=>"111011000",
  49259=>"100000000",
  49260=>"101100111",
  49261=>"001001011",
  49262=>"110101010",
  49263=>"111000000",
  49264=>"110101001",
  49265=>"011100011",
  49266=>"111110011",
  49267=>"000011000",
  49268=>"111100001",
  49269=>"100101010",
  49270=>"111000001",
  49271=>"110100101",
  49272=>"101100110",
  49273=>"110000011",
  49274=>"001011001",
  49275=>"111110000",
  49276=>"111001001",
  49277=>"000110011",
  49278=>"101100111",
  49279=>"001001001",
  49280=>"100001111",
  49281=>"100100011",
  49282=>"110011001",
  49283=>"101111101",
  49284=>"111011011",
  49285=>"001111000",
  49286=>"100011111",
  49287=>"100000001",
  49288=>"001010011",
  49289=>"101010111",
  49290=>"011000010",
  49291=>"000001100",
  49292=>"100100000",
  49293=>"010011110",
  49294=>"100000000",
  49295=>"011110010",
  49296=>"010100110",
  49297=>"001100100",
  49298=>"010110110",
  49299=>"100010001",
  49300=>"000111001",
  49301=>"110111101",
  49302=>"010011111",
  49303=>"000111100",
  49304=>"001110001",
  49305=>"100100111",
  49306=>"111000111",
  49307=>"000011010",
  49308=>"010011000",
  49309=>"100010000",
  49310=>"011000110",
  49311=>"011011110",
  49312=>"000111001",
  49313=>"010000001",
  49314=>"100011110",
  49315=>"110101000",
  49316=>"100010110",
  49317=>"000101000",
  49318=>"100111100",
  49319=>"010101010",
  49320=>"001011100",
  49321=>"010110111",
  49322=>"110001110",
  49323=>"011010101",
  49324=>"110111000",
  49325=>"000001001",
  49326=>"111010000",
  49327=>"000000101",
  49328=>"000110010",
  49329=>"010010110",
  49330=>"110000111",
  49331=>"001011010",
  49332=>"011110010",
  49333=>"000100110",
  49334=>"001110101",
  49335=>"011110101",
  49336=>"001010001",
  49337=>"100001001",
  49338=>"001100000",
  49339=>"110011011",
  49340=>"000110000",
  49341=>"001101100",
  49342=>"000001100",
  49343=>"110011011",
  49344=>"001001101",
  49345=>"000101101",
  49346=>"110100010",
  49347=>"000100111",
  49348=>"000010100",
  49349=>"001101110",
  49350=>"011111010",
  49351=>"100000010",
  49352=>"000100101",
  49353=>"010000000",
  49354=>"001011001",
  49355=>"111111010",
  49356=>"010000011",
  49357=>"111111011",
  49358=>"000100010",
  49359=>"010000100",
  49360=>"111000000",
  49361=>"010100100",
  49362=>"000110000",
  49363=>"011011011",
  49364=>"111111110",
  49365=>"010100111",
  49366=>"111011000",
  49367=>"001111111",
  49368=>"100100010",
  49369=>"111011000",
  49370=>"101111110",
  49371=>"001000001",
  49372=>"000110001",
  49373=>"001100001",
  49374=>"110000000",
  49375=>"010101011",
  49376=>"001100010",
  49377=>"110011000",
  49378=>"001010101",
  49379=>"011111110",
  49380=>"110100011",
  49381=>"011010101",
  49382=>"011100010",
  49383=>"010101111",
  49384=>"010010000",
  49385=>"001100100",
  49386=>"100011001",
  49387=>"101101111",
  49388=>"011101000",
  49389=>"110111010",
  49390=>"010010110",
  49391=>"001001010",
  49392=>"010000101",
  49393=>"001011110",
  49394=>"101110100",
  49395=>"101100010",
  49396=>"101001001",
  49397=>"110001000",
  49398=>"001011110",
  49399=>"111001111",
  49400=>"101011010",
  49401=>"000100000",
  49402=>"001001110",
  49403=>"100000010",
  49404=>"000000100",
  49405=>"011010000",
  49406=>"101010100",
  49407=>"110111111",
  49408=>"010101001",
  49409=>"010110011",
  49410=>"110110000",
  49411=>"000001111",
  49412=>"000111001",
  49413=>"100011110",
  49414=>"111000011",
  49415=>"100111100",
  49416=>"110001110",
  49417=>"101011111",
  49418=>"111000111",
  49419=>"010001110",
  49420=>"010000001",
  49421=>"100001001",
  49422=>"001011000",
  49423=>"001001010",
  49424=>"101011011",
  49425=>"000001100",
  49426=>"111011010",
  49427=>"011110011",
  49428=>"001011110",
  49429=>"010001000",
  49430=>"101111100",
  49431=>"110111000",
  49432=>"011000010",
  49433=>"011000001",
  49434=>"000111101",
  49435=>"111011010",
  49436=>"001101110",
  49437=>"101000010",
  49438=>"010110111",
  49439=>"111001000",
  49440=>"000001110",
  49441=>"000110001",
  49442=>"011110101",
  49443=>"011010010",
  49444=>"111000011",
  49445=>"010010011",
  49446=>"101010010",
  49447=>"111111111",
  49448=>"001000000",
  49449=>"000010100",
  49450=>"011011000",
  49451=>"100110011",
  49452=>"111101001",
  49453=>"101110111",
  49454=>"001100101",
  49455=>"100100001",
  49456=>"000011110",
  49457=>"110011001",
  49458=>"101000110",
  49459=>"000110000",
  49460=>"110000100",
  49461=>"011010100",
  49462=>"010011110",
  49463=>"010111100",
  49464=>"011100100",
  49465=>"100000011",
  49466=>"111010001",
  49467=>"001010110",
  49468=>"001110111",
  49469=>"100101101",
  49470=>"111110111",
  49471=>"011110101",
  49472=>"010000101",
  49473=>"110001001",
  49474=>"000000101",
  49475=>"100001110",
  49476=>"010000010",
  49477=>"011101000",
  49478=>"000000010",
  49479=>"010011110",
  49480=>"011010100",
  49481=>"001001100",
  49482=>"011110001",
  49483=>"011010101",
  49484=>"001110101",
  49485=>"100111011",
  49486=>"011011001",
  49487=>"111001001",
  49488=>"111000110",
  49489=>"101011101",
  49490=>"101001001",
  49491=>"010101111",
  49492=>"001111010",
  49493=>"010001011",
  49494=>"110100110",
  49495=>"001110011",
  49496=>"000100001",
  49497=>"001001111",
  49498=>"000100100",
  49499=>"111100011",
  49500=>"101110011",
  49501=>"100010110",
  49502=>"111011001",
  49503=>"101001010",
  49504=>"010110010",
  49505=>"011001000",
  49506=>"000100100",
  49507=>"001001000",
  49508=>"110111111",
  49509=>"010101101",
  49510=>"011000001",
  49511=>"000001111",
  49512=>"010000111",
  49513=>"000100111",
  49514=>"000101011",
  49515=>"101110001",
  49516=>"110011110",
  49517=>"010110011",
  49518=>"110110110",
  49519=>"011100000",
  49520=>"000000101",
  49521=>"001000000",
  49522=>"111000100",
  49523=>"001001110",
  49524=>"001000010",
  49525=>"101101001",
  49526=>"101001110",
  49527=>"111010111",
  49528=>"100111010",
  49529=>"010000101",
  49530=>"100001000",
  49531=>"000001110",
  49532=>"111101010",
  49533=>"100001001",
  49534=>"010110000",
  49535=>"110001100",
  49536=>"101111010",
  49537=>"011010000",
  49538=>"110110111",
  49539=>"101101010",
  49540=>"000110110",
  49541=>"101100111",
  49542=>"010111000",
  49543=>"000110001",
  49544=>"001011000",
  49545=>"000001011",
  49546=>"001000000",
  49547=>"110110001",
  49548=>"000011011",
  49549=>"001100111",
  49550=>"010101110",
  49551=>"101101110",
  49552=>"001000000",
  49553=>"011001011",
  49554=>"001000010",
  49555=>"110001010",
  49556=>"000110011",
  49557=>"100111111",
  49558=>"110010111",
  49559=>"001101110",
  49560=>"010101101",
  49561=>"011001101",
  49562=>"110000111",
  49563=>"010111100",
  49564=>"000000000",
  49565=>"001111001",
  49566=>"100001000",
  49567=>"010000110",
  49568=>"111011101",
  49569=>"001101001",
  49570=>"100110001",
  49571=>"010010011",
  49572=>"110101001",
  49573=>"001100001",
  49574=>"110011101",
  49575=>"101000111",
  49576=>"001010110",
  49577=>"000011001",
  49578=>"011101011",
  49579=>"110001000",
  49580=>"101111111",
  49581=>"100001001",
  49582=>"110110000",
  49583=>"100010000",
  49584=>"011110101",
  49585=>"101000110",
  49586=>"100000101",
  49587=>"001001000",
  49588=>"001101111",
  49589=>"011011011",
  49590=>"101110011",
  49591=>"000111011",
  49592=>"100101010",
  49593=>"010101110",
  49594=>"000110001",
  49595=>"100000111",
  49596=>"100001000",
  49597=>"110010010",
  49598=>"010011100",
  49599=>"100010101",
  49600=>"011010010",
  49601=>"110110001",
  49602=>"011001011",
  49603=>"101010101",
  49604=>"011000100",
  49605=>"110101010",
  49606=>"010001000",
  49607=>"101000111",
  49608=>"011000000",
  49609=>"011010100",
  49610=>"101111000",
  49611=>"000100001",
  49612=>"101100110",
  49613=>"000010000",
  49614=>"010101001",
  49615=>"011100101",
  49616=>"110011100",
  49617=>"010010100",
  49618=>"000010000",
  49619=>"111010110",
  49620=>"000111001",
  49621=>"000101010",
  49622=>"011101010",
  49623=>"100101001",
  49624=>"001111100",
  49625=>"110100010",
  49626=>"000010101",
  49627=>"110011010",
  49628=>"110001011",
  49629=>"001100010",
  49630=>"111011010",
  49631=>"110011101",
  49632=>"110010011",
  49633=>"010100111",
  49634=>"010110110",
  49635=>"000011011",
  49636=>"101011101",
  49637=>"110100000",
  49638=>"111000101",
  49639=>"111100011",
  49640=>"100101000",
  49641=>"010110110",
  49642=>"100100001",
  49643=>"010001010",
  49644=>"000001110",
  49645=>"110101010",
  49646=>"001111011",
  49647=>"001001100",
  49648=>"100010011",
  49649=>"110001000",
  49650=>"010010000",
  49651=>"101000000",
  49652=>"111100111",
  49653=>"001100100",
  49654=>"010110111",
  49655=>"101111000",
  49656=>"101110000",
  49657=>"111010010",
  49658=>"001101111",
  49659=>"001110001",
  49660=>"100111101",
  49661=>"011010000",
  49662=>"100100010",
  49663=>"101010100",
  49664=>"010001000",
  49665=>"001101010",
  49666=>"000100101",
  49667=>"000001001",
  49668=>"100011011",
  49669=>"001100100",
  49670=>"001101101",
  49671=>"101100111",
  49672=>"110001010",
  49673=>"000101001",
  49674=>"110110101",
  49675=>"000010101",
  49676=>"110011111",
  49677=>"010110011",
  49678=>"100010000",
  49679=>"100010010",
  49680=>"001010011",
  49681=>"100011101",
  49682=>"010010100",
  49683=>"110111000",
  49684=>"111000111",
  49685=>"000011010",
  49686=>"010001101",
  49687=>"010001100",
  49688=>"110100111",
  49689=>"011010101",
  49690=>"101100000",
  49691=>"001001010",
  49692=>"101010000",
  49693=>"101001000",
  49694=>"101001101",
  49695=>"111110100",
  49696=>"011000011",
  49697=>"000010011",
  49698=>"010010110",
  49699=>"000000011",
  49700=>"100111100",
  49701=>"001001100",
  49702=>"001011000",
  49703=>"010010111",
  49704=>"101001010",
  49705=>"111110111",
  49706=>"101110110",
  49707=>"101111001",
  49708=>"000110011",
  49709=>"110001010",
  49710=>"001001001",
  49711=>"111000100",
  49712=>"110101001",
  49713=>"111000111",
  49714=>"111101101",
  49715=>"101101011",
  49716=>"100111001",
  49717=>"010010000",
  49718=>"100111111",
  49719=>"011010001",
  49720=>"101011101",
  49721=>"000000100",
  49722=>"111100000",
  49723=>"100101110",
  49724=>"010110001",
  49725=>"001011001",
  49726=>"101100100",
  49727=>"010001110",
  49728=>"001101010",
  49729=>"110000010",
  49730=>"100010000",
  49731=>"010110001",
  49732=>"010001101",
  49733=>"100100011",
  49734=>"001100000",
  49735=>"011100111",
  49736=>"111000001",
  49737=>"010101110",
  49738=>"010001100",
  49739=>"100010000",
  49740=>"001100001",
  49741=>"010000100",
  49742=>"101111000",
  49743=>"110111111",
  49744=>"010110000",
  49745=>"011101001",
  49746=>"000011110",
  49747=>"001010000",
  49748=>"010010010",
  49749=>"001100010",
  49750=>"101110100",
  49751=>"001110110",
  49752=>"010101011",
  49753=>"101110110",
  49754=>"000111001",
  49755=>"100000110",
  49756=>"100010011",
  49757=>"011110101",
  49758=>"101011000",
  49759=>"000001101",
  49760=>"000011101",
  49761=>"001111110",
  49762=>"110101000",
  49763=>"110001001",
  49764=>"001110001",
  49765=>"010000110",
  49766=>"111100101",
  49767=>"000000111",
  49768=>"100101100",
  49769=>"001010010",
  49770=>"110101100",
  49771=>"101100110",
  49772=>"101011101",
  49773=>"100001111",
  49774=>"001111111",
  49775=>"111100001",
  49776=>"000001001",
  49777=>"010100100",
  49778=>"110110001",
  49779=>"010001001",
  49780=>"010011000",
  49781=>"100010011",
  49782=>"110100110",
  49783=>"101010111",
  49784=>"010110110",
  49785=>"111101110",
  49786=>"111110111",
  49787=>"100110101",
  49788=>"001001001",
  49789=>"001010011",
  49790=>"001110001",
  49791=>"011000110",
  49792=>"110101000",
  49793=>"111111001",
  49794=>"001111111",
  49795=>"011001111",
  49796=>"100101100",
  49797=>"000001001",
  49798=>"011010111",
  49799=>"010100111",
  49800=>"110101100",
  49801=>"110011010",
  49802=>"010110010",
  49803=>"110101111",
  49804=>"000000010",
  49805=>"001100001",
  49806=>"001110100",
  49807=>"011111111",
  49808=>"011101000",
  49809=>"000010100",
  49810=>"010110110",
  49811=>"101111111",
  49812=>"010000100",
  49813=>"010110000",
  49814=>"001110011",
  49815=>"000000010",
  49816=>"111101010",
  49817=>"111000110",
  49818=>"101001100",
  49819=>"110001111",
  49820=>"001000101",
  49821=>"001010110",
  49822=>"101100001",
  49823=>"101111110",
  49824=>"010010110",
  49825=>"101000000",
  49826=>"001101001",
  49827=>"010001001",
  49828=>"111110100",
  49829=>"110011001",
  49830=>"011111011",
  49831=>"001111010",
  49832=>"110011011",
  49833=>"010000011",
  49834=>"101001101",
  49835=>"001001000",
  49836=>"011010010",
  49837=>"110011001",
  49838=>"111111111",
  49839=>"111100100",
  49840=>"000110001",
  49841=>"100000011",
  49842=>"110000011",
  49843=>"100100001",
  49844=>"001011001",
  49845=>"011101011",
  49846=>"010101100",
  49847=>"010100100",
  49848=>"100111010",
  49849=>"011101000",
  49850=>"001000110",
  49851=>"111001011",
  49852=>"000101011",
  49853=>"001110010",
  49854=>"100001101",
  49855=>"111001011",
  49856=>"001000011",
  49857=>"001010001",
  49858=>"000010100",
  49859=>"110000001",
  49860=>"001011101",
  49861=>"010110010",
  49862=>"011100100",
  49863=>"001110110",
  49864=>"110001000",
  49865=>"100111001",
  49866=>"100001100",
  49867=>"010001010",
  49868=>"100011110",
  49869=>"101110110",
  49870=>"111011000",
  49871=>"101101011",
  49872=>"010000010",
  49873=>"110100111",
  49874=>"111110100",
  49875=>"110011101",
  49876=>"111000001",
  49877=>"000011010",
  49878=>"011101011",
  49879=>"110111010",
  49880=>"010000000",
  49881=>"111011011",
  49882=>"011100101",
  49883=>"100111110",
  49884=>"001000011",
  49885=>"101001010",
  49886=>"110100011",
  49887=>"110111101",
  49888=>"000011011",
  49889=>"111101101",
  49890=>"001101001",
  49891=>"111111011",
  49892=>"110101100",
  49893=>"000000011",
  49894=>"100011011",
  49895=>"010101000",
  49896=>"010001011",
  49897=>"111011101",
  49898=>"100001100",
  49899=>"101010110",
  49900=>"001001100",
  49901=>"110100011",
  49902=>"011010110",
  49903=>"001110110",
  49904=>"011110101",
  49905=>"000100111",
  49906=>"010001010",
  49907=>"111101110",
  49908=>"110011111",
  49909=>"001110011",
  49910=>"100110010",
  49911=>"001010001",
  49912=>"010001110",
  49913=>"010100000",
  49914=>"010010010",
  49915=>"100000100",
  49916=>"100101100",
  49917=>"101010001",
  49918=>"010101111",
  49919=>"010000011",
  49920=>"001100011",
  49921=>"010001010",
  49922=>"010011010",
  49923=>"100000101",
  49924=>"000101010",
  49925=>"101000011",
  49926=>"010011010",
  49927=>"110111011",
  49928=>"000001101",
  49929=>"111110110",
  49930=>"001100110",
  49931=>"111110001",
  49932=>"110111000",
  49933=>"100111101",
  49934=>"010110010",
  49935=>"100111111",
  49936=>"111100011",
  49937=>"101001100",
  49938=>"100100010",
  49939=>"101110011",
  49940=>"111001010",
  49941=>"100001011",
  49942=>"010011001",
  49943=>"100010001",
  49944=>"000001111",
  49945=>"001011101",
  49946=>"000100011",
  49947=>"011100001",
  49948=>"110111010",
  49949=>"001110011",
  49950=>"000000001",
  49951=>"111011000",
  49952=>"010101111",
  49953=>"101101111",
  49954=>"010101000",
  49955=>"011000001",
  49956=>"000100011",
  49957=>"110110010",
  49958=>"100010111",
  49959=>"000111100",
  49960=>"010010110",
  49961=>"111100001",
  49962=>"000101010",
  49963=>"011001100",
  49964=>"101011001",
  49965=>"000100001",
  49966=>"001110001",
  49967=>"110010101",
  49968=>"000001100",
  49969=>"000000101",
  49970=>"001001001",
  49971=>"011010000",
  49972=>"111001101",
  49973=>"101110011",
  49974=>"000011001",
  49975=>"010010110",
  49976=>"101100011",
  49977=>"001100011",
  49978=>"100011100",
  49979=>"100001011",
  49980=>"010000000",
  49981=>"001111010",
  49982=>"100001001",
  49983=>"100111010",
  49984=>"110110010",
  49985=>"001011000",
  49986=>"100000101",
  49987=>"101111101",
  49988=>"101101111",
  49989=>"011011010",
  49990=>"110100110",
  49991=>"010011111",
  49992=>"111011100",
  49993=>"110111000",
  49994=>"101111010",
  49995=>"101100100",
  49996=>"011000100",
  49997=>"111101110",
  49998=>"001000000",
  49999=>"011001110",
  50000=>"111000100",
  50001=>"111111001",
  50002=>"100000110",
  50003=>"010000111",
  50004=>"010000100",
  50005=>"001101100",
  50006=>"010100011",
  50007=>"010110000",
  50008=>"110111011",
  50009=>"011101101",
  50010=>"100011001",
  50011=>"001111010",
  50012=>"000101111",
  50013=>"110100101",
  50014=>"110101000",
  50015=>"100001000",
  50016=>"100111110",
  50017=>"010000010",
  50018=>"100001100",
  50019=>"100011011",
  50020=>"000010011",
  50021=>"101101000",
  50022=>"110100000",
  50023=>"101000001",
  50024=>"111101001",
  50025=>"000010101",
  50026=>"110001000",
  50027=>"011111010",
  50028=>"110000110",
  50029=>"011010010",
  50030=>"001001111",
  50031=>"110110101",
  50032=>"011000111",
  50033=>"011000001",
  50034=>"101011100",
  50035=>"101001111",
  50036=>"110010100",
  50037=>"111000011",
  50038=>"000100011",
  50039=>"001000110",
  50040=>"101011000",
  50041=>"001010001",
  50042=>"100110011",
  50043=>"100011111",
  50044=>"010001001",
  50045=>"011000010",
  50046=>"001110111",
  50047=>"100110011",
  50048=>"101111101",
  50049=>"011011001",
  50050=>"001010111",
  50051=>"011101101",
  50052=>"011110111",
  50053=>"000011000",
  50054=>"011110110",
  50055=>"000001100",
  50056=>"011001000",
  50057=>"000010110",
  50058=>"001010011",
  50059=>"010111010",
  50060=>"101000100",
  50061=>"010010000",
  50062=>"000111001",
  50063=>"010010001",
  50064=>"110000000",
  50065=>"110111110",
  50066=>"100010001",
  50067=>"100101111",
  50068=>"110101100",
  50069=>"000011010",
  50070=>"001100010",
  50071=>"100111110",
  50072=>"111101110",
  50073=>"110011010",
  50074=>"001110110",
  50075=>"101010110",
  50076=>"010111011",
  50077=>"001011111",
  50078=>"010001011",
  50079=>"100011010",
  50080=>"000000101",
  50081=>"100000110",
  50082=>"100010010",
  50083=>"100000010",
  50084=>"110100011",
  50085=>"111101101",
  50086=>"000001110",
  50087=>"111110011",
  50088=>"110101011",
  50089=>"010010101",
  50090=>"010010001",
  50091=>"110010101",
  50092=>"000001111",
  50093=>"010111100",
  50094=>"001110001",
  50095=>"110000100",
  50096=>"011011010",
  50097=>"011111010",
  50098=>"111111011",
  50099=>"100110100",
  50100=>"111100010",
  50101=>"101011101",
  50102=>"010010010",
  50103=>"010011110",
  50104=>"000000001",
  50105=>"101011011",
  50106=>"111011101",
  50107=>"001001011",
  50108=>"110000001",
  50109=>"110101011",
  50110=>"010000001",
  50111=>"011000001",
  50112=>"000010011",
  50113=>"101001101",
  50114=>"000001110",
  50115=>"011001001",
  50116=>"100001011",
  50117=>"010111001",
  50118=>"110001101",
  50119=>"110000111",
  50120=>"011011011",
  50121=>"111111111",
  50122=>"101101101",
  50123=>"100101000",
  50124=>"111110101",
  50125=>"011001101",
  50126=>"010010001",
  50127=>"000000001",
  50128=>"111111000",
  50129=>"010001000",
  50130=>"111011100",
  50131=>"110101101",
  50132=>"011101000",
  50133=>"011110010",
  50134=>"000101110",
  50135=>"101101011",
  50136=>"000000100",
  50137=>"011001011",
  50138=>"011100010",
  50139=>"000000001",
  50140=>"100101001",
  50141=>"111110011",
  50142=>"000000101",
  50143=>"100110111",
  50144=>"101111011",
  50145=>"110000011",
  50146=>"110100100",
  50147=>"001110111",
  50148=>"001111011",
  50149=>"111100011",
  50150=>"100100100",
  50151=>"111101011",
  50152=>"110101100",
  50153=>"001110011",
  50154=>"001001011",
  50155=>"001101001",
  50156=>"010010010",
  50157=>"010000010",
  50158=>"110010011",
  50159=>"111100100",
  50160=>"100011010",
  50161=>"111001001",
  50162=>"101000000",
  50163=>"001100111",
  50164=>"110100101",
  50165=>"011110000",
  50166=>"110110110",
  50167=>"111000101",
  50168=>"010100100",
  50169=>"110001001",
  50170=>"111100010",
  50171=>"111010111",
  50172=>"000011010",
  50173=>"000001100",
  50174=>"110010100",
  50175=>"001000001",
  50176=>"011010001",
  50177=>"001100100",
  50178=>"001011111",
  50179=>"100111111",
  50180=>"111000010",
  50181=>"110111010",
  50182=>"111100100",
  50183=>"111111101",
  50184=>"101110001",
  50185=>"110000000",
  50186=>"001110001",
  50187=>"010010100",
  50188=>"111110111",
  50189=>"011010100",
  50190=>"011011000",
  50191=>"110101010",
  50192=>"111010000",
  50193=>"000000010",
  50194=>"110101000",
  50195=>"000011001",
  50196=>"000000000",
  50197=>"000001110",
  50198=>"100111111",
  50199=>"111000101",
  50200=>"100010111",
  50201=>"000011011",
  50202=>"101011000",
  50203=>"101111110",
  50204=>"010101011",
  50205=>"110110100",
  50206=>"000010000",
  50207=>"101001111",
  50208=>"000100011",
  50209=>"000001101",
  50210=>"001101100",
  50211=>"000000100",
  50212=>"100010010",
  50213=>"010100110",
  50214=>"100100010",
  50215=>"001111100",
  50216=>"010011111",
  50217=>"001101011",
  50218=>"110100010",
  50219=>"010100111",
  50220=>"100101001",
  50221=>"111101001",
  50222=>"011101110",
  50223=>"111110111",
  50224=>"010000000",
  50225=>"101111111",
  50226=>"001100111",
  50227=>"100110000",
  50228=>"001100100",
  50229=>"010101000",
  50230=>"010001100",
  50231=>"100011110",
  50232=>"000001100",
  50233=>"100110100",
  50234=>"010001100",
  50235=>"100100111",
  50236=>"101000110",
  50237=>"110011100",
  50238=>"101011011",
  50239=>"001000010",
  50240=>"100101100",
  50241=>"101101001",
  50242=>"001000001",
  50243=>"111010000",
  50244=>"100011101",
  50245=>"110111001",
  50246=>"111101001",
  50247=>"110100001",
  50248=>"000111110",
  50249=>"111110101",
  50250=>"010001011",
  50251=>"000100000",
  50252=>"101011001",
  50253=>"100011010",
  50254=>"100100100",
  50255=>"111111110",
  50256=>"001010011",
  50257=>"001000010",
  50258=>"111000011",
  50259=>"101001001",
  50260=>"111010001",
  50261=>"111110000",
  50262=>"001000111",
  50263=>"111000110",
  50264=>"111010110",
  50265=>"000010110",
  50266=>"011001010",
  50267=>"000010110",
  50268=>"000000001",
  50269=>"101001110",
  50270=>"011000011",
  50271=>"111011101",
  50272=>"000000011",
  50273=>"110110011",
  50274=>"100110011",
  50275=>"000100101",
  50276=>"000011111",
  50277=>"000001000",
  50278=>"100110100",
  50279=>"100110110",
  50280=>"111000100",
  50281=>"111100011",
  50282=>"101100111",
  50283=>"011000110",
  50284=>"111100100",
  50285=>"101010010",
  50286=>"000001100",
  50287=>"001101100",
  50288=>"100001011",
  50289=>"010111100",
  50290=>"011100101",
  50291=>"011001111",
  50292=>"110111001",
  50293=>"101011100",
  50294=>"100000011",
  50295=>"010000001",
  50296=>"000001001",
  50297=>"100100001",
  50298=>"011011010",
  50299=>"101100010",
  50300=>"001001101",
  50301=>"100111010",
  50302=>"001001010",
  50303=>"011000111",
  50304=>"100001110",
  50305=>"000000010",
  50306=>"010011000",
  50307=>"101011000",
  50308=>"000001011",
  50309=>"101011001",
  50310=>"001011101",
  50311=>"110110101",
  50312=>"000000100",
  50313=>"011111101",
  50314=>"011001100",
  50315=>"110111001",
  50316=>"010101011",
  50317=>"001011101",
  50318=>"000101111",
  50319=>"011101001",
  50320=>"111111011",
  50321=>"110100101",
  50322=>"100101101",
  50323=>"000000110",
  50324=>"100011011",
  50325=>"110101011",
  50326=>"100111101",
  50327=>"011001111",
  50328=>"000101101",
  50329=>"101010110",
  50330=>"001010001",
  50331=>"000001011",
  50332=>"001001011",
  50333=>"010001111",
  50334=>"100100111",
  50335=>"101000010",
  50336=>"000100111",
  50337=>"010010001",
  50338=>"100110111",
  50339=>"000011110",
  50340=>"000100110",
  50341=>"000001101",
  50342=>"110001000",
  50343=>"000000100",
  50344=>"101010111",
  50345=>"001010011",
  50346=>"000101111",
  50347=>"001000001",
  50348=>"011101001",
  50349=>"111111001",
  50350=>"001001011",
  50351=>"011100110",
  50352=>"001111101",
  50353=>"010011000",
  50354=>"010100100",
  50355=>"110010111",
  50356=>"100001001",
  50357=>"110000010",
  50358=>"011101101",
  50359=>"101111100",
  50360=>"111111111",
  50361=>"010000100",
  50362=>"101111001",
  50363=>"111000101",
  50364=>"000100010",
  50365=>"101111000",
  50366=>"111111010",
  50367=>"000100000",
  50368=>"010000110",
  50369=>"111110001",
  50370=>"110001001",
  50371=>"000001011",
  50372=>"101101010",
  50373=>"100001111",
  50374=>"111110101",
  50375=>"110100001",
  50376=>"011101110",
  50377=>"111110000",
  50378=>"111100111",
  50379=>"001111000",
  50380=>"000011101",
  50381=>"000111000",
  50382=>"010001111",
  50383=>"000100111",
  50384=>"001000000",
  50385=>"011001111",
  50386=>"001001001",
  50387=>"010011001",
  50388=>"001000011",
  50389=>"000101100",
  50390=>"000000000",
  50391=>"110110101",
  50392=>"100100100",
  50393=>"011110100",
  50394=>"001010010",
  50395=>"110010001",
  50396=>"001101000",
  50397=>"001101101",
  50398=>"100100001",
  50399=>"001011100",
  50400=>"000100011",
  50401=>"011110010",
  50402=>"001101000",
  50403=>"000011110",
  50404=>"000100100",
  50405=>"101001100",
  50406=>"111010100",
  50407=>"001100110",
  50408=>"111100111",
  50409=>"111010010",
  50410=>"001011001",
  50411=>"001110111",
  50412=>"110000011",
  50413=>"110100111",
  50414=>"000000010",
  50415=>"110111100",
  50416=>"100111010",
  50417=>"000110000",
  50418=>"001111101",
  50419=>"111111100",
  50420=>"100100001",
  50421=>"011100110",
  50422=>"110000011",
  50423=>"110000001",
  50424=>"000001001",
  50425=>"011010100",
  50426=>"100011010",
  50427=>"000111011",
  50428=>"110100101",
  50429=>"011111000",
  50430=>"010010111",
  50431=>"001111011",
  50432=>"000101001",
  50433=>"001100101",
  50434=>"010101000",
  50435=>"101001010",
  50436=>"000100011",
  50437=>"011001001",
  50438=>"001001110",
  50439=>"101101100",
  50440=>"101011011",
  50441=>"000001110",
  50442=>"101101110",
  50443=>"111111111",
  50444=>"000011111",
  50445=>"000000001",
  50446=>"010001100",
  50447=>"101111000",
  50448=>"111001110",
  50449=>"110000110",
  50450=>"111011110",
  50451=>"010001111",
  50452=>"100111011",
  50453=>"001100111",
  50454=>"000010001",
  50455=>"100101010",
  50456=>"111000111",
  50457=>"101111011",
  50458=>"110111011",
  50459=>"101111111",
  50460=>"011101011",
  50461=>"001011011",
  50462=>"011010111",
  50463=>"110011001",
  50464=>"010000100",
  50465=>"110001000",
  50466=>"010101001",
  50467=>"000100000",
  50468=>"101101101",
  50469=>"011111001",
  50470=>"011111110",
  50471=>"111010000",
  50472=>"111000111",
  50473=>"100000111",
  50474=>"110001001",
  50475=>"010000100",
  50476=>"010011111",
  50477=>"111011000",
  50478=>"001010010",
  50479=>"010001100",
  50480=>"011000100",
  50481=>"100101100",
  50482=>"110100110",
  50483=>"000010111",
  50484=>"110100001",
  50485=>"110000110",
  50486=>"000001100",
  50487=>"010011010",
  50488=>"110010011",
  50489=>"110111001",
  50490=>"111001111",
  50491=>"110000101",
  50492=>"001010101",
  50493=>"011011110",
  50494=>"100010101",
  50495=>"101100011",
  50496=>"001110100",
  50497=>"000000100",
  50498=>"010110100",
  50499=>"100110011",
  50500=>"111011000",
  50501=>"100100000",
  50502=>"110011001",
  50503=>"010011011",
  50504=>"101010000",
  50505=>"110110001",
  50506=>"010100011",
  50507=>"111111010",
  50508=>"101011110",
  50509=>"001001101",
  50510=>"100110000",
  50511=>"111000010",
  50512=>"011100010",
  50513=>"111110001",
  50514=>"000100011",
  50515=>"110111000",
  50516=>"011101101",
  50517=>"110001111",
  50518=>"110110111",
  50519=>"000001000",
  50520=>"010011000",
  50521=>"100010000",
  50522=>"000010010",
  50523=>"101101000",
  50524=>"011010000",
  50525=>"000011011",
  50526=>"010100101",
  50527=>"110110101",
  50528=>"011011110",
  50529=>"001111001",
  50530=>"000110110",
  50531=>"000010010",
  50532=>"001001101",
  50533=>"000010000",
  50534=>"111100101",
  50535=>"111111110",
  50536=>"010001011",
  50537=>"101011100",
  50538=>"101110000",
  50539=>"000100010",
  50540=>"101000000",
  50541=>"111011011",
  50542=>"000011010",
  50543=>"011110100",
  50544=>"100101011",
  50545=>"010010111",
  50546=>"010010001",
  50547=>"000011001",
  50548=>"110010101",
  50549=>"110110100",
  50550=>"001001111",
  50551=>"010111011",
  50552=>"000111011",
  50553=>"001101111",
  50554=>"100000011",
  50555=>"010001011",
  50556=>"011100001",
  50557=>"111111010",
  50558=>"110110000",
  50559=>"111011011",
  50560=>"010010001",
  50561=>"011010000",
  50562=>"000101101",
  50563=>"001010001",
  50564=>"100000101",
  50565=>"110001001",
  50566=>"001000011",
  50567=>"110110111",
  50568=>"011011111",
  50569=>"010110101",
  50570=>"110110101",
  50571=>"000010011",
  50572=>"010110000",
  50573=>"011011001",
  50574=>"001000110",
  50575=>"100001110",
  50576=>"110000101",
  50577=>"111010001",
  50578=>"111111101",
  50579=>"111111111",
  50580=>"000101011",
  50581=>"101111110",
  50582=>"111001001",
  50583=>"111111100",
  50584=>"111011011",
  50585=>"010000000",
  50586=>"101010110",
  50587=>"100100111",
  50588=>"011111000",
  50589=>"001111001",
  50590=>"110011111",
  50591=>"101110111",
  50592=>"011100011",
  50593=>"010111011",
  50594=>"110100000",
  50595=>"000111111",
  50596=>"101101010",
  50597=>"101011010",
  50598=>"011011011",
  50599=>"010110111",
  50600=>"011011111",
  50601=>"100011101",
  50602=>"100100100",
  50603=>"111110011",
  50604=>"111000100",
  50605=>"000011001",
  50606=>"010011101",
  50607=>"010101101",
  50608=>"010000100",
  50609=>"010011010",
  50610=>"111111011",
  50611=>"110110110",
  50612=>"001010010",
  50613=>"010110001",
  50614=>"000101000",
  50615=>"100110110",
  50616=>"101000110",
  50617=>"111010111",
  50618=>"101010011",
  50619=>"100100010",
  50620=>"101001011",
  50621=>"111001011",
  50622=>"011101100",
  50623=>"111110110",
  50624=>"001000011",
  50625=>"011011100",
  50626=>"101110111",
  50627=>"001100110",
  50628=>"100100001",
  50629=>"000010111",
  50630=>"111110001",
  50631=>"010011110",
  50632=>"001101001",
  50633=>"111110110",
  50634=>"010100010",
  50635=>"011010010",
  50636=>"111001100",
  50637=>"001001101",
  50638=>"010010000",
  50639=>"001110111",
  50640=>"001110111",
  50641=>"011010100",
  50642=>"001011000",
  50643=>"011001011",
  50644=>"110011110",
  50645=>"001100100",
  50646=>"111101010",
  50647=>"001110010",
  50648=>"110101010",
  50649=>"000011100",
  50650=>"111100111",
  50651=>"111110010",
  50652=>"111101101",
  50653=>"000101110",
  50654=>"110000111",
  50655=>"010010001",
  50656=>"001000010",
  50657=>"001010000",
  50658=>"111001101",
  50659=>"111100101",
  50660=>"100010010",
  50661=>"111110100",
  50662=>"101000011",
  50663=>"001110011",
  50664=>"101010001",
  50665=>"010100000",
  50666=>"100001010",
  50667=>"101101100",
  50668=>"110110000",
  50669=>"011100110",
  50670=>"110000101",
  50671=>"111100000",
  50672=>"000011000",
  50673=>"010101010",
  50674=>"010001100",
  50675=>"111100010",
  50676=>"001111110",
  50677=>"101110011",
  50678=>"110000111",
  50679=>"101101110",
  50680=>"111111101",
  50681=>"001001001",
  50682=>"001001110",
  50683=>"111100001",
  50684=>"000000101",
  50685=>"010000101",
  50686=>"100100110",
  50687=>"101110110",
  50688=>"011011111",
  50689=>"001000100",
  50690=>"110000100",
  50691=>"000111010",
  50692=>"100010010",
  50693=>"011010001",
  50694=>"010011111",
  50695=>"011111001",
  50696=>"011110001",
  50697=>"010111101",
  50698=>"111011101",
  50699=>"001000000",
  50700=>"101001111",
  50701=>"111000000",
  50702=>"100111000",
  50703=>"000010000",
  50704=>"000111110",
  50705=>"011111100",
  50706=>"000000110",
  50707=>"000101000",
  50708=>"010101011",
  50709=>"110000001",
  50710=>"101101000",
  50711=>"110010000",
  50712=>"110101111",
  50713=>"010000111",
  50714=>"001010010",
  50715=>"111110011",
  50716=>"100111010",
  50717=>"110000001",
  50718=>"011011100",
  50719=>"110010000",
  50720=>"010101000",
  50721=>"110100000",
  50722=>"010010101",
  50723=>"010111101",
  50724=>"110101011",
  50725=>"100100000",
  50726=>"110111001",
  50727=>"001101000",
  50728=>"111100100",
  50729=>"011010010",
  50730=>"011111110",
  50731=>"010001010",
  50732=>"110010111",
  50733=>"000001111",
  50734=>"100111001",
  50735=>"111101010",
  50736=>"010010000",
  50737=>"000100010",
  50738=>"100110011",
  50739=>"010100100",
  50740=>"001011110",
  50741=>"010110101",
  50742=>"111110111",
  50743=>"001100100",
  50744=>"011001110",
  50745=>"100111011",
  50746=>"100011000",
  50747=>"010001001",
  50748=>"111111101",
  50749=>"100101101",
  50750=>"111110101",
  50751=>"100110101",
  50752=>"001110000",
  50753=>"001110111",
  50754=>"010110110",
  50755=>"100000000",
  50756=>"011101011",
  50757=>"000011000",
  50758=>"101101000",
  50759=>"110010100",
  50760=>"110111100",
  50761=>"111001100",
  50762=>"111100010",
  50763=>"111100100",
  50764=>"011010011",
  50765=>"100001000",
  50766=>"110001110",
  50767=>"010010101",
  50768=>"101100101",
  50769=>"111111011",
  50770=>"111010000",
  50771=>"011011100",
  50772=>"100110111",
  50773=>"011010110",
  50774=>"000100000",
  50775=>"101111001",
  50776=>"011010110",
  50777=>"011101010",
  50778=>"011011111",
  50779=>"110101001",
  50780=>"100000001",
  50781=>"000100010",
  50782=>"010011010",
  50783=>"001111100",
  50784=>"101111001",
  50785=>"110100000",
  50786=>"111011111",
  50787=>"000111010",
  50788=>"010100000",
  50789=>"101100101",
  50790=>"110011111",
  50791=>"010001100",
  50792=>"110000001",
  50793=>"111101011",
  50794=>"010010000",
  50795=>"101101100",
  50796=>"010011010",
  50797=>"110101101",
  50798=>"011000000",
  50799=>"100100100",
  50800=>"101001101",
  50801=>"100001001",
  50802=>"011100010",
  50803=>"011010000",
  50804=>"110010011",
  50805=>"001010100",
  50806=>"111010000",
  50807=>"000010101",
  50808=>"111100101",
  50809=>"010111010",
  50810=>"111111001",
  50811=>"000011011",
  50812=>"000001001",
  50813=>"011110100",
  50814=>"100010010",
  50815=>"010001000",
  50816=>"011101000",
  50817=>"110101111",
  50818=>"001100101",
  50819=>"001101101",
  50820=>"001101101",
  50821=>"110000010",
  50822=>"010100101",
  50823=>"011000110",
  50824=>"011001111",
  50825=>"101100011",
  50826=>"000101100",
  50827=>"001111111",
  50828=>"000001101",
  50829=>"011111110",
  50830=>"111101101",
  50831=>"110001100",
  50832=>"010010110",
  50833=>"101101001",
  50834=>"010101011",
  50835=>"001111011",
  50836=>"001000010",
  50837=>"000000000",
  50838=>"101100101",
  50839=>"000100000",
  50840=>"110011110",
  50841=>"000110111",
  50842=>"111010011",
  50843=>"001100001",
  50844=>"101001011",
  50845=>"101110100",
  50846=>"001010010",
  50847=>"011010000",
  50848=>"010110000",
  50849=>"110011011",
  50850=>"010101110",
  50851=>"110110111",
  50852=>"001001000",
  50853=>"000100100",
  50854=>"110001001",
  50855=>"000100110",
  50856=>"100111000",
  50857=>"000110100",
  50858=>"111010011",
  50859=>"000100011",
  50860=>"101110010",
  50861=>"010101101",
  50862=>"111000000",
  50863=>"001100100",
  50864=>"010011010",
  50865=>"001000101",
  50866=>"010111111",
  50867=>"100001011",
  50868=>"101010110",
  50869=>"011011000",
  50870=>"110100111",
  50871=>"111111010",
  50872=>"010111100",
  50873=>"101000011",
  50874=>"110000000",
  50875=>"101011001",
  50876=>"001110000",
  50877=>"100100011",
  50878=>"111010001",
  50879=>"010110010",
  50880=>"010111101",
  50881=>"000110110",
  50882=>"010011011",
  50883=>"010010100",
  50884=>"000001101",
  50885=>"100100010",
  50886=>"011000110",
  50887=>"001010100",
  50888=>"111100101",
  50889=>"011110001",
  50890=>"111101110",
  50891=>"000001010",
  50892=>"000010101",
  50893=>"011001001",
  50894=>"110101111",
  50895=>"000111011",
  50896=>"001011001",
  50897=>"101111111",
  50898=>"000000000",
  50899=>"001101100",
  50900=>"000101110",
  50901=>"010100100",
  50902=>"011111011",
  50903=>"110000101",
  50904=>"110010010",
  50905=>"111000110",
  50906=>"000101101",
  50907=>"001011101",
  50908=>"100010000",
  50909=>"001001101",
  50910=>"100111011",
  50911=>"111110110",
  50912=>"111100111",
  50913=>"010000111",
  50914=>"011110101",
  50915=>"101111011",
  50916=>"011010000",
  50917=>"110110110",
  50918=>"000110110",
  50919=>"010001110",
  50920=>"001100010",
  50921=>"111110111",
  50922=>"001111111",
  50923=>"011101001",
  50924=>"001000010",
  50925=>"111010001",
  50926=>"101101011",
  50927=>"000011001",
  50928=>"110101010",
  50929=>"101011101",
  50930=>"111011011",
  50931=>"111001101",
  50932=>"011101111",
  50933=>"000011011",
  50934=>"101101010",
  50935=>"111100001",
  50936=>"010101100",
  50937=>"100100011",
  50938=>"111000101",
  50939=>"010111010",
  50940=>"100001111",
  50941=>"001100100",
  50942=>"000001000",
  50943=>"011011011",
  50944=>"001001100",
  50945=>"000000011",
  50946=>"111010011",
  50947=>"000001001",
  50948=>"110000001",
  50949=>"110011011",
  50950=>"000000101",
  50951=>"000000100",
  50952=>"000100011",
  50953=>"110000110",
  50954=>"010110110",
  50955=>"001000100",
  50956=>"101001101",
  50957=>"001001001",
  50958=>"101000101",
  50959=>"100011101",
  50960=>"010010010",
  50961=>"001001100",
  50962=>"100010001",
  50963=>"111101100",
  50964=>"110000101",
  50965=>"000010000",
  50966=>"010110100",
  50967=>"011111011",
  50968=>"110110000",
  50969=>"101100001",
  50970=>"000111111",
  50971=>"110100000",
  50972=>"110111001",
  50973=>"011011000",
  50974=>"011110001",
  50975=>"001101010",
  50976=>"001000111",
  50977=>"100011110",
  50978=>"111110000",
  50979=>"000011011",
  50980=>"011001111",
  50981=>"100110111",
  50982=>"111000001",
  50983=>"101010011",
  50984=>"101010110",
  50985=>"001111001",
  50986=>"111100011",
  50987=>"001011000",
  50988=>"001000110",
  50989=>"010100001",
  50990=>"000010111",
  50991=>"000100000",
  50992=>"000111010",
  50993=>"101100011",
  50994=>"001011001",
  50995=>"010111110",
  50996=>"111100110",
  50997=>"100101010",
  50998=>"111101010",
  50999=>"010101100",
  51000=>"100010001",
  51001=>"100001111",
  51002=>"101111110",
  51003=>"100110100",
  51004=>"111110010",
  51005=>"010000101",
  51006=>"000111100",
  51007=>"001010001",
  51008=>"011111111",
  51009=>"100000000",
  51010=>"101011101",
  51011=>"001011110",
  51012=>"001100111",
  51013=>"011011111",
  51014=>"110010011",
  51015=>"101100110",
  51016=>"000111010",
  51017=>"110101110",
  51018=>"001110111",
  51019=>"100101110",
  51020=>"101101111",
  51021=>"110110100",
  51022=>"111000111",
  51023=>"010001111",
  51024=>"011110011",
  51025=>"101111101",
  51026=>"011110000",
  51027=>"000010101",
  51028=>"110101101",
  51029=>"000101111",
  51030=>"000000110",
  51031=>"010111100",
  51032=>"011010011",
  51033=>"000011000",
  51034=>"101001000",
  51035=>"011110100",
  51036=>"101100111",
  51037=>"011001010",
  51038=>"101101111",
  51039=>"001010110",
  51040=>"000000011",
  51041=>"001000101",
  51042=>"000101101",
  51043=>"100011011",
  51044=>"101101111",
  51045=>"000000101",
  51046=>"001100011",
  51047=>"101111110",
  51048=>"001010101",
  51049=>"111011011",
  51050=>"010001000",
  51051=>"011010100",
  51052=>"110101111",
  51053=>"000010101",
  51054=>"001110100",
  51055=>"000000101",
  51056=>"000100000",
  51057=>"000110110",
  51058=>"000111000",
  51059=>"011001100",
  51060=>"001011010",
  51061=>"101101110",
  51062=>"111100100",
  51063=>"000101010",
  51064=>"011110111",
  51065=>"001001101",
  51066=>"110100011",
  51067=>"010111101",
  51068=>"000101000",
  51069=>"000010000",
  51070=>"110101101",
  51071=>"111011110",
  51072=>"000111010",
  51073=>"001100110",
  51074=>"100100010",
  51075=>"000011100",
  51076=>"011000010",
  51077=>"010011010",
  51078=>"001001101",
  51079=>"000011111",
  51080=>"011001100",
  51081=>"000100001",
  51082=>"001000011",
  51083=>"100110101",
  51084=>"011110101",
  51085=>"000110011",
  51086=>"110010111",
  51087=>"111110000",
  51088=>"010011000",
  51089=>"110010111",
  51090=>"101100010",
  51091=>"011000011",
  51092=>"111001011",
  51093=>"011001111",
  51094=>"000000111",
  51095=>"110000000",
  51096=>"000011110",
  51097=>"110010001",
  51098=>"111110100",
  51099=>"110011111",
  51100=>"110110000",
  51101=>"100111001",
  51102=>"001111100",
  51103=>"100011001",
  51104=>"111100111",
  51105=>"101001001",
  51106=>"100010101",
  51107=>"110000111",
  51108=>"110000011",
  51109=>"110010100",
  51110=>"110101000",
  51111=>"010111000",
  51112=>"101011000",
  51113=>"111011011",
  51114=>"011001010",
  51115=>"010001011",
  51116=>"101001101",
  51117=>"000110110",
  51118=>"100100000",
  51119=>"000000100",
  51120=>"001001110",
  51121=>"111001011",
  51122=>"001110011",
  51123=>"111011101",
  51124=>"111010100",
  51125=>"010011111",
  51126=>"110000001",
  51127=>"000011100",
  51128=>"111110100",
  51129=>"111010100",
  51130=>"101101101",
  51131=>"101110000",
  51132=>"000010101",
  51133=>"010111000",
  51134=>"111101011",
  51135=>"011001100",
  51136=>"100000111",
  51137=>"000000100",
  51138=>"110000110",
  51139=>"101101010",
  51140=>"000110000",
  51141=>"101011101",
  51142=>"100111111",
  51143=>"011100100",
  51144=>"010000000",
  51145=>"000101010",
  51146=>"101110010",
  51147=>"110110101",
  51148=>"010011101",
  51149=>"011000110",
  51150=>"001010101",
  51151=>"100011100",
  51152=>"011001100",
  51153=>"100100111",
  51154=>"010111100",
  51155=>"011100101",
  51156=>"100000011",
  51157=>"000000010",
  51158=>"011101010",
  51159=>"110101111",
  51160=>"101110001",
  51161=>"000110110",
  51162=>"100110101",
  51163=>"110001001",
  51164=>"110010101",
  51165=>"110010100",
  51166=>"111010001",
  51167=>"100010111",
  51168=>"110100011",
  51169=>"101011110",
  51170=>"100001111",
  51171=>"000101100",
  51172=>"111001000",
  51173=>"111111001",
  51174=>"000101010",
  51175=>"101001110",
  51176=>"010110000",
  51177=>"110100000",
  51178=>"000001100",
  51179=>"111111000",
  51180=>"001110011",
  51181=>"111111100",
  51182=>"110110001",
  51183=>"101001101",
  51184=>"000111001",
  51185=>"001010110",
  51186=>"000000100",
  51187=>"100000101",
  51188=>"100000100",
  51189=>"010010110",
  51190=>"110011011",
  51191=>"111100011",
  51192=>"010100101",
  51193=>"111011001",
  51194=>"101110111",
  51195=>"111100101",
  51196=>"111011110",
  51197=>"000010010",
  51198=>"001111101",
  51199=>"111001011",
  51200=>"111111101",
  51201=>"100110110",
  51202=>"001010000",
  51203=>"011100010",
  51204=>"001111011",
  51205=>"001111001",
  51206=>"100101101",
  51207=>"101001100",
  51208=>"110110100",
  51209=>"010101000",
  51210=>"111111000",
  51211=>"101011000",
  51212=>"001111110",
  51213=>"110011100",
  51214=>"011111100",
  51215=>"111111101",
  51216=>"101100000",
  51217=>"100000101",
  51218=>"001110010",
  51219=>"011010110",
  51220=>"111011000",
  51221=>"100110100",
  51222=>"011011000",
  51223=>"010010010",
  51224=>"110001111",
  51225=>"101100110",
  51226=>"011110000",
  51227=>"011101011",
  51228=>"101010010",
  51229=>"010100011",
  51230=>"111100111",
  51231=>"010110000",
  51232=>"001111001",
  51233=>"011111111",
  51234=>"000100110",
  51235=>"000010001",
  51236=>"110011011",
  51237=>"100110101",
  51238=>"001011110",
  51239=>"101100100",
  51240=>"111010101",
  51241=>"111110011",
  51242=>"101011111",
  51243=>"000110011",
  51244=>"101100000",
  51245=>"100111101",
  51246=>"010000010",
  51247=>"100011100",
  51248=>"010110010",
  51249=>"110110111",
  51250=>"001000011",
  51251=>"110101011",
  51252=>"010000100",
  51253=>"111110100",
  51254=>"100100101",
  51255=>"101010110",
  51256=>"000100100",
  51257=>"010111110",
  51258=>"100000110",
  51259=>"110000101",
  51260=>"101001000",
  51261=>"010011111",
  51262=>"001000000",
  51263=>"010111111",
  51264=>"100011111",
  51265=>"000000111",
  51266=>"100000001",
  51267=>"001010001",
  51268=>"001110111",
  51269=>"001000011",
  51270=>"111111011",
  51271=>"100100101",
  51272=>"101110101",
  51273=>"111011100",
  51274=>"110101101",
  51275=>"010000100",
  51276=>"000111101",
  51277=>"000111110",
  51278=>"111111011",
  51279=>"111000111",
  51280=>"110010100",
  51281=>"101100000",
  51282=>"010101110",
  51283=>"101110100",
  51284=>"011001001",
  51285=>"001100111",
  51286=>"100101111",
  51287=>"011001111",
  51288=>"010110100",
  51289=>"111000101",
  51290=>"011110001",
  51291=>"111011010",
  51292=>"011000011",
  51293=>"001011010",
  51294=>"001000010",
  51295=>"110011011",
  51296=>"110001001",
  51297=>"001101011",
  51298=>"111000010",
  51299=>"001110001",
  51300=>"000100000",
  51301=>"011001110",
  51302=>"110010010",
  51303=>"100101101",
  51304=>"011110101",
  51305=>"000110010",
  51306=>"100100010",
  51307=>"111000100",
  51308=>"010000001",
  51309=>"111001011",
  51310=>"111010101",
  51311=>"100011110",
  51312=>"010010001",
  51313=>"000011111",
  51314=>"111010011",
  51315=>"110010101",
  51316=>"011110110",
  51317=>"110001000",
  51318=>"000100101",
  51319=>"111111100",
  51320=>"011000000",
  51321=>"010100101",
  51322=>"101011111",
  51323=>"110010101",
  51324=>"110010010",
  51325=>"110000000",
  51326=>"111011111",
  51327=>"011100011",
  51328=>"010101110",
  51329=>"001001110",
  51330=>"110001101",
  51331=>"111111100",
  51332=>"100000111",
  51333=>"001100101",
  51334=>"000111111",
  51335=>"111001011",
  51336=>"101110000",
  51337=>"111001100",
  51338=>"001110110",
  51339=>"001011001",
  51340=>"000000010",
  51341=>"101011111",
  51342=>"100000100",
  51343=>"111000110",
  51344=>"111000000",
  51345=>"100101011",
  51346=>"100111001",
  51347=>"010000000",
  51348=>"001000000",
  51349=>"000110100",
  51350=>"100010100",
  51351=>"111011000",
  51352=>"010010010",
  51353=>"111100011",
  51354=>"110110000",
  51355=>"001010101",
  51356=>"000011110",
  51357=>"110100110",
  51358=>"001011101",
  51359=>"011111101",
  51360=>"111110101",
  51361=>"100001110",
  51362=>"110100010",
  51363=>"010100010",
  51364=>"111011000",
  51365=>"010111001",
  51366=>"000001100",
  51367=>"010000011",
  51368=>"001011100",
  51369=>"000111100",
  51370=>"000000011",
  51371=>"110011000",
  51372=>"101010101",
  51373=>"010000110",
  51374=>"100010101",
  51375=>"000101000",
  51376=>"000001010",
  51377=>"101001101",
  51378=>"101100100",
  51379=>"111011000",
  51380=>"011001010",
  51381=>"000101110",
  51382=>"111010110",
  51383=>"110100111",
  51384=>"010111010",
  51385=>"000101000",
  51386=>"100100010",
  51387=>"001011000",
  51388=>"010101111",
  51389=>"110101001",
  51390=>"010101001",
  51391=>"010001110",
  51392=>"001100101",
  51393=>"001010100",
  51394=>"111000100",
  51395=>"101100001",
  51396=>"101010000",
  51397=>"000000110",
  51398=>"011100101",
  51399=>"110010000",
  51400=>"100110101",
  51401=>"101000101",
  51402=>"001110000",
  51403=>"100110111",
  51404=>"100000101",
  51405=>"100111000",
  51406=>"100010110",
  51407=>"101010110",
  51408=>"011001010",
  51409=>"100110000",
  51410=>"011010101",
  51411=>"110000110",
  51412=>"000001110",
  51413=>"000110110",
  51414=>"110110001",
  51415=>"010111001",
  51416=>"100100000",
  51417=>"011110010",
  51418=>"110000111",
  51419=>"001110010",
  51420=>"001011111",
  51421=>"010111111",
  51422=>"010111111",
  51423=>"111010000",
  51424=>"001001010",
  51425=>"000111110",
  51426=>"000011001",
  51427=>"000001010",
  51428=>"100010011",
  51429=>"000111111",
  51430=>"100100100",
  51431=>"000100000",
  51432=>"011001100",
  51433=>"000010011",
  51434=>"100000001",
  51435=>"100100110",
  51436=>"001010110",
  51437=>"001110111",
  51438=>"010010111",
  51439=>"101001011",
  51440=>"000111000",
  51441=>"001001110",
  51442=>"100010010",
  51443=>"000101100",
  51444=>"001001000",
  51445=>"000001101",
  51446=>"100010101",
  51447=>"010000001",
  51448=>"110111000",
  51449=>"110011110",
  51450=>"001100010",
  51451=>"111011100",
  51452=>"011101000",
  51453=>"100000100",
  51454=>"000110111",
  51455=>"000111010",
  51456=>"111000011",
  51457=>"001000010",
  51458=>"111111101",
  51459=>"110011010",
  51460=>"011001000",
  51461=>"110101110",
  51462=>"001010000",
  51463=>"111011110",
  51464=>"011100101",
  51465=>"110001001",
  51466=>"100100101",
  51467=>"000100000",
  51468=>"110110010",
  51469=>"010000001",
  51470=>"101011111",
  51471=>"111011111",
  51472=>"110100001",
  51473=>"011001101",
  51474=>"011011011",
  51475=>"000110000",
  51476=>"110110100",
  51477=>"110000000",
  51478=>"111010011",
  51479=>"000101001",
  51480=>"001001100",
  51481=>"001110000",
  51482=>"001010001",
  51483=>"010111101",
  51484=>"110100110",
  51485=>"100010100",
  51486=>"011101100",
  51487=>"110000000",
  51488=>"110001011",
  51489=>"111011101",
  51490=>"111111110",
  51491=>"100000101",
  51492=>"110001011",
  51493=>"100111000",
  51494=>"001000001",
  51495=>"101000111",
  51496=>"010110000",
  51497=>"010011011",
  51498=>"000010011",
  51499=>"101110001",
  51500=>"010011101",
  51501=>"000111011",
  51502=>"010011110",
  51503=>"111101101",
  51504=>"111000100",
  51505=>"011101000",
  51506=>"000000010",
  51507=>"011110111",
  51508=>"011010110",
  51509=>"011111011",
  51510=>"111111010",
  51511=>"110011110",
  51512=>"010111001",
  51513=>"000111101",
  51514=>"011110110",
  51515=>"001101111",
  51516=>"010001100",
  51517=>"110100111",
  51518=>"001011000",
  51519=>"101111101",
  51520=>"011011001",
  51521=>"111001100",
  51522=>"011001010",
  51523=>"011001000",
  51524=>"111101011",
  51525=>"011111001",
  51526=>"111010101",
  51527=>"001010001",
  51528=>"110111001",
  51529=>"100111011",
  51530=>"100010001",
  51531=>"111000111",
  51532=>"000000010",
  51533=>"000001001",
  51534=>"001000100",
  51535=>"001010010",
  51536=>"100011001",
  51537=>"011000010",
  51538=>"011111110",
  51539=>"101010010",
  51540=>"100000110",
  51541=>"100111100",
  51542=>"110110111",
  51543=>"101010011",
  51544=>"111101110",
  51545=>"000000010",
  51546=>"001001001",
  51547=>"110000000",
  51548=>"101010100",
  51549=>"111110101",
  51550=>"111001100",
  51551=>"101001101",
  51552=>"111010000",
  51553=>"011100101",
  51554=>"000001110",
  51555=>"100001010",
  51556=>"100011110",
  51557=>"011111110",
  51558=>"100111101",
  51559=>"000100000",
  51560=>"001001100",
  51561=>"111101111",
  51562=>"001000111",
  51563=>"100101000",
  51564=>"110110001",
  51565=>"101001010",
  51566=>"011000100",
  51567=>"110101111",
  51568=>"000110010",
  51569=>"011001110",
  51570=>"010100010",
  51571=>"110001111",
  51572=>"010000111",
  51573=>"010010110",
  51574=>"110010110",
  51575=>"100001101",
  51576=>"110000110",
  51577=>"001101100",
  51578=>"000011001",
  51579=>"011100000",
  51580=>"100100110",
  51581=>"011110101",
  51582=>"101011100",
  51583=>"010010001",
  51584=>"110101100",
  51585=>"110001010",
  51586=>"011000100",
  51587=>"101000011",
  51588=>"000100001",
  51589=>"010010010",
  51590=>"000110100",
  51591=>"011010000",
  51592=>"010000000",
  51593=>"011011011",
  51594=>"100100110",
  51595=>"111000110",
  51596=>"101000111",
  51597=>"001011010",
  51598=>"001000001",
  51599=>"101111110",
  51600=>"101111011",
  51601=>"010000000",
  51602=>"001111111",
  51603=>"011010000",
  51604=>"111110111",
  51605=>"001110110",
  51606=>"011100001",
  51607=>"110101011",
  51608=>"110010111",
  51609=>"110110110",
  51610=>"001010011",
  51611=>"111110100",
  51612=>"011001101",
  51613=>"110110100",
  51614=>"000000111",
  51615=>"010110011",
  51616=>"010010010",
  51617=>"011101100",
  51618=>"101010000",
  51619=>"111001111",
  51620=>"001101100",
  51621=>"111111101",
  51622=>"000110010",
  51623=>"010110101",
  51624=>"101001000",
  51625=>"110101000",
  51626=>"000101011",
  51627=>"011110000",
  51628=>"100000010",
  51629=>"010001100",
  51630=>"100010001",
  51631=>"011010101",
  51632=>"000100010",
  51633=>"100011000",
  51634=>"101111011",
  51635=>"001100001",
  51636=>"010111111",
  51637=>"010110111",
  51638=>"100100101",
  51639=>"110011110",
  51640=>"000111110",
  51641=>"100100101",
  51642=>"011000110",
  51643=>"000010010",
  51644=>"001000011",
  51645=>"010101101",
  51646=>"000100100",
  51647=>"010110010",
  51648=>"110001101",
  51649=>"010000111",
  51650=>"111110101",
  51651=>"101110111",
  51652=>"111001000",
  51653=>"100001001",
  51654=>"101100001",
  51655=>"100111011",
  51656=>"111001010",
  51657=>"010101101",
  51658=>"101101011",
  51659=>"011110100",
  51660=>"110100001",
  51661=>"111110011",
  51662=>"011000010",
  51663=>"100000001",
  51664=>"100100010",
  51665=>"001101101",
  51666=>"001010100",
  51667=>"001100011",
  51668=>"010000001",
  51669=>"100110110",
  51670=>"110001001",
  51671=>"000111001",
  51672=>"001011100",
  51673=>"000000101",
  51674=>"110100011",
  51675=>"101110110",
  51676=>"000100111",
  51677=>"011111101",
  51678=>"000011011",
  51679=>"000001000",
  51680=>"011100001",
  51681=>"001010111",
  51682=>"110001110",
  51683=>"100100010",
  51684=>"001000010",
  51685=>"011101110",
  51686=>"011001000",
  51687=>"011010111",
  51688=>"011001001",
  51689=>"010011100",
  51690=>"111110101",
  51691=>"001001111",
  51692=>"111110101",
  51693=>"111010110",
  51694=>"000101000",
  51695=>"001010000",
  51696=>"101101000",
  51697=>"110101111",
  51698=>"000010110",
  51699=>"110011100",
  51700=>"000000010",
  51701=>"101100101",
  51702=>"100110011",
  51703=>"110111001",
  51704=>"101101100",
  51705=>"101000111",
  51706=>"100110111",
  51707=>"010111001",
  51708=>"000000010",
  51709=>"000010111",
  51710=>"100100101",
  51711=>"110101001",
  51712=>"100100100",
  51713=>"001010101",
  51714=>"001111000",
  51715=>"100010111",
  51716=>"100010000",
  51717=>"111110111",
  51718=>"000111111",
  51719=>"000101100",
  51720=>"100110100",
  51721=>"000000001",
  51722=>"001100001",
  51723=>"100001010",
  51724=>"001101100",
  51725=>"010010011",
  51726=>"111011001",
  51727=>"001100001",
  51728=>"000001111",
  51729=>"011100000",
  51730=>"110100001",
  51731=>"011110100",
  51732=>"111010001",
  51733=>"100111100",
  51734=>"010111111",
  51735=>"111111101",
  51736=>"000001010",
  51737=>"010011101",
  51738=>"101000101",
  51739=>"000010111",
  51740=>"011001111",
  51741=>"100000010",
  51742=>"011011001",
  51743=>"110000000",
  51744=>"100001000",
  51745=>"100101010",
  51746=>"101110001",
  51747=>"010100101",
  51748=>"111111100",
  51749=>"010100100",
  51750=>"001110101",
  51751=>"110101111",
  51752=>"010111110",
  51753=>"010111010",
  51754=>"101001010",
  51755=>"001111000",
  51756=>"001011100",
  51757=>"110000110",
  51758=>"000010001",
  51759=>"110011100",
  51760=>"010101010",
  51761=>"100110000",
  51762=>"001000101",
  51763=>"100111111",
  51764=>"110000000",
  51765=>"101110001",
  51766=>"100111101",
  51767=>"101110010",
  51768=>"101011111",
  51769=>"010101010",
  51770=>"001111011",
  51771=>"010111011",
  51772=>"101101001",
  51773=>"010110000",
  51774=>"011011100",
  51775=>"000001000",
  51776=>"111111111",
  51777=>"100111111",
  51778=>"100100111",
  51779=>"101001000",
  51780=>"010100110",
  51781=>"101100111",
  51782=>"010100101",
  51783=>"001001000",
  51784=>"101110111",
  51785=>"101011100",
  51786=>"000001000",
  51787=>"000010010",
  51788=>"111001010",
  51789=>"010100011",
  51790=>"101101011",
  51791=>"010000011",
  51792=>"001010001",
  51793=>"111111010",
  51794=>"111011000",
  51795=>"101100001",
  51796=>"100000010",
  51797=>"011010100",
  51798=>"000000000",
  51799=>"001001101",
  51800=>"111001110",
  51801=>"000100011",
  51802=>"101010000",
  51803=>"011001110",
  51804=>"000100000",
  51805=>"000000010",
  51806=>"000101000",
  51807=>"110001110",
  51808=>"000011010",
  51809=>"110110000",
  51810=>"011110110",
  51811=>"100100000",
  51812=>"011111100",
  51813=>"011010101",
  51814=>"000000001",
  51815=>"000011100",
  51816=>"011010000",
  51817=>"010110001",
  51818=>"111000011",
  51819=>"000101111",
  51820=>"011001001",
  51821=>"101011111",
  51822=>"101111100",
  51823=>"100000000",
  51824=>"110101111",
  51825=>"100101010",
  51826=>"111100010",
  51827=>"011001111",
  51828=>"001100000",
  51829=>"100011010",
  51830=>"010101000",
  51831=>"010001110",
  51832=>"100010000",
  51833=>"010110100",
  51834=>"111110011",
  51835=>"111101100",
  51836=>"011000111",
  51837=>"100011111",
  51838=>"010110001",
  51839=>"100010000",
  51840=>"011010001",
  51841=>"011110111",
  51842=>"110110100",
  51843=>"100000101",
  51844=>"111111001",
  51845=>"000111101",
  51846=>"000011101",
  51847=>"001000101",
  51848=>"000111100",
  51849=>"100000101",
  51850=>"111111000",
  51851=>"100011100",
  51852=>"001000011",
  51853=>"100000111",
  51854=>"000010101",
  51855=>"010001011",
  51856=>"010001010",
  51857=>"100000110",
  51858=>"110100110",
  51859=>"110101010",
  51860=>"000001100",
  51861=>"011101111",
  51862=>"010100101",
  51863=>"101010101",
  51864=>"110101111",
  51865=>"100010000",
  51866=>"000101101",
  51867=>"001011011",
  51868=>"100001000",
  51869=>"111100010",
  51870=>"101011001",
  51871=>"100011101",
  51872=>"010010010",
  51873=>"110011101",
  51874=>"101011111",
  51875=>"110011101",
  51876=>"000101100",
  51877=>"010011101",
  51878=>"111001101",
  51879=>"011000000",
  51880=>"010100110",
  51881=>"010100010",
  51882=>"000000000",
  51883=>"000000101",
  51884=>"101110001",
  51885=>"010000010",
  51886=>"001010010",
  51887=>"000001101",
  51888=>"100000100",
  51889=>"110010010",
  51890=>"100001010",
  51891=>"001000111",
  51892=>"000101100",
  51893=>"010100001",
  51894=>"110001001",
  51895=>"000010000",
  51896=>"001110101",
  51897=>"111101010",
  51898=>"111100101",
  51899=>"000100111",
  51900=>"110010001",
  51901=>"000010000",
  51902=>"011011110",
  51903=>"100001110",
  51904=>"110100000",
  51905=>"111100110",
  51906=>"100001001",
  51907=>"111110010",
  51908=>"101011010",
  51909=>"001100010",
  51910=>"101111111",
  51911=>"000000100",
  51912=>"001000001",
  51913=>"100010110",
  51914=>"101001111",
  51915=>"010001010",
  51916=>"000100000",
  51917=>"111101010",
  51918=>"001100001",
  51919=>"100011011",
  51920=>"101111100",
  51921=>"111111100",
  51922=>"111110110",
  51923=>"101001010",
  51924=>"001010101",
  51925=>"000100111",
  51926=>"111101110",
  51927=>"101000001",
  51928=>"010000101",
  51929=>"010111000",
  51930=>"101101101",
  51931=>"110100011",
  51932=>"000001110",
  51933=>"011000000",
  51934=>"000000101",
  51935=>"101000010",
  51936=>"001110001",
  51937=>"110101001",
  51938=>"101110010",
  51939=>"001100011",
  51940=>"001011001",
  51941=>"010010100",
  51942=>"010100101",
  51943=>"101011000",
  51944=>"111100001",
  51945=>"111101111",
  51946=>"001110001",
  51947=>"001111001",
  51948=>"001001001",
  51949=>"101001011",
  51950=>"001000001",
  51951=>"100111010",
  51952=>"010010110",
  51953=>"100001010",
  51954=>"110011000",
  51955=>"001011110",
  51956=>"000111111",
  51957=>"001110101",
  51958=>"100011000",
  51959=>"100110100",
  51960=>"000010101",
  51961=>"111010010",
  51962=>"111010001",
  51963=>"101100111",
  51964=>"010110100",
  51965=>"100001001",
  51966=>"000000001",
  51967=>"001000011",
  51968=>"000000010",
  51969=>"001011011",
  51970=>"111111111",
  51971=>"000000001",
  51972=>"000001100",
  51973=>"001001110",
  51974=>"010011010",
  51975=>"001010110",
  51976=>"111111111",
  51977=>"111110101",
  51978=>"001010011",
  51979=>"011001001",
  51980=>"001101101",
  51981=>"010011101",
  51982=>"100111000",
  51983=>"000111000",
  51984=>"001101000",
  51985=>"111010000",
  51986=>"001101011",
  51987=>"101001100",
  51988=>"001101000",
  51989=>"001101010",
  51990=>"010110101",
  51991=>"001111000",
  51992=>"100110011",
  51993=>"101011000",
  51994=>"000101111",
  51995=>"111111101",
  51996=>"000001101",
  51997=>"101011011",
  51998=>"010010101",
  51999=>"100000111",
  52000=>"101100010",
  52001=>"110101100",
  52002=>"000000011",
  52003=>"101000011",
  52004=>"011110101",
  52005=>"111111001",
  52006=>"110010000",
  52007=>"101011100",
  52008=>"100111111",
  52009=>"010001011",
  52010=>"101010000",
  52011=>"101111111",
  52012=>"111111011",
  52013=>"111100001",
  52014=>"010000111",
  52015=>"101001101",
  52016=>"010010010",
  52017=>"010110011",
  52018=>"000101110",
  52019=>"001001101",
  52020=>"000100001",
  52021=>"001100101",
  52022=>"101010100",
  52023=>"111011110",
  52024=>"101000010",
  52025=>"110000110",
  52026=>"000010110",
  52027=>"101011101",
  52028=>"111001110",
  52029=>"001000100",
  52030=>"110100100",
  52031=>"011010010",
  52032=>"111011001",
  52033=>"101100100",
  52034=>"010110000",
  52035=>"001000110",
  52036=>"111100000",
  52037=>"010011001",
  52038=>"010000001",
  52039=>"111000011",
  52040=>"011001011",
  52041=>"110101011",
  52042=>"000011101",
  52043=>"000100100",
  52044=>"110011010",
  52045=>"111101101",
  52046=>"001000100",
  52047=>"000010010",
  52048=>"101001010",
  52049=>"011000011",
  52050=>"010001110",
  52051=>"010010010",
  52052=>"100001110",
  52053=>"110011000",
  52054=>"010011101",
  52055=>"000100101",
  52056=>"110101000",
  52057=>"111111100",
  52058=>"111001010",
  52059=>"110000001",
  52060=>"001111001",
  52061=>"110001101",
  52062=>"110100000",
  52063=>"001010111",
  52064=>"000000000",
  52065=>"000011101",
  52066=>"100000010",
  52067=>"010001111",
  52068=>"101100101",
  52069=>"100011000",
  52070=>"000000110",
  52071=>"001111110",
  52072=>"111111011",
  52073=>"111010101",
  52074=>"110011110",
  52075=>"110011110",
  52076=>"000001010",
  52077=>"001000001",
  52078=>"011010010",
  52079=>"100001010",
  52080=>"100010111",
  52081=>"100110001",
  52082=>"100101001",
  52083=>"000100000",
  52084=>"111000110",
  52085=>"000010000",
  52086=>"111100110",
  52087=>"000110010",
  52088=>"000011001",
  52089=>"000101111",
  52090=>"011111100",
  52091=>"110010100",
  52092=>"000001001",
  52093=>"000001111",
  52094=>"101000010",
  52095=>"100011011",
  52096=>"000100101",
  52097=>"100101110",
  52098=>"100000001",
  52099=>"000011000",
  52100=>"011010000",
  52101=>"010010010",
  52102=>"001000001",
  52103=>"011001101",
  52104=>"111001111",
  52105=>"100001000",
  52106=>"111111111",
  52107=>"010110010",
  52108=>"100110111",
  52109=>"110001110",
  52110=>"111011100",
  52111=>"111010001",
  52112=>"010000100",
  52113=>"111111010",
  52114=>"100010100",
  52115=>"100111111",
  52116=>"101111100",
  52117=>"011111111",
  52118=>"001001101",
  52119=>"110000000",
  52120=>"010001100",
  52121=>"111011100",
  52122=>"101111101",
  52123=>"000000110",
  52124=>"011000000",
  52125=>"000000110",
  52126=>"010101000",
  52127=>"010101110",
  52128=>"001001100",
  52129=>"001101001",
  52130=>"000000010",
  52131=>"111101010",
  52132=>"100110111",
  52133=>"111101111",
  52134=>"110010100",
  52135=>"111100000",
  52136=>"101111101",
  52137=>"000110001",
  52138=>"010110001",
  52139=>"100110010",
  52140=>"100010010",
  52141=>"101111101",
  52142=>"010101110",
  52143=>"000010000",
  52144=>"110000000",
  52145=>"110111010",
  52146=>"011110101",
  52147=>"000001101",
  52148=>"000000100",
  52149=>"111101110",
  52150=>"100110100",
  52151=>"101100110",
  52152=>"100110100",
  52153=>"010100010",
  52154=>"001111100",
  52155=>"110100100",
  52156=>"001001110",
  52157=>"110000000",
  52158=>"011110100",
  52159=>"011011110",
  52160=>"011101111",
  52161=>"000100101",
  52162=>"100001111",
  52163=>"111100111",
  52164=>"010000100",
  52165=>"010000111",
  52166=>"111100101",
  52167=>"110110100",
  52168=>"000110001",
  52169=>"100101010",
  52170=>"000111101",
  52171=>"100010110",
  52172=>"011110000",
  52173=>"001001101",
  52174=>"010011001",
  52175=>"100000001",
  52176=>"010110001",
  52177=>"011001111",
  52178=>"011010000",
  52179=>"010000010",
  52180=>"100111000",
  52181=>"011111111",
  52182=>"110011101",
  52183=>"101101010",
  52184=>"001000000",
  52185=>"101010000",
  52186=>"010011010",
  52187=>"111011100",
  52188=>"000100110",
  52189=>"111110010",
  52190=>"001010000",
  52191=>"101010111",
  52192=>"011101000",
  52193=>"110111001",
  52194=>"101001111",
  52195=>"000101011",
  52196=>"101000100",
  52197=>"000110100",
  52198=>"011011010",
  52199=>"010100101",
  52200=>"010000000",
  52201=>"000000000",
  52202=>"101100100",
  52203=>"010000011",
  52204=>"101001111",
  52205=>"100110110",
  52206=>"000010001",
  52207=>"010101111",
  52208=>"101010110",
  52209=>"000101101",
  52210=>"001101010",
  52211=>"111111101",
  52212=>"010110001",
  52213=>"000111101",
  52214=>"011111010",
  52215=>"111000011",
  52216=>"101110111",
  52217=>"000111111",
  52218=>"101000101",
  52219=>"010001010",
  52220=>"001001001",
  52221=>"110000001",
  52222=>"001101010",
  52223=>"001010111",
  52224=>"111111010",
  52225=>"101011010",
  52226=>"011010101",
  52227=>"011110000",
  52228=>"010110001",
  52229=>"110010010",
  52230=>"010000101",
  52231=>"010011000",
  52232=>"110001100",
  52233=>"010011100",
  52234=>"011000010",
  52235=>"111000111",
  52236=>"111110100",
  52237=>"100000101",
  52238=>"000101000",
  52239=>"110100011",
  52240=>"010010110",
  52241=>"100011011",
  52242=>"001100010",
  52243=>"011000010",
  52244=>"111111010",
  52245=>"100110000",
  52246=>"101001100",
  52247=>"010001001",
  52248=>"001000001",
  52249=>"000001010",
  52250=>"011100111",
  52251=>"000011010",
  52252=>"010101010",
  52253=>"110101110",
  52254=>"011011001",
  52255=>"100000000",
  52256=>"011000001",
  52257=>"000000000",
  52258=>"010001100",
  52259=>"111010101",
  52260=>"110010000",
  52261=>"000111100",
  52262=>"101001101",
  52263=>"010011001",
  52264=>"100111100",
  52265=>"001110010",
  52266=>"011100100",
  52267=>"110011010",
  52268=>"101011001",
  52269=>"011011110",
  52270=>"011001101",
  52271=>"010110010",
  52272=>"010011101",
  52273=>"110101100",
  52274=>"110001000",
  52275=>"000000101",
  52276=>"100010110",
  52277=>"101111011",
  52278=>"011000000",
  52279=>"101110000",
  52280=>"000011000",
  52281=>"110100101",
  52282=>"000000110",
  52283=>"010011100",
  52284=>"101000111",
  52285=>"111111110",
  52286=>"011010101",
  52287=>"000011001",
  52288=>"111011010",
  52289=>"001011111",
  52290=>"001101001",
  52291=>"111101001",
  52292=>"100001100",
  52293=>"101000000",
  52294=>"101010001",
  52295=>"000111011",
  52296=>"110000010",
  52297=>"000001001",
  52298=>"110010010",
  52299=>"010010001",
  52300=>"100001100",
  52301=>"001000010",
  52302=>"100100001",
  52303=>"011100001",
  52304=>"011000000",
  52305=>"001101101",
  52306=>"100111111",
  52307=>"110110000",
  52308=>"101110011",
  52309=>"010011000",
  52310=>"100101011",
  52311=>"100011001",
  52312=>"110011000",
  52313=>"101001000",
  52314=>"011001000",
  52315=>"111000010",
  52316=>"010111000",
  52317=>"000000110",
  52318=>"111100011",
  52319=>"100101011",
  52320=>"001101011",
  52321=>"010101100",
  52322=>"000000011",
  52323=>"011111111",
  52324=>"010111010",
  52325=>"100011111",
  52326=>"110100001",
  52327=>"010101101",
  52328=>"100101100",
  52329=>"010011100",
  52330=>"110100111",
  52331=>"111001101",
  52332=>"010101100",
  52333=>"111110010",
  52334=>"000101010",
  52335=>"110110110",
  52336=>"101011111",
  52337=>"010001111",
  52338=>"001100011",
  52339=>"111111111",
  52340=>"101001011",
  52341=>"001001111",
  52342=>"101101000",
  52343=>"111101000",
  52344=>"100101001",
  52345=>"110111000",
  52346=>"100100111",
  52347=>"000100110",
  52348=>"111110011",
  52349=>"001000000",
  52350=>"110100101",
  52351=>"000000000",
  52352=>"011011111",
  52353=>"100001001",
  52354=>"100000111",
  52355=>"111111111",
  52356=>"111111111",
  52357=>"000000000",
  52358=>"000111111",
  52359=>"000000110",
  52360=>"100111011",
  52361=>"000000000",
  52362=>"111100001",
  52363=>"100111000",
  52364=>"110000001",
  52365=>"100100110",
  52366=>"001111011",
  52367=>"110101011",
  52368=>"001010110",
  52369=>"111011111",
  52370=>"000000001",
  52371=>"101111100",
  52372=>"011000110",
  52373=>"101011111",
  52374=>"011010100",
  52375=>"010100111",
  52376=>"011001001",
  52377=>"100110100",
  52378=>"101100001",
  52379=>"110101011",
  52380=>"110111100",
  52381=>"001001110",
  52382=>"000100000",
  52383=>"111101111",
  52384=>"000110111",
  52385=>"010111111",
  52386=>"010011000",
  52387=>"000111010",
  52388=>"110111001",
  52389=>"000100011",
  52390=>"010001110",
  52391=>"000011111",
  52392=>"010001101",
  52393=>"101111001",
  52394=>"010010001",
  52395=>"111100111",
  52396=>"001000111",
  52397=>"011100010",
  52398=>"111101001",
  52399=>"110001101",
  52400=>"101001001",
  52401=>"100000000",
  52402=>"101110101",
  52403=>"110110101",
  52404=>"110110001",
  52405=>"000011011",
  52406=>"101101111",
  52407=>"000100001",
  52408=>"000000100",
  52409=>"101000000",
  52410=>"010110110",
  52411=>"100110110",
  52412=>"000111100",
  52413=>"000001001",
  52414=>"000101000",
  52415=>"011011001",
  52416=>"101000011",
  52417=>"010100011",
  52418=>"110010101",
  52419=>"100000001",
  52420=>"110010010",
  52421=>"100001101",
  52422=>"110111111",
  52423=>"110001111",
  52424=>"101011001",
  52425=>"001011000",
  52426=>"111111101",
  52427=>"111010101",
  52428=>"100110010",
  52429=>"010010001",
  52430=>"000010000",
  52431=>"000011000",
  52432=>"011011000",
  52433=>"001001111",
  52434=>"100100110",
  52435=>"001101010",
  52436=>"000001000",
  52437=>"010110011",
  52438=>"011100100",
  52439=>"010110001",
  52440=>"000110101",
  52441=>"000111011",
  52442=>"111110110",
  52443=>"101000111",
  52444=>"110011111",
  52445=>"100111001",
  52446=>"000100011",
  52447=>"000110101",
  52448=>"000111001",
  52449=>"000010000",
  52450=>"010100010",
  52451=>"010001101",
  52452=>"110111111",
  52453=>"110010000",
  52454=>"100110110",
  52455=>"011000011",
  52456=>"101010100",
  52457=>"110001000",
  52458=>"001100111",
  52459=>"010111111",
  52460=>"101100000",
  52461=>"101101100",
  52462=>"010100011",
  52463=>"100000011",
  52464=>"111110011",
  52465=>"000110010",
  52466=>"010011000",
  52467=>"100011011",
  52468=>"100000100",
  52469=>"001000100",
  52470=>"100011000",
  52471=>"011111110",
  52472=>"001010101",
  52473=>"010110010",
  52474=>"111000111",
  52475=>"111010001",
  52476=>"011100000",
  52477=>"001101001",
  52478=>"101100100",
  52479=>"000110111",
  52480=>"010011101",
  52481=>"111011001",
  52482=>"100111111",
  52483=>"000100100",
  52484=>"101011000",
  52485=>"000011000",
  52486=>"000100100",
  52487=>"011110101",
  52488=>"000000010",
  52489=>"011101110",
  52490=>"110110011",
  52491=>"001000001",
  52492=>"110110110",
  52493=>"000100110",
  52494=>"111101001",
  52495=>"110101001",
  52496=>"000110001",
  52497=>"001011011",
  52498=>"100111110",
  52499=>"111001100",
  52500=>"001111101",
  52501=>"000110010",
  52502=>"101011111",
  52503=>"101100111",
  52504=>"101010000",
  52505=>"111110110",
  52506=>"000011011",
  52507=>"001010011",
  52508=>"010001000",
  52509=>"010011101",
  52510=>"000000101",
  52511=>"101010001",
  52512=>"000100000",
  52513=>"001101100",
  52514=>"001010110",
  52515=>"000110111",
  52516=>"000100011",
  52517=>"110110011",
  52518=>"111110010",
  52519=>"111011001",
  52520=>"101010111",
  52521=>"101110010",
  52522=>"100101110",
  52523=>"100110000",
  52524=>"011010000",
  52525=>"111010011",
  52526=>"111011001",
  52527=>"100100101",
  52528=>"110110110",
  52529=>"111110010",
  52530=>"011110110",
  52531=>"101101000",
  52532=>"001001010",
  52533=>"011111010",
  52534=>"000110001",
  52535=>"111111101",
  52536=>"111100110",
  52537=>"011000011",
  52538=>"100011111",
  52539=>"111010100",
  52540=>"100001100",
  52541=>"011001001",
  52542=>"000111001",
  52543=>"111011000",
  52544=>"000001110",
  52545=>"111101111",
  52546=>"100000001",
  52547=>"110010111",
  52548=>"010000010",
  52549=>"011010000",
  52550=>"001000001",
  52551=>"010100011",
  52552=>"011001000",
  52553=>"000101110",
  52554=>"111100000",
  52555=>"110100110",
  52556=>"001011110",
  52557=>"100110000",
  52558=>"101010111",
  52559=>"111010101",
  52560=>"110010000",
  52561=>"011110010",
  52562=>"000011000",
  52563=>"010110011",
  52564=>"110010000",
  52565=>"110100100",
  52566=>"010010111",
  52567=>"000111000",
  52568=>"001110100",
  52569=>"011010100",
  52570=>"111010010",
  52571=>"010101010",
  52572=>"011110010",
  52573=>"000110101",
  52574=>"111111101",
  52575=>"001110100",
  52576=>"010000000",
  52577=>"011010001",
  52578=>"100110100",
  52579=>"011001010",
  52580=>"101010100",
  52581=>"111101100",
  52582=>"011010001",
  52583=>"000010000",
  52584=>"010111100",
  52585=>"111000100",
  52586=>"010111101",
  52587=>"101011100",
  52588=>"100110111",
  52589=>"110010111",
  52590=>"010010110",
  52591=>"001001101",
  52592=>"010101100",
  52593=>"100111111",
  52594=>"000010000",
  52595=>"110000010",
  52596=>"010110111",
  52597=>"000011000",
  52598=>"001001101",
  52599=>"111010001",
  52600=>"100011110",
  52601=>"010101011",
  52602=>"000101101",
  52603=>"111101000",
  52604=>"100001000",
  52605=>"001110100",
  52606=>"000010110",
  52607=>"111011000",
  52608=>"010011100",
  52609=>"100110010",
  52610=>"011111011",
  52611=>"110110101",
  52612=>"100111111",
  52613=>"101110001",
  52614=>"000110010",
  52615=>"011011010",
  52616=>"000100010",
  52617=>"000101011",
  52618=>"000101000",
  52619=>"111000110",
  52620=>"010000100",
  52621=>"100010011",
  52622=>"100000000",
  52623=>"011101111",
  52624=>"110000100",
  52625=>"001000010",
  52626=>"111110111",
  52627=>"100100110",
  52628=>"110111100",
  52629=>"101010010",
  52630=>"100111000",
  52631=>"011000110",
  52632=>"000001101",
  52633=>"010010100",
  52634=>"111110011",
  52635=>"000100111",
  52636=>"011111111",
  52637=>"000011110",
  52638=>"010101110",
  52639=>"001110101",
  52640=>"101000010",
  52641=>"011010111",
  52642=>"000011000",
  52643=>"001000100",
  52644=>"101100010",
  52645=>"111010101",
  52646=>"111111110",
  52647=>"111011100",
  52648=>"010001111",
  52649=>"000100001",
  52650=>"100000111",
  52651=>"101001010",
  52652=>"001010011",
  52653=>"101000100",
  52654=>"001100000",
  52655=>"010011010",
  52656=>"000010110",
  52657=>"010101111",
  52658=>"100001011",
  52659=>"100011000",
  52660=>"000011111",
  52661=>"111101100",
  52662=>"111000101",
  52663=>"000010010",
  52664=>"010001111",
  52665=>"110111101",
  52666=>"110101100",
  52667=>"011010010",
  52668=>"111110100",
  52669=>"110010100",
  52670=>"001000010",
  52671=>"000001010",
  52672=>"110100010",
  52673=>"000000011",
  52674=>"011011011",
  52675=>"010000100",
  52676=>"101000111",
  52677=>"010000100",
  52678=>"000000011",
  52679=>"001001000",
  52680=>"110001101",
  52681=>"100111100",
  52682=>"100111101",
  52683=>"010110100",
  52684=>"111111111",
  52685=>"101100111",
  52686=>"100111111",
  52687=>"011101001",
  52688=>"110000001",
  52689=>"000011000",
  52690=>"000111001",
  52691=>"001101100",
  52692=>"000011010",
  52693=>"010110100",
  52694=>"001001010",
  52695=>"010100000",
  52696=>"101001001",
  52697=>"000010101",
  52698=>"000110000",
  52699=>"001000010",
  52700=>"001111011",
  52701=>"101010111",
  52702=>"110000001",
  52703=>"010111000",
  52704=>"011100001",
  52705=>"010010010",
  52706=>"011001010",
  52707=>"011010001",
  52708=>"011011010",
  52709=>"100110000",
  52710=>"001001111",
  52711=>"010101100",
  52712=>"010110011",
  52713=>"001001010",
  52714=>"000010000",
  52715=>"000000001",
  52716=>"000000001",
  52717=>"111000001",
  52718=>"010110101",
  52719=>"010000110",
  52720=>"010010010",
  52721=>"110000111",
  52722=>"111010001",
  52723=>"110100000",
  52724=>"000000000",
  52725=>"011010111",
  52726=>"100010110",
  52727=>"010001111",
  52728=>"011110001",
  52729=>"111001011",
  52730=>"000010101",
  52731=>"010001101",
  52732=>"011101001",
  52733=>"110010101",
  52734=>"001110001",
  52735=>"000101101",
  52736=>"010011111",
  52737=>"110111111",
  52738=>"011010111",
  52739=>"111100101",
  52740=>"101001110",
  52741=>"010111100",
  52742=>"111111100",
  52743=>"101011000",
  52744=>"101011100",
  52745=>"000101010",
  52746=>"000011101",
  52747=>"010110101",
  52748=>"001010110",
  52749=>"111011101",
  52750=>"011001000",
  52751=>"010011001",
  52752=>"000000000",
  52753=>"100110101",
  52754=>"011100100",
  52755=>"110111110",
  52756=>"011011111",
  52757=>"011000110",
  52758=>"011000000",
  52759=>"100000100",
  52760=>"000010100",
  52761=>"010111010",
  52762=>"000110011",
  52763=>"111100100",
  52764=>"000001111",
  52765=>"001001000",
  52766=>"110111100",
  52767=>"010010001",
  52768=>"001110100",
  52769=>"011110001",
  52770=>"001001101",
  52771=>"110100001",
  52772=>"110011111",
  52773=>"010011001",
  52774=>"110111100",
  52775=>"010001011",
  52776=>"100010100",
  52777=>"100001011",
  52778=>"001011111",
  52779=>"011010010",
  52780=>"110101001",
  52781=>"010000000",
  52782=>"011000001",
  52783=>"111001100",
  52784=>"001101001",
  52785=>"100111100",
  52786=>"100100111",
  52787=>"101110101",
  52788=>"001000011",
  52789=>"001001100",
  52790=>"100010111",
  52791=>"000110111",
  52792=>"101001110",
  52793=>"001011010",
  52794=>"101110100",
  52795=>"110010101",
  52796=>"100110011",
  52797=>"001010001",
  52798=>"100110011",
  52799=>"001010011",
  52800=>"100100000",
  52801=>"111010101",
  52802=>"101110100",
  52803=>"101000110",
  52804=>"011111000",
  52805=>"000000111",
  52806=>"010000011",
  52807=>"111111101",
  52808=>"000100000",
  52809=>"001000011",
  52810=>"100011111",
  52811=>"001011001",
  52812=>"100101101",
  52813=>"011101011",
  52814=>"100011000",
  52815=>"110111001",
  52816=>"000000000",
  52817=>"001100010",
  52818=>"111111010",
  52819=>"100111000",
  52820=>"000100101",
  52821=>"100000111",
  52822=>"001010110",
  52823=>"110100001",
  52824=>"110111111",
  52825=>"111101001",
  52826=>"110100001",
  52827=>"111100110",
  52828=>"111011111",
  52829=>"010111001",
  52830=>"001110001",
  52831=>"101111111",
  52832=>"101000001",
  52833=>"001111101",
  52834=>"010111110",
  52835=>"000110001",
  52836=>"011110101",
  52837=>"100100101",
  52838=>"010011000",
  52839=>"100011010",
  52840=>"101011101",
  52841=>"110001101",
  52842=>"100111000",
  52843=>"010000010",
  52844=>"000100110",
  52845=>"111101101",
  52846=>"000111010",
  52847=>"011010110",
  52848=>"110110101",
  52849=>"010001011",
  52850=>"000010110",
  52851=>"001100010",
  52852=>"000001000",
  52853=>"101001110",
  52854=>"110111101",
  52855=>"011011001",
  52856=>"001100011",
  52857=>"001100101",
  52858=>"110011001",
  52859=>"111000100",
  52860=>"100111001",
  52861=>"101111111",
  52862=>"001001001",
  52863=>"001100011",
  52864=>"100110000",
  52865=>"000110100",
  52866=>"001111110",
  52867=>"011100101",
  52868=>"010110111",
  52869=>"111000001",
  52870=>"010010111",
  52871=>"011110110",
  52872=>"001101101",
  52873=>"101101000",
  52874=>"100000001",
  52875=>"100010100",
  52876=>"101010011",
  52877=>"001110111",
  52878=>"110111010",
  52879=>"011101001",
  52880=>"010011101",
  52881=>"100101100",
  52882=>"000011001",
  52883=>"110100111",
  52884=>"100101000",
  52885=>"000111000",
  52886=>"001101011",
  52887=>"110101111",
  52888=>"000111110",
  52889=>"110011110",
  52890=>"101111000",
  52891=>"100110001",
  52892=>"100110001",
  52893=>"001001011",
  52894=>"111011011",
  52895=>"000001110",
  52896=>"111110000",
  52897=>"000001001",
  52898=>"100011111",
  52899=>"111101001",
  52900=>"001100000",
  52901=>"000101010",
  52902=>"110101110",
  52903=>"000110110",
  52904=>"100000111",
  52905=>"101000010",
  52906=>"100111111",
  52907=>"100100101",
  52908=>"111010010",
  52909=>"001111111",
  52910=>"110101011",
  52911=>"000101010",
  52912=>"110000100",
  52913=>"101001001",
  52914=>"101110101",
  52915=>"011100111",
  52916=>"010000001",
  52917=>"111101010",
  52918=>"001010101",
  52919=>"001000010",
  52920=>"000101111",
  52921=>"011101110",
  52922=>"001011100",
  52923=>"111100010",
  52924=>"001111110",
  52925=>"101010110",
  52926=>"100001101",
  52927=>"101000000",
  52928=>"110011110",
  52929=>"111110010",
  52930=>"000000101",
  52931=>"000100101",
  52932=>"100111110",
  52933=>"101101101",
  52934=>"001010000",
  52935=>"000000010",
  52936=>"000010100",
  52937=>"101010001",
  52938=>"000011001",
  52939=>"011111101",
  52940=>"100111001",
  52941=>"101001111",
  52942=>"110101111",
  52943=>"101000111",
  52944=>"101111111",
  52945=>"000011000",
  52946=>"101000011",
  52947=>"000011010",
  52948=>"101000011",
  52949=>"001010000",
  52950=>"101010110",
  52951=>"110010101",
  52952=>"000011100",
  52953=>"111100111",
  52954=>"000101101",
  52955=>"001110110",
  52956=>"001110101",
  52957=>"110000000",
  52958=>"110010010",
  52959=>"001110100",
  52960=>"001111100",
  52961=>"010001111",
  52962=>"111001001",
  52963=>"010110010",
  52964=>"101100011",
  52965=>"000100011",
  52966=>"010110110",
  52967=>"101001011",
  52968=>"000101110",
  52969=>"101111100",
  52970=>"100100101",
  52971=>"100110010",
  52972=>"100111110",
  52973=>"111111101",
  52974=>"111000100",
  52975=>"001111111",
  52976=>"010111011",
  52977=>"101101101",
  52978=>"101000110",
  52979=>"110101111",
  52980=>"010010100",
  52981=>"011011010",
  52982=>"111111101",
  52983=>"010110111",
  52984=>"100010110",
  52985=>"110000111",
  52986=>"001101000",
  52987=>"011010101",
  52988=>"100010000",
  52989=>"000100101",
  52990=>"101011111",
  52991=>"101101001",
  52992=>"001101100",
  52993=>"001000001",
  52994=>"101101010",
  52995=>"010001101",
  52996=>"110001101",
  52997=>"000100110",
  52998=>"100100110",
  52999=>"000000011",
  53000=>"001000001",
  53001=>"010001010",
  53002=>"001110111",
  53003=>"000100101",
  53004=>"010101110",
  53005=>"110101110",
  53006=>"010100000",
  53007=>"111001001",
  53008=>"110100101",
  53009=>"000100100",
  53010=>"001100000",
  53011=>"110101010",
  53012=>"000110011",
  53013=>"110010001",
  53014=>"111011100",
  53015=>"111111110",
  53016=>"110011001",
  53017=>"011001010",
  53018=>"101010011",
  53019=>"110111110",
  53020=>"101010011",
  53021=>"111010110",
  53022=>"111101101",
  53023=>"101010110",
  53024=>"111011011",
  53025=>"000000101",
  53026=>"011111011",
  53027=>"101110101",
  53028=>"101000011",
  53029=>"100010010",
  53030=>"000100000",
  53031=>"010001101",
  53032=>"010110001",
  53033=>"111011000",
  53034=>"010101010",
  53035=>"101111000",
  53036=>"010000111",
  53037=>"111110011",
  53038=>"101000110",
  53039=>"101100101",
  53040=>"000000101",
  53041=>"100001100",
  53042=>"111010010",
  53043=>"111000110",
  53044=>"000001001",
  53045=>"010011001",
  53046=>"001110000",
  53047=>"110001101",
  53048=>"010010101",
  53049=>"010110110",
  53050=>"100100000",
  53051=>"010001011",
  53052=>"000010010",
  53053=>"000000111",
  53054=>"000011010",
  53055=>"100111100",
  53056=>"110101111",
  53057=>"010011101",
  53058=>"110111100",
  53059=>"010101011",
  53060=>"111001111",
  53061=>"111000010",
  53062=>"110001100",
  53063=>"000000011",
  53064=>"101100000",
  53065=>"010010111",
  53066=>"010101111",
  53067=>"110011101",
  53068=>"000001010",
  53069=>"100001011",
  53070=>"111100011",
  53071=>"111110000",
  53072=>"110000101",
  53073=>"010010100",
  53074=>"010011011",
  53075=>"011110110",
  53076=>"101011101",
  53077=>"110101100",
  53078=>"101000100",
  53079=>"010110111",
  53080=>"001001001",
  53081=>"110000111",
  53082=>"011111111",
  53083=>"110110010",
  53084=>"110110111",
  53085=>"011110101",
  53086=>"110011000",
  53087=>"001100101",
  53088=>"011010111",
  53089=>"101010100",
  53090=>"000010101",
  53091=>"101011111",
  53092=>"000111100",
  53093=>"001001010",
  53094=>"101011010",
  53095=>"111000110",
  53096=>"000000001",
  53097=>"110001010",
  53098=>"111010000",
  53099=>"010011100",
  53100=>"111001110",
  53101=>"000100010",
  53102=>"110000010",
  53103=>"100011110",
  53104=>"000011001",
  53105=>"111101011",
  53106=>"010011101",
  53107=>"110001100",
  53108=>"011011111",
  53109=>"111111000",
  53110=>"001110010",
  53111=>"101111010",
  53112=>"000101010",
  53113=>"110000110",
  53114=>"000011011",
  53115=>"100000000",
  53116=>"010110000",
  53117=>"110000001",
  53118=>"011100001",
  53119=>"010111111",
  53120=>"111001011",
  53121=>"000001000",
  53122=>"001100000",
  53123=>"111111010",
  53124=>"111011000",
  53125=>"000010101",
  53126=>"001000010",
  53127=>"000010000",
  53128=>"000011011",
  53129=>"100101000",
  53130=>"110110100",
  53131=>"100101010",
  53132=>"111111100",
  53133=>"101010010",
  53134=>"100101000",
  53135=>"111101111",
  53136=>"000001001",
  53137=>"110011110",
  53138=>"111100100",
  53139=>"110101000",
  53140=>"001101010",
  53141=>"101101100",
  53142=>"110000101",
  53143=>"111111010",
  53144=>"111000000",
  53145=>"100100011",
  53146=>"001011101",
  53147=>"110100111",
  53148=>"110001101",
  53149=>"101111110",
  53150=>"001100000",
  53151=>"011110001",
  53152=>"111110100",
  53153=>"101000100",
  53154=>"011110110",
  53155=>"110111011",
  53156=>"010100010",
  53157=>"111010101",
  53158=>"010011000",
  53159=>"000110101",
  53160=>"001110010",
  53161=>"001001011",
  53162=>"000100101",
  53163=>"100101010",
  53164=>"111101100",
  53165=>"010000010",
  53166=>"111100000",
  53167=>"000110010",
  53168=>"011101101",
  53169=>"110111011",
  53170=>"001111111",
  53171=>"111000110",
  53172=>"011111000",
  53173=>"001111011",
  53174=>"100110000",
  53175=>"000100001",
  53176=>"010010100",
  53177=>"001001011",
  53178=>"101100000",
  53179=>"111110110",
  53180=>"110000100",
  53181=>"110000101",
  53182=>"111000010",
  53183=>"010111111",
  53184=>"100001000",
  53185=>"110010010",
  53186=>"110100111",
  53187=>"100000011",
  53188=>"010000111",
  53189=>"111011101",
  53190=>"100111100",
  53191=>"101101010",
  53192=>"110000011",
  53193=>"010111101",
  53194=>"011000000",
  53195=>"001011001",
  53196=>"011010011",
  53197=>"101000000",
  53198=>"110111110",
  53199=>"001011101",
  53200=>"000001010",
  53201=>"110100101",
  53202=>"001100100",
  53203=>"100000101",
  53204=>"100000001",
  53205=>"101111010",
  53206=>"010001001",
  53207=>"000011011",
  53208=>"101000010",
  53209=>"011010101",
  53210=>"011000100",
  53211=>"001010110",
  53212=>"110111101",
  53213=>"011110101",
  53214=>"111101101",
  53215=>"110010100",
  53216=>"000000110",
  53217=>"010101111",
  53218=>"100000011",
  53219=>"100110011",
  53220=>"000011011",
  53221=>"111111110",
  53222=>"111010110",
  53223=>"111101011",
  53224=>"011110101",
  53225=>"010110111",
  53226=>"100100111",
  53227=>"110011111",
  53228=>"000111010",
  53229=>"000111010",
  53230=>"010001110",
  53231=>"010011110",
  53232=>"011111011",
  53233=>"011101101",
  53234=>"101010011",
  53235=>"101010101",
  53236=>"110100111",
  53237=>"111101111",
  53238=>"110111010",
  53239=>"111111011",
  53240=>"010110111",
  53241=>"111000100",
  53242=>"011101111",
  53243=>"010100000",
  53244=>"001010101",
  53245=>"111110100",
  53246=>"110010011",
  53247=>"011000011",
  53248=>"101011010",
  53249=>"111001011",
  53250=>"101010001",
  53251=>"001000011",
  53252=>"101010000",
  53253=>"101110001",
  53254=>"101000001",
  53255=>"010010000",
  53256=>"100101101",
  53257=>"101001001",
  53258=>"000000000",
  53259=>"111011001",
  53260=>"111010001",
  53261=>"101101010",
  53262=>"001101000",
  53263=>"111100111",
  53264=>"101011010",
  53265=>"011110000",
  53266=>"010010001",
  53267=>"100111111",
  53268=>"000110101",
  53269=>"110010011",
  53270=>"000000110",
  53271=>"000001100",
  53272=>"111100001",
  53273=>"001111000",
  53274=>"000111111",
  53275=>"000001000",
  53276=>"001100011",
  53277=>"000010001",
  53278=>"010111011",
  53279=>"111011010",
  53280=>"011001011",
  53281=>"010010010",
  53282=>"010011110",
  53283=>"101100111",
  53284=>"110001001",
  53285=>"111111011",
  53286=>"011111110",
  53287=>"011101110",
  53288=>"101110010",
  53289=>"010111001",
  53290=>"100001110",
  53291=>"111111001",
  53292=>"111100101",
  53293=>"101101001",
  53294=>"101010110",
  53295=>"110000100",
  53296=>"000101110",
  53297=>"010111010",
  53298=>"010010001",
  53299=>"100101001",
  53300=>"011010010",
  53301=>"000101100",
  53302=>"011101000",
  53303=>"110110011",
  53304=>"101001010",
  53305=>"011100011",
  53306=>"001010101",
  53307=>"110110011",
  53308=>"001101111",
  53309=>"101001001",
  53310=>"000110001",
  53311=>"111111111",
  53312=>"011001110",
  53313=>"011000000",
  53314=>"001000100",
  53315=>"001011100",
  53316=>"011101000",
  53317=>"100000000",
  53318=>"101101101",
  53319=>"000011000",
  53320=>"100100000",
  53321=>"001101000",
  53322=>"010001011",
  53323=>"101011011",
  53324=>"000111001",
  53325=>"111011111",
  53326=>"101000000",
  53327=>"001011011",
  53328=>"011110110",
  53329=>"010000011",
  53330=>"011000010",
  53331=>"001101100",
  53332=>"010100110",
  53333=>"011101010",
  53334=>"111111010",
  53335=>"110011100",
  53336=>"110011010",
  53337=>"011000110",
  53338=>"100101011",
  53339=>"011101010",
  53340=>"011111000",
  53341=>"110010111",
  53342=>"010011100",
  53343=>"001001000",
  53344=>"000111110",
  53345=>"000110011",
  53346=>"010000000",
  53347=>"101010011",
  53348=>"100110001",
  53349=>"010010100",
  53350=>"000000000",
  53351=>"000111110",
  53352=>"111101001",
  53353=>"110111000",
  53354=>"100001000",
  53355=>"010010000",
  53356=>"011101100",
  53357=>"110100011",
  53358=>"000101111",
  53359=>"000100001",
  53360=>"001011011",
  53361=>"011100111",
  53362=>"110101111",
  53363=>"111111001",
  53364=>"110110011",
  53365=>"111011001",
  53366=>"011110010",
  53367=>"010111011",
  53368=>"100110111",
  53369=>"000010011",
  53370=>"000000100",
  53371=>"011000101",
  53372=>"011011001",
  53373=>"000011111",
  53374=>"100011000",
  53375=>"000101001",
  53376=>"001001000",
  53377=>"101010100",
  53378=>"000100001",
  53379=>"001111010",
  53380=>"001011001",
  53381=>"111000000",
  53382=>"100001101",
  53383=>"100011000",
  53384=>"111111010",
  53385=>"100110001",
  53386=>"101000100",
  53387=>"011111000",
  53388=>"110011010",
  53389=>"110101111",
  53390=>"110011100",
  53391=>"001100000",
  53392=>"010100001",
  53393=>"110000011",
  53394=>"000011110",
  53395=>"011100101",
  53396=>"000111000",
  53397=>"110000000",
  53398=>"000010101",
  53399=>"001011011",
  53400=>"110010010",
  53401=>"101010100",
  53402=>"100001100",
  53403=>"101100101",
  53404=>"101000100",
  53405=>"110100100",
  53406=>"101011000",
  53407=>"010001011",
  53408=>"010001100",
  53409=>"001111011",
  53410=>"001010100",
  53411=>"001111001",
  53412=>"110111111",
  53413=>"011111100",
  53414=>"011011011",
  53415=>"101001001",
  53416=>"010011101",
  53417=>"111000001",
  53418=>"001100101",
  53419=>"010011000",
  53420=>"011011101",
  53421=>"000101101",
  53422=>"110111101",
  53423=>"000110111",
  53424=>"010011011",
  53425=>"100101111",
  53426=>"111110101",
  53427=>"111101100",
  53428=>"011110100",
  53429=>"000111000",
  53430=>"001011111",
  53431=>"010000011",
  53432=>"000110101",
  53433=>"000110000",
  53434=>"100101010",
  53435=>"111000111",
  53436=>"111110100",
  53437=>"110010011",
  53438=>"011000101",
  53439=>"111100111",
  53440=>"000001110",
  53441=>"011011111",
  53442=>"010011100",
  53443=>"011110000",
  53444=>"001111111",
  53445=>"001010010",
  53446=>"010010110",
  53447=>"101101011",
  53448=>"011110101",
  53449=>"101101001",
  53450=>"100100111",
  53451=>"010000111",
  53452=>"001000100",
  53453=>"011111110",
  53454=>"001111001",
  53455=>"001101100",
  53456=>"001111011",
  53457=>"111111001",
  53458=>"101000100",
  53459=>"101000111",
  53460=>"000001010",
  53461=>"001010100",
  53462=>"001100000",
  53463=>"110000011",
  53464=>"001101000",
  53465=>"001101101",
  53466=>"110001000",
  53467=>"011001010",
  53468=>"001110011",
  53469=>"001000000",
  53470=>"111001111",
  53471=>"001100000",
  53472=>"110100101",
  53473=>"100001001",
  53474=>"111101101",
  53475=>"110010011",
  53476=>"101111100",
  53477=>"110100001",
  53478=>"011111010",
  53479=>"111011101",
  53480=>"100011101",
  53481=>"111011110",
  53482=>"101111101",
  53483=>"100101001",
  53484=>"110100111",
  53485=>"001100010",
  53486=>"010000101",
  53487=>"001001011",
  53488=>"001010000",
  53489=>"011001100",
  53490=>"011100100",
  53491=>"111010111",
  53492=>"100001011",
  53493=>"100010111",
  53494=>"111110100",
  53495=>"101110000",
  53496=>"101100001",
  53497=>"011111111",
  53498=>"100101100",
  53499=>"101001000",
  53500=>"000010110",
  53501=>"101100100",
  53502=>"101110001",
  53503=>"000011110",
  53504=>"000000011",
  53505=>"001111111",
  53506=>"011101111",
  53507=>"000101111",
  53508=>"000111000",
  53509=>"000111001",
  53510=>"010100000",
  53511=>"110010111",
  53512=>"010101110",
  53513=>"100110101",
  53514=>"000000100",
  53515=>"010000000",
  53516=>"101111000",
  53517=>"011100010",
  53518=>"100010010",
  53519=>"000100100",
  53520=>"101100101",
  53521=>"010011111",
  53522=>"000111010",
  53523=>"100000101",
  53524=>"000101000",
  53525=>"111001111",
  53526=>"001011000",
  53527=>"111111110",
  53528=>"111110000",
  53529=>"000000110",
  53530=>"001110100",
  53531=>"011001110",
  53532=>"000111011",
  53533=>"100010100",
  53534=>"011010010",
  53535=>"110000100",
  53536=>"000011110",
  53537=>"011111000",
  53538=>"010101000",
  53539=>"111101011",
  53540=>"001111111",
  53541=>"011100101",
  53542=>"000110000",
  53543=>"110101011",
  53544=>"100000010",
  53545=>"100111111",
  53546=>"001011001",
  53547=>"001000010",
  53548=>"000110000",
  53549=>"110101101",
  53550=>"111110011",
  53551=>"001111001",
  53552=>"101011011",
  53553=>"111000001",
  53554=>"101111010",
  53555=>"000101111",
  53556=>"001011100",
  53557=>"111111000",
  53558=>"001010011",
  53559=>"000110100",
  53560=>"011011010",
  53561=>"000001001",
  53562=>"110111011",
  53563=>"011111010",
  53564=>"000010110",
  53565=>"000000000",
  53566=>"011000101",
  53567=>"111011011",
  53568=>"000101001",
  53569=>"011000000",
  53570=>"000011110",
  53571=>"100010000",
  53572=>"011101111",
  53573=>"111100101",
  53574=>"011011010",
  53575=>"101001000",
  53576=>"100011001",
  53577=>"010000111",
  53578=>"100001010",
  53579=>"011100101",
  53580=>"100110111",
  53581=>"110010100",
  53582=>"111001111",
  53583=>"111100000",
  53584=>"110010011",
  53585=>"110110110",
  53586=>"111111110",
  53587=>"110000011",
  53588=>"001011010",
  53589=>"010111011",
  53590=>"000001110",
  53591=>"010100101",
  53592=>"011010101",
  53593=>"111111100",
  53594=>"101001001",
  53595=>"011010110",
  53596=>"000100010",
  53597=>"011011000",
  53598=>"100011100",
  53599=>"100001011",
  53600=>"101100010",
  53601=>"010001110",
  53602=>"001001001",
  53603=>"011110000",
  53604=>"110001100",
  53605=>"110111101",
  53606=>"001100101",
  53607=>"111010010",
  53608=>"011100100",
  53609=>"110011010",
  53610=>"100100001",
  53611=>"010010001",
  53612=>"101110001",
  53613=>"111000111",
  53614=>"101001110",
  53615=>"111110000",
  53616=>"111110010",
  53617=>"000010011",
  53618=>"101001010",
  53619=>"100100110",
  53620=>"110010011",
  53621=>"111110001",
  53622=>"110100001",
  53623=>"011111011",
  53624=>"000011101",
  53625=>"011101000",
  53626=>"111110010",
  53627=>"011001101",
  53628=>"100000101",
  53629=>"111100110",
  53630=>"000011010",
  53631=>"110101000",
  53632=>"001110100",
  53633=>"100011000",
  53634=>"000000110",
  53635=>"101110000",
  53636=>"010011111",
  53637=>"001010110",
  53638=>"110010010",
  53639=>"011010101",
  53640=>"000001000",
  53641=>"000111101",
  53642=>"000110000",
  53643=>"001011101",
  53644=>"100010000",
  53645=>"001011101",
  53646=>"101011101",
  53647=>"011010110",
  53648=>"001010000",
  53649=>"110001011",
  53650=>"011101000",
  53651=>"010010000",
  53652=>"100101111",
  53653=>"101000011",
  53654=>"100011011",
  53655=>"000101000",
  53656=>"100110001",
  53657=>"111010001",
  53658=>"000011110",
  53659=>"010111001",
  53660=>"111001101",
  53661=>"111110011",
  53662=>"111000110",
  53663=>"010000000",
  53664=>"101000111",
  53665=>"101100101",
  53666=>"000000111",
  53667=>"110010101",
  53668=>"001101111",
  53669=>"110010010",
  53670=>"100111111",
  53671=>"011111111",
  53672=>"001100111",
  53673=>"001001110",
  53674=>"010011111",
  53675=>"100101101",
  53676=>"000000101",
  53677=>"111100100",
  53678=>"000000101",
  53679=>"111100100",
  53680=>"000011101",
  53681=>"010000101",
  53682=>"111101101",
  53683=>"100111010",
  53684=>"100111101",
  53685=>"010010101",
  53686=>"100110001",
  53687=>"010001101",
  53688=>"101101111",
  53689=>"100000010",
  53690=>"110100101",
  53691=>"111000111",
  53692=>"000001001",
  53693=>"111111000",
  53694=>"000110100",
  53695=>"110101100",
  53696=>"010000011",
  53697=>"101101001",
  53698=>"010110001",
  53699=>"100001010",
  53700=>"010010010",
  53701=>"100110100",
  53702=>"000111100",
  53703=>"011100110",
  53704=>"001001110",
  53705=>"010010010",
  53706=>"100010101",
  53707=>"011011111",
  53708=>"110110000",
  53709=>"001100000",
  53710=>"101000000",
  53711=>"100010010",
  53712=>"011101000",
  53713=>"011001010",
  53714=>"010111001",
  53715=>"110110011",
  53716=>"011000011",
  53717=>"011011110",
  53718=>"111110110",
  53719=>"011010101",
  53720=>"000101010",
  53721=>"101110010",
  53722=>"111111111",
  53723=>"001100101",
  53724=>"111001001",
  53725=>"010100101",
  53726=>"000011110",
  53727=>"001000101",
  53728=>"001010011",
  53729=>"100101000",
  53730=>"100001101",
  53731=>"011100100",
  53732=>"111110110",
  53733=>"111110111",
  53734=>"111011000",
  53735=>"011011000",
  53736=>"011101111",
  53737=>"010101111",
  53738=>"111111001",
  53739=>"101001001",
  53740=>"101001101",
  53741=>"100011011",
  53742=>"111000011",
  53743=>"110110000",
  53744=>"100011110",
  53745=>"001110101",
  53746=>"001101111",
  53747=>"011011100",
  53748=>"011101011",
  53749=>"111110010",
  53750=>"011111000",
  53751=>"100010100",
  53752=>"010111111",
  53753=>"101001111",
  53754=>"111010111",
  53755=>"111000000",
  53756=>"011011111",
  53757=>"000000101",
  53758=>"011110011",
  53759=>"001100001",
  53760=>"100111110",
  53761=>"110110010",
  53762=>"101101000",
  53763=>"100001010",
  53764=>"010011101",
  53765=>"100111110",
  53766=>"100111001",
  53767=>"100001000",
  53768=>"000011111",
  53769=>"000000110",
  53770=>"100011010",
  53771=>"101001111",
  53772=>"010110000",
  53773=>"110011100",
  53774=>"000111010",
  53775=>"001100000",
  53776=>"111010110",
  53777=>"000111111",
  53778=>"110100101",
  53779=>"000101010",
  53780=>"101110000",
  53781=>"001110101",
  53782=>"101100100",
  53783=>"100110111",
  53784=>"010010111",
  53785=>"000101010",
  53786=>"100010010",
  53787=>"111111110",
  53788=>"111110000",
  53789=>"001010000",
  53790=>"101001110",
  53791=>"000111110",
  53792=>"001000001",
  53793=>"011010011",
  53794=>"111000000",
  53795=>"001001001",
  53796=>"000010001",
  53797=>"101001001",
  53798=>"001000010",
  53799=>"100111000",
  53800=>"000001101",
  53801=>"011010001",
  53802=>"000001100",
  53803=>"000111001",
  53804=>"110111011",
  53805=>"100101111",
  53806=>"000011110",
  53807=>"110111101",
  53808=>"101111111",
  53809=>"001101101",
  53810=>"001101000",
  53811=>"110111000",
  53812=>"001001100",
  53813=>"110101101",
  53814=>"111100011",
  53815=>"000100100",
  53816=>"110100001",
  53817=>"101111011",
  53818=>"111000000",
  53819=>"011101100",
  53820=>"101101101",
  53821=>"000110101",
  53822=>"111011000",
  53823=>"100101011",
  53824=>"000111111",
  53825=>"101100100",
  53826=>"111101001",
  53827=>"100101101",
  53828=>"010111111",
  53829=>"101010010",
  53830=>"010011110",
  53831=>"011000000",
  53832=>"011111110",
  53833=>"000100010",
  53834=>"011000111",
  53835=>"011110111",
  53836=>"000001111",
  53837=>"101101101",
  53838=>"001110001",
  53839=>"000011110",
  53840=>"010110100",
  53841=>"011100000",
  53842=>"111111010",
  53843=>"100011000",
  53844=>"000100101",
  53845=>"111111111",
  53846=>"000000110",
  53847=>"110010111",
  53848=>"000110101",
  53849=>"000011101",
  53850=>"000111111",
  53851=>"111111110",
  53852=>"111110100",
  53853=>"010011010",
  53854=>"110111001",
  53855=>"000100011",
  53856=>"010101101",
  53857=>"010110100",
  53858=>"101011110",
  53859=>"011001011",
  53860=>"010100011",
  53861=>"011100011",
  53862=>"010010010",
  53863=>"110110011",
  53864=>"010100100",
  53865=>"101110001",
  53866=>"000110001",
  53867=>"111011110",
  53868=>"110110100",
  53869=>"110101000",
  53870=>"010000100",
  53871=>"011001100",
  53872=>"011011101",
  53873=>"010111110",
  53874=>"001010111",
  53875=>"100100111",
  53876=>"000011000",
  53877=>"000101001",
  53878=>"100010111",
  53879=>"100111010",
  53880=>"100010101",
  53881=>"001111101",
  53882=>"100011100",
  53883=>"001110111",
  53884=>"011110011",
  53885=>"010011110",
  53886=>"011110101",
  53887=>"111000001",
  53888=>"011000111",
  53889=>"111000110",
  53890=>"000000000",
  53891=>"111001110",
  53892=>"001101111",
  53893=>"101110010",
  53894=>"011101001",
  53895=>"000011011",
  53896=>"110111001",
  53897=>"001000000",
  53898=>"111010111",
  53899=>"000010001",
  53900=>"010111100",
  53901=>"101101000",
  53902=>"010000010",
  53903=>"010010010",
  53904=>"100001111",
  53905=>"000110110",
  53906=>"001011111",
  53907=>"010010110",
  53908=>"010000101",
  53909=>"101001011",
  53910=>"110110010",
  53911=>"001111110",
  53912=>"111101100",
  53913=>"101000111",
  53914=>"110100110",
  53915=>"101000101",
  53916=>"011100010",
  53917=>"000001000",
  53918=>"101111110",
  53919=>"010111100",
  53920=>"011111101",
  53921=>"101100001",
  53922=>"001010000",
  53923=>"001000110",
  53924=>"110101100",
  53925=>"100110110",
  53926=>"100000101",
  53927=>"001100011",
  53928=>"111111010",
  53929=>"101101000",
  53930=>"100101100",
  53931=>"001100101",
  53932=>"000001001",
  53933=>"010010100",
  53934=>"110101111",
  53935=>"111110001",
  53936=>"101100101",
  53937=>"100000110",
  53938=>"000111101",
  53939=>"101101100",
  53940=>"101100011",
  53941=>"010111111",
  53942=>"001010110",
  53943=>"101101100",
  53944=>"100011101",
  53945=>"100011010",
  53946=>"000111010",
  53947=>"101100011",
  53948=>"111011110",
  53949=>"011000010",
  53950=>"011010001",
  53951=>"011000110",
  53952=>"001011100",
  53953=>"101001110",
  53954=>"011001110",
  53955=>"001000001",
  53956=>"000000000",
  53957=>"100010010",
  53958=>"100110101",
  53959=>"010000000",
  53960=>"001100100",
  53961=>"000000000",
  53962=>"111000000",
  53963=>"111010011",
  53964=>"010111101",
  53965=>"010100000",
  53966=>"101000010",
  53967=>"111011110",
  53968=>"010110111",
  53969=>"101100101",
  53970=>"100101001",
  53971=>"011000110",
  53972=>"001010010",
  53973=>"000000010",
  53974=>"111001111",
  53975=>"011010011",
  53976=>"001000011",
  53977=>"001100011",
  53978=>"000010011",
  53979=>"000000011",
  53980=>"000010101",
  53981=>"100110111",
  53982=>"111000010",
  53983=>"000000010",
  53984=>"111101011",
  53985=>"000010001",
  53986=>"010000101",
  53987=>"100011111",
  53988=>"011011001",
  53989=>"001110000",
  53990=>"011111011",
  53991=>"100001001",
  53992=>"001011100",
  53993=>"000010001",
  53994=>"001000110",
  53995=>"011000001",
  53996=>"000110110",
  53997=>"011101100",
  53998=>"111011101",
  53999=>"100111101",
  54000=>"001001001",
  54001=>"000001011",
  54002=>"111111100",
  54003=>"110010000",
  54004=>"101100111",
  54005=>"010100100",
  54006=>"011111001",
  54007=>"101010101",
  54008=>"011110011",
  54009=>"000011101",
  54010=>"101011001",
  54011=>"011001111",
  54012=>"001011111",
  54013=>"000110100",
  54014=>"000100110",
  54015=>"000010111",
  54016=>"101110110",
  54017=>"110000001",
  54018=>"000111010",
  54019=>"010101010",
  54020=>"001000001",
  54021=>"000000100",
  54022=>"100011000",
  54023=>"000001000",
  54024=>"100000100",
  54025=>"011001000",
  54026=>"100011101",
  54027=>"000011101",
  54028=>"000001000",
  54029=>"100001110",
  54030=>"000000010",
  54031=>"110110010",
  54032=>"011001010",
  54033=>"011011000",
  54034=>"100000100",
  54035=>"111010000",
  54036=>"001000110",
  54037=>"100001000",
  54038=>"110111001",
  54039=>"101100101",
  54040=>"001101101",
  54041=>"111100000",
  54042=>"100001001",
  54043=>"110011101",
  54044=>"101010101",
  54045=>"000001111",
  54046=>"101011000",
  54047=>"000100000",
  54048=>"101111111",
  54049=>"110000010",
  54050=>"010000111",
  54051=>"000000111",
  54052=>"011101011",
  54053=>"000100000",
  54054=>"100101101",
  54055=>"111000100",
  54056=>"000010010",
  54057=>"000111001",
  54058=>"111011001",
  54059=>"000100100",
  54060=>"111011101",
  54061=>"001001010",
  54062=>"111101010",
  54063=>"001001000",
  54064=>"001011000",
  54065=>"001100000",
  54066=>"110011100",
  54067=>"011010010",
  54068=>"100111001",
  54069=>"110010111",
  54070=>"010000010",
  54071=>"111100011",
  54072=>"101001000",
  54073=>"110101100",
  54074=>"011000100",
  54075=>"111101011",
  54076=>"110001000",
  54077=>"000000101",
  54078=>"000011001",
  54079=>"000000011",
  54080=>"011111011",
  54081=>"010100111",
  54082=>"010001000",
  54083=>"101000101",
  54084=>"101110100",
  54085=>"001110111",
  54086=>"110110011",
  54087=>"011000101",
  54088=>"010100100",
  54089=>"010100000",
  54090=>"000111100",
  54091=>"010101010",
  54092=>"110110101",
  54093=>"010111111",
  54094=>"111010010",
  54095=>"110100001",
  54096=>"100010000",
  54097=>"101010110",
  54098=>"000001000",
  54099=>"000110011",
  54100=>"110010001",
  54101=>"111111111",
  54102=>"001010011",
  54103=>"101101110",
  54104=>"100101001",
  54105=>"001100001",
  54106=>"010011101",
  54107=>"001100110",
  54108=>"101001101",
  54109=>"110100000",
  54110=>"101111001",
  54111=>"111111101",
  54112=>"001011110",
  54113=>"011010100",
  54114=>"111000011",
  54115=>"101111101",
  54116=>"011011100",
  54117=>"111000011",
  54118=>"111110001",
  54119=>"001001110",
  54120=>"111110001",
  54121=>"100100011",
  54122=>"001000011",
  54123=>"111011110",
  54124=>"000110110",
  54125=>"001101000",
  54126=>"111000001",
  54127=>"101101011",
  54128=>"010110000",
  54129=>"011000100",
  54130=>"101110010",
  54131=>"011000110",
  54132=>"101001100",
  54133=>"110000111",
  54134=>"000000111",
  54135=>"000010010",
  54136=>"101001000",
  54137=>"001101100",
  54138=>"001101011",
  54139=>"011101011",
  54140=>"000000001",
  54141=>"101001110",
  54142=>"111111100",
  54143=>"010001011",
  54144=>"110010010",
  54145=>"000100001",
  54146=>"010100100",
  54147=>"111101110",
  54148=>"011100111",
  54149=>"011011000",
  54150=>"010110100",
  54151=>"101001111",
  54152=>"010010011",
  54153=>"000111100",
  54154=>"110011111",
  54155=>"111000100",
  54156=>"111110100",
  54157=>"011111000",
  54158=>"110101110",
  54159=>"110100111",
  54160=>"100010001",
  54161=>"101011000",
  54162=>"111111001",
  54163=>"101000010",
  54164=>"000010001",
  54165=>"100001001",
  54166=>"000110001",
  54167=>"111101001",
  54168=>"001101011",
  54169=>"101100100",
  54170=>"000100010",
  54171=>"010101000",
  54172=>"100100110",
  54173=>"011110010",
  54174=>"000000111",
  54175=>"001110110",
  54176=>"010101011",
  54177=>"111011001",
  54178=>"111101101",
  54179=>"100000000",
  54180=>"011101001",
  54181=>"110110110",
  54182=>"010100011",
  54183=>"011100101",
  54184=>"001100000",
  54185=>"000001100",
  54186=>"001101100",
  54187=>"010100101",
  54188=>"011110111",
  54189=>"001100100",
  54190=>"000100101",
  54191=>"001100011",
  54192=>"001010100",
  54193=>"010101110",
  54194=>"000101101",
  54195=>"010100100",
  54196=>"000000011",
  54197=>"010011110",
  54198=>"001000000",
  54199=>"111001001",
  54200=>"111010100",
  54201=>"001000101",
  54202=>"111011111",
  54203=>"001001001",
  54204=>"101000111",
  54205=>"011101011",
  54206=>"001010000",
  54207=>"101000100",
  54208=>"111001010",
  54209=>"001110110",
  54210=>"000101011",
  54211=>"100100100",
  54212=>"001010000",
  54213=>"110100000",
  54214=>"000001001",
  54215=>"011100111",
  54216=>"100111011",
  54217=>"101100010",
  54218=>"101000001",
  54219=>"110000000",
  54220=>"101111110",
  54221=>"000110011",
  54222=>"111000011",
  54223=>"101110111",
  54224=>"100101110",
  54225=>"111101000",
  54226=>"010010011",
  54227=>"100001100",
  54228=>"101001010",
  54229=>"001011010",
  54230=>"010000011",
  54231=>"000000000",
  54232=>"111011101",
  54233=>"000100111",
  54234=>"011010010",
  54235=>"000101101",
  54236=>"011100000",
  54237=>"000011111",
  54238=>"011111111",
  54239=>"111101000",
  54240=>"100011000",
  54241=>"111100010",
  54242=>"111101111",
  54243=>"001111010",
  54244=>"101001111",
  54245=>"010110011",
  54246=>"110000010",
  54247=>"110010110",
  54248=>"101111110",
  54249=>"111001110",
  54250=>"011001101",
  54251=>"100010001",
  54252=>"111011010",
  54253=>"000000010",
  54254=>"101101100",
  54255=>"111111010",
  54256=>"001000011",
  54257=>"010111101",
  54258=>"110111100",
  54259=>"011010000",
  54260=>"001011010",
  54261=>"100110111",
  54262=>"001001011",
  54263=>"011100101",
  54264=>"010111001",
  54265=>"011111101",
  54266=>"001010001",
  54267=>"011011110",
  54268=>"011000110",
  54269=>"010001100",
  54270=>"010110110",
  54271=>"011111001",
  54272=>"111000110",
  54273=>"001000110",
  54274=>"001010100",
  54275=>"110000101",
  54276=>"000001000",
  54277=>"100101101",
  54278=>"101000110",
  54279=>"011011010",
  54280=>"000011001",
  54281=>"101001101",
  54282=>"100101101",
  54283=>"010011100",
  54284=>"011111000",
  54285=>"000111111",
  54286=>"010101001",
  54287=>"110010110",
  54288=>"111111110",
  54289=>"010100010",
  54290=>"101100100",
  54291=>"101111110",
  54292=>"000000101",
  54293=>"100001000",
  54294=>"101100110",
  54295=>"010001101",
  54296=>"100000000",
  54297=>"111101101",
  54298=>"111111011",
  54299=>"110100100",
  54300=>"110111000",
  54301=>"111110010",
  54302=>"010101111",
  54303=>"110101001",
  54304=>"000111011",
  54305=>"000100101",
  54306=>"011110011",
  54307=>"101111001",
  54308=>"100110101",
  54309=>"011101101",
  54310=>"100010111",
  54311=>"001100000",
  54312=>"000000100",
  54313=>"000000000",
  54314=>"110110111",
  54315=>"010001000",
  54316=>"100011100",
  54317=>"110101001",
  54318=>"001101100",
  54319=>"011011011",
  54320=>"010101100",
  54321=>"110111011",
  54322=>"001011110",
  54323=>"000100110",
  54324=>"011000111",
  54325=>"000101100",
  54326=>"001101110",
  54327=>"000010100",
  54328=>"010110011",
  54329=>"100101101",
  54330=>"000001111",
  54331=>"101110000",
  54332=>"011101100",
  54333=>"000111101",
  54334=>"111010111",
  54335=>"000111011",
  54336=>"110111000",
  54337=>"100110000",
  54338=>"001000001",
  54339=>"011110011",
  54340=>"110111001",
  54341=>"111111100",
  54342=>"101111011",
  54343=>"111100100",
  54344=>"111000100",
  54345=>"110011010",
  54346=>"011001111",
  54347=>"001011101",
  54348=>"111010010",
  54349=>"001001011",
  54350=>"101110110",
  54351=>"010100111",
  54352=>"100001110",
  54353=>"000010001",
  54354=>"001001010",
  54355=>"001000000",
  54356=>"001000010",
  54357=>"000000011",
  54358=>"111101100",
  54359=>"110011011",
  54360=>"011000111",
  54361=>"110100011",
  54362=>"011001100",
  54363=>"000000100",
  54364=>"111100100",
  54365=>"001100011",
  54366=>"000010100",
  54367=>"000100011",
  54368=>"101010111",
  54369=>"011110110",
  54370=>"000000010",
  54371=>"000011001",
  54372=>"101001011",
  54373=>"010010111",
  54374=>"101001011",
  54375=>"011101000",
  54376=>"000111110",
  54377=>"001001100",
  54378=>"100000111",
  54379=>"101000001",
  54380=>"110001100",
  54381=>"101001110",
  54382=>"010010011",
  54383=>"010100011",
  54384=>"100000101",
  54385=>"110110011",
  54386=>"010110111",
  54387=>"011010011",
  54388=>"110110011",
  54389=>"111001111",
  54390=>"111010000",
  54391=>"111011010",
  54392=>"000011101",
  54393=>"011110010",
  54394=>"100111101",
  54395=>"100100111",
  54396=>"000001101",
  54397=>"000010110",
  54398=>"000001000",
  54399=>"100111111",
  54400=>"111010000",
  54401=>"011001101",
  54402=>"111000001",
  54403=>"011001100",
  54404=>"000101111",
  54405=>"000001100",
  54406=>"110101000",
  54407=>"111011011",
  54408=>"100011101",
  54409=>"000100101",
  54410=>"111110100",
  54411=>"010001000",
  54412=>"110100110",
  54413=>"011110001",
  54414=>"101100011",
  54415=>"101001101",
  54416=>"111001000",
  54417=>"101001100",
  54418=>"001000011",
  54419=>"001101101",
  54420=>"110100001",
  54421=>"000010101",
  54422=>"010110111",
  54423=>"011111100",
  54424=>"111110110",
  54425=>"111010001",
  54426=>"011100110",
  54427=>"111100000",
  54428=>"101101011",
  54429=>"010010110",
  54430=>"101111011",
  54431=>"111000111",
  54432=>"010101100",
  54433=>"100011101",
  54434=>"000100110",
  54435=>"000100001",
  54436=>"011110111",
  54437=>"111000011",
  54438=>"010111110",
  54439=>"010110000",
  54440=>"101111101",
  54441=>"001000000",
  54442=>"011001100",
  54443=>"101110111",
  54444=>"110000001",
  54445=>"101111111",
  54446=>"000101101",
  54447=>"100001011",
  54448=>"110000001",
  54449=>"000000100",
  54450=>"001011000",
  54451=>"000010110",
  54452=>"111001101",
  54453=>"011101000",
  54454=>"001010010",
  54455=>"000110000",
  54456=>"101101010",
  54457=>"001101010",
  54458=>"111000101",
  54459=>"010100101",
  54460=>"110111001",
  54461=>"110000111",
  54462=>"111111010",
  54463=>"000011100",
  54464=>"001000101",
  54465=>"000101100",
  54466=>"100101100",
  54467=>"111111001",
  54468=>"110010001",
  54469=>"101010101",
  54470=>"000111011",
  54471=>"101101011",
  54472=>"100000010",
  54473=>"111111000",
  54474=>"010111111",
  54475=>"110000011",
  54476=>"110101000",
  54477=>"100011010",
  54478=>"111101101",
  54479=>"011100110",
  54480=>"000110000",
  54481=>"001110111",
  54482=>"110010100",
  54483=>"001001001",
  54484=>"001110000",
  54485=>"111010001",
  54486=>"000000111",
  54487=>"100100101",
  54488=>"110110011",
  54489=>"100100001",
  54490=>"000011001",
  54491=>"100111100",
  54492=>"100110100",
  54493=>"011011101",
  54494=>"011101101",
  54495=>"110010110",
  54496=>"001110100",
  54497=>"000000000",
  54498=>"011011100",
  54499=>"101010000",
  54500=>"010011100",
  54501=>"100010101",
  54502=>"001101101",
  54503=>"101100111",
  54504=>"000101110",
  54505=>"101111111",
  54506=>"110000111",
  54507=>"110101111",
  54508=>"010010010",
  54509=>"100100100",
  54510=>"100001111",
  54511=>"011100110",
  54512=>"011100000",
  54513=>"010111101",
  54514=>"111010011",
  54515=>"000011010",
  54516=>"010011111",
  54517=>"001001111",
  54518=>"000001101",
  54519=>"011111011",
  54520=>"000011010",
  54521=>"001100000",
  54522=>"011010110",
  54523=>"001010100",
  54524=>"100101000",
  54525=>"001010011",
  54526=>"100011111",
  54527=>"011000100",
  54528=>"010011000",
  54529=>"011010111",
  54530=>"110111000",
  54531=>"010100110",
  54532=>"010100001",
  54533=>"000001010",
  54534=>"111101000",
  54535=>"011000101",
  54536=>"110100100",
  54537=>"000000000",
  54538=>"110000111",
  54539=>"001001010",
  54540=>"001011000",
  54541=>"000000100",
  54542=>"001100101",
  54543=>"000101001",
  54544=>"100100010",
  54545=>"101111111",
  54546=>"000111001",
  54547=>"111000010",
  54548=>"101000001",
  54549=>"000011111",
  54550=>"011000000",
  54551=>"011110101",
  54552=>"110101010",
  54553=>"101001111",
  54554=>"100110100",
  54555=>"111001100",
  54556=>"000101000",
  54557=>"011110011",
  54558=>"001100111",
  54559=>"101110010",
  54560=>"100000001",
  54561=>"011110110",
  54562=>"010000100",
  54563=>"011001110",
  54564=>"110111001",
  54565=>"010101100",
  54566=>"100101110",
  54567=>"111100010",
  54568=>"111010111",
  54569=>"110101010",
  54570=>"111010101",
  54571=>"001001111",
  54572=>"000101001",
  54573=>"101100101",
  54574=>"000000001",
  54575=>"100101100",
  54576=>"100100000",
  54577=>"101101111",
  54578=>"110010101",
  54579=>"100111111",
  54580=>"001101010",
  54581=>"010000111",
  54582=>"100000110",
  54583=>"010010011",
  54584=>"111011111",
  54585=>"000011111",
  54586=>"101001011",
  54587=>"110010100",
  54588=>"001111011",
  54589=>"111101101",
  54590=>"110100110",
  54591=>"010011011",
  54592=>"010100111",
  54593=>"100111010",
  54594=>"111110001",
  54595=>"101000101",
  54596=>"011001001",
  54597=>"101110011",
  54598=>"110000011",
  54599=>"000011111",
  54600=>"110110000",
  54601=>"010010011",
  54602=>"100000011",
  54603=>"011011000",
  54604=>"011010001",
  54605=>"011001111",
  54606=>"110010011",
  54607=>"000111001",
  54608=>"100000011",
  54609=>"101111010",
  54610=>"011001110",
  54611=>"010011000",
  54612=>"111000101",
  54613=>"000010010",
  54614=>"100010011",
  54615=>"000100011",
  54616=>"011000111",
  54617=>"010111111",
  54618=>"110001111",
  54619=>"001110101",
  54620=>"100100001",
  54621=>"110010100",
  54622=>"101101011",
  54623=>"101001110",
  54624=>"100111111",
  54625=>"111101101",
  54626=>"101100101",
  54627=>"101101101",
  54628=>"101011111",
  54629=>"000100000",
  54630=>"101000010",
  54631=>"111101111",
  54632=>"000111100",
  54633=>"111110000",
  54634=>"101101110",
  54635=>"001000111",
  54636=>"011011110",
  54637=>"001001000",
  54638=>"110000101",
  54639=>"110011001",
  54640=>"100101111",
  54641=>"110010110",
  54642=>"111000100",
  54643=>"010010010",
  54644=>"111001110",
  54645=>"111110101",
  54646=>"010111110",
  54647=>"000001100",
  54648=>"011011000",
  54649=>"101000011",
  54650=>"101110010",
  54651=>"011011100",
  54652=>"010100101",
  54653=>"010100100",
  54654=>"100000011",
  54655=>"111011101",
  54656=>"100001111",
  54657=>"000001010",
  54658=>"001110101",
  54659=>"011110000",
  54660=>"100110011",
  54661=>"101111000",
  54662=>"110000011",
  54663=>"000100111",
  54664=>"101111110",
  54665=>"100000110",
  54666=>"000010000",
  54667=>"110111110",
  54668=>"001001110",
  54669=>"110111111",
  54670=>"001111111",
  54671=>"011011110",
  54672=>"111000011",
  54673=>"111111000",
  54674=>"010011000",
  54675=>"001001001",
  54676=>"001000100",
  54677=>"100000110",
  54678=>"110111001",
  54679=>"101110011",
  54680=>"000110000",
  54681=>"011001001",
  54682=>"111000011",
  54683=>"110010100",
  54684=>"000000100",
  54685=>"000010000",
  54686=>"010110001",
  54687=>"001100011",
  54688=>"100110010",
  54689=>"011100010",
  54690=>"000001011",
  54691=>"001110011",
  54692=>"000001101",
  54693=>"001001111",
  54694=>"011110011",
  54695=>"011101100",
  54696=>"000000111",
  54697=>"111101001",
  54698=>"100001000",
  54699=>"001101000",
  54700=>"000111001",
  54701=>"010101110",
  54702=>"101100111",
  54703=>"010111111",
  54704=>"100110001",
  54705=>"100010011",
  54706=>"000110011",
  54707=>"000001100",
  54708=>"100000001",
  54709=>"101111100",
  54710=>"111000000",
  54711=>"100111001",
  54712=>"010000111",
  54713=>"110100101",
  54714=>"100100000",
  54715=>"110111110",
  54716=>"111100100",
  54717=>"010100001",
  54718=>"101100111",
  54719=>"101100101",
  54720=>"101011001",
  54721=>"111100110",
  54722=>"110101000",
  54723=>"110011000",
  54724=>"100000110",
  54725=>"100001000",
  54726=>"010001111",
  54727=>"101110101",
  54728=>"111011011",
  54729=>"101101001",
  54730=>"110101011",
  54731=>"101011100",
  54732=>"100101001",
  54733=>"000100111",
  54734=>"000000000",
  54735=>"100001111",
  54736=>"001000001",
  54737=>"100011111",
  54738=>"110001111",
  54739=>"001011010",
  54740=>"000111000",
  54741=>"010001001",
  54742=>"000001101",
  54743=>"110111110",
  54744=>"001101100",
  54745=>"111011100",
  54746=>"011111000",
  54747=>"110011111",
  54748=>"110010100",
  54749=>"110001001",
  54750=>"110000111",
  54751=>"111111101",
  54752=>"011011010",
  54753=>"010101100",
  54754=>"011111111",
  54755=>"101001011",
  54756=>"110110001",
  54757=>"000001000",
  54758=>"010111100",
  54759=>"100001101",
  54760=>"100001010",
  54761=>"010110011",
  54762=>"010000010",
  54763=>"100001100",
  54764=>"000010110",
  54765=>"011111101",
  54766=>"110101001",
  54767=>"110100111",
  54768=>"110111110",
  54769=>"111001100",
  54770=>"000000101",
  54771=>"010010010",
  54772=>"110001010",
  54773=>"101011010",
  54774=>"100010100",
  54775=>"111001110",
  54776=>"110111110",
  54777=>"111100000",
  54778=>"010010001",
  54779=>"110010000",
  54780=>"110001101",
  54781=>"000011011",
  54782=>"000000100",
  54783=>"010111110",
  54784=>"111011010",
  54785=>"000111011",
  54786=>"000011101",
  54787=>"100011101",
  54788=>"011101100",
  54789=>"000011001",
  54790=>"100000101",
  54791=>"100010100",
  54792=>"000111001",
  54793=>"100101111",
  54794=>"100101111",
  54795=>"100011001",
  54796=>"001001001",
  54797=>"111111100",
  54798=>"000000000",
  54799=>"101010111",
  54800=>"001000101",
  54801=>"110100100",
  54802=>"110000101",
  54803=>"101010100",
  54804=>"011010001",
  54805=>"100000011",
  54806=>"110000001",
  54807=>"001111010",
  54808=>"011000000",
  54809=>"110001011",
  54810=>"100001010",
  54811=>"101010111",
  54812=>"110001111",
  54813=>"000000011",
  54814=>"001001100",
  54815=>"100001000",
  54816=>"000000111",
  54817=>"011111111",
  54818=>"000011011",
  54819=>"000111000",
  54820=>"000101000",
  54821=>"010101000",
  54822=>"101110101",
  54823=>"100100001",
  54824=>"110110010",
  54825=>"101011100",
  54826=>"001110111",
  54827=>"010101001",
  54828=>"001001101",
  54829=>"100000100",
  54830=>"101000101",
  54831=>"001000000",
  54832=>"001001110",
  54833=>"000000011",
  54834=>"001101100",
  54835=>"011110010",
  54836=>"001011100",
  54837=>"011111000",
  54838=>"100001100",
  54839=>"000011100",
  54840=>"110110101",
  54841=>"010100101",
  54842=>"101000110",
  54843=>"010110000",
  54844=>"001110110",
  54845=>"000001000",
  54846=>"010100011",
  54847=>"110111110",
  54848=>"001011001",
  54849=>"101111111",
  54850=>"110110110",
  54851=>"001100010",
  54852=>"101011011",
  54853=>"110000101",
  54854=>"100000011",
  54855=>"101011101",
  54856=>"001000001",
  54857=>"001011010",
  54858=>"110110110",
  54859=>"010001101",
  54860=>"011101101",
  54861=>"111000000",
  54862=>"010101000",
  54863=>"001000000",
  54864=>"000100000",
  54865=>"110101101",
  54866=>"100110001",
  54867=>"000100001",
  54868=>"100000001",
  54869=>"000010010",
  54870=>"010100011",
  54871=>"100110000",
  54872=>"001011001",
  54873=>"111110111",
  54874=>"001111111",
  54875=>"111001011",
  54876=>"101010100",
  54877=>"100000110",
  54878=>"011111100",
  54879=>"000010111",
  54880=>"010100111",
  54881=>"111000101",
  54882=>"110101111",
  54883=>"010101010",
  54884=>"010111011",
  54885=>"101101110",
  54886=>"011110110",
  54887=>"111111011",
  54888=>"110001011",
  54889=>"001010001",
  54890=>"111101111",
  54891=>"000111000",
  54892=>"010111011",
  54893=>"110101001",
  54894=>"111101101",
  54895=>"110011000",
  54896=>"111010001",
  54897=>"011011100",
  54898=>"110001011",
  54899=>"001101000",
  54900=>"111001001",
  54901=>"110011010",
  54902=>"001001110",
  54903=>"111001001",
  54904=>"001101101",
  54905=>"010110010",
  54906=>"101101101",
  54907=>"010111110",
  54908=>"101011100",
  54909=>"001100000",
  54910=>"001010111",
  54911=>"010100010",
  54912=>"100111100",
  54913=>"100101110",
  54914=>"000101110",
  54915=>"011100010",
  54916=>"011001100",
  54917=>"011101000",
  54918=>"111101110",
  54919=>"011001000",
  54920=>"110000101",
  54921=>"001001001",
  54922=>"010110110",
  54923=>"111011110",
  54924=>"011101010",
  54925=>"011110111",
  54926=>"101001101",
  54927=>"111110011",
  54928=>"001110111",
  54929=>"000011001",
  54930=>"100111001",
  54931=>"111100011",
  54932=>"000011110",
  54933=>"011000000",
  54934=>"111011101",
  54935=>"100111110",
  54936=>"001110011",
  54937=>"111101110",
  54938=>"010111100",
  54939=>"100011001",
  54940=>"010100101",
  54941=>"010010111",
  54942=>"010101010",
  54943=>"111100001",
  54944=>"001000010",
  54945=>"110111010",
  54946=>"110110010",
  54947=>"111011110",
  54948=>"001101110",
  54949=>"100111100",
  54950=>"110001001",
  54951=>"000001000",
  54952=>"001000101",
  54953=>"111101111",
  54954=>"000101110",
  54955=>"110100101",
  54956=>"111000110",
  54957=>"101001110",
  54958=>"101001000",
  54959=>"010100001",
  54960=>"110101101",
  54961=>"111010111",
  54962=>"101001100",
  54963=>"100000100",
  54964=>"110011111",
  54965=>"011101100",
  54966=>"010111100",
  54967=>"010110110",
  54968=>"111001011",
  54969=>"111000110",
  54970=>"010110100",
  54971=>"010000010",
  54972=>"110111011",
  54973=>"000100100",
  54974=>"100010110",
  54975=>"100111110",
  54976=>"010100000",
  54977=>"110011110",
  54978=>"110000000",
  54979=>"100010001",
  54980=>"011010110",
  54981=>"100111010",
  54982=>"010010010",
  54983=>"010001110",
  54984=>"011001001",
  54985=>"000000100",
  54986=>"101110011",
  54987=>"010111110",
  54988=>"000001101",
  54989=>"010010111",
  54990=>"101000111",
  54991=>"000011001",
  54992=>"010110100",
  54993=>"101111011",
  54994=>"001010111",
  54995=>"001011001",
  54996=>"101111000",
  54997=>"010011011",
  54998=>"001010001",
  54999=>"110100000",
  55000=>"011110000",
  55001=>"000001001",
  55002=>"100100111",
  55003=>"001100000",
  55004=>"100101000",
  55005=>"111000011",
  55006=>"111001110",
  55007=>"100011110",
  55008=>"001100111",
  55009=>"110000000",
  55010=>"100000100",
  55011=>"010100000",
  55012=>"001011110",
  55013=>"001101101",
  55014=>"011111101",
  55015=>"001111000",
  55016=>"010001000",
  55017=>"101110110",
  55018=>"100111101",
  55019=>"011111001",
  55020=>"100001000",
  55021=>"111111011",
  55022=>"110000111",
  55023=>"111111111",
  55024=>"000100000",
  55025=>"001111001",
  55026=>"000000011",
  55027=>"000011110",
  55028=>"110100100",
  55029=>"100110001",
  55030=>"011000111",
  55031=>"010010110",
  55032=>"000010001",
  55033=>"111101001",
  55034=>"100010101",
  55035=>"010001100",
  55036=>"110111000",
  55037=>"011001000",
  55038=>"010000000",
  55039=>"000111010",
  55040=>"000010011",
  55041=>"100111011",
  55042=>"110111001",
  55043=>"111101010",
  55044=>"110011100",
  55045=>"000001011",
  55046=>"101110110",
  55047=>"000100111",
  55048=>"100011101",
  55049=>"001100000",
  55050=>"111000010",
  55051=>"001000001",
  55052=>"010000001",
  55053=>"111111111",
  55054=>"101110100",
  55055=>"111101110",
  55056=>"010100111",
  55057=>"011010100",
  55058=>"100110000",
  55059=>"001011111",
  55060=>"100110011",
  55061=>"100100010",
  55062=>"111110111",
  55063=>"010100001",
  55064=>"001001111",
  55065=>"110101000",
  55066=>"111010001",
  55067=>"001010001",
  55068=>"111000101",
  55069=>"111000101",
  55070=>"100101011",
  55071=>"001000000",
  55072=>"111010110",
  55073=>"001100010",
  55074=>"110101000",
  55075=>"100010111",
  55076=>"111000100",
  55077=>"000001000",
  55078=>"000011010",
  55079=>"111100001",
  55080=>"010001010",
  55081=>"110101110",
  55082=>"100011001",
  55083=>"100001110",
  55084=>"001111100",
  55085=>"000000010",
  55086=>"100111110",
  55087=>"111111110",
  55088=>"001010110",
  55089=>"110110101",
  55090=>"010000000",
  55091=>"101011011",
  55092=>"000110111",
  55093=>"101111000",
  55094=>"000001110",
  55095=>"111100100",
  55096=>"010111000",
  55097=>"001010101",
  55098=>"101111111",
  55099=>"011111101",
  55100=>"100001001",
  55101=>"100100000",
  55102=>"101100101",
  55103=>"110110000",
  55104=>"001001000",
  55105=>"001001110",
  55106=>"100100100",
  55107=>"100011011",
  55108=>"010101101",
  55109=>"101011111",
  55110=>"000111110",
  55111=>"011001010",
  55112=>"110000101",
  55113=>"010000000",
  55114=>"111100110",
  55115=>"100011000",
  55116=>"100111110",
  55117=>"000110011",
  55118=>"110000110",
  55119=>"000111100",
  55120=>"100110001",
  55121=>"000100011",
  55122=>"000111110",
  55123=>"100000001",
  55124=>"100010111",
  55125=>"111001111",
  55126=>"011000001",
  55127=>"111100111",
  55128=>"111110000",
  55129=>"111011001",
  55130=>"111010101",
  55131=>"101111010",
  55132=>"100001011",
  55133=>"001010100",
  55134=>"010011011",
  55135=>"000010000",
  55136=>"101101001",
  55137=>"101011110",
  55138=>"110000010",
  55139=>"011001011",
  55140=>"000100011",
  55141=>"100011111",
  55142=>"101010101",
  55143=>"101000010",
  55144=>"101001000",
  55145=>"001000001",
  55146=>"101011110",
  55147=>"001000000",
  55148=>"000101111",
  55149=>"101110010",
  55150=>"111010000",
  55151=>"011111110",
  55152=>"000110111",
  55153=>"111010110",
  55154=>"100000101",
  55155=>"111111110",
  55156=>"100111001",
  55157=>"111111110",
  55158=>"000001001",
  55159=>"111111000",
  55160=>"110100000",
  55161=>"010001010",
  55162=>"010000101",
  55163=>"110110000",
  55164=>"111010010",
  55165=>"000000000",
  55166=>"101110001",
  55167=>"010011011",
  55168=>"010101011",
  55169=>"100101000",
  55170=>"101101100",
  55171=>"100010010",
  55172=>"100110001",
  55173=>"111000000",
  55174=>"001110000",
  55175=>"000100011",
  55176=>"111010001",
  55177=>"001110000",
  55178=>"110011010",
  55179=>"111000110",
  55180=>"010111110",
  55181=>"001000000",
  55182=>"100110000",
  55183=>"100100000",
  55184=>"100001111",
  55185=>"011000110",
  55186=>"010010010",
  55187=>"011001011",
  55188=>"010111110",
  55189=>"001011110",
  55190=>"001111100",
  55191=>"010011011",
  55192=>"011011001",
  55193=>"100000001",
  55194=>"110000110",
  55195=>"001000110",
  55196=>"110010111",
  55197=>"111111011",
  55198=>"111101100",
  55199=>"011011110",
  55200=>"010110101",
  55201=>"001010010",
  55202=>"101101010",
  55203=>"011111011",
  55204=>"000000000",
  55205=>"011100100",
  55206=>"010011111",
  55207=>"010011001",
  55208=>"101110111",
  55209=>"101111111",
  55210=>"101000010",
  55211=>"100000000",
  55212=>"000011100",
  55213=>"011101001",
  55214=>"111000000",
  55215=>"101110001",
  55216=>"001111000",
  55217=>"101100001",
  55218=>"010001001",
  55219=>"011001010",
  55220=>"110001100",
  55221=>"011010001",
  55222=>"100010010",
  55223=>"001010101",
  55224=>"100101111",
  55225=>"101111010",
  55226=>"000100000",
  55227=>"100000101",
  55228=>"011111000",
  55229=>"100010000",
  55230=>"111101000",
  55231=>"111000111",
  55232=>"000101000",
  55233=>"111001000",
  55234=>"001111001",
  55235=>"011001101",
  55236=>"000000101",
  55237=>"111110001",
  55238=>"101110001",
  55239=>"010111111",
  55240=>"010011000",
  55241=>"000100100",
  55242=>"000001000",
  55243=>"110000111",
  55244=>"111110010",
  55245=>"110101100",
  55246=>"100000110",
  55247=>"101001011",
  55248=>"000100010",
  55249=>"101000010",
  55250=>"100111111",
  55251=>"011000010",
  55252=>"000000101",
  55253=>"110010000",
  55254=>"100110010",
  55255=>"100100010",
  55256=>"111001011",
  55257=>"000111111",
  55258=>"000011010",
  55259=>"011100011",
  55260=>"011001001",
  55261=>"000001010",
  55262=>"010011000",
  55263=>"110010111",
  55264=>"100010011",
  55265=>"000000011",
  55266=>"010001110",
  55267=>"111001000",
  55268=>"000100001",
  55269=>"111110101",
  55270=>"001011001",
  55271=>"010110111",
  55272=>"011110000",
  55273=>"011001001",
  55274=>"011111000",
  55275=>"111110000",
  55276=>"001100101",
  55277=>"110011111",
  55278=>"011101000",
  55279=>"000010011",
  55280=>"110110110",
  55281=>"100000100",
  55282=>"110111111",
  55283=>"010000101",
  55284=>"011010001",
  55285=>"101110111",
  55286=>"001100011",
  55287=>"010000001",
  55288=>"010111101",
  55289=>"111001100",
  55290=>"000010000",
  55291=>"000000001",
  55292=>"101001110",
  55293=>"110101000",
  55294=>"011011011",
  55295=>"101010010",
  55296=>"010011001",
  55297=>"110011111",
  55298=>"000101101",
  55299=>"001111110",
  55300=>"101100000",
  55301=>"101100000",
  55302=>"011110100",
  55303=>"010101001",
  55304=>"101100000",
  55305=>"110010111",
  55306=>"010111000",
  55307=>"010000110",
  55308=>"101011001",
  55309=>"000100011",
  55310=>"110100000",
  55311=>"001101011",
  55312=>"001111000",
  55313=>"010000101",
  55314=>"111110111",
  55315=>"100000000",
  55316=>"001010010",
  55317=>"011100100",
  55318=>"110111111",
  55319=>"001000001",
  55320=>"011110111",
  55321=>"100100011",
  55322=>"110000011",
  55323=>"011001010",
  55324=>"000010011",
  55325=>"010100010",
  55326=>"110000010",
  55327=>"111000001",
  55328=>"110000101",
  55329=>"100000010",
  55330=>"111110111",
  55331=>"110010100",
  55332=>"110011101",
  55333=>"110000010",
  55334=>"101011101",
  55335=>"111111110",
  55336=>"100000100",
  55337=>"001010001",
  55338=>"010100111",
  55339=>"011000110",
  55340=>"100000101",
  55341=>"001010001",
  55342=>"001110111",
  55343=>"110011010",
  55344=>"110011010",
  55345=>"111000011",
  55346=>"011101000",
  55347=>"111001010",
  55348=>"000100010",
  55349=>"010001010",
  55350=>"101001000",
  55351=>"110010010",
  55352=>"110101101",
  55353=>"101100100",
  55354=>"010000010",
  55355=>"101011010",
  55356=>"000111111",
  55357=>"100110001",
  55358=>"100100000",
  55359=>"100011011",
  55360=>"101101000",
  55361=>"001100010",
  55362=>"101100001",
  55363=>"011011101",
  55364=>"111011111",
  55365=>"110011100",
  55366=>"111100001",
  55367=>"000011011",
  55368=>"111001000",
  55369=>"100000110",
  55370=>"100110000",
  55371=>"100001000",
  55372=>"101100000",
  55373=>"001000111",
  55374=>"001010000",
  55375=>"011110011",
  55376=>"110000011",
  55377=>"000011100",
  55378=>"011001010",
  55379=>"011011000",
  55380=>"111011100",
  55381=>"111001011",
  55382=>"110010100",
  55383=>"110101001",
  55384=>"011001101",
  55385=>"100101001",
  55386=>"010011111",
  55387=>"000011000",
  55388=>"000011001",
  55389=>"001001011",
  55390=>"100000100",
  55391=>"110010000",
  55392=>"010111100",
  55393=>"111000001",
  55394=>"100101001",
  55395=>"011110010",
  55396=>"110100101",
  55397=>"001011011",
  55398=>"001011011",
  55399=>"111100001",
  55400=>"111010100",
  55401=>"000000010",
  55402=>"100111010",
  55403=>"101111110",
  55404=>"011001100",
  55405=>"010000100",
  55406=>"101010111",
  55407=>"111111111",
  55408=>"000100111",
  55409=>"001010000",
  55410=>"010001011",
  55411=>"100110110",
  55412=>"000110100",
  55413=>"000000011",
  55414=>"111010000",
  55415=>"000100001",
  55416=>"011110001",
  55417=>"110010111",
  55418=>"100111110",
  55419=>"111100111",
  55420=>"100011101",
  55421=>"110111010",
  55422=>"001000011",
  55423=>"111101101",
  55424=>"001111011",
  55425=>"100101101",
  55426=>"001010100",
  55427=>"101001001",
  55428=>"100110011",
  55429=>"110100001",
  55430=>"100111101",
  55431=>"001000101",
  55432=>"001100111",
  55433=>"110100110",
  55434=>"011011000",
  55435=>"010010111",
  55436=>"011100100",
  55437=>"010101001",
  55438=>"111011100",
  55439=>"010101001",
  55440=>"111101010",
  55441=>"001100100",
  55442=>"010100110",
  55443=>"001011011",
  55444=>"101010100",
  55445=>"010000000",
  55446=>"110000100",
  55447=>"110000011",
  55448=>"011111100",
  55449=>"010000101",
  55450=>"100011100",
  55451=>"010001010",
  55452=>"011010100",
  55453=>"000001110",
  55454=>"111101101",
  55455=>"010100111",
  55456=>"001100001",
  55457=>"011100101",
  55458=>"000011100",
  55459=>"001001011",
  55460=>"001001100",
  55461=>"011101000",
  55462=>"011000110",
  55463=>"010100101",
  55464=>"011000111",
  55465=>"101101000",
  55466=>"111101101",
  55467=>"010100010",
  55468=>"110000110",
  55469=>"111000001",
  55470=>"001101100",
  55471=>"011000000",
  55472=>"000111011",
  55473=>"101001000",
  55474=>"101000111",
  55475=>"111001001",
  55476=>"000101100",
  55477=>"100101001",
  55478=>"100000000",
  55479=>"011110000",
  55480=>"110001000",
  55481=>"110100111",
  55482=>"001000000",
  55483=>"001100101",
  55484=>"111110001",
  55485=>"000101110",
  55486=>"010001110",
  55487=>"011001001",
  55488=>"100010100",
  55489=>"001001101",
  55490=>"111100101",
  55491=>"011011010",
  55492=>"111111111",
  55493=>"110000000",
  55494=>"100000000",
  55495=>"000000000",
  55496=>"000011110",
  55497=>"111101111",
  55498=>"010001010",
  55499=>"100100011",
  55500=>"100011100",
  55501=>"101101111",
  55502=>"110011011",
  55503=>"110111000",
  55504=>"001010000",
  55505=>"001001100",
  55506=>"010000101",
  55507=>"100000011",
  55508=>"000000001",
  55509=>"000101101",
  55510=>"101110100",
  55511=>"110110100",
  55512=>"011011000",
  55513=>"000101101",
  55514=>"101000010",
  55515=>"010100000",
  55516=>"011000101",
  55517=>"011001111",
  55518=>"001111001",
  55519=>"111111111",
  55520=>"100011010",
  55521=>"111100001",
  55522=>"011000101",
  55523=>"011010001",
  55524=>"001101101",
  55525=>"111000011",
  55526=>"001000000",
  55527=>"000001111",
  55528=>"010001011",
  55529=>"010100010",
  55530=>"011011100",
  55531=>"000010010",
  55532=>"101100111",
  55533=>"000111011",
  55534=>"011010001",
  55535=>"000100101",
  55536=>"001101110",
  55537=>"110011001",
  55538=>"010100000",
  55539=>"110110001",
  55540=>"000010110",
  55541=>"000000100",
  55542=>"110010101",
  55543=>"010010011",
  55544=>"011001110",
  55545=>"101001010",
  55546=>"010011000",
  55547=>"100110000",
  55548=>"000111000",
  55549=>"011011001",
  55550=>"010101101",
  55551=>"110000100",
  55552=>"010001001",
  55553=>"111010101",
  55554=>"000000001",
  55555=>"001011000",
  55556=>"000101101",
  55557=>"110000000",
  55558=>"100010001",
  55559=>"010001011",
  55560=>"001000011",
  55561=>"010101000",
  55562=>"001000010",
  55563=>"111000000",
  55564=>"100110011",
  55565=>"111010001",
  55566=>"111001111",
  55567=>"011000000",
  55568=>"010111111",
  55569=>"011000001",
  55570=>"101111110",
  55571=>"011110111",
  55572=>"001001000",
  55573=>"111111100",
  55574=>"011111100",
  55575=>"101110111",
  55576=>"011101001",
  55577=>"101011011",
  55578=>"000000011",
  55579=>"000110100",
  55580=>"000001000",
  55581=>"010110001",
  55582=>"000000011",
  55583=>"010001000",
  55584=>"011010111",
  55585=>"001111010",
  55586=>"010010110",
  55587=>"000101011",
  55588=>"001111101",
  55589=>"000001111",
  55590=>"111001011",
  55591=>"011000101",
  55592=>"111011100",
  55593=>"101001010",
  55594=>"111001100",
  55595=>"010111111",
  55596=>"110110101",
  55597=>"000010001",
  55598=>"001000010",
  55599=>"000100011",
  55600=>"011001001",
  55601=>"111001001",
  55602=>"111100000",
  55603=>"000111111",
  55604=>"001100101",
  55605=>"001001101",
  55606=>"001111101",
  55607=>"110101111",
  55608=>"101010010",
  55609=>"110111001",
  55610=>"100001011",
  55611=>"101010001",
  55612=>"001100010",
  55613=>"111110110",
  55614=>"100111011",
  55615=>"111001011",
  55616=>"101010100",
  55617=>"001000001",
  55618=>"011001000",
  55619=>"000000101",
  55620=>"101101111",
  55621=>"100100111",
  55622=>"101100100",
  55623=>"011011001",
  55624=>"000000010",
  55625=>"110100101",
  55626=>"001001111",
  55627=>"001000010",
  55628=>"000101010",
  55629=>"011111100",
  55630=>"001100111",
  55631=>"100011001",
  55632=>"000010000",
  55633=>"100010011",
  55634=>"000100011",
  55635=>"100001011",
  55636=>"010010100",
  55637=>"101011110",
  55638=>"011111000",
  55639=>"011111101",
  55640=>"001010101",
  55641=>"100000000",
  55642=>"000001101",
  55643=>"100000010",
  55644=>"110111011",
  55645=>"001001101",
  55646=>"101101100",
  55647=>"100011110",
  55648=>"011111001",
  55649=>"010110000",
  55650=>"011011111",
  55651=>"101000100",
  55652=>"000100101",
  55653=>"000011001",
  55654=>"000011110",
  55655=>"110111011",
  55656=>"011011011",
  55657=>"010011001",
  55658=>"111010100",
  55659=>"011011011",
  55660=>"100101011",
  55661=>"001001001",
  55662=>"011110111",
  55663=>"011000000",
  55664=>"010100100",
  55665=>"111110110",
  55666=>"110100001",
  55667=>"111111001",
  55668=>"110001100",
  55669=>"011001100",
  55670=>"011100101",
  55671=>"100000101",
  55672=>"001100101",
  55673=>"101100000",
  55674=>"110001111",
  55675=>"100010101",
  55676=>"011101000",
  55677=>"110010100",
  55678=>"010010001",
  55679=>"100100001",
  55680=>"010000001",
  55681=>"011101100",
  55682=>"011011000",
  55683=>"110011100",
  55684=>"111101010",
  55685=>"011100000",
  55686=>"010010010",
  55687=>"011001010",
  55688=>"101101001",
  55689=>"100101010",
  55690=>"110111100",
  55691=>"100101100",
  55692=>"000001000",
  55693=>"101010000",
  55694=>"010111011",
  55695=>"101100110",
  55696=>"110101010",
  55697=>"111010000",
  55698=>"111001011",
  55699=>"010101110",
  55700=>"110000111",
  55701=>"010001101",
  55702=>"010010000",
  55703=>"001001001",
  55704=>"111010111",
  55705=>"000001111",
  55706=>"100001001",
  55707=>"111101110",
  55708=>"010101011",
  55709=>"000100000",
  55710=>"101000011",
  55711=>"101011011",
  55712=>"010111111",
  55713=>"010100010",
  55714=>"010011110",
  55715=>"001000010",
  55716=>"011101111",
  55717=>"000100011",
  55718=>"111011101",
  55719=>"001011010",
  55720=>"101110010",
  55721=>"011010110",
  55722=>"100001010",
  55723=>"011010000",
  55724=>"001010001",
  55725=>"101111001",
  55726=>"011110110",
  55727=>"100111000",
  55728=>"011101000",
  55729=>"001001010",
  55730=>"101101001",
  55731=>"100001101",
  55732=>"111100001",
  55733=>"011000100",
  55734=>"001001000",
  55735=>"000011011",
  55736=>"000001100",
  55737=>"110000010",
  55738=>"001000000",
  55739=>"110110111",
  55740=>"010001100",
  55741=>"011110111",
  55742=>"101011010",
  55743=>"110001010",
  55744=>"001000001",
  55745=>"101001101",
  55746=>"111100001",
  55747=>"000011100",
  55748=>"011001111",
  55749=>"110111011",
  55750=>"111011010",
  55751=>"110000100",
  55752=>"001000111",
  55753=>"010000011",
  55754=>"011111111",
  55755=>"110010000",
  55756=>"001011110",
  55757=>"111101110",
  55758=>"110011010",
  55759=>"111001000",
  55760=>"010110011",
  55761=>"010001010",
  55762=>"100010110",
  55763=>"100000110",
  55764=>"000101110",
  55765=>"101010011",
  55766=>"111101011",
  55767=>"101101000",
  55768=>"101100100",
  55769=>"110011000",
  55770=>"100100110",
  55771=>"111111011",
  55772=>"110000011",
  55773=>"011010100",
  55774=>"110000111",
  55775=>"001100100",
  55776=>"001100011",
  55777=>"101100100",
  55778=>"010110101",
  55779=>"111001001",
  55780=>"001001111",
  55781=>"111111110",
  55782=>"001100010",
  55783=>"110101001",
  55784=>"101110000",
  55785=>"100001100",
  55786=>"101000001",
  55787=>"010011100",
  55788=>"011111010",
  55789=>"010001010",
  55790=>"101100000",
  55791=>"101010110",
  55792=>"100111010",
  55793=>"111011101",
  55794=>"111100000",
  55795=>"011100101",
  55796=>"000001001",
  55797=>"001110000",
  55798=>"000010011",
  55799=>"001010001",
  55800=>"000111100",
  55801=>"110011101",
  55802=>"000110111",
  55803=>"011100111",
  55804=>"000100100",
  55805=>"110001100",
  55806=>"000100111",
  55807=>"110101110",
  55808=>"010110101",
  55809=>"011011010",
  55810=>"110110000",
  55811=>"101110000",
  55812=>"000110111",
  55813=>"101110010",
  55814=>"001010111",
  55815=>"001000111",
  55816=>"101100100",
  55817=>"100000111",
  55818=>"111011000",
  55819=>"011110000",
  55820=>"110110110",
  55821=>"110101100",
  55822=>"101110100",
  55823=>"110001000",
  55824=>"110011110",
  55825=>"010101111",
  55826=>"001000101",
  55827=>"111101000",
  55828=>"100001001",
  55829=>"111000000",
  55830=>"110000000",
  55831=>"111001100",
  55832=>"111010000",
  55833=>"001001000",
  55834=>"011000001",
  55835=>"001101010",
  55836=>"010111000",
  55837=>"100111000",
  55838=>"111101110",
  55839=>"101111101",
  55840=>"111110011",
  55841=>"000001001",
  55842=>"001001010",
  55843=>"111010000",
  55844=>"011101110",
  55845=>"011001010",
  55846=>"000101011",
  55847=>"110100010",
  55848=>"001010100",
  55849=>"100111101",
  55850=>"100000000",
  55851=>"101110111",
  55852=>"111000111",
  55853=>"011010000",
  55854=>"110111110",
  55855=>"101010011",
  55856=>"100010110",
  55857=>"111001110",
  55858=>"011011001",
  55859=>"100000001",
  55860=>"101110100",
  55861=>"010011000",
  55862=>"110010000",
  55863=>"001001100",
  55864=>"111010000",
  55865=>"101001111",
  55866=>"111100111",
  55867=>"001101000",
  55868=>"101100100",
  55869=>"000110110",
  55870=>"001101010",
  55871=>"101111110",
  55872=>"101001011",
  55873=>"011001010",
  55874=>"110000100",
  55875=>"110111011",
  55876=>"011001011",
  55877=>"000010011",
  55878=>"001111011",
  55879=>"100100111",
  55880=>"000101110",
  55881=>"111110100",
  55882=>"010110101",
  55883=>"101001000",
  55884=>"011011000",
  55885=>"111100001",
  55886=>"110110111",
  55887=>"101101100",
  55888=>"111101101",
  55889=>"101110111",
  55890=>"110011111",
  55891=>"100111000",
  55892=>"110011000",
  55893=>"110000001",
  55894=>"110101100",
  55895=>"111100110",
  55896=>"100000011",
  55897=>"101001111",
  55898=>"010111011",
  55899=>"111010000",
  55900=>"110000010",
  55901=>"100111110",
  55902=>"000010001",
  55903=>"000101011",
  55904=>"010111001",
  55905=>"000000000",
  55906=>"111100100",
  55907=>"001101000",
  55908=>"010110001",
  55909=>"110000010",
  55910=>"010010011",
  55911=>"100101001",
  55912=>"100000111",
  55913=>"111000001",
  55914=>"111111011",
  55915=>"001100000",
  55916=>"100010110",
  55917=>"101100011",
  55918=>"110101011",
  55919=>"010010010",
  55920=>"100000100",
  55921=>"000100000",
  55922=>"001001101",
  55923=>"001000000",
  55924=>"111011010",
  55925=>"010011001",
  55926=>"111110001",
  55927=>"000100010",
  55928=>"111100010",
  55929=>"111010001",
  55930=>"111101111",
  55931=>"010110011",
  55932=>"011101010",
  55933=>"010000000",
  55934=>"111101000",
  55935=>"001010110",
  55936=>"011001001",
  55937=>"011111110",
  55938=>"110010100",
  55939=>"111101111",
  55940=>"010000011",
  55941=>"000001101",
  55942=>"011001000",
  55943=>"111101010",
  55944=>"001101111",
  55945=>"101010001",
  55946=>"101101100",
  55947=>"111111000",
  55948=>"000101000",
  55949=>"001101100",
  55950=>"101100011",
  55951=>"000001101",
  55952=>"100001110",
  55953=>"101101101",
  55954=>"101110001",
  55955=>"010011001",
  55956=>"000010111",
  55957=>"101100110",
  55958=>"110111011",
  55959=>"100100010",
  55960=>"011010000",
  55961=>"011111111",
  55962=>"010001010",
  55963=>"101111011",
  55964=>"011111001",
  55965=>"110001101",
  55966=>"011101000",
  55967=>"000100100",
  55968=>"111010000",
  55969=>"101101101",
  55970=>"110011011",
  55971=>"000111011",
  55972=>"010110001",
  55973=>"001110010",
  55974=>"001000001",
  55975=>"001011000",
  55976=>"010010010",
  55977=>"010000001",
  55978=>"001010011",
  55979=>"111100110",
  55980=>"101010010",
  55981=>"111000001",
  55982=>"010011100",
  55983=>"011110011",
  55984=>"100110100",
  55985=>"101010010",
  55986=>"110100011",
  55987=>"011011101",
  55988=>"001110100",
  55989=>"010001110",
  55990=>"111101001",
  55991=>"011100101",
  55992=>"011000101",
  55993=>"110100100",
  55994=>"100010011",
  55995=>"011011001",
  55996=>"100011010",
  55997=>"010001011",
  55998=>"100001000",
  55999=>"011001001",
  56000=>"001010000",
  56001=>"010110111",
  56002=>"001111010",
  56003=>"000101111",
  56004=>"101001000",
  56005=>"111001110",
  56006=>"111111011",
  56007=>"000110101",
  56008=>"111111000",
  56009=>"100111101",
  56010=>"010010110",
  56011=>"110001011",
  56012=>"101011011",
  56013=>"011110100",
  56014=>"011010110",
  56015=>"010111111",
  56016=>"100101110",
  56017=>"010011001",
  56018=>"110100001",
  56019=>"101011010",
  56020=>"001111111",
  56021=>"101000100",
  56022=>"001101001",
  56023=>"010011010",
  56024=>"110010101",
  56025=>"010111111",
  56026=>"001101101",
  56027=>"110101000",
  56028=>"000011000",
  56029=>"010000000",
  56030=>"001110011",
  56031=>"101010111",
  56032=>"000001110",
  56033=>"100010001",
  56034=>"000101111",
  56035=>"101001010",
  56036=>"000001100",
  56037=>"011010111",
  56038=>"000000111",
  56039=>"101010100",
  56040=>"001000010",
  56041=>"000111111",
  56042=>"011101001",
  56043=>"010100111",
  56044=>"010010110",
  56045=>"000101100",
  56046=>"110110110",
  56047=>"101100110",
  56048=>"100110001",
  56049=>"110000011",
  56050=>"100010101",
  56051=>"000111101",
  56052=>"000010010",
  56053=>"100010110",
  56054=>"110101110",
  56055=>"011010100",
  56056=>"101011000",
  56057=>"110011101",
  56058=>"011101110",
  56059=>"001011111",
  56060=>"001101000",
  56061=>"110100110",
  56062=>"111010111",
  56063=>"111010011",
  56064=>"110000000",
  56065=>"111011000",
  56066=>"010001011",
  56067=>"010110001",
  56068=>"110001111",
  56069=>"001000011",
  56070=>"010101001",
  56071=>"011011010",
  56072=>"011010110",
  56073=>"001001101",
  56074=>"001010111",
  56075=>"101110010",
  56076=>"011010001",
  56077=>"111101100",
  56078=>"000011010",
  56079=>"100101110",
  56080=>"111010001",
  56081=>"100010000",
  56082=>"001010111",
  56083=>"000101001",
  56084=>"110111110",
  56085=>"101101111",
  56086=>"001110000",
  56087=>"010100110",
  56088=>"111100010",
  56089=>"011000001",
  56090=>"000001100",
  56091=>"000011011",
  56092=>"001011001",
  56093=>"001000011",
  56094=>"000110110",
  56095=>"010110101",
  56096=>"011110100",
  56097=>"101000111",
  56098=>"110010110",
  56099=>"111110111",
  56100=>"101010101",
  56101=>"011110111",
  56102=>"011001100",
  56103=>"101110101",
  56104=>"100001110",
  56105=>"110111111",
  56106=>"000100100",
  56107=>"110110111",
  56108=>"000000010",
  56109=>"010101010",
  56110=>"000000000",
  56111=>"000101001",
  56112=>"001001001",
  56113=>"001001110",
  56114=>"110110001",
  56115=>"010010100",
  56116=>"111101010",
  56117=>"100001101",
  56118=>"010111111",
  56119=>"010100010",
  56120=>"101000010",
  56121=>"000100111",
  56122=>"011011110",
  56123=>"111010010",
  56124=>"001100000",
  56125=>"010001001",
  56126=>"100101100",
  56127=>"011001011",
  56128=>"110101000",
  56129=>"100110111",
  56130=>"100001001",
  56131=>"100100110",
  56132=>"111010010",
  56133=>"111000001",
  56134=>"001010100",
  56135=>"000110110",
  56136=>"111100111",
  56137=>"111111010",
  56138=>"111001011",
  56139=>"111101000",
  56140=>"011100100",
  56141=>"010111010",
  56142=>"001100011",
  56143=>"001011110",
  56144=>"010001010",
  56145=>"100001001",
  56146=>"111101101",
  56147=>"100101010",
  56148=>"000110001",
  56149=>"110111001",
  56150=>"010110010",
  56151=>"010000110",
  56152=>"001110110",
  56153=>"110100100",
  56154=>"111111101",
  56155=>"101001101",
  56156=>"111110000",
  56157=>"010011001",
  56158=>"010010011",
  56159=>"011101000",
  56160=>"010100011",
  56161=>"010000001",
  56162=>"111000001",
  56163=>"010001100",
  56164=>"100111011",
  56165=>"010011000",
  56166=>"111111101",
  56167=>"110111100",
  56168=>"111011001",
  56169=>"001000010",
  56170=>"110101110",
  56171=>"110101011",
  56172=>"011110000",
  56173=>"000000110",
  56174=>"111001111",
  56175=>"000110100",
  56176=>"111100010",
  56177=>"010000010",
  56178=>"100111011",
  56179=>"101110000",
  56180=>"000111110",
  56181=>"000101110",
  56182=>"100010111",
  56183=>"001010001",
  56184=>"111110000",
  56185=>"110011011",
  56186=>"010110100",
  56187=>"010101101",
  56188=>"101011000",
  56189=>"100011001",
  56190=>"111101001",
  56191=>"001011011",
  56192=>"101001001",
  56193=>"101010000",
  56194=>"001001001",
  56195=>"001001100",
  56196=>"100001010",
  56197=>"011000011",
  56198=>"101000000",
  56199=>"000001011",
  56200=>"010110111",
  56201=>"100000001",
  56202=>"000001100",
  56203=>"011010000",
  56204=>"110011000",
  56205=>"010101110",
  56206=>"000010110",
  56207=>"001011101",
  56208=>"010111010",
  56209=>"001000110",
  56210=>"010110100",
  56211=>"000010011",
  56212=>"101101010",
  56213=>"111011011",
  56214=>"000011111",
  56215=>"111110101",
  56216=>"010011111",
  56217=>"111101011",
  56218=>"000001110",
  56219=>"001000110",
  56220=>"101001010",
  56221=>"101001011",
  56222=>"001000000",
  56223=>"110111101",
  56224=>"101101000",
  56225=>"011000111",
  56226=>"101011010",
  56227=>"100100010",
  56228=>"001001001",
  56229=>"001001111",
  56230=>"010111101",
  56231=>"111111000",
  56232=>"101110110",
  56233=>"001110000",
  56234=>"111010100",
  56235=>"100101010",
  56236=>"100111100",
  56237=>"001101010",
  56238=>"100001111",
  56239=>"010101100",
  56240=>"111100111",
  56241=>"000011111",
  56242=>"001010111",
  56243=>"001110011",
  56244=>"111111111",
  56245=>"011100101",
  56246=>"100011011",
  56247=>"100000001",
  56248=>"101101001",
  56249=>"100000111",
  56250=>"000000101",
  56251=>"100100101",
  56252=>"010110000",
  56253=>"011100000",
  56254=>"101000010",
  56255=>"000001001",
  56256=>"011011011",
  56257=>"000000100",
  56258=>"100011110",
  56259=>"001000010",
  56260=>"111100010",
  56261=>"000101011",
  56262=>"111001000",
  56263=>"001001010",
  56264=>"010001000",
  56265=>"100001111",
  56266=>"010100111",
  56267=>"001001111",
  56268=>"110011000",
  56269=>"001111100",
  56270=>"010000111",
  56271=>"001001010",
  56272=>"001001010",
  56273=>"011000111",
  56274=>"010111011",
  56275=>"001101011",
  56276=>"011011000",
  56277=>"011111111",
  56278=>"001000000",
  56279=>"100010001",
  56280=>"100100001",
  56281=>"001011110",
  56282=>"110111101",
  56283=>"000001100",
  56284=>"111101000",
  56285=>"000000101",
  56286=>"110001100",
  56287=>"010110011",
  56288=>"001000110",
  56289=>"100100101",
  56290=>"001101001",
  56291=>"010110100",
  56292=>"100101001",
  56293=>"010100111",
  56294=>"100001001",
  56295=>"010101101",
  56296=>"000000011",
  56297=>"010001111",
  56298=>"001010000",
  56299=>"011101001",
  56300=>"111001110",
  56301=>"001010000",
  56302=>"110110010",
  56303=>"001010101",
  56304=>"001010011",
  56305=>"110101001",
  56306=>"101001101",
  56307=>"000010111",
  56308=>"100000101",
  56309=>"000101001",
  56310=>"000011011",
  56311=>"001111000",
  56312=>"100111001",
  56313=>"100110111",
  56314=>"010000000",
  56315=>"100000110",
  56316=>"000011111",
  56317=>"100110010",
  56318=>"010110010",
  56319=>"010100010",
  56320=>"100101101",
  56321=>"001111000",
  56322=>"011111000",
  56323=>"011000111",
  56324=>"111100011",
  56325=>"101000001",
  56326=>"000110001",
  56327=>"101100110",
  56328=>"011110110",
  56329=>"111100110",
  56330=>"001111000",
  56331=>"011111110",
  56332=>"100101000",
  56333=>"110010100",
  56334=>"110111010",
  56335=>"000101100",
  56336=>"110110011",
  56337=>"000111100",
  56338=>"110000110",
  56339=>"100001100",
  56340=>"101010101",
  56341=>"010010100",
  56342=>"010111110",
  56343=>"100101111",
  56344=>"101100010",
  56345=>"000000001",
  56346=>"011000101",
  56347=>"000100000",
  56348=>"000000101",
  56349=>"111101000",
  56350=>"111011000",
  56351=>"000010001",
  56352=>"000001111",
  56353=>"000101001",
  56354=>"011000100",
  56355=>"011111100",
  56356=>"110111101",
  56357=>"100001010",
  56358=>"101101000",
  56359=>"010010100",
  56360=>"010000001",
  56361=>"100011111",
  56362=>"010100111",
  56363=>"100011011",
  56364=>"111010010",
  56365=>"101111001",
  56366=>"000101010",
  56367=>"111000000",
  56368=>"011110011",
  56369=>"100110001",
  56370=>"010100000",
  56371=>"111011100",
  56372=>"001001000",
  56373=>"111010001",
  56374=>"000101100",
  56375=>"001110111",
  56376=>"000011011",
  56377=>"101000110",
  56378=>"101000100",
  56379=>"001000001",
  56380=>"010010100",
  56381=>"000111111",
  56382=>"111011001",
  56383=>"000111111",
  56384=>"111111000",
  56385=>"010011011",
  56386=>"011100000",
  56387=>"000001110",
  56388=>"111011011",
  56389=>"001011011",
  56390=>"111110100",
  56391=>"100111011",
  56392=>"001101110",
  56393=>"011101111",
  56394=>"111000000",
  56395=>"011010010",
  56396=>"101100101",
  56397=>"101100101",
  56398=>"110111111",
  56399=>"110000011",
  56400=>"100010110",
  56401=>"000111111",
  56402=>"001101011",
  56403=>"011010001",
  56404=>"101100010",
  56405=>"111111111",
  56406=>"011000100",
  56407=>"100101111",
  56408=>"101010100",
  56409=>"110100000",
  56410=>"111010000",
  56411=>"000000110",
  56412=>"011111111",
  56413=>"100000001",
  56414=>"000100100",
  56415=>"101001100",
  56416=>"001001001",
  56417=>"111110101",
  56418=>"000001001",
  56419=>"100000000",
  56420=>"000101011",
  56421=>"010010000",
  56422=>"011111110",
  56423=>"000000100",
  56424=>"110101101",
  56425=>"010101010",
  56426=>"011110000",
  56427=>"000110101",
  56428=>"110010000",
  56429=>"110101111",
  56430=>"111001111",
  56431=>"000110001",
  56432=>"001000010",
  56433=>"010110110",
  56434=>"110111110",
  56435=>"100111011",
  56436=>"101101010",
  56437=>"010111100",
  56438=>"011101000",
  56439=>"000110100",
  56440=>"000111110",
  56441=>"110010000",
  56442=>"100111100",
  56443=>"100111000",
  56444=>"100011110",
  56445=>"110011000",
  56446=>"101110011",
  56447=>"010111010",
  56448=>"001000001",
  56449=>"011000001",
  56450=>"001011100",
  56451=>"100101111",
  56452=>"111111000",
  56453=>"110101011",
  56454=>"110110100",
  56455=>"011111011",
  56456=>"011001111",
  56457=>"010101001",
  56458=>"101100100",
  56459=>"000000011",
  56460=>"100110111",
  56461=>"111101000",
  56462=>"110000111",
  56463=>"111001111",
  56464=>"100000011",
  56465=>"001001110",
  56466=>"001101010",
  56467=>"001100011",
  56468=>"001100111",
  56469=>"110111011",
  56470=>"010001101",
  56471=>"000010001",
  56472=>"001110000",
  56473=>"111011110",
  56474=>"110110100",
  56475=>"111011101",
  56476=>"011000111",
  56477=>"010110000",
  56478=>"000110000",
  56479=>"011110101",
  56480=>"011010100",
  56481=>"011000001",
  56482=>"111010100",
  56483=>"000100001",
  56484=>"101000110",
  56485=>"111111011",
  56486=>"100010001",
  56487=>"110110000",
  56488=>"010001110",
  56489=>"111111000",
  56490=>"010110001",
  56491=>"101000010",
  56492=>"110010010",
  56493=>"100101110",
  56494=>"010100001",
  56495=>"111111000",
  56496=>"001011011",
  56497=>"011011101",
  56498=>"010101101",
  56499=>"011110110",
  56500=>"000011010",
  56501=>"000010000",
  56502=>"001000001",
  56503=>"011011100",
  56504=>"100001110",
  56505=>"100100011",
  56506=>"011110000",
  56507=>"100011010",
  56508=>"101000110",
  56509=>"010011001",
  56510=>"001001001",
  56511=>"111011000",
  56512=>"101010010",
  56513=>"111110010",
  56514=>"000111000",
  56515=>"010011010",
  56516=>"110110101",
  56517=>"100100100",
  56518=>"000000010",
  56519=>"111001100",
  56520=>"010011000",
  56521=>"111101110",
  56522=>"011111010",
  56523=>"011111110",
  56524=>"100000101",
  56525=>"010101101",
  56526=>"000111101",
  56527=>"001011110",
  56528=>"010110011",
  56529=>"101010101",
  56530=>"100110100",
  56531=>"110101001",
  56532=>"000111001",
  56533=>"001010001",
  56534=>"110000000",
  56535=>"000101010",
  56536=>"100001011",
  56537=>"101000001",
  56538=>"001110011",
  56539=>"010111010",
  56540=>"100011001",
  56541=>"101010011",
  56542=>"011100110",
  56543=>"010011000",
  56544=>"101010011",
  56545=>"001111111",
  56546=>"011011101",
  56547=>"000101110",
  56548=>"000010111",
  56549=>"100100110",
  56550=>"110110100",
  56551=>"001010100",
  56552=>"110110011",
  56553=>"111110100",
  56554=>"000011001",
  56555=>"111101101",
  56556=>"010101100",
  56557=>"000010111",
  56558=>"010001011",
  56559=>"111000001",
  56560=>"101011011",
  56561=>"111111101",
  56562=>"100001100",
  56563=>"011100001",
  56564=>"111010001",
  56565=>"110100000",
  56566=>"000000011",
  56567=>"110010100",
  56568=>"100100110",
  56569=>"001001111",
  56570=>"010000110",
  56571=>"100010010",
  56572=>"000000110",
  56573=>"110011110",
  56574=>"001101000",
  56575=>"000001101",
  56576=>"011100110",
  56577=>"101100011",
  56578=>"000101010",
  56579=>"000110010",
  56580=>"101110111",
  56581=>"000001001",
  56582=>"000011011",
  56583=>"110100100",
  56584=>"001101110",
  56585=>"111101011",
  56586=>"000111110",
  56587=>"000111001",
  56588=>"110010111",
  56589=>"010010111",
  56590=>"011010101",
  56591=>"000110111",
  56592=>"110001111",
  56593=>"110101011",
  56594=>"110101010",
  56595=>"001011001",
  56596=>"010110000",
  56597=>"110100110",
  56598=>"000100000",
  56599=>"111011110",
  56600=>"110010100",
  56601=>"100110001",
  56602=>"101010000",
  56603=>"111010000",
  56604=>"010111100",
  56605=>"010100110",
  56606=>"001010010",
  56607=>"100011000",
  56608=>"100010011",
  56609=>"101001110",
  56610=>"101111101",
  56611=>"110001101",
  56612=>"110110010",
  56613=>"111101001",
  56614=>"010110011",
  56615=>"000101101",
  56616=>"100000011",
  56617=>"101001000",
  56618=>"110111100",
  56619=>"000011001",
  56620=>"111111000",
  56621=>"000101110",
  56622=>"001101100",
  56623=>"001001111",
  56624=>"101110101",
  56625=>"010111001",
  56626=>"110111000",
  56627=>"011110011",
  56628=>"011001110",
  56629=>"110011101",
  56630=>"011111110",
  56631=>"110110010",
  56632=>"001001011",
  56633=>"110111101",
  56634=>"010110101",
  56635=>"011010001",
  56636=>"001011001",
  56637=>"010000001",
  56638=>"000001001",
  56639=>"011110010",
  56640=>"010100000",
  56641=>"000100011",
  56642=>"101110110",
  56643=>"001001101",
  56644=>"001100001",
  56645=>"101100010",
  56646=>"101001010",
  56647=>"010110101",
  56648=>"011110100",
  56649=>"101000110",
  56650=>"110100001",
  56651=>"000111101",
  56652=>"101100000",
  56653=>"000110111",
  56654=>"010111100",
  56655=>"111011010",
  56656=>"010000100",
  56657=>"101101111",
  56658=>"010111011",
  56659=>"010011100",
  56660=>"110010101",
  56661=>"001100111",
  56662=>"100010000",
  56663=>"101110011",
  56664=>"100101000",
  56665=>"111110101",
  56666=>"010111100",
  56667=>"111100110",
  56668=>"001101010",
  56669=>"000000111",
  56670=>"101110100",
  56671=>"000111001",
  56672=>"101001001",
  56673=>"111011111",
  56674=>"100111100",
  56675=>"001000101",
  56676=>"111001010",
  56677=>"110101110",
  56678=>"000010110",
  56679=>"110010001",
  56680=>"100001000",
  56681=>"001010111",
  56682=>"101000100",
  56683=>"011110000",
  56684=>"000010000",
  56685=>"111111011",
  56686=>"110110010",
  56687=>"000000001",
  56688=>"001001101",
  56689=>"100101111",
  56690=>"001011111",
  56691=>"100000011",
  56692=>"101000000",
  56693=>"010000001",
  56694=>"001011100",
  56695=>"101101110",
  56696=>"100010011",
  56697=>"100110011",
  56698=>"000110001",
  56699=>"111111000",
  56700=>"101011001",
  56701=>"010001010",
  56702=>"001011111",
  56703=>"100001100",
  56704=>"111000000",
  56705=>"011111110",
  56706=>"011011111",
  56707=>"010000010",
  56708=>"101111110",
  56709=>"100110011",
  56710=>"001011101",
  56711=>"010000010",
  56712=>"101001101",
  56713=>"001110000",
  56714=>"010011110",
  56715=>"011010101",
  56716=>"101100010",
  56717=>"000011101",
  56718=>"111100100",
  56719=>"111101010",
  56720=>"101110111",
  56721=>"100110000",
  56722=>"101100110",
  56723=>"001001011",
  56724=>"010011111",
  56725=>"000100001",
  56726=>"101010111",
  56727=>"100111001",
  56728=>"110000100",
  56729=>"100000101",
  56730=>"011000111",
  56731=>"011010111",
  56732=>"010010110",
  56733=>"111110100",
  56734=>"101110110",
  56735=>"010110000",
  56736=>"010011001",
  56737=>"100110011",
  56738=>"101100100",
  56739=>"011111010",
  56740=>"100000000",
  56741=>"111000001",
  56742=>"011100011",
  56743=>"001011101",
  56744=>"101000111",
  56745=>"010101000",
  56746=>"100100110",
  56747=>"010110010",
  56748=>"011011000",
  56749=>"011010000",
  56750=>"111000110",
  56751=>"101111110",
  56752=>"010000101",
  56753=>"000010000",
  56754=>"101001010",
  56755=>"000000110",
  56756=>"101101011",
  56757=>"101000110",
  56758=>"000011111",
  56759=>"101101110",
  56760=>"000001001",
  56761=>"000101100",
  56762=>"111001100",
  56763=>"110000011",
  56764=>"011001001",
  56765=>"101010001",
  56766=>"011011000",
  56767=>"111011000",
  56768=>"011100100",
  56769=>"000100110",
  56770=>"000001010",
  56771=>"000010001",
  56772=>"111100011",
  56773=>"011101111",
  56774=>"101101110",
  56775=>"111101000",
  56776=>"100000100",
  56777=>"110110010",
  56778=>"001000100",
  56779=>"111001100",
  56780=>"110110101",
  56781=>"101010100",
  56782=>"011110010",
  56783=>"101010110",
  56784=>"100101001",
  56785=>"001000001",
  56786=>"001100000",
  56787=>"011011000",
  56788=>"001010111",
  56789=>"001101100",
  56790=>"110010100",
  56791=>"110001000",
  56792=>"010010111",
  56793=>"111111010",
  56794=>"110101011",
  56795=>"000010001",
  56796=>"101011010",
  56797=>"100011110",
  56798=>"110111110",
  56799=>"000111100",
  56800=>"010100110",
  56801=>"100111001",
  56802=>"111010000",
  56803=>"011110000",
  56804=>"001111011",
  56805=>"111000100",
  56806=>"000101101",
  56807=>"101111000",
  56808=>"001101000",
  56809=>"011001011",
  56810=>"000010111",
  56811=>"001111101",
  56812=>"001000100",
  56813=>"000000000",
  56814=>"100100010",
  56815=>"101101110",
  56816=>"111001110",
  56817=>"111010001",
  56818=>"000001011",
  56819=>"101100100",
  56820=>"100111000",
  56821=>"101010101",
  56822=>"111101011",
  56823=>"110001011",
  56824=>"001111000",
  56825=>"100110011",
  56826=>"110101111",
  56827=>"001101001",
  56828=>"000100000",
  56829=>"000100000",
  56830=>"001011111",
  56831=>"111111000",
  56832=>"000011111",
  56833=>"110000101",
  56834=>"000101010",
  56835=>"110010110",
  56836=>"011111011",
  56837=>"000100111",
  56838=>"100011001",
  56839=>"010000101",
  56840=>"001000000",
  56841=>"110011010",
  56842=>"000110010",
  56843=>"010011000",
  56844=>"001101000",
  56845=>"101110001",
  56846=>"111000111",
  56847=>"001110010",
  56848=>"100101100",
  56849=>"011111101",
  56850=>"101111001",
  56851=>"110001000",
  56852=>"010111100",
  56853=>"000011110",
  56854=>"101101110",
  56855=>"101011000",
  56856=>"001100010",
  56857=>"111111101",
  56858=>"000000001",
  56859=>"110011101",
  56860=>"101000001",
  56861=>"110000010",
  56862=>"100100101",
  56863=>"010011111",
  56864=>"000001010",
  56865=>"101111011",
  56866=>"001011111",
  56867=>"010001000",
  56868=>"011001011",
  56869=>"111110111",
  56870=>"001001110",
  56871=>"010000000",
  56872=>"100001000",
  56873=>"110000001",
  56874=>"111101001",
  56875=>"010111100",
  56876=>"010101011",
  56877=>"000001011",
  56878=>"111010001",
  56879=>"011000010",
  56880=>"010100111",
  56881=>"111101011",
  56882=>"010100111",
  56883=>"111010111",
  56884=>"110000100",
  56885=>"101011001",
  56886=>"011110100",
  56887=>"111000011",
  56888=>"010000000",
  56889=>"111001000",
  56890=>"101110111",
  56891=>"001001001",
  56892=>"000000111",
  56893=>"110010010",
  56894=>"101001010",
  56895=>"100001101",
  56896=>"110100101",
  56897=>"110001111",
  56898=>"110001001",
  56899=>"010011001",
  56900=>"110111000",
  56901=>"011110010",
  56902=>"100100001",
  56903=>"000010110",
  56904=>"110100011",
  56905=>"100101000",
  56906=>"011110000",
  56907=>"011001111",
  56908=>"101110111",
  56909=>"110110010",
  56910=>"100001101",
  56911=>"001001010",
  56912=>"010100000",
  56913=>"011000001",
  56914=>"001111101",
  56915=>"000100010",
  56916=>"011000010",
  56917=>"011110110",
  56918=>"011111011",
  56919=>"110100111",
  56920=>"100011111",
  56921=>"001100000",
  56922=>"010101100",
  56923=>"010101101",
  56924=>"101100000",
  56925=>"111111101",
  56926=>"101101000",
  56927=>"000111100",
  56928=>"000110011",
  56929=>"110101101",
  56930=>"101101101",
  56931=>"001001101",
  56932=>"111110011",
  56933=>"001100111",
  56934=>"101111000",
  56935=>"001000010",
  56936=>"001010111",
  56937=>"100011110",
  56938=>"111111001",
  56939=>"010000000",
  56940=>"100010101",
  56941=>"011011111",
  56942=>"101001110",
  56943=>"100111100",
  56944=>"010011101",
  56945=>"001011000",
  56946=>"100111011",
  56947=>"001101010",
  56948=>"001010110",
  56949=>"110100110",
  56950=>"011100000",
  56951=>"100010011",
  56952=>"011001010",
  56953=>"110100111",
  56954=>"101010001",
  56955=>"000011000",
  56956=>"110001000",
  56957=>"001110110",
  56958=>"110101100",
  56959=>"111110011",
  56960=>"100010001",
  56961=>"001010100",
  56962=>"001101000",
  56963=>"000000001",
  56964=>"000110110",
  56965=>"110101101",
  56966=>"010100100",
  56967=>"011011001",
  56968=>"100110010",
  56969=>"110100110",
  56970=>"111011111",
  56971=>"110001101",
  56972=>"000010010",
  56973=>"110001110",
  56974=>"110001100",
  56975=>"000010101",
  56976=>"010101100",
  56977=>"101100101",
  56978=>"110001111",
  56979=>"001111000",
  56980=>"101000000",
  56981=>"000010001",
  56982=>"000101001",
  56983=>"000001001",
  56984=>"011001101",
  56985=>"110010101",
  56986=>"000011001",
  56987=>"100101010",
  56988=>"100010000",
  56989=>"110100100",
  56990=>"110000011",
  56991=>"010010000",
  56992=>"011000011",
  56993=>"100101010",
  56994=>"000000000",
  56995=>"100101111",
  56996=>"011000100",
  56997=>"100110111",
  56998=>"110111001",
  56999=>"100100011",
  57000=>"001001100",
  57001=>"100001101",
  57002=>"001000110",
  57003=>"001000001",
  57004=>"010000111",
  57005=>"101011011",
  57006=>"111100100",
  57007=>"110000011",
  57008=>"100001111",
  57009=>"101111001",
  57010=>"011010100",
  57011=>"110001010",
  57012=>"010110001",
  57013=>"000110101",
  57014=>"011111010",
  57015=>"000011000",
  57016=>"010001010",
  57017=>"011100111",
  57018=>"001100011",
  57019=>"000000110",
  57020=>"010000110",
  57021=>"000000100",
  57022=>"101101100",
  57023=>"001011110",
  57024=>"001110110",
  57025=>"111111101",
  57026=>"000101110",
  57027=>"000111111",
  57028=>"110001111",
  57029=>"011010010",
  57030=>"010111111",
  57031=>"110010010",
  57032=>"000101000",
  57033=>"100001011",
  57034=>"110000011",
  57035=>"011100011",
  57036=>"100110111",
  57037=>"101111100",
  57038=>"101110001",
  57039=>"011010000",
  57040=>"100110000",
  57041=>"100100011",
  57042=>"101111011",
  57043=>"110010000",
  57044=>"100100111",
  57045=>"001001110",
  57046=>"001011011",
  57047=>"001000111",
  57048=>"000001111",
  57049=>"001101000",
  57050=>"001100100",
  57051=>"010101001",
  57052=>"101101001",
  57053=>"111100001",
  57054=>"011001010",
  57055=>"001011000",
  57056=>"111000010",
  57057=>"010010000",
  57058=>"011011101",
  57059=>"010010101",
  57060=>"000010001",
  57061=>"110011111",
  57062=>"001100110",
  57063=>"100101101",
  57064=>"011110001",
  57065=>"110001101",
  57066=>"000011111",
  57067=>"010100000",
  57068=>"100100101",
  57069=>"100001110",
  57070=>"000001010",
  57071=>"101110011",
  57072=>"011010101",
  57073=>"000111111",
  57074=>"001110010",
  57075=>"111111001",
  57076=>"010010101",
  57077=>"011000010",
  57078=>"011010000",
  57079=>"001001110",
  57080=>"101010010",
  57081=>"011100000",
  57082=>"100010001",
  57083=>"010000111",
  57084=>"001001011",
  57085=>"100011010",
  57086=>"001000011",
  57087=>"111111101",
  57088=>"011001000",
  57089=>"100010100",
  57090=>"011001100",
  57091=>"111101000",
  57092=>"100101110",
  57093=>"010001001",
  57094=>"101011100",
  57095=>"101111110",
  57096=>"010111001",
  57097=>"010100011",
  57098=>"111001111",
  57099=>"111001011",
  57100=>"001010001",
  57101=>"010110011",
  57102=>"110000000",
  57103=>"010111110",
  57104=>"011001111",
  57105=>"100001010",
  57106=>"101000000",
  57107=>"011101101",
  57108=>"001110100",
  57109=>"011010010",
  57110=>"100000000",
  57111=>"110011001",
  57112=>"000100100",
  57113=>"100010001",
  57114=>"111111111",
  57115=>"000011011",
  57116=>"001000011",
  57117=>"100110111",
  57118=>"110010010",
  57119=>"001000011",
  57120=>"001111111",
  57121=>"001111000",
  57122=>"110100101",
  57123=>"100000000",
  57124=>"101000101",
  57125=>"100110000",
  57126=>"011110101",
  57127=>"001001010",
  57128=>"010100000",
  57129=>"101111100",
  57130=>"111001000",
  57131=>"001100100",
  57132=>"001111010",
  57133=>"110011101",
  57134=>"000100000",
  57135=>"110000111",
  57136=>"111101001",
  57137=>"111010101",
  57138=>"100010101",
  57139=>"101111111",
  57140=>"000110011",
  57141=>"111100100",
  57142=>"000010010",
  57143=>"001111100",
  57144=>"000111011",
  57145=>"000000100",
  57146=>"000011010",
  57147=>"010111111",
  57148=>"000000101",
  57149=>"001110110",
  57150=>"111100100",
  57151=>"001011001",
  57152=>"011000011",
  57153=>"010101011",
  57154=>"000010010",
  57155=>"001110111",
  57156=>"101101011",
  57157=>"100010000",
  57158=>"101001101",
  57159=>"110010011",
  57160=>"110001110",
  57161=>"010011100",
  57162=>"101011010",
  57163=>"101010101",
  57164=>"000100000",
  57165=>"110010010",
  57166=>"000010000",
  57167=>"110000100",
  57168=>"001100000",
  57169=>"111001011",
  57170=>"010000110",
  57171=>"110000001",
  57172=>"111111011",
  57173=>"010100100",
  57174=>"000100010",
  57175=>"010000001",
  57176=>"011100001",
  57177=>"011111001",
  57178=>"111100110",
  57179=>"100101111",
  57180=>"011100111",
  57181=>"110101101",
  57182=>"010001100",
  57183=>"010100110",
  57184=>"110100000",
  57185=>"111010101",
  57186=>"000001010",
  57187=>"100101111",
  57188=>"010111000",
  57189=>"111000011",
  57190=>"010100110",
  57191=>"010100010",
  57192=>"101010000",
  57193=>"010000010",
  57194=>"110000100",
  57195=>"011100111",
  57196=>"010101000",
  57197=>"010011100",
  57198=>"101100111",
  57199=>"111100101",
  57200=>"101111000",
  57201=>"010100101",
  57202=>"000110000",
  57203=>"000111100",
  57204=>"000010110",
  57205=>"001101001",
  57206=>"001110011",
  57207=>"011110000",
  57208=>"001001100",
  57209=>"110100101",
  57210=>"010100110",
  57211=>"011011000",
  57212=>"100110110",
  57213=>"111011101",
  57214=>"100000110",
  57215=>"110111010",
  57216=>"100011110",
  57217=>"001101010",
  57218=>"001000111",
  57219=>"010101111",
  57220=>"000111010",
  57221=>"000101010",
  57222=>"111101111",
  57223=>"010100010",
  57224=>"100110101",
  57225=>"001101000",
  57226=>"100001100",
  57227=>"011100100",
  57228=>"011010111",
  57229=>"001100010",
  57230=>"001111011",
  57231=>"001111111",
  57232=>"010000100",
  57233=>"011110101",
  57234=>"001000111",
  57235=>"000110011",
  57236=>"111110101",
  57237=>"111100000",
  57238=>"010100001",
  57239=>"000101101",
  57240=>"001101110",
  57241=>"100100101",
  57242=>"001100001",
  57243=>"000110100",
  57244=>"010000101",
  57245=>"111001010",
  57246=>"001000001",
  57247=>"111011010",
  57248=>"110100000",
  57249=>"110100000",
  57250=>"001011110",
  57251=>"100101010",
  57252=>"100000001",
  57253=>"110101110",
  57254=>"000101111",
  57255=>"101111011",
  57256=>"100101100",
  57257=>"010001001",
  57258=>"011110011",
  57259=>"001100110",
  57260=>"000010000",
  57261=>"011001110",
  57262=>"001111110",
  57263=>"101010010",
  57264=>"010010110",
  57265=>"011011010",
  57266=>"001000000",
  57267=>"011000110",
  57268=>"010111001",
  57269=>"100111110",
  57270=>"111100011",
  57271=>"111011001",
  57272=>"001001100",
  57273=>"100110100",
  57274=>"110010101",
  57275=>"101010101",
  57276=>"110000101",
  57277=>"010110100",
  57278=>"000011011",
  57279=>"010100110",
  57280=>"011111001",
  57281=>"111101101",
  57282=>"000000100",
  57283=>"110001100",
  57284=>"100000111",
  57285=>"101011100",
  57286=>"100010000",
  57287=>"000011111",
  57288=>"100001011",
  57289=>"101101101",
  57290=>"101100001",
  57291=>"110110000",
  57292=>"010101111",
  57293=>"100100111",
  57294=>"011111001",
  57295=>"001110100",
  57296=>"110101100",
  57297=>"001101110",
  57298=>"001001010",
  57299=>"011110100",
  57300=>"101000101",
  57301=>"010000011",
  57302=>"010001011",
  57303=>"110000111",
  57304=>"000010101",
  57305=>"001110110",
  57306=>"100111100",
  57307=>"000010110",
  57308=>"000010100",
  57309=>"001111111",
  57310=>"101000101",
  57311=>"000001010",
  57312=>"010100010",
  57313=>"001110100",
  57314=>"010101110",
  57315=>"100100100",
  57316=>"011010101",
  57317=>"101000001",
  57318=>"001110101",
  57319=>"011110000",
  57320=>"110010011",
  57321=>"100110001",
  57322=>"101001111",
  57323=>"110100111",
  57324=>"111111001",
  57325=>"011101111",
  57326=>"100100101",
  57327=>"110111010",
  57328=>"011100111",
  57329=>"010011101",
  57330=>"001101001",
  57331=>"000110010",
  57332=>"010100001",
  57333=>"010111110",
  57334=>"010110000",
  57335=>"000100000",
  57336=>"011010000",
  57337=>"001001000",
  57338=>"101111001",
  57339=>"100111010",
  57340=>"100100111",
  57341=>"001011100",
  57342=>"111000111",
  57343=>"010111110",
  57344=>"011110011",
  57345=>"011000111",
  57346=>"101100010",
  57347=>"111010011",
  57348=>"010011000",
  57349=>"000000110",
  57350=>"100011001",
  57351=>"111000001",
  57352=>"010100101",
  57353=>"110010010",
  57354=>"010001100",
  57355=>"111100100",
  57356=>"000001100",
  57357=>"010111010",
  57358=>"101111001",
  57359=>"111111011",
  57360=>"000110101",
  57361=>"110100001",
  57362=>"001011011",
  57363=>"100111000",
  57364=>"001100111",
  57365=>"101111111",
  57366=>"110011010",
  57367=>"111000010",
  57368=>"110010100",
  57369=>"101101001",
  57370=>"110010101",
  57371=>"000010001",
  57372=>"001000100",
  57373=>"011011000",
  57374=>"000001101",
  57375=>"110100110",
  57376=>"111011101",
  57377=>"000101011",
  57378=>"001011011",
  57379=>"000100101",
  57380=>"000100000",
  57381=>"001111111",
  57382=>"000100100",
  57383=>"011111110",
  57384=>"000001111",
  57385=>"011011010",
  57386=>"011110000",
  57387=>"001010110",
  57388=>"110101001",
  57389=>"111001111",
  57390=>"101111100",
  57391=>"100000110",
  57392=>"111011111",
  57393=>"110001100",
  57394=>"010111001",
  57395=>"011000110",
  57396=>"000011111",
  57397=>"011010100",
  57398=>"110010010",
  57399=>"011110011",
  57400=>"101110110",
  57401=>"001000000",
  57402=>"010101111",
  57403=>"100111001",
  57404=>"100011001",
  57405=>"110111111",
  57406=>"101101011",
  57407=>"000000001",
  57408=>"110101110",
  57409=>"111010000",
  57410=>"001100000",
  57411=>"011010011",
  57412=>"100011100",
  57413=>"110100111",
  57414=>"000001011",
  57415=>"101000000",
  57416=>"111011011",
  57417=>"110110000",
  57418=>"010101100",
  57419=>"100000100",
  57420=>"011111010",
  57421=>"010010010",
  57422=>"111101011",
  57423=>"111110110",
  57424=>"001011011",
  57425=>"000101010",
  57426=>"001010110",
  57427=>"100000010",
  57428=>"010111111",
  57429=>"011001001",
  57430=>"110011000",
  57431=>"110001001",
  57432=>"101001000",
  57433=>"010010000",
  57434=>"000010011",
  57435=>"011100000",
  57436=>"100110011",
  57437=>"011001101",
  57438=>"101110001",
  57439=>"000000001",
  57440=>"000010001",
  57441=>"011010111",
  57442=>"100100101",
  57443=>"111001111",
  57444=>"100000001",
  57445=>"010110100",
  57446=>"011111001",
  57447=>"000101011",
  57448=>"010110010",
  57449=>"011110010",
  57450=>"010011010",
  57451=>"011011011",
  57452=>"110110100",
  57453=>"011001101",
  57454=>"010101101",
  57455=>"010011111",
  57456=>"101000110",
  57457=>"101001101",
  57458=>"111111110",
  57459=>"001000101",
  57460=>"000100111",
  57461=>"001111100",
  57462=>"111101100",
  57463=>"000101100",
  57464=>"111101110",
  57465=>"011000010",
  57466=>"010011111",
  57467=>"100100010",
  57468=>"000011001",
  57469=>"101001000",
  57470=>"000100000",
  57471=>"010111001",
  57472=>"110110001",
  57473=>"000000001",
  57474=>"001010010",
  57475=>"100100111",
  57476=>"111011010",
  57477=>"001100111",
  57478=>"011010100",
  57479=>"100001110",
  57480=>"000110011",
  57481=>"001100110",
  57482=>"100011000",
  57483=>"101111000",
  57484=>"100000101",
  57485=>"110000011",
  57486=>"101000011",
  57487=>"001111100",
  57488=>"000000011",
  57489=>"010110111",
  57490=>"100110000",
  57491=>"000001111",
  57492=>"000001101",
  57493=>"111111100",
  57494=>"110010011",
  57495=>"101111000",
  57496=>"010110001",
  57497=>"111110111",
  57498=>"101001110",
  57499=>"011010101",
  57500=>"111001010",
  57501=>"111001101",
  57502=>"101000010",
  57503=>"101111000",
  57504=>"001001010",
  57505=>"001101100",
  57506=>"111110001",
  57507=>"010011011",
  57508=>"000001001",
  57509=>"111111110",
  57510=>"111100101",
  57511=>"101011010",
  57512=>"110011010",
  57513=>"101100000",
  57514=>"001000011",
  57515=>"000011000",
  57516=>"111000000",
  57517=>"111001011",
  57518=>"100100000",
  57519=>"000000011",
  57520=>"000011000",
  57521=>"111110100",
  57522=>"011110101",
  57523=>"001101001",
  57524=>"101100110",
  57525=>"111011111",
  57526=>"000001000",
  57527=>"100101101",
  57528=>"001000000",
  57529=>"101100001",
  57530=>"000001110",
  57531=>"000010000",
  57532=>"111001001",
  57533=>"000010001",
  57534=>"011000011",
  57535=>"100011101",
  57536=>"001000100",
  57537=>"000001110",
  57538=>"011110000",
  57539=>"111100100",
  57540=>"010001000",
  57541=>"001001010",
  57542=>"001111101",
  57543=>"111011001",
  57544=>"101100010",
  57545=>"000110101",
  57546=>"000000000",
  57547=>"100101110",
  57548=>"101100011",
  57549=>"011011001",
  57550=>"000000100",
  57551=>"000110011",
  57552=>"110100000",
  57553=>"001011010",
  57554=>"111001011",
  57555=>"101101011",
  57556=>"001010100",
  57557=>"111000110",
  57558=>"100010101",
  57559=>"111011101",
  57560=>"001011001",
  57561=>"010111101",
  57562=>"011110111",
  57563=>"010110101",
  57564=>"100110101",
  57565=>"001001000",
  57566=>"001010010",
  57567=>"100101100",
  57568=>"101111001",
  57569=>"001110100",
  57570=>"010100011",
  57571=>"111001111",
  57572=>"011110101",
  57573=>"000101100",
  57574=>"001110010",
  57575=>"000011110",
  57576=>"111101110",
  57577=>"010010001",
  57578=>"111010111",
  57579=>"010101001",
  57580=>"101100110",
  57581=>"100100000",
  57582=>"011001110",
  57583=>"000010000",
  57584=>"110111101",
  57585=>"111111110",
  57586=>"000110010",
  57587=>"111110101",
  57588=>"011101001",
  57589=>"010101010",
  57590=>"111111100",
  57591=>"001100100",
  57592=>"110100110",
  57593=>"001001010",
  57594=>"111011100",
  57595=>"111110001",
  57596=>"000000011",
  57597=>"100100111",
  57598=>"000110010",
  57599=>"101011111",
  57600=>"101011111",
  57601=>"010111010",
  57602=>"000010101",
  57603=>"001101011",
  57604=>"111110010",
  57605=>"011101011",
  57606=>"011001101",
  57607=>"111000000",
  57608=>"101111000",
  57609=>"010001100",
  57610=>"101010101",
  57611=>"011000001",
  57612=>"000011111",
  57613=>"010100000",
  57614=>"101001011",
  57615=>"001001110",
  57616=>"100110111",
  57617=>"011110101",
  57618=>"000000000",
  57619=>"110010001",
  57620=>"110010100",
  57621=>"101110100",
  57622=>"000100100",
  57623=>"010100100",
  57624=>"101001111",
  57625=>"101011101",
  57626=>"000101101",
  57627=>"111001100",
  57628=>"001101001",
  57629=>"011011001",
  57630=>"111110001",
  57631=>"010001000",
  57632=>"100010111",
  57633=>"100010100",
  57634=>"010110110",
  57635=>"010111010",
  57636=>"011000000",
  57637=>"111110001",
  57638=>"001011100",
  57639=>"100001110",
  57640=>"111011111",
  57641=>"111111000",
  57642=>"101001000",
  57643=>"101101010",
  57644=>"001101011",
  57645=>"110111010",
  57646=>"001000010",
  57647=>"111000011",
  57648=>"100000000",
  57649=>"000111101",
  57650=>"100110111",
  57651=>"000010001",
  57652=>"110100100",
  57653=>"110111100",
  57654=>"110010010",
  57655=>"110100111",
  57656=>"111101111",
  57657=>"011011001",
  57658=>"110110011",
  57659=>"110110000",
  57660=>"001001011",
  57661=>"001101010",
  57662=>"010001010",
  57663=>"000110011",
  57664=>"001100110",
  57665=>"011101110",
  57666=>"000000011",
  57667=>"111001010",
  57668=>"100111100",
  57669=>"000101101",
  57670=>"110000010",
  57671=>"001010011",
  57672=>"000011101",
  57673=>"010100011",
  57674=>"001001001",
  57675=>"010010010",
  57676=>"110110111",
  57677=>"010100001",
  57678=>"001110010",
  57679=>"010111001",
  57680=>"011110010",
  57681=>"101100001",
  57682=>"100010011",
  57683=>"111101011",
  57684=>"101001110",
  57685=>"001111101",
  57686=>"101110111",
  57687=>"010001111",
  57688=>"110111000",
  57689=>"000001111",
  57690=>"000111010",
  57691=>"101001100",
  57692=>"011101000",
  57693=>"011100101",
  57694=>"100010000",
  57695=>"100010111",
  57696=>"111100111",
  57697=>"111111001",
  57698=>"101000101",
  57699=>"100000011",
  57700=>"000100101",
  57701=>"110000001",
  57702=>"011010001",
  57703=>"111110010",
  57704=>"001010011",
  57705=>"110000001",
  57706=>"000000101",
  57707=>"100011000",
  57708=>"110100110",
  57709=>"110111100",
  57710=>"100100000",
  57711=>"111010001",
  57712=>"010001100",
  57713=>"111111001",
  57714=>"110111010",
  57715=>"011100001",
  57716=>"011100010",
  57717=>"111111110",
  57718=>"010000100",
  57719=>"101111001",
  57720=>"101101110",
  57721=>"011101110",
  57722=>"000101010",
  57723=>"001000111",
  57724=>"110001010",
  57725=>"111111100",
  57726=>"101110110",
  57727=>"010111111",
  57728=>"110110000",
  57729=>"000011000",
  57730=>"001100101",
  57731=>"010011000",
  57732=>"011011101",
  57733=>"001000010",
  57734=>"110000110",
  57735=>"110010001",
  57736=>"001110000",
  57737=>"111000110",
  57738=>"000001001",
  57739=>"110111110",
  57740=>"100001110",
  57741=>"011110110",
  57742=>"101000110",
  57743=>"000001011",
  57744=>"000011010",
  57745=>"000111001",
  57746=>"111010001",
  57747=>"100111110",
  57748=>"111100101",
  57749=>"000001011",
  57750=>"001110011",
  57751=>"111001011",
  57752=>"011010011",
  57753=>"001001001",
  57754=>"010101011",
  57755=>"011001100",
  57756=>"000010101",
  57757=>"000000101",
  57758=>"000000100",
  57759=>"101110111",
  57760=>"011100010",
  57761=>"111001001",
  57762=>"011111110",
  57763=>"000001000",
  57764=>"010100100",
  57765=>"100000010",
  57766=>"111000000",
  57767=>"101000000",
  57768=>"011111100",
  57769=>"110010000",
  57770=>"110011110",
  57771=>"100011010",
  57772=>"011011010",
  57773=>"101001000",
  57774=>"110111101",
  57775=>"100101010",
  57776=>"011011001",
  57777=>"101001001",
  57778=>"001110111",
  57779=>"110010101",
  57780=>"010011011",
  57781=>"101001011",
  57782=>"010111111",
  57783=>"100111010",
  57784=>"111011001",
  57785=>"101000011",
  57786=>"111010011",
  57787=>"011001011",
  57788=>"111111100",
  57789=>"010101101",
  57790=>"010000001",
  57791=>"010101011",
  57792=>"011010010",
  57793=>"101010001",
  57794=>"011110001",
  57795=>"000000001",
  57796=>"001010011",
  57797=>"100101001",
  57798=>"001111101",
  57799=>"100110101",
  57800=>"101111000",
  57801=>"100011000",
  57802=>"100001000",
  57803=>"111110000",
  57804=>"001000101",
  57805=>"110100000",
  57806=>"111100011",
  57807=>"001110000",
  57808=>"001000000",
  57809=>"100001111",
  57810=>"001111101",
  57811=>"001011010",
  57812=>"111101100",
  57813=>"000000100",
  57814=>"111011110",
  57815=>"110111011",
  57816=>"011010011",
  57817=>"011001110",
  57818=>"010100001",
  57819=>"011110110",
  57820=>"011001110",
  57821=>"110000101",
  57822=>"101110111",
  57823=>"101100000",
  57824=>"001111011",
  57825=>"111101100",
  57826=>"001000010",
  57827=>"000010001",
  57828=>"111100011",
  57829=>"011110000",
  57830=>"101010001",
  57831=>"010010000",
  57832=>"010001111",
  57833=>"100110110",
  57834=>"100100010",
  57835=>"111011011",
  57836=>"001001001",
  57837=>"111111110",
  57838=>"001001100",
  57839=>"010110011",
  57840=>"001011101",
  57841=>"101100110",
  57842=>"100001001",
  57843=>"111001001",
  57844=>"001011110",
  57845=>"101100001",
  57846=>"010000100",
  57847=>"111110001",
  57848=>"010001000",
  57849=>"111000101",
  57850=>"101010000",
  57851=>"000010100",
  57852=>"000101000",
  57853=>"100000000",
  57854=>"100011111",
  57855=>"101101111",
  57856=>"100111011",
  57857=>"001000101",
  57858=>"101100110",
  57859=>"000100001",
  57860=>"100001001",
  57861=>"000010101",
  57862=>"001000000",
  57863=>"001001100",
  57864=>"000010110",
  57865=>"011101000",
  57866=>"010101101",
  57867=>"000101010",
  57868=>"000100100",
  57869=>"111100010",
  57870=>"100010101",
  57871=>"000000101",
  57872=>"111000100",
  57873=>"100000111",
  57874=>"000111100",
  57875=>"110111010",
  57876=>"110001101",
  57877=>"101101000",
  57878=>"011010000",
  57879=>"000111000",
  57880=>"001100011",
  57881=>"000001101",
  57882=>"010000010",
  57883=>"011101100",
  57884=>"110110000",
  57885=>"111110100",
  57886=>"010100010",
  57887=>"000001011",
  57888=>"010100011",
  57889=>"110001011",
  57890=>"000101110",
  57891=>"111101100",
  57892=>"110111110",
  57893=>"111011100",
  57894=>"001111100",
  57895=>"001000011",
  57896=>"010000001",
  57897=>"000010001",
  57898=>"001111011",
  57899=>"111000100",
  57900=>"101101111",
  57901=>"000001010",
  57902=>"110000000",
  57903=>"010101111",
  57904=>"100101011",
  57905=>"010010101",
  57906=>"110010110",
  57907=>"100010110",
  57908=>"010010101",
  57909=>"000001101",
  57910=>"000011001",
  57911=>"110011111",
  57912=>"001000110",
  57913=>"010000100",
  57914=>"111001101",
  57915=>"000111100",
  57916=>"111100001",
  57917=>"100010001",
  57918=>"000110110",
  57919=>"000100111",
  57920=>"100100100",
  57921=>"110111010",
  57922=>"110111001",
  57923=>"010111001",
  57924=>"101110010",
  57925=>"111000000",
  57926=>"111000000",
  57927=>"001011101",
  57928=>"000000001",
  57929=>"100001101",
  57930=>"001011100",
  57931=>"010011101",
  57932=>"110001001",
  57933=>"001100110",
  57934=>"100010111",
  57935=>"111111001",
  57936=>"010111010",
  57937=>"100000100",
  57938=>"101010000",
  57939=>"110111001",
  57940=>"110011011",
  57941=>"000000000",
  57942=>"010011000",
  57943=>"010101001",
  57944=>"111100110",
  57945=>"001111111",
  57946=>"110001011",
  57947=>"110010100",
  57948=>"100011001",
  57949=>"000111101",
  57950=>"001001100",
  57951=>"011111100",
  57952=>"000011100",
  57953=>"001001111",
  57954=>"100001101",
  57955=>"011100011",
  57956=>"101001110",
  57957=>"011110111",
  57958=>"011001110",
  57959=>"000001010",
  57960=>"101110100",
  57961=>"100101001",
  57962=>"001011101",
  57963=>"000101000",
  57964=>"000000100",
  57965=>"011100000",
  57966=>"101110000",
  57967=>"110000111",
  57968=>"101011011",
  57969=>"111010101",
  57970=>"100000001",
  57971=>"000001100",
  57972=>"111111011",
  57973=>"000010001",
  57974=>"000010010",
  57975=>"110010111",
  57976=>"101110110",
  57977=>"000111010",
  57978=>"010010111",
  57979=>"111100011",
  57980=>"001001000",
  57981=>"101010010",
  57982=>"111100111",
  57983=>"101001110",
  57984=>"000000010",
  57985=>"100100001",
  57986=>"111111000",
  57987=>"000011000",
  57988=>"001100010",
  57989=>"111101111",
  57990=>"001100001",
  57991=>"001000000",
  57992=>"000000101",
  57993=>"010011100",
  57994=>"001100110",
  57995=>"010100100",
  57996=>"101110111",
  57997=>"010111010",
  57998=>"011111100",
  57999=>"011011001",
  58000=>"001101111",
  58001=>"000001010",
  58002=>"111110100",
  58003=>"101111011",
  58004=>"001101101",
  58005=>"001110111",
  58006=>"101010100",
  58007=>"001010110",
  58008=>"101101110",
  58009=>"101101011",
  58010=>"110110100",
  58011=>"001010110",
  58012=>"010011010",
  58013=>"011100100",
  58014=>"001001001",
  58015=>"011100100",
  58016=>"111111000",
  58017=>"100010111",
  58018=>"100111001",
  58019=>"110101100",
  58020=>"011110111",
  58021=>"010100101",
  58022=>"010100001",
  58023=>"111000000",
  58024=>"011101000",
  58025=>"111100000",
  58026=>"000000001",
  58027=>"111101100",
  58028=>"011111011",
  58029=>"111110000",
  58030=>"111001011",
  58031=>"010111000",
  58032=>"111101000",
  58033=>"010111001",
  58034=>"011100110",
  58035=>"001100010",
  58036=>"000000011",
  58037=>"100101100",
  58038=>"100000100",
  58039=>"000100101",
  58040=>"100111100",
  58041=>"100000000",
  58042=>"101001000",
  58043=>"110011100",
  58044=>"101001101",
  58045=>"110000101",
  58046=>"111000100",
  58047=>"111000101",
  58048=>"100101101",
  58049=>"000111110",
  58050=>"000000001",
  58051=>"000000001",
  58052=>"001111001",
  58053=>"010111100",
  58054=>"111010101",
  58055=>"011010010",
  58056=>"101001111",
  58057=>"100001110",
  58058=>"000100010",
  58059=>"000010000",
  58060=>"011100101",
  58061=>"100110011",
  58062=>"101110111",
  58063=>"101101111",
  58064=>"110101110",
  58065=>"101111000",
  58066=>"010000111",
  58067=>"000000010",
  58068=>"100100100",
  58069=>"000011011",
  58070=>"111100001",
  58071=>"010111010",
  58072=>"011111101",
  58073=>"111010101",
  58074=>"100010110",
  58075=>"111010111",
  58076=>"111000100",
  58077=>"100000010",
  58078=>"101101101",
  58079=>"101110110",
  58080=>"010111010",
  58081=>"001010001",
  58082=>"100110111",
  58083=>"011101111",
  58084=>"011101000",
  58085=>"101101101",
  58086=>"110010000",
  58087=>"100110100",
  58088=>"010001001",
  58089=>"111011111",
  58090=>"101111001",
  58091=>"111101101",
  58092=>"010011011",
  58093=>"000001100",
  58094=>"110000101",
  58095=>"010000000",
  58096=>"000100000",
  58097=>"001100101",
  58098=>"011001000",
  58099=>"101000100",
  58100=>"110011101",
  58101=>"100011010",
  58102=>"001001110",
  58103=>"101010110",
  58104=>"000001010",
  58105=>"010010000",
  58106=>"001011111",
  58107=>"011110001",
  58108=>"100001011",
  58109=>"100100010",
  58110=>"000011111",
  58111=>"010111100",
  58112=>"100101011",
  58113=>"011010100",
  58114=>"001111000",
  58115=>"000111010",
  58116=>"110100010",
  58117=>"100101011",
  58118=>"001111001",
  58119=>"101011011",
  58120=>"110001111",
  58121=>"001000011",
  58122=>"001111011",
  58123=>"000110010",
  58124=>"000011001",
  58125=>"011111011",
  58126=>"101001110",
  58127=>"010100110",
  58128=>"110111111",
  58129=>"011001111",
  58130=>"011111100",
  58131=>"001011111",
  58132=>"010101100",
  58133=>"010001011",
  58134=>"010011010",
  58135=>"111011001",
  58136=>"000110100",
  58137=>"110011101",
  58138=>"011011000",
  58139=>"000010111",
  58140=>"000101010",
  58141=>"011110010",
  58142=>"000111111",
  58143=>"100111010",
  58144=>"101100011",
  58145=>"101001111",
  58146=>"011010000",
  58147=>"010010001",
  58148=>"100000000",
  58149=>"110101100",
  58150=>"111000011",
  58151=>"101010100",
  58152=>"011011001",
  58153=>"110111111",
  58154=>"000101010",
  58155=>"001111110",
  58156=>"000100011",
  58157=>"111000000",
  58158=>"110011000",
  58159=>"101000000",
  58160=>"000001110",
  58161=>"011111110",
  58162=>"011011010",
  58163=>"101111001",
  58164=>"101001010",
  58165=>"111011110",
  58166=>"110010000",
  58167=>"000101001",
  58168=>"001100100",
  58169=>"001111000",
  58170=>"111100011",
  58171=>"110101011",
  58172=>"110110100",
  58173=>"100100110",
  58174=>"001000111",
  58175=>"100111110",
  58176=>"101010010",
  58177=>"010110001",
  58178=>"100000010",
  58179=>"011000000",
  58180=>"010011000",
  58181=>"100011010",
  58182=>"100000111",
  58183=>"011111000",
  58184=>"110001111",
  58185=>"010011011",
  58186=>"100000011",
  58187=>"100011110",
  58188=>"001111000",
  58189=>"100101011",
  58190=>"001001111",
  58191=>"000011111",
  58192=>"110010000",
  58193=>"110000010",
  58194=>"101001000",
  58195=>"101111111",
  58196=>"000110101",
  58197=>"110010100",
  58198=>"010100100",
  58199=>"111010101",
  58200=>"100111111",
  58201=>"001000111",
  58202=>"011101111",
  58203=>"010111100",
  58204=>"111110000",
  58205=>"100101010",
  58206=>"001010100",
  58207=>"001010000",
  58208=>"111001000",
  58209=>"001010000",
  58210=>"010111111",
  58211=>"000101001",
  58212=>"001010001",
  58213=>"110101011",
  58214=>"100010000",
  58215=>"111110001",
  58216=>"000001011",
  58217=>"010101010",
  58218=>"001101011",
  58219=>"001000010",
  58220=>"001011101",
  58221=>"000011111",
  58222=>"011111010",
  58223=>"101111101",
  58224=>"011100010",
  58225=>"111111010",
  58226=>"101110110",
  58227=>"101011100",
  58228=>"111001011",
  58229=>"111111101",
  58230=>"100011010",
  58231=>"011000111",
  58232=>"110010111",
  58233=>"100110100",
  58234=>"100100000",
  58235=>"000011101",
  58236=>"100000110",
  58237=>"000010111",
  58238=>"100011010",
  58239=>"000100011",
  58240=>"110111101",
  58241=>"110000111",
  58242=>"001010101",
  58243=>"010111001",
  58244=>"100011110",
  58245=>"111111010",
  58246=>"111011011",
  58247=>"100110101",
  58248=>"111110100",
  58249=>"111100001",
  58250=>"001101101",
  58251=>"101111001",
  58252=>"100111111",
  58253=>"101000110",
  58254=>"111011101",
  58255=>"010000001",
  58256=>"110111111",
  58257=>"100010111",
  58258=>"000001100",
  58259=>"100000111",
  58260=>"000100011",
  58261=>"000011010",
  58262=>"110010101",
  58263=>"001110101",
  58264=>"100111111",
  58265=>"011010100",
  58266=>"010010001",
  58267=>"011110001",
  58268=>"111101110",
  58269=>"010000110",
  58270=>"011100111",
  58271=>"100110110",
  58272=>"000001110",
  58273=>"101101111",
  58274=>"111111111",
  58275=>"101101111",
  58276=>"101111110",
  58277=>"001101011",
  58278=>"000011100",
  58279=>"111101001",
  58280=>"111011111",
  58281=>"101010010",
  58282=>"010011110",
  58283=>"110101111",
  58284=>"111001100",
  58285=>"000010111",
  58286=>"010110110",
  58287=>"100011011",
  58288=>"111100111",
  58289=>"011111001",
  58290=>"001111111",
  58291=>"010010101",
  58292=>"011111110",
  58293=>"100000110",
  58294=>"011000110",
  58295=>"010110110",
  58296=>"000010110",
  58297=>"111000100",
  58298=>"010011110",
  58299=>"011100100",
  58300=>"100001101",
  58301=>"000110111",
  58302=>"111100110",
  58303=>"101000011",
  58304=>"100100001",
  58305=>"011100111",
  58306=>"100001011",
  58307=>"111100001",
  58308=>"000000100",
  58309=>"010101000",
  58310=>"111110011",
  58311=>"011101100",
  58312=>"000101010",
  58313=>"111010110",
  58314=>"000100111",
  58315=>"101101100",
  58316=>"101110001",
  58317=>"111111110",
  58318=>"011001100",
  58319=>"100110100",
  58320=>"110000000",
  58321=>"100001110",
  58322=>"010000000",
  58323=>"111010101",
  58324=>"000100100",
  58325=>"000100100",
  58326=>"001001110",
  58327=>"001011010",
  58328=>"111110100",
  58329=>"100000100",
  58330=>"110110100",
  58331=>"111011010",
  58332=>"000100001",
  58333=>"000101111",
  58334=>"011000010",
  58335=>"001000010",
  58336=>"101111100",
  58337=>"000111110",
  58338=>"100100101",
  58339=>"110011101",
  58340=>"000100000",
  58341=>"101011010",
  58342=>"000100010",
  58343=>"110100101",
  58344=>"000000000",
  58345=>"000011011",
  58346=>"100001011",
  58347=>"000010111",
  58348=>"011110110",
  58349=>"110001001",
  58350=>"111110101",
  58351=>"000101100",
  58352=>"000111111",
  58353=>"100110010",
  58354=>"000001100",
  58355=>"111001101",
  58356=>"000100000",
  58357=>"110101011",
  58358=>"101001000",
  58359=>"110111010",
  58360=>"111111010",
  58361=>"111110000",
  58362=>"101100010",
  58363=>"110000010",
  58364=>"001000010",
  58365=>"100101101",
  58366=>"101100000",
  58367=>"010100000",
  58368=>"010001011",
  58369=>"110101001",
  58370=>"100100010",
  58371=>"001100100",
  58372=>"010111010",
  58373=>"110101111",
  58374=>"100001001",
  58375=>"000000100",
  58376=>"001110111",
  58377=>"010011111",
  58378=>"011001100",
  58379=>"010001111",
  58380=>"000111100",
  58381=>"001001011",
  58382=>"000101001",
  58383=>"110011100",
  58384=>"001111100",
  58385=>"011011010",
  58386=>"111110100",
  58387=>"110101010",
  58388=>"000010111",
  58389=>"111011100",
  58390=>"001010100",
  58391=>"000001100",
  58392=>"111111000",
  58393=>"100000011",
  58394=>"001100110",
  58395=>"111000101",
  58396=>"010010000",
  58397=>"101100011",
  58398=>"010100110",
  58399=>"001110011",
  58400=>"101111010",
  58401=>"001111000",
  58402=>"101010101",
  58403=>"001011101",
  58404=>"110000001",
  58405=>"000000001",
  58406=>"001000101",
  58407=>"100001000",
  58408=>"100111111",
  58409=>"000100111",
  58410=>"011000001",
  58411=>"011000000",
  58412=>"101101101",
  58413=>"100001101",
  58414=>"110011001",
  58415=>"011011000",
  58416=>"010101101",
  58417=>"000001011",
  58418=>"011101111",
  58419=>"001101000",
  58420=>"110001101",
  58421=>"111111011",
  58422=>"011000011",
  58423=>"110110000",
  58424=>"111101011",
  58425=>"100110110",
  58426=>"010000001",
  58427=>"100001011",
  58428=>"011110011",
  58429=>"000111110",
  58430=>"110001011",
  58431=>"101000100",
  58432=>"101110101",
  58433=>"101110001",
  58434=>"010101001",
  58435=>"110010000",
  58436=>"001011010",
  58437=>"000000100",
  58438=>"011011110",
  58439=>"011111000",
  58440=>"100000111",
  58441=>"101010011",
  58442=>"100010110",
  58443=>"110010001",
  58444=>"100100000",
  58445=>"011011101",
  58446=>"100111011",
  58447=>"001000001",
  58448=>"000010100",
  58449=>"111101101",
  58450=>"110101100",
  58451=>"010011111",
  58452=>"111011110",
  58453=>"111110000",
  58454=>"101000000",
  58455=>"011010011",
  58456=>"110000110",
  58457=>"001111000",
  58458=>"100110110",
  58459=>"010111011",
  58460=>"011001011",
  58461=>"101100011",
  58462=>"111101110",
  58463=>"001000111",
  58464=>"011001101",
  58465=>"111101111",
  58466=>"001101000",
  58467=>"000001111",
  58468=>"101001001",
  58469=>"110100110",
  58470=>"111111110",
  58471=>"101000001",
  58472=>"110111011",
  58473=>"101111000",
  58474=>"100001110",
  58475=>"000101010",
  58476=>"101110111",
  58477=>"010111110",
  58478=>"011011011",
  58479=>"111011001",
  58480=>"000100011",
  58481=>"101110010",
  58482=>"111010110",
  58483=>"110001111",
  58484=>"110110000",
  58485=>"111111000",
  58486=>"100110000",
  58487=>"011111100",
  58488=>"001010010",
  58489=>"110001101",
  58490=>"101101100",
  58491=>"110111101",
  58492=>"110011100",
  58493=>"110101111",
  58494=>"100101001",
  58495=>"010111111",
  58496=>"101110000",
  58497=>"110011011",
  58498=>"001001111",
  58499=>"011101001",
  58500=>"000110100",
  58501=>"011010100",
  58502=>"001101011",
  58503=>"000110110",
  58504=>"000010110",
  58505=>"010110011",
  58506=>"000000001",
  58507=>"011000110",
  58508=>"111101011",
  58509=>"000101011",
  58510=>"111101101",
  58511=>"111000001",
  58512=>"001011100",
  58513=>"011011001",
  58514=>"010000011",
  58515=>"101010001",
  58516=>"110001000",
  58517=>"110110111",
  58518=>"111001010",
  58519=>"010110010",
  58520=>"000011111",
  58521=>"101010110",
  58522=>"010101010",
  58523=>"000101111",
  58524=>"110110000",
  58525=>"110011111",
  58526=>"001001000",
  58527=>"011111100",
  58528=>"010010010",
  58529=>"001011111",
  58530=>"101011111",
  58531=>"010110101",
  58532=>"001111011",
  58533=>"010101110",
  58534=>"110101110",
  58535=>"110010011",
  58536=>"001100000",
  58537=>"001001011",
  58538=>"111010100",
  58539=>"100100001",
  58540=>"100100111",
  58541=>"001010100",
  58542=>"100011011",
  58543=>"010010001",
  58544=>"100110010",
  58545=>"001101101",
  58546=>"110010011",
  58547=>"100101111",
  58548=>"011100010",
  58549=>"111100110",
  58550=>"100100010",
  58551=>"111111101",
  58552=>"011110001",
  58553=>"000101111",
  58554=>"110011011",
  58555=>"110101010",
  58556=>"010111001",
  58557=>"110011001",
  58558=>"000000010",
  58559=>"011101000",
  58560=>"101110000",
  58561=>"010111001",
  58562=>"000110101",
  58563=>"111110010",
  58564=>"100101111",
  58565=>"011101000",
  58566=>"111001000",
  58567=>"000110110",
  58568=>"000010001",
  58569=>"111101111",
  58570=>"111000110",
  58571=>"111011100",
  58572=>"000100011",
  58573=>"011110111",
  58574=>"001000111",
  58575=>"110101001",
  58576=>"111010111",
  58577=>"110111001",
  58578=>"011011111",
  58579=>"111100101",
  58580=>"110010001",
  58581=>"111111111",
  58582=>"001101001",
  58583=>"110010010",
  58584=>"010010110",
  58585=>"100000001",
  58586=>"110100110",
  58587=>"111101000",
  58588=>"001111100",
  58589=>"100001100",
  58590=>"101111011",
  58591=>"111001111",
  58592=>"111111101",
  58593=>"110110111",
  58594=>"101011000",
  58595=>"011101110",
  58596=>"110000001",
  58597=>"100110110",
  58598=>"000001000",
  58599=>"111111110",
  58600=>"100001010",
  58601=>"101111101",
  58602=>"101011000",
  58603=>"010100010",
  58604=>"000110010",
  58605=>"110010011",
  58606=>"010001000",
  58607=>"110111101",
  58608=>"000011000",
  58609=>"111111110",
  58610=>"111001000",
  58611=>"101001001",
  58612=>"010101100",
  58613=>"100001101",
  58614=>"000110110",
  58615=>"000010001",
  58616=>"000110100",
  58617=>"010100100",
  58618=>"000011111",
  58619=>"000100111",
  58620=>"000010101",
  58621=>"110000011",
  58622=>"011101101",
  58623=>"000001011",
  58624=>"110000000",
  58625=>"110101011",
  58626=>"010011110",
  58627=>"001010010",
  58628=>"101110111",
  58629=>"110010001",
  58630=>"011000101",
  58631=>"100001111",
  58632=>"010001101",
  58633=>"010110001",
  58634=>"010010001",
  58635=>"011100000",
  58636=>"101010010",
  58637=>"110100101",
  58638=>"001101010",
  58639=>"111110001",
  58640=>"110110001",
  58641=>"010000000",
  58642=>"111001001",
  58643=>"000011111",
  58644=>"011101000",
  58645=>"000100001",
  58646=>"010001011",
  58647=>"000100100",
  58648=>"100111011",
  58649=>"010100100",
  58650=>"011100000",
  58651=>"111011100",
  58652=>"011111010",
  58653=>"000100101",
  58654=>"110000101",
  58655=>"111010010",
  58656=>"101000000",
  58657=>"101100011",
  58658=>"001001001",
  58659=>"100101100",
  58660=>"110001100",
  58661=>"011100110",
  58662=>"110001101",
  58663=>"010011100",
  58664=>"011101011",
  58665=>"111100111",
  58666=>"011001011",
  58667=>"001111011",
  58668=>"000000001",
  58669=>"101110100",
  58670=>"001010000",
  58671=>"000100101",
  58672=>"001100011",
  58673=>"101100110",
  58674=>"001001001",
  58675=>"010010010",
  58676=>"000010011",
  58677=>"100110011",
  58678=>"100111001",
  58679=>"101111111",
  58680=>"110101110",
  58681=>"100010010",
  58682=>"111001110",
  58683=>"110011100",
  58684=>"011011101",
  58685=>"010101000",
  58686=>"100001010",
  58687=>"001011001",
  58688=>"111100111",
  58689=>"111110100",
  58690=>"101111010",
  58691=>"110010000",
  58692=>"100000100",
  58693=>"000011001",
  58694=>"110010010",
  58695=>"101001101",
  58696=>"111011001",
  58697=>"100101000",
  58698=>"110110001",
  58699=>"111000101",
  58700=>"110111111",
  58701=>"000110110",
  58702=>"100000100",
  58703=>"101100110",
  58704=>"010000010",
  58705=>"100110101",
  58706=>"001010000",
  58707=>"100101011",
  58708=>"000110110",
  58709=>"110111010",
  58710=>"110000000",
  58711=>"010100011",
  58712=>"101001010",
  58713=>"001011110",
  58714=>"001000010",
  58715=>"110111011",
  58716=>"101001011",
  58717=>"001100100",
  58718=>"111010000",
  58719=>"111101001",
  58720=>"000101100",
  58721=>"111011000",
  58722=>"110111001",
  58723=>"010111010",
  58724=>"010000110",
  58725=>"110000111",
  58726=>"000001101",
  58727=>"000110001",
  58728=>"101110001",
  58729=>"011101101",
  58730=>"100101101",
  58731=>"001001111",
  58732=>"011010110",
  58733=>"110111111",
  58734=>"101000100",
  58735=>"100000010",
  58736=>"011010100",
  58737=>"111101000",
  58738=>"001100111",
  58739=>"110100101",
  58740=>"011011101",
  58741=>"000111001",
  58742=>"101100000",
  58743=>"011100000",
  58744=>"001010110",
  58745=>"001110111",
  58746=>"111011010",
  58747=>"100001111",
  58748=>"110010110",
  58749=>"001100110",
  58750=>"111100101",
  58751=>"101011011",
  58752=>"111110010",
  58753=>"101010000",
  58754=>"001101101",
  58755=>"111111010",
  58756=>"010110100",
  58757=>"101110100",
  58758=>"001011000",
  58759=>"110100110",
  58760=>"000001010",
  58761=>"101111101",
  58762=>"000011100",
  58763=>"011010101",
  58764=>"111111111",
  58765=>"111010111",
  58766=>"101111111",
  58767=>"111000100",
  58768=>"111101110",
  58769=>"110110000",
  58770=>"011111001",
  58771=>"100101110",
  58772=>"010010001",
  58773=>"100100101",
  58774=>"110100110",
  58775=>"000101010",
  58776=>"011010011",
  58777=>"011010010",
  58778=>"001110000",
  58779=>"110101111",
  58780=>"010100110",
  58781=>"111100000",
  58782=>"001110001",
  58783=>"000110110",
  58784=>"001011001",
  58785=>"011110001",
  58786=>"001111000",
  58787=>"000001000",
  58788=>"011101110",
  58789=>"001000001",
  58790=>"000110100",
  58791=>"001111010",
  58792=>"010110111",
  58793=>"100111100",
  58794=>"100001001",
  58795=>"010001011",
  58796=>"111001000",
  58797=>"111111000",
  58798=>"011110000",
  58799=>"010001101",
  58800=>"100000100",
  58801=>"100010100",
  58802=>"110011011",
  58803=>"010011011",
  58804=>"010001100",
  58805=>"110111001",
  58806=>"011111010",
  58807=>"111111101",
  58808=>"000001001",
  58809=>"011110110",
  58810=>"011111111",
  58811=>"101111110",
  58812=>"011011010",
  58813=>"100000111",
  58814=>"100100110",
  58815=>"111001111",
  58816=>"010111010",
  58817=>"110100101",
  58818=>"011010110",
  58819=>"101011110",
  58820=>"010100010",
  58821=>"010010111",
  58822=>"111001111",
  58823=>"100011000",
  58824=>"100111010",
  58825=>"000000100",
  58826=>"101010010",
  58827=>"101011011",
  58828=>"110001100",
  58829=>"110011101",
  58830=>"011011111",
  58831=>"110011100",
  58832=>"111111110",
  58833=>"010101000",
  58834=>"100011001",
  58835=>"001101101",
  58836=>"000010100",
  58837=>"011001111",
  58838=>"100111011",
  58839=>"111010001",
  58840=>"110001100",
  58841=>"010011000",
  58842=>"110101001",
  58843=>"110111100",
  58844=>"100011011",
  58845=>"001101111",
  58846=>"101010001",
  58847=>"010000010",
  58848=>"001100110",
  58849=>"000101101",
  58850=>"110100010",
  58851=>"001101100",
  58852=>"101111101",
  58853=>"000001011",
  58854=>"010000111",
  58855=>"110100111",
  58856=>"000000000",
  58857=>"010110010",
  58858=>"110101100",
  58859=>"111000111",
  58860=>"010111101",
  58861=>"101001100",
  58862=>"000001010",
  58863=>"000001001",
  58864=>"000011000",
  58865=>"110100001",
  58866=>"000001000",
  58867=>"011101111",
  58868=>"111111011",
  58869=>"010011101",
  58870=>"100011100",
  58871=>"001101111",
  58872=>"110000100",
  58873=>"011101101",
  58874=>"111100100",
  58875=>"100011100",
  58876=>"010111010",
  58877=>"000100111",
  58878=>"011001001",
  58879=>"001011000",
  58880=>"001010100",
  58881=>"010111100",
  58882=>"110001100",
  58883=>"010000010",
  58884=>"110010010",
  58885=>"001011110",
  58886=>"010101111",
  58887=>"000010100",
  58888=>"101100110",
  58889=>"101011001",
  58890=>"111101011",
  58891=>"101110111",
  58892=>"100101100",
  58893=>"010010000",
  58894=>"110000001",
  58895=>"010010011",
  58896=>"110101111",
  58897=>"001101111",
  58898=>"100111111",
  58899=>"010011000",
  58900=>"010110100",
  58901=>"000100111",
  58902=>"010000110",
  58903=>"000101100",
  58904=>"101111111",
  58905=>"000110011",
  58906=>"110100011",
  58907=>"111001011",
  58908=>"010110011",
  58909=>"001110110",
  58910=>"010111010",
  58911=>"010011011",
  58912=>"101010000",
  58913=>"001101111",
  58914=>"101100000",
  58915=>"100100101",
  58916=>"000011011",
  58917=>"011101110",
  58918=>"101010010",
  58919=>"001110000",
  58920=>"111100000",
  58921=>"010000010",
  58922=>"011101111",
  58923=>"101111101",
  58924=>"101000110",
  58925=>"111000000",
  58926=>"111011100",
  58927=>"110110101",
  58928=>"011011110",
  58929=>"011101000",
  58930=>"101011001",
  58931=>"101100001",
  58932=>"110001011",
  58933=>"001100101",
  58934=>"011000100",
  58935=>"011100010",
  58936=>"100100010",
  58937=>"100110011",
  58938=>"101011111",
  58939=>"000000110",
  58940=>"110001111",
  58941=>"101011000",
  58942=>"011101111",
  58943=>"000101000",
  58944=>"100110100",
  58945=>"100011101",
  58946=>"001111011",
  58947=>"010111111",
  58948=>"111110111",
  58949=>"111101000",
  58950=>"101110001",
  58951=>"111011110",
  58952=>"110100010",
  58953=>"000111111",
  58954=>"011011010",
  58955=>"110011100",
  58956=>"110010011",
  58957=>"101110101",
  58958=>"001100101",
  58959=>"011111110",
  58960=>"100010000",
  58961=>"010010110",
  58962=>"101111101",
  58963=>"010001000",
  58964=>"001010010",
  58965=>"111011001",
  58966=>"110001100",
  58967=>"100101000",
  58968=>"100011101",
  58969=>"101011001",
  58970=>"000110011",
  58971=>"001101100",
  58972=>"011101011",
  58973=>"001000010",
  58974=>"101101011",
  58975=>"101011110",
  58976=>"010110111",
  58977=>"100101101",
  58978=>"001100110",
  58979=>"101010110",
  58980=>"100011111",
  58981=>"001010001",
  58982=>"000001011",
  58983=>"110011001",
  58984=>"001100111",
  58985=>"111101000",
  58986=>"010100010",
  58987=>"110110011",
  58988=>"001001100",
  58989=>"000100000",
  58990=>"001101010",
  58991=>"111101000",
  58992=>"010000111",
  58993=>"111110010",
  58994=>"110110100",
  58995=>"100010000",
  58996=>"011111001",
  58997=>"001101110",
  58998=>"110011110",
  58999=>"100000101",
  59000=>"001110001",
  59001=>"000000101",
  59002=>"101000000",
  59003=>"000011001",
  59004=>"110100000",
  59005=>"110011100",
  59006=>"011101001",
  59007=>"011101101",
  59008=>"010010101",
  59009=>"001001111",
  59010=>"100111000",
  59011=>"010001001",
  59012=>"010000011",
  59013=>"101101110",
  59014=>"010011111",
  59015=>"000010000",
  59016=>"100101011",
  59017=>"000000111",
  59018=>"001010001",
  59019=>"010101010",
  59020=>"001010011",
  59021=>"111111111",
  59022=>"101111111",
  59023=>"011110111",
  59024=>"100000110",
  59025=>"111010000",
  59026=>"111111101",
  59027=>"010111001",
  59028=>"001011100",
  59029=>"000000011",
  59030=>"101001101",
  59031=>"111110011",
  59032=>"110101101",
  59033=>"000101100",
  59034=>"101010010",
  59035=>"010000010",
  59036=>"011110010",
  59037=>"011001111",
  59038=>"100011000",
  59039=>"010111001",
  59040=>"101000000",
  59041=>"111110100",
  59042=>"111100111",
  59043=>"100101001",
  59044=>"110110100",
  59045=>"000111011",
  59046=>"011011010",
  59047=>"001110110",
  59048=>"011011001",
  59049=>"101100001",
  59050=>"011011110",
  59051=>"100111010",
  59052=>"010011101",
  59053=>"100101011",
  59054=>"100001010",
  59055=>"001111000",
  59056=>"101101111",
  59057=>"110111110",
  59058=>"101111110",
  59059=>"010110110",
  59060=>"000001111",
  59061=>"111101000",
  59062=>"011111101",
  59063=>"000111110",
  59064=>"111000001",
  59065=>"011100010",
  59066=>"010001110",
  59067=>"000010011",
  59068=>"111010100",
  59069=>"010101000",
  59070=>"111101001",
  59071=>"010101001",
  59072=>"001010111",
  59073=>"001001001",
  59074=>"100111000",
  59075=>"111111000",
  59076=>"111101110",
  59077=>"111011000",
  59078=>"000001111",
  59079=>"101001101",
  59080=>"001111010",
  59081=>"001010111",
  59082=>"111011010",
  59083=>"101000011",
  59084=>"100001010",
  59085=>"110110011",
  59086=>"100100111",
  59087=>"110011100",
  59088=>"000101101",
  59089=>"101000111",
  59090=>"110001101",
  59091=>"101110010",
  59092=>"111100010",
  59093=>"000100111",
  59094=>"110100001",
  59095=>"001000010",
  59096=>"000111101",
  59097=>"110111100",
  59098=>"000011101",
  59099=>"011101011",
  59100=>"011001111",
  59101=>"010101001",
  59102=>"100100000",
  59103=>"000110000",
  59104=>"011001010",
  59105=>"110111100",
  59106=>"010100100",
  59107=>"000010000",
  59108=>"010000101",
  59109=>"100110000",
  59110=>"101110000",
  59111=>"011001110",
  59112=>"111100101",
  59113=>"001001000",
  59114=>"001011010",
  59115=>"101000010",
  59116=>"011010000",
  59117=>"001111000",
  59118=>"000001110",
  59119=>"010111101",
  59120=>"011110001",
  59121=>"011110011",
  59122=>"010000001",
  59123=>"010101111",
  59124=>"100101111",
  59125=>"011111111",
  59126=>"001011111",
  59127=>"001010011",
  59128=>"011110011",
  59129=>"101010011",
  59130=>"100101111",
  59131=>"110011111",
  59132=>"010000111",
  59133=>"010010101",
  59134=>"111110110",
  59135=>"101111010",
  59136=>"111011100",
  59137=>"110000011",
  59138=>"010101100",
  59139=>"101000010",
  59140=>"110101010",
  59141=>"110111101",
  59142=>"000000001",
  59143=>"100101101",
  59144=>"010100001",
  59145=>"111100110",
  59146=>"010101101",
  59147=>"111000100",
  59148=>"100101100",
  59149=>"111110011",
  59150=>"110100110",
  59151=>"011011000",
  59152=>"000010110",
  59153=>"011010001",
  59154=>"011110111",
  59155=>"000000100",
  59156=>"111111000",
  59157=>"111110111",
  59158=>"111101011",
  59159=>"001011011",
  59160=>"101000001",
  59161=>"001111001",
  59162=>"101011000",
  59163=>"100100011",
  59164=>"001110101",
  59165=>"000001111",
  59166=>"101100101",
  59167=>"010111010",
  59168=>"010100010",
  59169=>"110110110",
  59170=>"110100010",
  59171=>"111111011",
  59172=>"000111111",
  59173=>"100010111",
  59174=>"111010000",
  59175=>"001011011",
  59176=>"111111010",
  59177=>"000101001",
  59178=>"001110011",
  59179=>"010010001",
  59180=>"110011011",
  59181=>"110100110",
  59182=>"111101001",
  59183=>"110111110",
  59184=>"011111010",
  59185=>"001001011",
  59186=>"001100110",
  59187=>"001000000",
  59188=>"001110000",
  59189=>"000100111",
  59190=>"011011011",
  59191=>"100101010",
  59192=>"000001100",
  59193=>"000111010",
  59194=>"110111010",
  59195=>"100000101",
  59196=>"110100101",
  59197=>"100000101",
  59198=>"010001110",
  59199=>"001010010",
  59200=>"000100100",
  59201=>"111100111",
  59202=>"100110010",
  59203=>"011100010",
  59204=>"111111101",
  59205=>"100111110",
  59206=>"110101111",
  59207=>"001110011",
  59208=>"101001011",
  59209=>"000011011",
  59210=>"001001111",
  59211=>"010100100",
  59212=>"111000000",
  59213=>"000011111",
  59214=>"110111110",
  59215=>"100110000",
  59216=>"111110011",
  59217=>"111100011",
  59218=>"000011101",
  59219=>"111100001",
  59220=>"101111011",
  59221=>"011011000",
  59222=>"010010011",
  59223=>"101110001",
  59224=>"100011101",
  59225=>"111010100",
  59226=>"111100011",
  59227=>"110111111",
  59228=>"110111000",
  59229=>"101101111",
  59230=>"111110001",
  59231=>"101011001",
  59232=>"110000000",
  59233=>"011111010",
  59234=>"111000000",
  59235=>"011000011",
  59236=>"011001001",
  59237=>"100110010",
  59238=>"001000101",
  59239=>"011110100",
  59240=>"000100011",
  59241=>"101111010",
  59242=>"111111010",
  59243=>"000101101",
  59244=>"101111111",
  59245=>"001111110",
  59246=>"011110111",
  59247=>"100101111",
  59248=>"000010100",
  59249=>"010000100",
  59250=>"111100110",
  59251=>"001111110",
  59252=>"100010100",
  59253=>"110110101",
  59254=>"110110110",
  59255=>"001110100",
  59256=>"011000101",
  59257=>"111001101",
  59258=>"011000010",
  59259=>"110111000",
  59260=>"000011000",
  59261=>"010100101",
  59262=>"111110100",
  59263=>"000000110",
  59264=>"001000101",
  59265=>"011100001",
  59266=>"010100010",
  59267=>"110100111",
  59268=>"011010101",
  59269=>"100110011",
  59270=>"011010000",
  59271=>"100101001",
  59272=>"001011110",
  59273=>"010101111",
  59274=>"010011000",
  59275=>"000111110",
  59276=>"000110110",
  59277=>"101111011",
  59278=>"001011100",
  59279=>"000001010",
  59280=>"100100101",
  59281=>"001110011",
  59282=>"110010110",
  59283=>"000111110",
  59284=>"010010111",
  59285=>"111011101",
  59286=>"111001000",
  59287=>"000001001",
  59288=>"110110101",
  59289=>"011001100",
  59290=>"010111101",
  59291=>"110010111",
  59292=>"101000011",
  59293=>"000001101",
  59294=>"100011000",
  59295=>"011011001",
  59296=>"000010101",
  59297=>"101010000",
  59298=>"010110111",
  59299=>"011100100",
  59300=>"011101111",
  59301=>"101110011",
  59302=>"100010000",
  59303=>"110110011",
  59304=>"011100000",
  59305=>"010001111",
  59306=>"010001111",
  59307=>"000100111",
  59308=>"100011110",
  59309=>"111010100",
  59310=>"000000100",
  59311=>"000111110",
  59312=>"100101011",
  59313=>"110000011",
  59314=>"100010100",
  59315=>"000001010",
  59316=>"001010010",
  59317=>"110011010",
  59318=>"101110100",
  59319=>"110110011",
  59320=>"000010000",
  59321=>"111000001",
  59322=>"010000100",
  59323=>"100001101",
  59324=>"000000011",
  59325=>"010100110",
  59326=>"011100011",
  59327=>"110101101",
  59328=>"110100110",
  59329=>"100001000",
  59330=>"100001010",
  59331=>"100100110",
  59332=>"111001111",
  59333=>"011010110",
  59334=>"001010111",
  59335=>"001101101",
  59336=>"110110001",
  59337=>"110111101",
  59338=>"000101011",
  59339=>"101000100",
  59340=>"010101001",
  59341=>"101010100",
  59342=>"110001110",
  59343=>"000011110",
  59344=>"011011000",
  59345=>"010100000",
  59346=>"111100000",
  59347=>"101000010",
  59348=>"110111111",
  59349=>"010011011",
  59350=>"110110011",
  59351=>"110001011",
  59352=>"001000010",
  59353=>"000010011",
  59354=>"101100001",
  59355=>"000100001",
  59356=>"001111111",
  59357=>"001101111",
  59358=>"011110110",
  59359=>"001010100",
  59360=>"001001101",
  59361=>"101101001",
  59362=>"000110111",
  59363=>"000011010",
  59364=>"110111100",
  59365=>"111111010",
  59366=>"111010001",
  59367=>"000000101",
  59368=>"101000100",
  59369=>"000111101",
  59370=>"100000011",
  59371=>"010000100",
  59372=>"001110110",
  59373=>"000101110",
  59374=>"010111100",
  59375=>"011100011",
  59376=>"001001111",
  59377=>"001110110",
  59378=>"110010000",
  59379=>"001000111",
  59380=>"101011111",
  59381=>"110101100",
  59382=>"110001001",
  59383=>"111001110",
  59384=>"110001000",
  59385=>"001100100",
  59386=>"111101000",
  59387=>"101010010",
  59388=>"101101111",
  59389=>"110000010",
  59390=>"101011101",
  59391=>"001101010",
  59392=>"100101100",
  59393=>"110000000",
  59394=>"000101011",
  59395=>"010011011",
  59396=>"010101110",
  59397=>"111011110",
  59398=>"000000011",
  59399=>"100101010",
  59400=>"011010110",
  59401=>"101000011",
  59402=>"000010110",
  59403=>"110111000",
  59404=>"000011011",
  59405=>"101001101",
  59406=>"111101111",
  59407=>"000110000",
  59408=>"110100010",
  59409=>"001110000",
  59410=>"000111111",
  59411=>"010101011",
  59412=>"100001011",
  59413=>"000110001",
  59414=>"110101110",
  59415=>"011001110",
  59416=>"011000001",
  59417=>"000111010",
  59418=>"111101100",
  59419=>"100111110",
  59420=>"100000000",
  59421=>"001001011",
  59422=>"110000000",
  59423=>"010000010",
  59424=>"101110100",
  59425=>"000001110",
  59426=>"010011000",
  59427=>"010011011",
  59428=>"000101111",
  59429=>"100100101",
  59430=>"100001100",
  59431=>"101111101",
  59432=>"010010111",
  59433=>"001001011",
  59434=>"011101000",
  59435=>"001011110",
  59436=>"101000011",
  59437=>"000011111",
  59438=>"111010111",
  59439=>"001101100",
  59440=>"000010110",
  59441=>"111001001",
  59442=>"101110011",
  59443=>"001000010",
  59444=>"110001111",
  59445=>"000010000",
  59446=>"010010110",
  59447=>"000010010",
  59448=>"110100100",
  59449=>"001110110",
  59450=>"011110110",
  59451=>"100101100",
  59452=>"000000010",
  59453=>"110111100",
  59454=>"100101111",
  59455=>"101011111",
  59456=>"111000001",
  59457=>"000000110",
  59458=>"010001010",
  59459=>"011000101",
  59460=>"010111010",
  59461=>"110000011",
  59462=>"001000100",
  59463=>"001000001",
  59464=>"111000111",
  59465=>"100100010",
  59466=>"110010010",
  59467=>"001000100",
  59468=>"001110100",
  59469=>"010101000",
  59470=>"100111011",
  59471=>"000110100",
  59472=>"111000001",
  59473=>"101000111",
  59474=>"101100011",
  59475=>"011001001",
  59476=>"100101101",
  59477=>"100000011",
  59478=>"011000110",
  59479=>"100101101",
  59480=>"000101011",
  59481=>"111001010",
  59482=>"001100011",
  59483=>"000000000",
  59484=>"010000010",
  59485=>"101110100",
  59486=>"111011100",
  59487=>"111000011",
  59488=>"011101000",
  59489=>"010111101",
  59490=>"010110011",
  59491=>"000011111",
  59492=>"000010110",
  59493=>"111100100",
  59494=>"011101110",
  59495=>"110001111",
  59496=>"011110101",
  59497=>"100000101",
  59498=>"100010111",
  59499=>"110010101",
  59500=>"000110001",
  59501=>"001101001",
  59502=>"101010011",
  59503=>"000010110",
  59504=>"100010110",
  59505=>"001011111",
  59506=>"000001000",
  59507=>"011010101",
  59508=>"111101011",
  59509=>"010111111",
  59510=>"110111101",
  59511=>"001100110",
  59512=>"000100000",
  59513=>"111101101",
  59514=>"001000101",
  59515=>"011000110",
  59516=>"010010001",
  59517=>"100110010",
  59518=>"111110000",
  59519=>"000100010",
  59520=>"100000110",
  59521=>"001110011",
  59522=>"100111011",
  59523=>"000111001",
  59524=>"000000100",
  59525=>"011110101",
  59526=>"001111001",
  59527=>"110000011",
  59528=>"110111111",
  59529=>"001100100",
  59530=>"001000001",
  59531=>"111110111",
  59532=>"100011010",
  59533=>"100011111",
  59534=>"100011111",
  59535=>"001100101",
  59536=>"010001000",
  59537=>"011101101",
  59538=>"100111001",
  59539=>"010111010",
  59540=>"101000000",
  59541=>"110101110",
  59542=>"101010110",
  59543=>"000000000",
  59544=>"011000111",
  59545=>"111101010",
  59546=>"101000000",
  59547=>"001000101",
  59548=>"101011111",
  59549=>"001001111",
  59550=>"111001001",
  59551=>"001001011",
  59552=>"000011010",
  59553=>"111111011",
  59554=>"011100001",
  59555=>"000111010",
  59556=>"011110111",
  59557=>"011101111",
  59558=>"001110101",
  59559=>"001001001",
  59560=>"110100000",
  59561=>"110000110",
  59562=>"011101010",
  59563=>"101010110",
  59564=>"110000010",
  59565=>"110101100",
  59566=>"001110010",
  59567=>"000100000",
  59568=>"111101100",
  59569=>"100111111",
  59570=>"011001110",
  59571=>"010101100",
  59572=>"000001101",
  59573=>"010011110",
  59574=>"100100000",
  59575=>"011001001",
  59576=>"101001101",
  59577=>"101100100",
  59578=>"111110110",
  59579=>"100101111",
  59580=>"000001101",
  59581=>"000001000",
  59582=>"000100010",
  59583=>"100111110",
  59584=>"000010110",
  59585=>"011100100",
  59586=>"011000111",
  59587=>"010000110",
  59588=>"001110101",
  59589=>"100101111",
  59590=>"001100011",
  59591=>"010110011",
  59592=>"101111110",
  59593=>"111010010",
  59594=>"000001011",
  59595=>"000011101",
  59596=>"111100110",
  59597=>"000110111",
  59598=>"111001000",
  59599=>"011111110",
  59600=>"010010001",
  59601=>"101110110",
  59602=>"010110010",
  59603=>"000101110",
  59604=>"111100001",
  59605=>"000110011",
  59606=>"111110100",
  59607=>"110011100",
  59608=>"110001001",
  59609=>"011011111",
  59610=>"100010101",
  59611=>"010010010",
  59612=>"011110000",
  59613=>"011110110",
  59614=>"100100010",
  59615=>"001111011",
  59616=>"000000011",
  59617=>"111010111",
  59618=>"110111100",
  59619=>"001111111",
  59620=>"101110110",
  59621=>"101011000",
  59622=>"000110010",
  59623=>"001001101",
  59624=>"011110000",
  59625=>"111101011",
  59626=>"000111001",
  59627=>"001011101",
  59628=>"000011011",
  59629=>"001010000",
  59630=>"111101010",
  59631=>"001001001",
  59632=>"010000001",
  59633=>"100000101",
  59634=>"001110101",
  59635=>"001011111",
  59636=>"100111110",
  59637=>"000011000",
  59638=>"111010011",
  59639=>"000011010",
  59640=>"010011111",
  59641=>"011001000",
  59642=>"010100110",
  59643=>"101010010",
  59644=>"000100101",
  59645=>"000000100",
  59646=>"100111111",
  59647=>"101110111",
  59648=>"111110010",
  59649=>"011111000",
  59650=>"011101100",
  59651=>"101101111",
  59652=>"111101111",
  59653=>"011000110",
  59654=>"110001110",
  59655=>"001111101",
  59656=>"111011001",
  59657=>"111100000",
  59658=>"010011010",
  59659=>"110000010",
  59660=>"111100001",
  59661=>"010011011",
  59662=>"110110000",
  59663=>"100000111",
  59664=>"001011010",
  59665=>"110110011",
  59666=>"000111011",
  59667=>"111101100",
  59668=>"111000110",
  59669=>"111101111",
  59670=>"011000100",
  59671=>"011000110",
  59672=>"110000000",
  59673=>"010000111",
  59674=>"001001111",
  59675=>"111000111",
  59676=>"000000011",
  59677=>"010001100",
  59678=>"100100010",
  59679=>"000111001",
  59680=>"100111110",
  59681=>"011001111",
  59682=>"000110010",
  59683=>"000011001",
  59684=>"101101011",
  59685=>"101111010",
  59686=>"010000000",
  59687=>"010000011",
  59688=>"111111101",
  59689=>"011000001",
  59690=>"011001101",
  59691=>"100110011",
  59692=>"000111001",
  59693=>"001000000",
  59694=>"001010011",
  59695=>"010011011",
  59696=>"111111111",
  59697=>"111011101",
  59698=>"110001101",
  59699=>"010010001",
  59700=>"010001111",
  59701=>"001000011",
  59702=>"001011100",
  59703=>"101111110",
  59704=>"101111111",
  59705=>"101011001",
  59706=>"001000100",
  59707=>"110111001",
  59708=>"011010100",
  59709=>"110101111",
  59710=>"110001010",
  59711=>"111101101",
  59712=>"101011001",
  59713=>"111110010",
  59714=>"010011101",
  59715=>"010000010",
  59716=>"010100001",
  59717=>"101111110",
  59718=>"001010001",
  59719=>"101101101",
  59720=>"011000011",
  59721=>"001000000",
  59722=>"011001110",
  59723=>"000011011",
  59724=>"001011100",
  59725=>"101110101",
  59726=>"000001110",
  59727=>"110001001",
  59728=>"001011001",
  59729=>"111011000",
  59730=>"010110010",
  59731=>"010010000",
  59732=>"111100101",
  59733=>"010000011",
  59734=>"001100010",
  59735=>"101000001",
  59736=>"111010100",
  59737=>"110100001",
  59738=>"100000001",
  59739=>"011101110",
  59740=>"000101110",
  59741=>"000111001",
  59742=>"101001010",
  59743=>"101110111",
  59744=>"011101101",
  59745=>"111000111",
  59746=>"010010000",
  59747=>"010000000",
  59748=>"101111110",
  59749=>"101011000",
  59750=>"011111111",
  59751=>"011111101",
  59752=>"111100100",
  59753=>"000010001",
  59754=>"001001110",
  59755=>"101001001",
  59756=>"000000000",
  59757=>"011000000",
  59758=>"100001011",
  59759=>"111101111",
  59760=>"000100010",
  59761=>"110111110",
  59762=>"011000000",
  59763=>"111101111",
  59764=>"110100010",
  59765=>"010100111",
  59766=>"001001111",
  59767=>"000000101",
  59768=>"111011011",
  59769=>"000011100",
  59770=>"000011111",
  59771=>"111101000",
  59772=>"111010010",
  59773=>"010100101",
  59774=>"010011000",
  59775=>"010101011",
  59776=>"010110110",
  59777=>"000000000",
  59778=>"001010010",
  59779=>"011111000",
  59780=>"110011001",
  59781=>"100001111",
  59782=>"011011010",
  59783=>"110110010",
  59784=>"110101011",
  59785=>"101100010",
  59786=>"001110111",
  59787=>"110010011",
  59788=>"010010001",
  59789=>"111111011",
  59790=>"000010000",
  59791=>"011111101",
  59792=>"001010100",
  59793=>"000001101",
  59794=>"010101000",
  59795=>"111100111",
  59796=>"101110111",
  59797=>"010010000",
  59798=>"000000010",
  59799=>"101100100",
  59800=>"111101111",
  59801=>"100000001",
  59802=>"110001000",
  59803=>"010010111",
  59804=>"111111110",
  59805=>"000111010",
  59806=>"010000000",
  59807=>"111100100",
  59808=>"110101010",
  59809=>"000001100",
  59810=>"110111100",
  59811=>"000010010",
  59812=>"110010000",
  59813=>"101111000",
  59814=>"011111101",
  59815=>"110110101",
  59816=>"100000110",
  59817=>"111110000",
  59818=>"110000000",
  59819=>"111010101",
  59820=>"001010110",
  59821=>"010110100",
  59822=>"111000000",
  59823=>"110100010",
  59824=>"001111001",
  59825=>"010010111",
  59826=>"001011000",
  59827=>"011011101",
  59828=>"111001110",
  59829=>"010110100",
  59830=>"111111001",
  59831=>"010111111",
  59832=>"111110001",
  59833=>"000101011",
  59834=>"101101100",
  59835=>"100111010",
  59836=>"011010010",
  59837=>"010010101",
  59838=>"111001000",
  59839=>"100011011",
  59840=>"010101000",
  59841=>"000110001",
  59842=>"001111010",
  59843=>"111001001",
  59844=>"101010000",
  59845=>"000001100",
  59846=>"111101001",
  59847=>"000101110",
  59848=>"001001000",
  59849=>"001010110",
  59850=>"001000100",
  59851=>"111011111",
  59852=>"100100000",
  59853=>"100011110",
  59854=>"001001010",
  59855=>"001111101",
  59856=>"000110111",
  59857=>"010100110",
  59858=>"010000100",
  59859=>"111101100",
  59860=>"000010110",
  59861=>"000111100",
  59862=>"100110111",
  59863=>"000011111",
  59864=>"111000101",
  59865=>"101110011",
  59866=>"000111100",
  59867=>"110011110",
  59868=>"100001000",
  59869=>"101111111",
  59870=>"101011101",
  59871=>"110011000",
  59872=>"010101111",
  59873=>"010101101",
  59874=>"111011000",
  59875=>"001000010",
  59876=>"010101100",
  59877=>"110010111",
  59878=>"000110011",
  59879=>"001110101",
  59880=>"001010100",
  59881=>"000111000",
  59882=>"011000011",
  59883=>"000111000",
  59884=>"000101110",
  59885=>"001010010",
  59886=>"000000000",
  59887=>"111001100",
  59888=>"010100111",
  59889=>"111011010",
  59890=>"001110100",
  59891=>"100110100",
  59892=>"100010011",
  59893=>"100111010",
  59894=>"001111001",
  59895=>"100010100",
  59896=>"100101000",
  59897=>"111000101",
  59898=>"111001000",
  59899=>"101010000",
  59900=>"111000101",
  59901=>"101111011",
  59902=>"000111000",
  59903=>"001100000",
  59904=>"001111110",
  59905=>"110000110",
  59906=>"100011110",
  59907=>"110011010",
  59908=>"111101110",
  59909=>"100000000",
  59910=>"101110000",
  59911=>"001010000",
  59912=>"110010001",
  59913=>"010100000",
  59914=>"001110110",
  59915=>"110010010",
  59916=>"010101110",
  59917=>"010000110",
  59918=>"001001000",
  59919=>"101000111",
  59920=>"111111001",
  59921=>"011100101",
  59922=>"110000110",
  59923=>"110101011",
  59924=>"100110110",
  59925=>"100011100",
  59926=>"101010010",
  59927=>"010010000",
  59928=>"011001010",
  59929=>"001101101",
  59930=>"000000000",
  59931=>"010111100",
  59932=>"110001011",
  59933=>"100010111",
  59934=>"111100111",
  59935=>"101001111",
  59936=>"001000011",
  59937=>"111010100",
  59938=>"000000111",
  59939=>"001010110",
  59940=>"100101010",
  59941=>"100000011",
  59942=>"101001001",
  59943=>"111111000",
  59944=>"111010010",
  59945=>"101010000",
  59946=>"101110011",
  59947=>"110101101",
  59948=>"100011001",
  59949=>"000001000",
  59950=>"101000001",
  59951=>"010110000",
  59952=>"000101000",
  59953=>"000100011",
  59954=>"001011111",
  59955=>"101000111",
  59956=>"101110100",
  59957=>"011100101",
  59958=>"110000011",
  59959=>"001110101",
  59960=>"100110110",
  59961=>"010110001",
  59962=>"101000000",
  59963=>"111000001",
  59964=>"001100000",
  59965=>"000001111",
  59966=>"000010010",
  59967=>"001011010",
  59968=>"010000110",
  59969=>"011011100",
  59970=>"000110000",
  59971=>"101101111",
  59972=>"000111010",
  59973=>"111111010",
  59974=>"000100100",
  59975=>"011011010",
  59976=>"010011110",
  59977=>"010101111",
  59978=>"011010010",
  59979=>"101001010",
  59980=>"101000001",
  59981=>"110001011",
  59982=>"000010000",
  59983=>"100010100",
  59984=>"000100000",
  59985=>"110010100",
  59986=>"110111111",
  59987=>"010001011",
  59988=>"010111101",
  59989=>"110010000",
  59990=>"101001101",
  59991=>"100110100",
  59992=>"111111101",
  59993=>"010010010",
  59994=>"110001010",
  59995=>"011111011",
  59996=>"101100111",
  59997=>"100001100",
  59998=>"010101001",
  59999=>"111101010",
  60000=>"011100001",
  60001=>"010010000",
  60002=>"010010001",
  60003=>"011111110",
  60004=>"101110100",
  60005=>"111101001",
  60006=>"000111001",
  60007=>"001001010",
  60008=>"000101101",
  60009=>"111111100",
  60010=>"001101010",
  60011=>"110001000",
  60012=>"001011000",
  60013=>"100100001",
  60014=>"001101101",
  60015=>"010110000",
  60016=>"111101000",
  60017=>"110110011",
  60018=>"101110110",
  60019=>"000001101",
  60020=>"000011001",
  60021=>"010100000",
  60022=>"101001011",
  60023=>"000000000",
  60024=>"111100101",
  60025=>"011010011",
  60026=>"110111110",
  60027=>"001011111",
  60028=>"101110100",
  60029=>"001101010",
  60030=>"100001111",
  60031=>"000100110",
  60032=>"100110110",
  60033=>"000101100",
  60034=>"000110101",
  60035=>"000001101",
  60036=>"010100101",
  60037=>"111011000",
  60038=>"100011100",
  60039=>"001100011",
  60040=>"111000001",
  60041=>"010101001",
  60042=>"110000100",
  60043=>"001100011",
  60044=>"011000110",
  60045=>"111011001",
  60046=>"011010011",
  60047=>"111100010",
  60048=>"010101001",
  60049=>"111000010",
  60050=>"001010111",
  60051=>"010111100",
  60052=>"101011111",
  60053=>"000110010",
  60054=>"111001110",
  60055=>"100110111",
  60056=>"011110011",
  60057=>"111111001",
  60058=>"010011110",
  60059=>"110111101",
  60060=>"100110001",
  60061=>"011011101",
  60062=>"110111110",
  60063=>"000001000",
  60064=>"110101100",
  60065=>"011001000",
  60066=>"110101010",
  60067=>"101000010",
  60068=>"000100001",
  60069=>"111101000",
  60070=>"101100000",
  60071=>"000011101",
  60072=>"000111111",
  60073=>"010001001",
  60074=>"010101011",
  60075=>"101100100",
  60076=>"010100011",
  60077=>"010001010",
  60078=>"010111111",
  60079=>"100110000",
  60080=>"000111111",
  60081=>"101110000",
  60082=>"011110010",
  60083=>"011110111",
  60084=>"011001001",
  60085=>"111111111",
  60086=>"010000010",
  60087=>"001101011",
  60088=>"010100100",
  60089=>"101000000",
  60090=>"110111011",
  60091=>"100101100",
  60092=>"010001110",
  60093=>"001110100",
  60094=>"011101000",
  60095=>"011001010",
  60096=>"101111000",
  60097=>"101100101",
  60098=>"100110010",
  60099=>"011010111",
  60100=>"100010001",
  60101=>"001000101",
  60102=>"000000010",
  60103=>"010010100",
  60104=>"101101010",
  60105=>"110010001",
  60106=>"111110001",
  60107=>"110010100",
  60108=>"000100010",
  60109=>"010000101",
  60110=>"100101101",
  60111=>"011011100",
  60112=>"101001100",
  60113=>"011011011",
  60114=>"011111100",
  60115=>"101100100",
  60116=>"101001110",
  60117=>"011000011",
  60118=>"101000000",
  60119=>"100001001",
  60120=>"110000000",
  60121=>"101101110",
  60122=>"110111101",
  60123=>"101001001",
  60124=>"111110100",
  60125=>"001001111",
  60126=>"111111110",
  60127=>"000100000",
  60128=>"111100111",
  60129=>"110000111",
  60130=>"101100001",
  60131=>"000100101",
  60132=>"011110111",
  60133=>"111011110",
  60134=>"010101000",
  60135=>"000100011",
  60136=>"010110000",
  60137=>"111101001",
  60138=>"011001000",
  60139=>"111001001",
  60140=>"000001101",
  60141=>"001100000",
  60142=>"101101111",
  60143=>"011110010",
  60144=>"000010010",
  60145=>"010000011",
  60146=>"001100101",
  60147=>"101011111",
  60148=>"010100101",
  60149=>"010011110",
  60150=>"110010001",
  60151=>"101101011",
  60152=>"001011011",
  60153=>"010110111",
  60154=>"111110110",
  60155=>"100000001",
  60156=>"011110111",
  60157=>"001001000",
  60158=>"001000110",
  60159=>"101100000",
  60160=>"101100000",
  60161=>"110101000",
  60162=>"111100001",
  60163=>"000101111",
  60164=>"100011110",
  60165=>"101100111",
  60166=>"010111110",
  60167=>"011101101",
  60168=>"100110010",
  60169=>"000110000",
  60170=>"011000110",
  60171=>"011111101",
  60172=>"010110001",
  60173=>"011011100",
  60174=>"001111000",
  60175=>"100001100",
  60176=>"101101101",
  60177=>"101100111",
  60178=>"010010000",
  60179=>"011101101",
  60180=>"001110100",
  60181=>"011101111",
  60182=>"001110001",
  60183=>"100010011",
  60184=>"100110110",
  60185=>"000001100",
  60186=>"001100001",
  60187=>"011000001",
  60188=>"010100101",
  60189=>"000100001",
  60190=>"001111111",
  60191=>"000111100",
  60192=>"001000000",
  60193=>"101111100",
  60194=>"000000001",
  60195=>"001010011",
  60196=>"100010110",
  60197=>"000000010",
  60198=>"101001010",
  60199=>"001001101",
  60200=>"010010010",
  60201=>"101000100",
  60202=>"111111111",
  60203=>"111001000",
  60204=>"010000000",
  60205=>"001110011",
  60206=>"001111101",
  60207=>"011110011",
  60208=>"101011010",
  60209=>"111111011",
  60210=>"011000110",
  60211=>"001110010",
  60212=>"111001101",
  60213=>"111000000",
  60214=>"100000010",
  60215=>"001011011",
  60216=>"100000100",
  60217=>"011001110",
  60218=>"101101011",
  60219=>"111110111",
  60220=>"010111000",
  60221=>"110111111",
  60222=>"101110001",
  60223=>"100100101",
  60224=>"111010110",
  60225=>"000000110",
  60226=>"101101000",
  60227=>"010011010",
  60228=>"100111111",
  60229=>"011111000",
  60230=>"100100001",
  60231=>"101111010",
  60232=>"000011000",
  60233=>"100010111",
  60234=>"110110011",
  60235=>"000000000",
  60236=>"011000011",
  60237=>"101001010",
  60238=>"101100010",
  60239=>"001100101",
  60240=>"100101110",
  60241=>"010000000",
  60242=>"000110011",
  60243=>"101001100",
  60244=>"110100111",
  60245=>"010111111",
  60246=>"100001011",
  60247=>"110101001",
  60248=>"110111101",
  60249=>"111011010",
  60250=>"111110111",
  60251=>"010000100",
  60252=>"101110101",
  60253=>"001000011",
  60254=>"000110101",
  60255=>"000010000",
  60256=>"110101001",
  60257=>"000111111",
  60258=>"111100100",
  60259=>"010010110",
  60260=>"111010110",
  60261=>"111010110",
  60262=>"000100011",
  60263=>"111101111",
  60264=>"001000100",
  60265=>"000101000",
  60266=>"010011100",
  60267=>"011000110",
  60268=>"000011111",
  60269=>"110111111",
  60270=>"010110000",
  60271=>"000100010",
  60272=>"011000110",
  60273=>"111101101",
  60274=>"101011010",
  60275=>"110100111",
  60276=>"101110100",
  60277=>"101100000",
  60278=>"011100001",
  60279=>"001011111",
  60280=>"111110010",
  60281=>"001000111",
  60282=>"001011111",
  60283=>"001001010",
  60284=>"010010100",
  60285=>"001000011",
  60286=>"010000000",
  60287=>"000101111",
  60288=>"010010011",
  60289=>"011000010",
  60290=>"110001100",
  60291=>"101101111",
  60292=>"110000010",
  60293=>"000101010",
  60294=>"111111100",
  60295=>"000111010",
  60296=>"011100110",
  60297=>"100111010",
  60298=>"000010111",
  60299=>"110101111",
  60300=>"111110100",
  60301=>"111110010",
  60302=>"110000010",
  60303=>"000001100",
  60304=>"011000100",
  60305=>"010001111",
  60306=>"010100000",
  60307=>"100000001",
  60308=>"000111101",
  60309=>"111011101",
  60310=>"001001101",
  60311=>"100110101",
  60312=>"111011110",
  60313=>"000110000",
  60314=>"010010000",
  60315=>"101111110",
  60316=>"100111000",
  60317=>"111101101",
  60318=>"001001010",
  60319=>"001010011",
  60320=>"010110100",
  60321=>"111010100",
  60322=>"001000010",
  60323=>"001101011",
  60324=>"001111000",
  60325=>"101011000",
  60326=>"011111000",
  60327=>"001111001",
  60328=>"010001000",
  60329=>"011011011",
  60330=>"101001001",
  60331=>"100101011",
  60332=>"100011010",
  60333=>"100100001",
  60334=>"101100111",
  60335=>"010011101",
  60336=>"111111111",
  60337=>"011011100",
  60338=>"011100110",
  60339=>"111010110",
  60340=>"011101100",
  60341=>"100100001",
  60342=>"110101001",
  60343=>"111100000",
  60344=>"111101001",
  60345=>"001101101",
  60346=>"100010110",
  60347=>"100010111",
  60348=>"101100010",
  60349=>"010100010",
  60350=>"010110111",
  60351=>"011111000",
  60352=>"100101001",
  60353=>"100001010",
  60354=>"111011001",
  60355=>"000010011",
  60356=>"010000011",
  60357=>"100000001",
  60358=>"100000110",
  60359=>"111101111",
  60360=>"010010110",
  60361=>"010010001",
  60362=>"110111111",
  60363=>"001001100",
  60364=>"010110111",
  60365=>"100010110",
  60366=>"011011100",
  60367=>"001111010",
  60368=>"000010011",
  60369=>"100101101",
  60370=>"111111011",
  60371=>"101010010",
  60372=>"100110101",
  60373=>"100111100",
  60374=>"001100111",
  60375=>"001011001",
  60376=>"101101111",
  60377=>"110110111",
  60378=>"100101011",
  60379=>"101010000",
  60380=>"000111101",
  60381=>"100011101",
  60382=>"011111000",
  60383=>"111110011",
  60384=>"100110100",
  60385=>"111011000",
  60386=>"110000000",
  60387=>"000100010",
  60388=>"010111001",
  60389=>"000000000",
  60390=>"101010111",
  60391=>"111101000",
  60392=>"110111111",
  60393=>"100101001",
  60394=>"011010111",
  60395=>"111111100",
  60396=>"001001101",
  60397=>"110111011",
  60398=>"100111101",
  60399=>"000110000",
  60400=>"111100111",
  60401=>"110110100",
  60402=>"111110111",
  60403=>"111010011",
  60404=>"110110101",
  60405=>"001010000",
  60406=>"101001100",
  60407=>"010111000",
  60408=>"010100110",
  60409=>"111001001",
  60410=>"100001000",
  60411=>"101000000",
  60412=>"101100111",
  60413=>"000100000",
  60414=>"111001000",
  60415=>"010100100",
  60416=>"101000001",
  60417=>"001100001",
  60418=>"010001001",
  60419=>"100110111",
  60420=>"100111111",
  60421=>"100100101",
  60422=>"101000011",
  60423=>"111111101",
  60424=>"010011111",
  60425=>"101111101",
  60426=>"111100011",
  60427=>"000100001",
  60428=>"110101101",
  60429=>"111111101",
  60430=>"110010100",
  60431=>"011110010",
  60432=>"100010101",
  60433=>"010111010",
  60434=>"010111011",
  60435=>"101100001",
  60436=>"000111111",
  60437=>"001111001",
  60438=>"000001111",
  60439=>"101110000",
  60440=>"110001010",
  60441=>"010001001",
  60442=>"011110101",
  60443=>"101111100",
  60444=>"100011010",
  60445=>"000100101",
  60446=>"110111100",
  60447=>"110010010",
  60448=>"101101100",
  60449=>"111010101",
  60450=>"010111011",
  60451=>"101110001",
  60452=>"011111000",
  60453=>"011010000",
  60454=>"011110001",
  60455=>"110101011",
  60456=>"110000100",
  60457=>"001010010",
  60458=>"111110101",
  60459=>"000100101",
  60460=>"001000111",
  60461=>"110100110",
  60462=>"100111010",
  60463=>"111111010",
  60464=>"001001100",
  60465=>"010011101",
  60466=>"100101000",
  60467=>"010001011",
  60468=>"111011101",
  60469=>"011111010",
  60470=>"000101100",
  60471=>"000101111",
  60472=>"101101001",
  60473=>"000010100",
  60474=>"101100001",
  60475=>"001111111",
  60476=>"010110100",
  60477=>"111010100",
  60478=>"001111000",
  60479=>"111101110",
  60480=>"110000111",
  60481=>"100011110",
  60482=>"111111111",
  60483=>"111100001",
  60484=>"110111010",
  60485=>"110000101",
  60486=>"000011101",
  60487=>"111111100",
  60488=>"011000111",
  60489=>"100011100",
  60490=>"111000110",
  60491=>"000101000",
  60492=>"101110110",
  60493=>"000111011",
  60494=>"110100001",
  60495=>"000010000",
  60496=>"101100011",
  60497=>"100010100",
  60498=>"010101111",
  60499=>"010110101",
  60500=>"000000110",
  60501=>"101000101",
  60502=>"101011101",
  60503=>"001010011",
  60504=>"110000101",
  60505=>"001010011",
  60506=>"001111001",
  60507=>"111111010",
  60508=>"101101110",
  60509=>"001000101",
  60510=>"101010111",
  60511=>"111111100",
  60512=>"111001000",
  60513=>"000001001",
  60514=>"011111000",
  60515=>"101011101",
  60516=>"100001111",
  60517=>"111001000",
  60518=>"100000100",
  60519=>"000000101",
  60520=>"001111101",
  60521=>"011100010",
  60522=>"001100100",
  60523=>"001101101",
  60524=>"011100101",
  60525=>"100011001",
  60526=>"010101011",
  60527=>"001111111",
  60528=>"101010101",
  60529=>"111011101",
  60530=>"001010001",
  60531=>"100110100",
  60532=>"110001010",
  60533=>"101110001",
  60534=>"101100010",
  60535=>"100110101",
  60536=>"000101111",
  60537=>"101000010",
  60538=>"111100100",
  60539=>"110111110",
  60540=>"101100110",
  60541=>"101111100",
  60542=>"010011101",
  60543=>"100001001",
  60544=>"011001000",
  60545=>"000000011",
  60546=>"010100011",
  60547=>"011010101",
  60548=>"011110110",
  60549=>"111000011",
  60550=>"101100000",
  60551=>"110001011",
  60552=>"000000010",
  60553=>"100100011",
  60554=>"101111100",
  60555=>"101000000",
  60556=>"100100100",
  60557=>"100001010",
  60558=>"010011010",
  60559=>"000111111",
  60560=>"101000111",
  60561=>"000010111",
  60562=>"010001011",
  60563=>"111000011",
  60564=>"111001100",
  60565=>"100001110",
  60566=>"111010101",
  60567=>"111001111",
  60568=>"110000011",
  60569=>"000000001",
  60570=>"001001010",
  60571=>"110001010",
  60572=>"001000110",
  60573=>"101110100",
  60574=>"000011001",
  60575=>"010000001",
  60576=>"100111100",
  60577=>"110011001",
  60578=>"011110001",
  60579=>"111000111",
  60580=>"010101001",
  60581=>"110011001",
  60582=>"010001001",
  60583=>"001110101",
  60584=>"101101110",
  60585=>"011100000",
  60586=>"101001001",
  60587=>"011000110",
  60588=>"001110011",
  60589=>"111001110",
  60590=>"100000111",
  60591=>"011010001",
  60592=>"110000100",
  60593=>"110000011",
  60594=>"010111001",
  60595=>"001011011",
  60596=>"011110111",
  60597=>"000110001",
  60598=>"111010001",
  60599=>"101111011",
  60600=>"111011110",
  60601=>"101101111",
  60602=>"111110110",
  60603=>"000100011",
  60604=>"000001000",
  60605=>"010011110",
  60606=>"000000101",
  60607=>"110111110",
  60608=>"100110111",
  60609=>"110100111",
  60610=>"001101010",
  60611=>"100101010",
  60612=>"010010010",
  60613=>"110011001",
  60614=>"100010111",
  60615=>"010101000",
  60616=>"001000111",
  60617=>"110010100",
  60618=>"110100000",
  60619=>"000001001",
  60620=>"100110000",
  60621=>"001111010",
  60622=>"110110110",
  60623=>"101100011",
  60624=>"111111111",
  60625=>"100110011",
  60626=>"011001101",
  60627=>"101101110",
  60628=>"010110111",
  60629=>"001111000",
  60630=>"000111101",
  60631=>"001000011",
  60632=>"110111111",
  60633=>"010110111",
  60634=>"100111011",
  60635=>"001000110",
  60636=>"111010010",
  60637=>"000011101",
  60638=>"101101011",
  60639=>"100000100",
  60640=>"111111111",
  60641=>"001000101",
  60642=>"010110010",
  60643=>"110101111",
  60644=>"011000100",
  60645=>"011110111",
  60646=>"000100000",
  60647=>"011001101",
  60648=>"111011100",
  60649=>"110101011",
  60650=>"001011010",
  60651=>"101010001",
  60652=>"010111001",
  60653=>"111110111",
  60654=>"011000010",
  60655=>"010000000",
  60656=>"010011000",
  60657=>"010111100",
  60658=>"100110001",
  60659=>"111101011",
  60660=>"110011000",
  60661=>"011010110",
  60662=>"100010000",
  60663=>"101101100",
  60664=>"000100100",
  60665=>"010100011",
  60666=>"010110111",
  60667=>"001011110",
  60668=>"010111100",
  60669=>"111101000",
  60670=>"110000010",
  60671=>"100111100",
  60672=>"101100101",
  60673=>"001111111",
  60674=>"000010110",
  60675=>"011111100",
  60676=>"010100000",
  60677=>"000100010",
  60678=>"001110111",
  60679=>"100100000",
  60680=>"110100111",
  60681=>"101110110",
  60682=>"001010000",
  60683=>"111101011",
  60684=>"110101110",
  60685=>"011101001",
  60686=>"000111001",
  60687=>"011111001",
  60688=>"111011000",
  60689=>"001110110",
  60690=>"101000011",
  60691=>"101111000",
  60692=>"000101010",
  60693=>"111101001",
  60694=>"101101011",
  60695=>"111110010",
  60696=>"100110100",
  60697=>"010011111",
  60698=>"101010000",
  60699=>"111111001",
  60700=>"000011111",
  60701=>"011001010",
  60702=>"111100101",
  60703=>"100000001",
  60704=>"101100011",
  60705=>"111101001",
  60706=>"111110110",
  60707=>"101110010",
  60708=>"111100001",
  60709=>"010101110",
  60710=>"010111000",
  60711=>"111100101",
  60712=>"011010011",
  60713=>"111111100",
  60714=>"110100110",
  60715=>"011010110",
  60716=>"011010100",
  60717=>"100111111",
  60718=>"011100010",
  60719=>"010101001",
  60720=>"100100110",
  60721=>"110110010",
  60722=>"110101111",
  60723=>"100110111",
  60724=>"000110110",
  60725=>"011111110",
  60726=>"000000101",
  60727=>"100001001",
  60728=>"110100111",
  60729=>"101100111",
  60730=>"101101011",
  60731=>"100100100",
  60732=>"111100000",
  60733=>"011010110",
  60734=>"111010111",
  60735=>"001001010",
  60736=>"100100101",
  60737=>"111000011",
  60738=>"110111011",
  60739=>"100110111",
  60740=>"000100001",
  60741=>"111000111",
  60742=>"111011100",
  60743=>"000100101",
  60744=>"111010010",
  60745=>"010101010",
  60746=>"001001101",
  60747=>"100011100",
  60748=>"001000011",
  60749=>"010110000",
  60750=>"001011000",
  60751=>"100100110",
  60752=>"001111001",
  60753=>"110110110",
  60754=>"000110110",
  60755=>"000100101",
  60756=>"010011101",
  60757=>"010001111",
  60758=>"100001110",
  60759=>"100010001",
  60760=>"101101010",
  60761=>"101010100",
  60762=>"010101101",
  60763=>"011110100",
  60764=>"000010000",
  60765=>"111100000",
  60766=>"111010010",
  60767=>"000000110",
  60768=>"010101000",
  60769=>"101011001",
  60770=>"110110001",
  60771=>"100001100",
  60772=>"010111010",
  60773=>"001110111",
  60774=>"011101010",
  60775=>"101000010",
  60776=>"001010001",
  60777=>"001111111",
  60778=>"111000111",
  60779=>"101100010",
  60780=>"010011011",
  60781=>"110111010",
  60782=>"111101111",
  60783=>"000010001",
  60784=>"001100011",
  60785=>"111111100",
  60786=>"011010011",
  60787=>"001010110",
  60788=>"011011011",
  60789=>"001011001",
  60790=>"001010111",
  60791=>"111100100",
  60792=>"111010011",
  60793=>"000101110",
  60794=>"110101100",
  60795=>"001100011",
  60796=>"011000000",
  60797=>"110011111",
  60798=>"000000110",
  60799=>"001001111",
  60800=>"000101101",
  60801=>"110000011",
  60802=>"101111110",
  60803=>"111111110",
  60804=>"000101111",
  60805=>"001111011",
  60806=>"000000011",
  60807=>"010000001",
  60808=>"111101111",
  60809=>"100001001",
  60810=>"111010011",
  60811=>"101111001",
  60812=>"111111111",
  60813=>"001010101",
  60814=>"101100011",
  60815=>"101001111",
  60816=>"000101110",
  60817=>"100101111",
  60818=>"101111111",
  60819=>"000111111",
  60820=>"010101101",
  60821=>"110111000",
  60822=>"111010110",
  60823=>"001010101",
  60824=>"000101001",
  60825=>"110001111",
  60826=>"000001011",
  60827=>"101111111",
  60828=>"111110011",
  60829=>"100100011",
  60830=>"001010111",
  60831=>"101010011",
  60832=>"111010101",
  60833=>"111111111",
  60834=>"100010100",
  60835=>"001011100",
  60836=>"011111110",
  60837=>"111111101",
  60838=>"101100000",
  60839=>"010110111",
  60840=>"000101110",
  60841=>"001111111",
  60842=>"101001001",
  60843=>"111010111",
  60844=>"001011001",
  60845=>"110110111",
  60846=>"001010010",
  60847=>"011011010",
  60848=>"001111000",
  60849=>"110000111",
  60850=>"011010110",
  60851=>"101111011",
  60852=>"111101001",
  60853=>"000001111",
  60854=>"011100011",
  60855=>"100011110",
  60856=>"010001101",
  60857=>"000100100",
  60858=>"100110110",
  60859=>"111111001",
  60860=>"111110010",
  60861=>"010001110",
  60862=>"000001111",
  60863=>"100011111",
  60864=>"110110100",
  60865=>"100100001",
  60866=>"001011011",
  60867=>"110011101",
  60868=>"011011000",
  60869=>"110001000",
  60870=>"110110001",
  60871=>"001101110",
  60872=>"110101000",
  60873=>"100001110",
  60874=>"110010011",
  60875=>"101101010",
  60876=>"000101100",
  60877=>"101010100",
  60878=>"101101100",
  60879=>"110110010",
  60880=>"011011011",
  60881=>"011110110",
  60882=>"100011010",
  60883=>"000101010",
  60884=>"000011101",
  60885=>"111001001",
  60886=>"111111110",
  60887=>"101010010",
  60888=>"011100000",
  60889=>"011000100",
  60890=>"110110111",
  60891=>"100001101",
  60892=>"110011110",
  60893=>"000100111",
  60894=>"111101101",
  60895=>"001010111",
  60896=>"010101010",
  60897=>"001000111",
  60898=>"010010101",
  60899=>"011101011",
  60900=>"011000000",
  60901=>"000001011",
  60902=>"011011011",
  60903=>"111111111",
  60904=>"110011110",
  60905=>"010100101",
  60906=>"010011100",
  60907=>"100001100",
  60908=>"011001101",
  60909=>"110101100",
  60910=>"101111111",
  60911=>"100100111",
  60912=>"011110100",
  60913=>"001111000",
  60914=>"100101010",
  60915=>"100011111",
  60916=>"011100011",
  60917=>"010010011",
  60918=>"011110110",
  60919=>"010000110",
  60920=>"111010100",
  60921=>"011101111",
  60922=>"100110010",
  60923=>"111111101",
  60924=>"000001000",
  60925=>"011111101",
  60926=>"111001000",
  60927=>"001101001",
  60928=>"001011100",
  60929=>"100010001",
  60930=>"101000001",
  60931=>"111011111",
  60932=>"101111001",
  60933=>"111010001",
  60934=>"001100001",
  60935=>"010111110",
  60936=>"011101110",
  60937=>"110101011",
  60938=>"000000100",
  60939=>"011111010",
  60940=>"100001111",
  60941=>"101111111",
  60942=>"001000010",
  60943=>"101010000",
  60944=>"000000001",
  60945=>"011011000",
  60946=>"000000010",
  60947=>"010101100",
  60948=>"110010110",
  60949=>"100110111",
  60950=>"110000010",
  60951=>"001100011",
  60952=>"001011110",
  60953=>"100000110",
  60954=>"100011011",
  60955=>"010000011",
  60956=>"001110101",
  60957=>"101111101",
  60958=>"100111111",
  60959=>"000100000",
  60960=>"011001001",
  60961=>"001111100",
  60962=>"111110101",
  60963=>"100010100",
  60964=>"101011101",
  60965=>"101101110",
  60966=>"100001000",
  60967=>"111110111",
  60968=>"011100000",
  60969=>"110101101",
  60970=>"111001100",
  60971=>"110001010",
  60972=>"010111010",
  60973=>"100010110",
  60974=>"000101111",
  60975=>"111110010",
  60976=>"011000000",
  60977=>"000101111",
  60978=>"010010111",
  60979=>"011011001",
  60980=>"110101001",
  60981=>"011001100",
  60982=>"100100011",
  60983=>"100011111",
  60984=>"111000100",
  60985=>"100001011",
  60986=>"011011000",
  60987=>"110000110",
  60988=>"010101101",
  60989=>"110010111",
  60990=>"100111010",
  60991=>"000000010",
  60992=>"011100001",
  60993=>"101110111",
  60994=>"100000011",
  60995=>"000100000",
  60996=>"011000110",
  60997=>"110100010",
  60998=>"101010110",
  60999=>"111110110",
  61000=>"110111110",
  61001=>"100111001",
  61002=>"010001101",
  61003=>"011101100",
  61004=>"111111011",
  61005=>"101111101",
  61006=>"001000001",
  61007=>"101111011",
  61008=>"011001010",
  61009=>"100010000",
  61010=>"101111111",
  61011=>"010100100",
  61012=>"000101100",
  61013=>"011011001",
  61014=>"101111111",
  61015=>"111100010",
  61016=>"010110101",
  61017=>"110100011",
  61018=>"110010010",
  61019=>"100001001",
  61020=>"001000100",
  61021=>"000101011",
  61022=>"010100100",
  61023=>"111110001",
  61024=>"011110110",
  61025=>"111010011",
  61026=>"001110000",
  61027=>"110010010",
  61028=>"001000100",
  61029=>"001011001",
  61030=>"110101011",
  61031=>"100101101",
  61032=>"110111111",
  61033=>"001010011",
  61034=>"001101011",
  61035=>"001011110",
  61036=>"111010110",
  61037=>"000100000",
  61038=>"010010010",
  61039=>"000001001",
  61040=>"100111101",
  61041=>"111011100",
  61042=>"010011101",
  61043=>"100000101",
  61044=>"001101110",
  61045=>"101100011",
  61046=>"101100101",
  61047=>"001000101",
  61048=>"101110001",
  61049=>"000000000",
  61050=>"011001000",
  61051=>"000010011",
  61052=>"011100111",
  61053=>"111011000",
  61054=>"101111101",
  61055=>"000100110",
  61056=>"111110101",
  61057=>"001011011",
  61058=>"011111100",
  61059=>"101001010",
  61060=>"101001111",
  61061=>"101000001",
  61062=>"011011101",
  61063=>"001100000",
  61064=>"001001100",
  61065=>"110111010",
  61066=>"110101001",
  61067=>"001100100",
  61068=>"111110010",
  61069=>"001100011",
  61070=>"001111111",
  61071=>"110100100",
  61072=>"101001001",
  61073=>"101000001",
  61074=>"111110110",
  61075=>"001000100",
  61076=>"100101010",
  61077=>"100000110",
  61078=>"011000100",
  61079=>"100010110",
  61080=>"011100010",
  61081=>"011011001",
  61082=>"010110000",
  61083=>"011011010",
  61084=>"011010010",
  61085=>"010010011",
  61086=>"111100000",
  61087=>"100111100",
  61088=>"001010011",
  61089=>"001001001",
  61090=>"100001000",
  61091=>"111111011",
  61092=>"100000011",
  61093=>"101100100",
  61094=>"111000110",
  61095=>"101010111",
  61096=>"110101000",
  61097=>"101011100",
  61098=>"100101111",
  61099=>"111010101",
  61100=>"111110100",
  61101=>"101011111",
  61102=>"010110011",
  61103=>"000000011",
  61104=>"110100010",
  61105=>"101101111",
  61106=>"111111001",
  61107=>"010100111",
  61108=>"000011011",
  61109=>"101101101",
  61110=>"001111101",
  61111=>"000100010",
  61112=>"111110100",
  61113=>"011111100",
  61114=>"000100001",
  61115=>"000101000",
  61116=>"111010110",
  61117=>"011011111",
  61118=>"100101111",
  61119=>"101000100",
  61120=>"110101101",
  61121=>"010001000",
  61122=>"010101001",
  61123=>"110111110",
  61124=>"000010010",
  61125=>"101000101",
  61126=>"001011011",
  61127=>"011010011",
  61128=>"110011010",
  61129=>"110000000",
  61130=>"000110111",
  61131=>"100010111",
  61132=>"001010000",
  61133=>"110011110",
  61134=>"101011110",
  61135=>"111011101",
  61136=>"001000000",
  61137=>"011100111",
  61138=>"001100010",
  61139=>"000100111",
  61140=>"101111100",
  61141=>"111010000",
  61142=>"011011010",
  61143=>"111000011",
  61144=>"001011110",
  61145=>"011000110",
  61146=>"111111101",
  61147=>"110010011",
  61148=>"111011110",
  61149=>"011001000",
  61150=>"111101100",
  61151=>"011110100",
  61152=>"101100011",
  61153=>"001100111",
  61154=>"010010110",
  61155=>"000000011",
  61156=>"100111001",
  61157=>"000000101",
  61158=>"101101010",
  61159=>"000110000",
  61160=>"111111100",
  61161=>"010100001",
  61162=>"000011101",
  61163=>"001010000",
  61164=>"010001010",
  61165=>"001111110",
  61166=>"001101011",
  61167=>"111111101",
  61168=>"111111110",
  61169=>"000111000",
  61170=>"011111101",
  61171=>"001011011",
  61172=>"111011001",
  61173=>"010010011",
  61174=>"111111001",
  61175=>"101000001",
  61176=>"110101001",
  61177=>"010111100",
  61178=>"111111001",
  61179=>"110001110",
  61180=>"111110011",
  61181=>"100011100",
  61182=>"110101111",
  61183=>"101110000",
  61184=>"010011010",
  61185=>"111001111",
  61186=>"010000101",
  61187=>"011110001",
  61188=>"100000011",
  61189=>"100100100",
  61190=>"000011101",
  61191=>"101100101",
  61192=>"000101110",
  61193=>"011001100",
  61194=>"010011101",
  61195=>"001100010",
  61196=>"111110101",
  61197=>"010000100",
  61198=>"100000101",
  61199=>"100000101",
  61200=>"111000111",
  61201=>"000011101",
  61202=>"001100111",
  61203=>"101101001",
  61204=>"000101011",
  61205=>"101010001",
  61206=>"100011010",
  61207=>"000000000",
  61208=>"000110111",
  61209=>"000110010",
  61210=>"011001000",
  61211=>"110110111",
  61212=>"001001001",
  61213=>"010010110",
  61214=>"101100111",
  61215=>"001101000",
  61216=>"111010111",
  61217=>"011011110",
  61218=>"101101000",
  61219=>"111100111",
  61220=>"111111111",
  61221=>"000100010",
  61222=>"000010000",
  61223=>"010010000",
  61224=>"010101111",
  61225=>"001001100",
  61226=>"110001000",
  61227=>"111101110",
  61228=>"011000100",
  61229=>"101110011",
  61230=>"010100000",
  61231=>"001011000",
  61232=>"000010010",
  61233=>"110000011",
  61234=>"100111111",
  61235=>"101011011",
  61236=>"100010111",
  61237=>"100111110",
  61238=>"101011101",
  61239=>"001001111",
  61240=>"101111010",
  61241=>"101000101",
  61242=>"011000001",
  61243=>"010110001",
  61244=>"110111010",
  61245=>"110011010",
  61246=>"110010011",
  61247=>"000011110",
  61248=>"101111110",
  61249=>"110110100",
  61250=>"001100010",
  61251=>"101011011",
  61252=>"010100111",
  61253=>"110011010",
  61254=>"011011000",
  61255=>"000100000",
  61256=>"000001001",
  61257=>"000000010",
  61258=>"111001110",
  61259=>"100000010",
  61260=>"100100101",
  61261=>"000100010",
  61262=>"100100101",
  61263=>"001101010",
  61264=>"010001110",
  61265=>"101010001",
  61266=>"000000001",
  61267=>"101111011",
  61268=>"001001000",
  61269=>"111000001",
  61270=>"110110110",
  61271=>"000100111",
  61272=>"100011001",
  61273=>"010010001",
  61274=>"110110111",
  61275=>"111001001",
  61276=>"100111110",
  61277=>"111111000",
  61278=>"100011000",
  61279=>"111110111",
  61280=>"111101010",
  61281=>"111001011",
  61282=>"011011001",
  61283=>"011000100",
  61284=>"100100001",
  61285=>"111110111",
  61286=>"010101111",
  61287=>"100011111",
  61288=>"011010000",
  61289=>"111100111",
  61290=>"101100010",
  61291=>"011101101",
  61292=>"011001011",
  61293=>"001110111",
  61294=>"111110110",
  61295=>"000111111",
  61296=>"111101101",
  61297=>"110010100",
  61298=>"011000001",
  61299=>"001010111",
  61300=>"101001111",
  61301=>"110110110",
  61302=>"101111011",
  61303=>"110101011",
  61304=>"111100001",
  61305=>"010011101",
  61306=>"100000010",
  61307=>"001001110",
  61308=>"100100111",
  61309=>"010100001",
  61310=>"011100100",
  61311=>"010110010",
  61312=>"000111111",
  61313=>"110110000",
  61314=>"100110101",
  61315=>"100001000",
  61316=>"011100010",
  61317=>"011101100",
  61318=>"010100100",
  61319=>"111111110",
  61320=>"010011100",
  61321=>"111111100",
  61322=>"111111111",
  61323=>"000001011",
  61324=>"100111010",
  61325=>"110010010",
  61326=>"001100001",
  61327=>"100000010",
  61328=>"010011111",
  61329=>"000000000",
  61330=>"101001010",
  61331=>"101001010",
  61332=>"010111000",
  61333=>"111000010",
  61334=>"111110111",
  61335=>"000001111",
  61336=>"011000000",
  61337=>"000001010",
  61338=>"000110110",
  61339=>"100000110",
  61340=>"111000000",
  61341=>"010110111",
  61342=>"000111111",
  61343=>"101100111",
  61344=>"001110100",
  61345=>"100111010",
  61346=>"001010111",
  61347=>"011111101",
  61348=>"111110111",
  61349=>"000011100",
  61350=>"000111011",
  61351=>"101110000",
  61352=>"011101000",
  61353=>"101011100",
  61354=>"000101010",
  61355=>"101100001",
  61356=>"111000101",
  61357=>"000000101",
  61358=>"001101000",
  61359=>"100001001",
  61360=>"000000001",
  61361=>"101110111",
  61362=>"011010000",
  61363=>"000011001",
  61364=>"010111000",
  61365=>"110010001",
  61366=>"001000000",
  61367=>"110100011",
  61368=>"100000010",
  61369=>"000011001",
  61370=>"000010110",
  61371=>"010101001",
  61372=>"111111110",
  61373=>"111101011",
  61374=>"110111111",
  61375=>"111000001",
  61376=>"011110110",
  61377=>"111010011",
  61378=>"101101111",
  61379=>"010110100",
  61380=>"101111110",
  61381=>"111011000",
  61382=>"100101101",
  61383=>"011010001",
  61384=>"101111100",
  61385=>"111111100",
  61386=>"101000010",
  61387=>"110101111",
  61388=>"001111010",
  61389=>"010010111",
  61390=>"100111111",
  61391=>"101000011",
  61392=>"101100011",
  61393=>"111010100",
  61394=>"101111000",
  61395=>"011011100",
  61396=>"111010011",
  61397=>"010000011",
  61398=>"001000111",
  61399=>"110111101",
  61400=>"000010101",
  61401=>"000000110",
  61402=>"111010000",
  61403=>"110101010",
  61404=>"111111010",
  61405=>"111100011",
  61406=>"100110010",
  61407=>"000001100",
  61408=>"011101101",
  61409=>"110001101",
  61410=>"110011010",
  61411=>"111010001",
  61412=>"110001110",
  61413=>"100000101",
  61414=>"101100010",
  61415=>"111100111",
  61416=>"110111011",
  61417=>"010111110",
  61418=>"111101100",
  61419=>"111100101",
  61420=>"101110100",
  61421=>"000011010",
  61422=>"110110111",
  61423=>"011000101",
  61424=>"010100100",
  61425=>"100101000",
  61426=>"111000111",
  61427=>"000110110",
  61428=>"010001001",
  61429=>"111111110",
  61430=>"011110110",
  61431=>"111110011",
  61432=>"100010010",
  61433=>"001001001",
  61434=>"010100001",
  61435=>"111001000",
  61436=>"010101100",
  61437=>"010010011",
  61438=>"111000100",
  61439=>"111101011",
  61440=>"110001000",
  61441=>"110000010",
  61442=>"101111111",
  61443=>"001010110",
  61444=>"000010000",
  61445=>"001000110",
  61446=>"110000100",
  61447=>"011100000",
  61448=>"010101101",
  61449=>"101010011",
  61450=>"010011000",
  61451=>"011110110",
  61452=>"000011100",
  61453=>"000111011",
  61454=>"000011101",
  61455=>"000110110",
  61456=>"110101100",
  61457=>"100100010",
  61458=>"000100010",
  61459=>"111101001",
  61460=>"100110000",
  61461=>"110111011",
  61462=>"111100111",
  61463=>"011001001",
  61464=>"110000011",
  61465=>"010010100",
  61466=>"010110101",
  61467=>"000111010",
  61468=>"001011110",
  61469=>"111000010",
  61470=>"100100000",
  61471=>"000000101",
  61472=>"111011101",
  61473=>"011010101",
  61474=>"001001110",
  61475=>"001001000",
  61476=>"101100001",
  61477=>"011010101",
  61478=>"100101011",
  61479=>"010000101",
  61480=>"110100010",
  61481=>"000110010",
  61482=>"100101100",
  61483=>"001000000",
  61484=>"010111110",
  61485=>"110110101",
  61486=>"001100010",
  61487=>"101110110",
  61488=>"001101110",
  61489=>"100000011",
  61490=>"001001001",
  61491=>"010011000",
  61492=>"011011100",
  61493=>"010000111",
  61494=>"110000111",
  61495=>"010100100",
  61496=>"101101010",
  61497=>"001010001",
  61498=>"110010000",
  61499=>"101111000",
  61500=>"000010100",
  61501=>"000100000",
  61502=>"010011100",
  61503=>"000100010",
  61504=>"000011011",
  61505=>"110111000",
  61506=>"111111000",
  61507=>"111110101",
  61508=>"100011111",
  61509=>"011100011",
  61510=>"000111101",
  61511=>"101010100",
  61512=>"111001011",
  61513=>"101100101",
  61514=>"110000001",
  61515=>"010101001",
  61516=>"010011000",
  61517=>"100011000",
  61518=>"010000011",
  61519=>"001011110",
  61520=>"111101001",
  61521=>"001110011",
  61522=>"000110110",
  61523=>"001101000",
  61524=>"000101100",
  61525=>"100000000",
  61526=>"101110110",
  61527=>"111101111",
  61528=>"110111010",
  61529=>"100001100",
  61530=>"011100000",
  61531=>"000010010",
  61532=>"110111111",
  61533=>"111111010",
  61534=>"100001110",
  61535=>"110011101",
  61536=>"000001101",
  61537=>"110001110",
  61538=>"000100101",
  61539=>"110001100",
  61540=>"101110001",
  61541=>"010011111",
  61542=>"101101111",
  61543=>"100010100",
  61544=>"010110111",
  61545=>"111101111",
  61546=>"100001100",
  61547=>"101000100",
  61548=>"100111011",
  61549=>"110101001",
  61550=>"110010001",
  61551=>"110111110",
  61552=>"100001001",
  61553=>"010110010",
  61554=>"110100110",
  61555=>"000101100",
  61556=>"101000101",
  61557=>"100110000",
  61558=>"101110010",
  61559=>"101010100",
  61560=>"110111111",
  61561=>"000010011",
  61562=>"010110010",
  61563=>"001001111",
  61564=>"110011100",
  61565=>"010001010",
  61566=>"100000001",
  61567=>"011111001",
  61568=>"111011011",
  61569=>"001100111",
  61570=>"011101000",
  61571=>"100000010",
  61572=>"101100110",
  61573=>"011111101",
  61574=>"010100011",
  61575=>"100100100",
  61576=>"111110111",
  61577=>"101110111",
  61578=>"011100100",
  61579=>"110010110",
  61580=>"100101110",
  61581=>"001100111",
  61582=>"010111111",
  61583=>"000001011",
  61584=>"101101100",
  61585=>"110111111",
  61586=>"010000101",
  61587=>"000111010",
  61588=>"001001010",
  61589=>"101111000",
  61590=>"010101001",
  61591=>"000100000",
  61592=>"000100110",
  61593=>"100100000",
  61594=>"111001000",
  61595=>"110011011",
  61596=>"101011111",
  61597=>"001001110",
  61598=>"010011111",
  61599=>"000001001",
  61600=>"000101101",
  61601=>"110100011",
  61602=>"111001111",
  61603=>"011100001",
  61604=>"111010101",
  61605=>"110101001",
  61606=>"010010010",
  61607=>"111001110",
  61608=>"000101001",
  61609=>"110111111",
  61610=>"010101010",
  61611=>"101101101",
  61612=>"100111100",
  61613=>"100100010",
  61614=>"100010000",
  61615=>"111101110",
  61616=>"011111000",
  61617=>"000100110",
  61618=>"111000100",
  61619=>"010100100",
  61620=>"000101101",
  61621=>"010010101",
  61622=>"001101000",
  61623=>"010000101",
  61624=>"101001010",
  61625=>"111001111",
  61626=>"110100011",
  61627=>"110000011",
  61628=>"100011111",
  61629=>"011101001",
  61630=>"001011000",
  61631=>"000000000",
  61632=>"100101001",
  61633=>"101111111",
  61634=>"001110111",
  61635=>"000110100",
  61636=>"010100110",
  61637=>"101010011",
  61638=>"110011010",
  61639=>"001100101",
  61640=>"001010000",
  61641=>"001100000",
  61642=>"111111100",
  61643=>"001101000",
  61644=>"010001011",
  61645=>"100111011",
  61646=>"001001000",
  61647=>"000000110",
  61648=>"100110101",
  61649=>"110010001",
  61650=>"111101001",
  61651=>"101011000",
  61652=>"101000100",
  61653=>"010110111",
  61654=>"000010101",
  61655=>"110000111",
  61656=>"010011110",
  61657=>"000110011",
  61658=>"011000101",
  61659=>"101000111",
  61660=>"100001000",
  61661=>"000011110",
  61662=>"001011101",
  61663=>"110101001",
  61664=>"101001000",
  61665=>"000010110",
  61666=>"010001100",
  61667=>"001001010",
  61668=>"111011101",
  61669=>"101010101",
  61670=>"011100010",
  61671=>"111010100",
  61672=>"111111010",
  61673=>"000010101",
  61674=>"000000110",
  61675=>"000010101",
  61676=>"101110011",
  61677=>"010111010",
  61678=>"011111001",
  61679=>"001110111",
  61680=>"111111110",
  61681=>"100010001",
  61682=>"101100101",
  61683=>"100011001",
  61684=>"100101000",
  61685=>"011001000",
  61686=>"010100010",
  61687=>"001111010",
  61688=>"100101110",
  61689=>"000011101",
  61690=>"011111001",
  61691=>"011001100",
  61692=>"010000001",
  61693=>"100100010",
  61694=>"101000001",
  61695=>"100011111",
  61696=>"100010011",
  61697=>"101011100",
  61698=>"110011111",
  61699=>"000000100",
  61700=>"010011101",
  61701=>"011000100",
  61702=>"111000110",
  61703=>"111011000",
  61704=>"111000001",
  61705=>"111110000",
  61706=>"000010010",
  61707=>"110001110",
  61708=>"110000010",
  61709=>"100000110",
  61710=>"111101110",
  61711=>"101001111",
  61712=>"011011111",
  61713=>"101110101",
  61714=>"001001000",
  61715=>"111111000",
  61716=>"011111011",
  61717=>"001100110",
  61718=>"100100010",
  61719=>"000000001",
  61720=>"110011010",
  61721=>"101110000",
  61722=>"111110100",
  61723=>"100011101",
  61724=>"110100101",
  61725=>"100101101",
  61726=>"101101011",
  61727=>"100001010",
  61728=>"100001111",
  61729=>"111100010",
  61730=>"011010001",
  61731=>"010101110",
  61732=>"001100010",
  61733=>"000100110",
  61734=>"010100000",
  61735=>"000001101",
  61736=>"000111011",
  61737=>"000100010",
  61738=>"001100100",
  61739=>"000011000",
  61740=>"110110110",
  61741=>"010000011",
  61742=>"001100101",
  61743=>"101011010",
  61744=>"110011001",
  61745=>"110011010",
  61746=>"001101101",
  61747=>"010001011",
  61748=>"011010010",
  61749=>"011000110",
  61750=>"000010001",
  61751=>"110010001",
  61752=>"101101111",
  61753=>"011100011",
  61754=>"001010111",
  61755=>"101111010",
  61756=>"000101011",
  61757=>"001011100",
  61758=>"000100010",
  61759=>"000011101",
  61760=>"011010110",
  61761=>"010001011",
  61762=>"111011000",
  61763=>"110101001",
  61764=>"101101011",
  61765=>"100000101",
  61766=>"100100010",
  61767=>"000011000",
  61768=>"101000100",
  61769=>"000001001",
  61770=>"000011100",
  61771=>"101100110",
  61772=>"101111001",
  61773=>"111110000",
  61774=>"100010110",
  61775=>"101000111",
  61776=>"000010000",
  61777=>"100101101",
  61778=>"000101001",
  61779=>"111101011",
  61780=>"010001100",
  61781=>"111001111",
  61782=>"100000010",
  61783=>"001101010",
  61784=>"010000010",
  61785=>"011000010",
  61786=>"000100001",
  61787=>"010010001",
  61788=>"011110111",
  61789=>"001110100",
  61790=>"110110100",
  61791=>"001110010",
  61792=>"101111110",
  61793=>"101100110",
  61794=>"000110111",
  61795=>"010100000",
  61796=>"111011111",
  61797=>"000011000",
  61798=>"100101101",
  61799=>"011011111",
  61800=>"110010110",
  61801=>"101000010",
  61802=>"000011010",
  61803=>"111100100",
  61804=>"000010001",
  61805=>"010101000",
  61806=>"100011000",
  61807=>"011101111",
  61808=>"011111011",
  61809=>"101000011",
  61810=>"011101010",
  61811=>"111010000",
  61812=>"001111110",
  61813=>"110101001",
  61814=>"111101010",
  61815=>"110100110",
  61816=>"100010010",
  61817=>"001011111",
  61818=>"011000101",
  61819=>"010010110",
  61820=>"100110110",
  61821=>"101111001",
  61822=>"111110001",
  61823=>"111100001",
  61824=>"011101001",
  61825=>"010010101",
  61826=>"100111110",
  61827=>"110101100",
  61828=>"111011010",
  61829=>"100101100",
  61830=>"110010110",
  61831=>"000110100",
  61832=>"110001100",
  61833=>"010010110",
  61834=>"101000100",
  61835=>"111010011",
  61836=>"101100010",
  61837=>"001111000",
  61838=>"010011011",
  61839=>"010111011",
  61840=>"110101111",
  61841=>"111111100",
  61842=>"101001100",
  61843=>"001100001",
  61844=>"111010001",
  61845=>"100110111",
  61846=>"011110010",
  61847=>"111011100",
  61848=>"101111100",
  61849=>"000101111",
  61850=>"100011110",
  61851=>"011011011",
  61852=>"101011010",
  61853=>"000110100",
  61854=>"111001110",
  61855=>"011110111",
  61856=>"110100010",
  61857=>"110100000",
  61858=>"110100010",
  61859=>"111001100",
  61860=>"101110010",
  61861=>"000000101",
  61862=>"101000001",
  61863=>"011011100",
  61864=>"010111001",
  61865=>"111000010",
  61866=>"101001100",
  61867=>"101110000",
  61868=>"010110101",
  61869=>"000110011",
  61870=>"010000100",
  61871=>"010110111",
  61872=>"011111001",
  61873=>"010010101",
  61874=>"000011100",
  61875=>"100101010",
  61876=>"001111100",
  61877=>"011111000",
  61878=>"110010001",
  61879=>"101011010",
  61880=>"100000000",
  61881=>"010000001",
  61882=>"100000010",
  61883=>"111000111",
  61884=>"100101000",
  61885=>"011110011",
  61886=>"100110011",
  61887=>"111001101",
  61888=>"101101101",
  61889=>"101011111",
  61890=>"101111110",
  61891=>"100010010",
  61892=>"000011000",
  61893=>"000100110",
  61894=>"011001001",
  61895=>"100111000",
  61896=>"100010011",
  61897=>"101111110",
  61898=>"010100110",
  61899=>"010111110",
  61900=>"011110000",
  61901=>"001011111",
  61902=>"101111100",
  61903=>"001101101",
  61904=>"101001010",
  61905=>"111100000",
  61906=>"101010010",
  61907=>"101001010",
  61908=>"111100111",
  61909=>"001000001",
  61910=>"000101011",
  61911=>"110010111",
  61912=>"011111111",
  61913=>"111110101",
  61914=>"000010111",
  61915=>"101001100",
  61916=>"100011001",
  61917=>"100111010",
  61918=>"011110011",
  61919=>"111001011",
  61920=>"100010111",
  61921=>"010111000",
  61922=>"010110001",
  61923=>"011100010",
  61924=>"001011101",
  61925=>"110000101",
  61926=>"111101001",
  61927=>"000011010",
  61928=>"011100001",
  61929=>"010000010",
  61930=>"000101011",
  61931=>"101001101",
  61932=>"110001011",
  61933=>"010010011",
  61934=>"000110001",
  61935=>"011100100",
  61936=>"101011011",
  61937=>"111001110",
  61938=>"000110101",
  61939=>"001110111",
  61940=>"000010101",
  61941=>"010101010",
  61942=>"110000010",
  61943=>"110000100",
  61944=>"000001101",
  61945=>"011111001",
  61946=>"110101001",
  61947=>"010010001",
  61948=>"000010001",
  61949=>"101100000",
  61950=>"001011011",
  61951=>"101111110",
  61952=>"101100010",
  61953=>"111001000",
  61954=>"110100100",
  61955=>"001100010",
  61956=>"100010100",
  61957=>"100011010",
  61958=>"110110110",
  61959=>"000000000",
  61960=>"000110100",
  61961=>"100001001",
  61962=>"100001011",
  61963=>"000111000",
  61964=>"101100000",
  61965=>"111001000",
  61966=>"010100001",
  61967=>"100001101",
  61968=>"101010111",
  61969=>"100000000",
  61970=>"111011111",
  61971=>"011101010",
  61972=>"110010000",
  61973=>"001110110",
  61974=>"000101001",
  61975=>"101011111",
  61976=>"100001100",
  61977=>"110001110",
  61978=>"110011111",
  61979=>"011101011",
  61980=>"101001011",
  61981=>"010100111",
  61982=>"001110011",
  61983=>"110110001",
  61984=>"111001101",
  61985=>"001100100",
  61986=>"111001011",
  61987=>"110101101",
  61988=>"000000001",
  61989=>"001000000",
  61990=>"111111110",
  61991=>"010000010",
  61992=>"110110000",
  61993=>"101000010",
  61994=>"101100011",
  61995=>"000001011",
  61996=>"000110001",
  61997=>"000000011",
  61998=>"111001101",
  61999=>"101111101",
  62000=>"001111101",
  62001=>"010110000",
  62002=>"111110001",
  62003=>"010000011",
  62004=>"111011000",
  62005=>"010100101",
  62006=>"001010010",
  62007=>"010001100",
  62008=>"011101100",
  62009=>"110010110",
  62010=>"001101100",
  62011=>"100010000",
  62012=>"100110000",
  62013=>"000110100",
  62014=>"111100100",
  62015=>"010001101",
  62016=>"101010011",
  62017=>"100011001",
  62018=>"100100011",
  62019=>"111000010",
  62020=>"111110111",
  62021=>"100100001",
  62022=>"001000001",
  62023=>"000110000",
  62024=>"001001110",
  62025=>"011011101",
  62026=>"010000110",
  62027=>"101111101",
  62028=>"110010000",
  62029=>"001001000",
  62030=>"110110010",
  62031=>"011100000",
  62032=>"000010011",
  62033=>"000000011",
  62034=>"100101001",
  62035=>"110111000",
  62036=>"010011011",
  62037=>"111000100",
  62038=>"111101111",
  62039=>"011101010",
  62040=>"011001110",
  62041=>"001110100",
  62042=>"100000001",
  62043=>"100100100",
  62044=>"001010110",
  62045=>"101011110",
  62046=>"100101100",
  62047=>"010001001",
  62048=>"100100110",
  62049=>"100100011",
  62050=>"110010100",
  62051=>"111001000",
  62052=>"111111000",
  62053=>"000001111",
  62054=>"111000111",
  62055=>"101111110",
  62056=>"010101110",
  62057=>"101011110",
  62058=>"011101000",
  62059=>"010000101",
  62060=>"010100001",
  62061=>"101100010",
  62062=>"001101001",
  62063=>"011001011",
  62064=>"000110111",
  62065=>"100000100",
  62066=>"011001000",
  62067=>"100110010",
  62068=>"000110001",
  62069=>"101100111",
  62070=>"010101110",
  62071=>"001100100",
  62072=>"001011110",
  62073=>"111110111",
  62074=>"010010111",
  62075=>"100011110",
  62076=>"011000100",
  62077=>"111001101",
  62078=>"100111111",
  62079=>"010110000",
  62080=>"100100100",
  62081=>"111010100",
  62082=>"001011111",
  62083=>"101111010",
  62084=>"110000010",
  62085=>"000001000",
  62086=>"111000001",
  62087=>"111100001",
  62088=>"111101001",
  62089=>"111110111",
  62090=>"100101000",
  62091=>"101110011",
  62092=>"110101000",
  62093=>"100110100",
  62094=>"111111001",
  62095=>"110110011",
  62096=>"000111010",
  62097=>"111001110",
  62098=>"101101011",
  62099=>"010100100",
  62100=>"001100100",
  62101=>"010110100",
  62102=>"101111110",
  62103=>"010101011",
  62104=>"111011010",
  62105=>"101001010",
  62106=>"100001011",
  62107=>"001100000",
  62108=>"010101001",
  62109=>"000000111",
  62110=>"001000011",
  62111=>"111010011",
  62112=>"100001110",
  62113=>"001010000",
  62114=>"110001100",
  62115=>"000000010",
  62116=>"001010010",
  62117=>"000011011",
  62118=>"010000001",
  62119=>"011111101",
  62120=>"100110010",
  62121=>"111111010",
  62122=>"001110001",
  62123=>"001110011",
  62124=>"010010001",
  62125=>"111111011",
  62126=>"010010110",
  62127=>"011101111",
  62128=>"111101011",
  62129=>"010100000",
  62130=>"001101101",
  62131=>"011110101",
  62132=>"110110010",
  62133=>"111101101",
  62134=>"110000001",
  62135=>"010010100",
  62136=>"001111011",
  62137=>"111100010",
  62138=>"000010101",
  62139=>"011100111",
  62140=>"101100110",
  62141=>"001000001",
  62142=>"111011001",
  62143=>"001011101",
  62144=>"101101111",
  62145=>"010100101",
  62146=>"010110011",
  62147=>"010000101",
  62148=>"100100111",
  62149=>"101100100",
  62150=>"000001001",
  62151=>"101011101",
  62152=>"011110011",
  62153=>"100000010",
  62154=>"111010011",
  62155=>"100110101",
  62156=>"110001000",
  62157=>"011101100",
  62158=>"100101100",
  62159=>"110110001",
  62160=>"110001001",
  62161=>"110011010",
  62162=>"110110001",
  62163=>"011111011",
  62164=>"111111011",
  62165=>"110100001",
  62166=>"110011011",
  62167=>"110000001",
  62168=>"100000101",
  62169=>"000101001",
  62170=>"110010101",
  62171=>"000000111",
  62172=>"000100000",
  62173=>"100100110",
  62174=>"010011011",
  62175=>"011010110",
  62176=>"110111000",
  62177=>"000101111",
  62178=>"111100000",
  62179=>"111111000",
  62180=>"000000111",
  62181=>"010001000",
  62182=>"101100000",
  62183=>"000001100",
  62184=>"111001110",
  62185=>"100111001",
  62186=>"111100001",
  62187=>"111011111",
  62188=>"000000100",
  62189=>"001001011",
  62190=>"111011110",
  62191=>"000001110",
  62192=>"010100100",
  62193=>"000000100",
  62194=>"100101100",
  62195=>"100110111",
  62196=>"001100010",
  62197=>"010101110",
  62198=>"111110101",
  62199=>"011101000",
  62200=>"001010100",
  62201=>"010001010",
  62202=>"010011001",
  62203=>"011100001",
  62204=>"001111111",
  62205=>"101101000",
  62206=>"100111001",
  62207=>"000010101",
  62208=>"001011010",
  62209=>"011111100",
  62210=>"111100001",
  62211=>"000110101",
  62212=>"010111010",
  62213=>"011100000",
  62214=>"001000110",
  62215=>"100110000",
  62216=>"111000101",
  62217=>"010100001",
  62218=>"111110010",
  62219=>"011011001",
  62220=>"001000010",
  62221=>"101101011",
  62222=>"010000110",
  62223=>"010000010",
  62224=>"010101100",
  62225=>"001011011",
  62226=>"010100111",
  62227=>"111011110",
  62228=>"100110111",
  62229=>"001011111",
  62230=>"110000010",
  62231=>"110101000",
  62232=>"111001000",
  62233=>"100011000",
  62234=>"110001010",
  62235=>"111010101",
  62236=>"001111111",
  62237=>"100111010",
  62238=>"100010101",
  62239=>"000000000",
  62240=>"010010000",
  62241=>"100000100",
  62242=>"101101000",
  62243=>"110100001",
  62244=>"001100111",
  62245=>"101100000",
  62246=>"001011101",
  62247=>"110110011",
  62248=>"000010001",
  62249=>"001011000",
  62250=>"110011001",
  62251=>"110101101",
  62252=>"001101111",
  62253=>"001010000",
  62254=>"111001100",
  62255=>"010001010",
  62256=>"111000000",
  62257=>"100000111",
  62258=>"001101001",
  62259=>"000001111",
  62260=>"110010011",
  62261=>"111001101",
  62262=>"000000011",
  62263=>"000011111",
  62264=>"110101110",
  62265=>"010011001",
  62266=>"100110101",
  62267=>"110010111",
  62268=>"100001111",
  62269=>"001110000",
  62270=>"110100101",
  62271=>"110100011",
  62272=>"100101001",
  62273=>"111111011",
  62274=>"000000000",
  62275=>"101110001",
  62276=>"111001100",
  62277=>"111010101",
  62278=>"111101111",
  62279=>"100101000",
  62280=>"001110100",
  62281=>"110101001",
  62282=>"011111100",
  62283=>"010100010",
  62284=>"110100100",
  62285=>"011011100",
  62286=>"111101000",
  62287=>"110101010",
  62288=>"001001011",
  62289=>"101001101",
  62290=>"100111111",
  62291=>"110111000",
  62292=>"001101001",
  62293=>"101110110",
  62294=>"101001010",
  62295=>"000001001",
  62296=>"001110111",
  62297=>"010001110",
  62298=>"011101010",
  62299=>"001001001",
  62300=>"011111111",
  62301=>"111101110",
  62302=>"001000001",
  62303=>"010110011",
  62304=>"010000110",
  62305=>"100110101",
  62306=>"000001000",
  62307=>"001001100",
  62308=>"100010011",
  62309=>"111000101",
  62310=>"101100100",
  62311=>"111011001",
  62312=>"000000011",
  62313=>"110000110",
  62314=>"011011100",
  62315=>"000111000",
  62316=>"100101101",
  62317=>"001100011",
  62318=>"011000100",
  62319=>"111100110",
  62320=>"110001111",
  62321=>"011100111",
  62322=>"111010101",
  62323=>"100111000",
  62324=>"100100010",
  62325=>"100001000",
  62326=>"110001001",
  62327=>"001001110",
  62328=>"101010011",
  62329=>"001000101",
  62330=>"110001111",
  62331=>"100101100",
  62332=>"001110000",
  62333=>"101011011",
  62334=>"111101111",
  62335=>"011110101",
  62336=>"101011010",
  62337=>"100011101",
  62338=>"001101101",
  62339=>"111010011",
  62340=>"011101110",
  62341=>"111111000",
  62342=>"011111010",
  62343=>"101101000",
  62344=>"001110001",
  62345=>"110010101",
  62346=>"011000011",
  62347=>"001100011",
  62348=>"001100000",
  62349=>"101000001",
  62350=>"001111110",
  62351=>"100000100",
  62352=>"011001110",
  62353=>"011111111",
  62354=>"010001010",
  62355=>"111010101",
  62356=>"110011111",
  62357=>"101010010",
  62358=>"101011110",
  62359=>"010110100",
  62360=>"101000101",
  62361=>"111111111",
  62362=>"111110000",
  62363=>"000010010",
  62364=>"111001100",
  62365=>"101010100",
  62366=>"001100011",
  62367=>"001000011",
  62368=>"111111110",
  62369=>"010001010",
  62370=>"011101010",
  62371=>"101010011",
  62372=>"011110000",
  62373=>"101111010",
  62374=>"001110101",
  62375=>"011110000",
  62376=>"010001000",
  62377=>"100010110",
  62378=>"011110100",
  62379=>"100011010",
  62380=>"010010110",
  62381=>"111010110",
  62382=>"011011110",
  62383=>"010100010",
  62384=>"010001111",
  62385=>"001110110",
  62386=>"101011001",
  62387=>"010110101",
  62388=>"100101110",
  62389=>"111100111",
  62390=>"000111011",
  62391=>"101111000",
  62392=>"111000001",
  62393=>"001000100",
  62394=>"001011011",
  62395=>"001001000",
  62396=>"101001110",
  62397=>"000001001",
  62398=>"111011001",
  62399=>"001011000",
  62400=>"101001001",
  62401=>"000100001",
  62402=>"000001100",
  62403=>"111011011",
  62404=>"100101100",
  62405=>"100111011",
  62406=>"111011100",
  62407=>"000000001",
  62408=>"011110011",
  62409=>"100010010",
  62410=>"111010111",
  62411=>"001111100",
  62412=>"111101010",
  62413=>"111110000",
  62414=>"011111011",
  62415=>"101010100",
  62416=>"010000001",
  62417=>"101011100",
  62418=>"010010000",
  62419=>"001101111",
  62420=>"001100111",
  62421=>"100000001",
  62422=>"110110111",
  62423=>"011011010",
  62424=>"011000000",
  62425=>"010010100",
  62426=>"101111100",
  62427=>"000111110",
  62428=>"101011110",
  62429=>"100001000",
  62430=>"111001001",
  62431=>"110100011",
  62432=>"101100010",
  62433=>"011111101",
  62434=>"000101000",
  62435=>"110100001",
  62436=>"111000100",
  62437=>"000010010",
  62438=>"001000111",
  62439=>"000110011",
  62440=>"011000110",
  62441=>"110000010",
  62442=>"100100010",
  62443=>"000111000",
  62444=>"001111101",
  62445=>"110000000",
  62446=>"000011010",
  62447=>"011001000",
  62448=>"111110001",
  62449=>"110111010",
  62450=>"001111000",
  62451=>"100001110",
  62452=>"010000001",
  62453=>"001110000",
  62454=>"001001000",
  62455=>"000111010",
  62456=>"010011110",
  62457=>"100101001",
  62458=>"010010001",
  62459=>"000111111",
  62460=>"010110000",
  62461=>"100100110",
  62462=>"001001010",
  62463=>"000111010",
  62464=>"111101101",
  62465=>"001111011",
  62466=>"010111111",
  62467=>"010100111",
  62468=>"101101001",
  62469=>"111010110",
  62470=>"000011101",
  62471=>"111001100",
  62472=>"000001100",
  62473=>"000100110",
  62474=>"100011000",
  62475=>"100100111",
  62476=>"010000011",
  62477=>"111111101",
  62478=>"001001110",
  62479=>"110111111",
  62480=>"000011101",
  62481=>"000101111",
  62482=>"111100010",
  62483=>"111100000",
  62484=>"011001000",
  62485=>"110000101",
  62486=>"100000010",
  62487=>"001100010",
  62488=>"010110111",
  62489=>"001000111",
  62490=>"110101010",
  62491=>"001110011",
  62492=>"001010010",
  62493=>"000111010",
  62494=>"100111111",
  62495=>"111100110",
  62496=>"110010010",
  62497=>"111001000",
  62498=>"100011010",
  62499=>"001110110",
  62500=>"000001000",
  62501=>"001100101",
  62502=>"100111100",
  62503=>"000100110",
  62504=>"110011101",
  62505=>"101110011",
  62506=>"100111101",
  62507=>"000110101",
  62508=>"110110000",
  62509=>"101011110",
  62510=>"010010000",
  62511=>"110100111",
  62512=>"000010000",
  62513=>"111000100",
  62514=>"011100000",
  62515=>"000110101",
  62516=>"001101111",
  62517=>"101001000",
  62518=>"101011010",
  62519=>"010000111",
  62520=>"100001000",
  62521=>"010001001",
  62522=>"100010010",
  62523=>"111001011",
  62524=>"100100010",
  62525=>"011010110",
  62526=>"101011101",
  62527=>"110111010",
  62528=>"001101000",
  62529=>"110010110",
  62530=>"010010000",
  62531=>"101111100",
  62532=>"101001000",
  62533=>"110111111",
  62534=>"001011111",
  62535=>"110000110",
  62536=>"011110101",
  62537=>"110110001",
  62538=>"011010011",
  62539=>"000010010",
  62540=>"101010110",
  62541=>"101011110",
  62542=>"110101111",
  62543=>"111101011",
  62544=>"100111010",
  62545=>"100001110",
  62546=>"111011100",
  62547=>"111010101",
  62548=>"001000011",
  62549=>"011100010",
  62550=>"011010000",
  62551=>"000011000",
  62552=>"110001010",
  62553=>"111101010",
  62554=>"111111011",
  62555=>"011001011",
  62556=>"011000111",
  62557=>"000011011",
  62558=>"001101100",
  62559=>"011010010",
  62560=>"110000010",
  62561=>"010010100",
  62562=>"000011001",
  62563=>"111001001",
  62564=>"010000000",
  62565=>"111000110",
  62566=>"001010110",
  62567=>"011010110",
  62568=>"101011101",
  62569=>"011011110",
  62570=>"011001101",
  62571=>"010111110",
  62572=>"011010100",
  62573=>"100001001",
  62574=>"101111000",
  62575=>"000001111",
  62576=>"011001001",
  62577=>"000100101",
  62578=>"000100001",
  62579=>"000100111",
  62580=>"100101000",
  62581=>"110010100",
  62582=>"011011110",
  62583=>"010100100",
  62584=>"101110100",
  62585=>"001100110",
  62586=>"111111111",
  62587=>"000110101",
  62588=>"000000001",
  62589=>"010101010",
  62590=>"110110100",
  62591=>"000110001",
  62592=>"001011101",
  62593=>"011010100",
  62594=>"001000100",
  62595=>"000001110",
  62596=>"000000111",
  62597=>"000101110",
  62598=>"111001000",
  62599=>"000001110",
  62600=>"000110011",
  62601=>"101010000",
  62602=>"000101011",
  62603=>"011111111",
  62604=>"011111111",
  62605=>"001010101",
  62606=>"010010101",
  62607=>"010011110",
  62608=>"101100101",
  62609=>"111101000",
  62610=>"000111111",
  62611=>"111110101",
  62612=>"101001011",
  62613=>"110100010",
  62614=>"111111000",
  62615=>"111001011",
  62616=>"111111011",
  62617=>"011111000",
  62618=>"010000010",
  62619=>"100110111",
  62620=>"010001010",
  62621=>"001000011",
  62622=>"110110000",
  62623=>"000111000",
  62624=>"001110010",
  62625=>"101010111",
  62626=>"110000000",
  62627=>"000101100",
  62628=>"100010100",
  62629=>"011011011",
  62630=>"101110011",
  62631=>"101000100",
  62632=>"100001010",
  62633=>"100101101",
  62634=>"100001001",
  62635=>"101000101",
  62636=>"000101001",
  62637=>"011010100",
  62638=>"001110100",
  62639=>"001110110",
  62640=>"001000111",
  62641=>"001000000",
  62642=>"101100011",
  62643=>"110000000",
  62644=>"110110110",
  62645=>"101011010",
  62646=>"001111010",
  62647=>"111100111",
  62648=>"001001011",
  62649=>"010001010",
  62650=>"101000101",
  62651=>"000101011",
  62652=>"011110111",
  62653=>"000000001",
  62654=>"100000011",
  62655=>"000000111",
  62656=>"011000110",
  62657=>"000010011",
  62658=>"000101010",
  62659=>"001001011",
  62660=>"011010110",
  62661=>"010101100",
  62662=>"001001011",
  62663=>"111100011",
  62664=>"001010011",
  62665=>"101001110",
  62666=>"010011110",
  62667=>"101100011",
  62668=>"100101000",
  62669=>"011101101",
  62670=>"101101110",
  62671=>"101001110",
  62672=>"000101010",
  62673=>"011101111",
  62674=>"001100110",
  62675=>"111001100",
  62676=>"111100001",
  62677=>"010000110",
  62678=>"110001111",
  62679=>"111111111",
  62680=>"011000001",
  62681=>"100001000",
  62682=>"001011110",
  62683=>"011001101",
  62684=>"011001011",
  62685=>"110110010",
  62686=>"101011011",
  62687=>"011101100",
  62688=>"110100110",
  62689=>"110000110",
  62690=>"000110101",
  62691=>"011111111",
  62692=>"110000100",
  62693=>"011110011",
  62694=>"001111100",
  62695=>"010001111",
  62696=>"100111111",
  62697=>"100001000",
  62698=>"011000000",
  62699=>"110010010",
  62700=>"010010001",
  62701=>"101000111",
  62702=>"001001111",
  62703=>"101010110",
  62704=>"000000111",
  62705=>"010111100",
  62706=>"000001111",
  62707=>"001011010",
  62708=>"011110011",
  62709=>"000011110",
  62710=>"111000110",
  62711=>"100101000",
  62712=>"110010001",
  62713=>"010000001",
  62714=>"110001000",
  62715=>"101011001",
  62716=>"110010100",
  62717=>"011111010",
  62718=>"010001111",
  62719=>"011100000",
  62720=>"100001000",
  62721=>"101010011",
  62722=>"100010000",
  62723=>"010100101",
  62724=>"101100101",
  62725=>"010111000",
  62726=>"001010100",
  62727=>"001110010",
  62728=>"111010011",
  62729=>"111000101",
  62730=>"000100011",
  62731=>"111100010",
  62732=>"001011101",
  62733=>"100100110",
  62734=>"100111100",
  62735=>"001011111",
  62736=>"110010001",
  62737=>"100111010",
  62738=>"011011000",
  62739=>"001110011",
  62740=>"001111011",
  62741=>"101101100",
  62742=>"000100100",
  62743=>"101000000",
  62744=>"010110111",
  62745=>"101010111",
  62746=>"100110101",
  62747=>"000001000",
  62748=>"110011001",
  62749=>"010010010",
  62750=>"111110101",
  62751=>"101001111",
  62752=>"001110011",
  62753=>"101110111",
  62754=>"100001010",
  62755=>"101000101",
  62756=>"001001111",
  62757=>"110101110",
  62758=>"111111110",
  62759=>"111000000",
  62760=>"101100111",
  62761=>"110100011",
  62762=>"011111011",
  62763=>"010010000",
  62764=>"110111100",
  62765=>"100111111",
  62766=>"001101010",
  62767=>"010100110",
  62768=>"110101100",
  62769=>"101100101",
  62770=>"111111001",
  62771=>"100100011",
  62772=>"111010001",
  62773=>"001010110",
  62774=>"011011100",
  62775=>"001101110",
  62776=>"111011001",
  62777=>"011011100",
  62778=>"111110111",
  62779=>"000101011",
  62780=>"011101101",
  62781=>"111000100",
  62782=>"010100101",
  62783=>"110100010",
  62784=>"011100000",
  62785=>"000111100",
  62786=>"110010110",
  62787=>"100001100",
  62788=>"001000011",
  62789=>"101111001",
  62790=>"010010011",
  62791=>"011110100",
  62792=>"010100010",
  62793=>"111000000",
  62794=>"101011010",
  62795=>"001010000",
  62796=>"100100000",
  62797=>"011001000",
  62798=>"101000101",
  62799=>"111010000",
  62800=>"111111001",
  62801=>"001100000",
  62802=>"101000011",
  62803=>"110110100",
  62804=>"000011100",
  62805=>"111000100",
  62806=>"111111110",
  62807=>"000111111",
  62808=>"111110010",
  62809=>"011100110",
  62810=>"110011000",
  62811=>"100000001",
  62812=>"111001100",
  62813=>"001011001",
  62814=>"010001110",
  62815=>"110001000",
  62816=>"100100110",
  62817=>"101001110",
  62818=>"000000011",
  62819=>"000001101",
  62820=>"011101111",
  62821=>"101001110",
  62822=>"000010101",
  62823=>"011010101",
  62824=>"001011101",
  62825=>"110111111",
  62826=>"111010001",
  62827=>"011100011",
  62828=>"000110110",
  62829=>"000111111",
  62830=>"001011011",
  62831=>"010011011",
  62832=>"011111111",
  62833=>"101000011",
  62834=>"110111011",
  62835=>"100101011",
  62836=>"011111000",
  62837=>"001001000",
  62838=>"011111001",
  62839=>"001010110",
  62840=>"101111000",
  62841=>"000111101",
  62842=>"110011110",
  62843=>"011100111",
  62844=>"001100101",
  62845=>"000001010",
  62846=>"001010000",
  62847=>"000011110",
  62848=>"000010001",
  62849=>"110011001",
  62850=>"001101100",
  62851=>"001111110",
  62852=>"001000000",
  62853=>"000111110",
  62854=>"001110010",
  62855=>"010110000",
  62856=>"101000000",
  62857=>"110101101",
  62858=>"010011010",
  62859=>"010110100",
  62860=>"111111101",
  62861=>"010111100",
  62862=>"001111001",
  62863=>"000100000",
  62864=>"111011001",
  62865=>"001000011",
  62866=>"101000011",
  62867=>"011100010",
  62868=>"101000010",
  62869=>"000110011",
  62870=>"101010001",
  62871=>"100111110",
  62872=>"111010111",
  62873=>"000111010",
  62874=>"010101000",
  62875=>"001001101",
  62876=>"100101101",
  62877=>"110101000",
  62878=>"011011011",
  62879=>"110110101",
  62880=>"100011011",
  62881=>"111010101",
  62882=>"011100101",
  62883=>"001111110",
  62884=>"111011000",
  62885=>"111010111",
  62886=>"011101010",
  62887=>"110000100",
  62888=>"010101111",
  62889=>"101111101",
  62890=>"001100100",
  62891=>"001010010",
  62892=>"111110011",
  62893=>"001010100",
  62894=>"101011010",
  62895=>"101110101",
  62896=>"111111100",
  62897=>"111110011",
  62898=>"111001101",
  62899=>"010100100",
  62900=>"110001100",
  62901=>"100101000",
  62902=>"010110000",
  62903=>"000010010",
  62904=>"011100100",
  62905=>"101000001",
  62906=>"101011101",
  62907=>"110100011",
  62908=>"111110110",
  62909=>"101110011",
  62910=>"000011011",
  62911=>"001010110",
  62912=>"001100111",
  62913=>"101110111",
  62914=>"100011110",
  62915=>"011010010",
  62916=>"000001011",
  62917=>"010101011",
  62918=>"010000010",
  62919=>"011010100",
  62920=>"000101000",
  62921=>"111111101",
  62922=>"000001001",
  62923=>"010110101",
  62924=>"000101111",
  62925=>"011101001",
  62926=>"101101110",
  62927=>"011101110",
  62928=>"100010110",
  62929=>"011110110",
  62930=>"000001101",
  62931=>"101110011",
  62932=>"011001111",
  62933=>"010100111",
  62934=>"000000000",
  62935=>"110111011",
  62936=>"101011001",
  62937=>"000011000",
  62938=>"100111010",
  62939=>"111110100",
  62940=>"110010111",
  62941=>"100110011",
  62942=>"011111000",
  62943=>"100010001",
  62944=>"000111110",
  62945=>"101101010",
  62946=>"111010111",
  62947=>"110110000",
  62948=>"110100101",
  62949=>"001100001",
  62950=>"010010001",
  62951=>"101110110",
  62952=>"000111001",
  62953=>"000010111",
  62954=>"110000110",
  62955=>"101110001",
  62956=>"110100111",
  62957=>"001011000",
  62958=>"111010101",
  62959=>"000101100",
  62960=>"010000100",
  62961=>"010010010",
  62962=>"011010010",
  62963=>"011111011",
  62964=>"101111000",
  62965=>"101110110",
  62966=>"101101010",
  62967=>"000011111",
  62968=>"111110100",
  62969=>"000110001",
  62970=>"010100101",
  62971=>"100010110",
  62972=>"010001010",
  62973=>"000100110",
  62974=>"100101101",
  62975=>"110101000",
  62976=>"101011110",
  62977=>"111010100",
  62978=>"010110100",
  62979=>"111010011",
  62980=>"001000111",
  62981=>"100010001",
  62982=>"100101000",
  62983=>"110001011",
  62984=>"000101110",
  62985=>"001110111",
  62986=>"110001010",
  62987=>"011000010",
  62988=>"000110101",
  62989=>"000000001",
  62990=>"111110111",
  62991=>"100111111",
  62992=>"111110000",
  62993=>"101000101",
  62994=>"010111000",
  62995=>"010111101",
  62996=>"011110100",
  62997=>"011100000",
  62998=>"100000000",
  62999=>"000101111",
  63000=>"110011110",
  63001=>"000000100",
  63002=>"001011110",
  63003=>"101011010",
  63004=>"100111111",
  63005=>"010010101",
  63006=>"000000010",
  63007=>"000110100",
  63008=>"011001101",
  63009=>"100000100",
  63010=>"010111110",
  63011=>"011001011",
  63012=>"100010111",
  63013=>"111010111",
  63014=>"000001100",
  63015=>"010001011",
  63016=>"000001111",
  63017=>"101101010",
  63018=>"011000100",
  63019=>"110000100",
  63020=>"100110111",
  63021=>"110111011",
  63022=>"010101100",
  63023=>"011100101",
  63024=>"000000101",
  63025=>"011011010",
  63026=>"000110011",
  63027=>"001001011",
  63028=>"111011001",
  63029=>"100110101",
  63030=>"010111000",
  63031=>"110011011",
  63032=>"111010001",
  63033=>"000001100",
  63034=>"111100101",
  63035=>"100010110",
  63036=>"101111100",
  63037=>"000010100",
  63038=>"001111011",
  63039=>"110111001",
  63040=>"001111010",
  63041=>"101000101",
  63042=>"111011100",
  63043=>"111010011",
  63044=>"010101100",
  63045=>"101000001",
  63046=>"100111100",
  63047=>"111010111",
  63048=>"000001001",
  63049=>"010000010",
  63050=>"100000001",
  63051=>"110101011",
  63052=>"111111010",
  63053=>"111110001",
  63054=>"011001100",
  63055=>"101111000",
  63056=>"111011111",
  63057=>"010001010",
  63058=>"001001011",
  63059=>"010011011",
  63060=>"010101010",
  63061=>"000000010",
  63062=>"110100100",
  63063=>"110011110",
  63064=>"000011000",
  63065=>"000000010",
  63066=>"001000001",
  63067=>"011100110",
  63068=>"100000010",
  63069=>"100110001",
  63070=>"010100101",
  63071=>"001011011",
  63072=>"100010000",
  63073=>"110001111",
  63074=>"110010101",
  63075=>"001001000",
  63076=>"011001111",
  63077=>"001000000",
  63078=>"000001101",
  63079=>"010111100",
  63080=>"101000110",
  63081=>"000001000",
  63082=>"110100010",
  63083=>"010101011",
  63084=>"010010010",
  63085=>"101001111",
  63086=>"001000110",
  63087=>"010111101",
  63088=>"110011111",
  63089=>"101001001",
  63090=>"000100010",
  63091=>"111100111",
  63092=>"011101010",
  63093=>"011001100",
  63094=>"100101010",
  63095=>"111010110",
  63096=>"101101000",
  63097=>"010011110",
  63098=>"001011100",
  63099=>"100110110",
  63100=>"001001110",
  63101=>"100110011",
  63102=>"010010010",
  63103=>"101011111",
  63104=>"000000011",
  63105=>"001000010",
  63106=>"001010101",
  63107=>"011000010",
  63108=>"001100000",
  63109=>"100000010",
  63110=>"110000011",
  63111=>"011111110",
  63112=>"110011100",
  63113=>"001011111",
  63114=>"110101111",
  63115=>"010000110",
  63116=>"000000011",
  63117=>"101101101",
  63118=>"101100011",
  63119=>"011010101",
  63120=>"010110101",
  63121=>"000000011",
  63122=>"110100010",
  63123=>"100000101",
  63124=>"111100100",
  63125=>"110111001",
  63126=>"010001111",
  63127=>"100001000",
  63128=>"011110100",
  63129=>"000010101",
  63130=>"111110100",
  63131=>"100110101",
  63132=>"010001110",
  63133=>"011111000",
  63134=>"010101000",
  63135=>"001001110",
  63136=>"011001000",
  63137=>"000100001",
  63138=>"100000000",
  63139=>"010001011",
  63140=>"110001000",
  63141=>"001000010",
  63142=>"011111001",
  63143=>"000000101",
  63144=>"111011110",
  63145=>"001101101",
  63146=>"001000010",
  63147=>"001100100",
  63148=>"110110101",
  63149=>"010100111",
  63150=>"110101000",
  63151=>"010001000",
  63152=>"010000000",
  63153=>"111010101",
  63154=>"101101010",
  63155=>"100000110",
  63156=>"110101111",
  63157=>"000011010",
  63158=>"111111011",
  63159=>"000011010",
  63160=>"010011111",
  63161=>"100110111",
  63162=>"110111011",
  63163=>"000010111",
  63164=>"011001001",
  63165=>"011001001",
  63166=>"001111111",
  63167=>"111100100",
  63168=>"101010111",
  63169=>"101000100",
  63170=>"110011010",
  63171=>"000011000",
  63172=>"000111001",
  63173=>"110111001",
  63174=>"000010100",
  63175=>"000100000",
  63176=>"010100111",
  63177=>"100011011",
  63178=>"101110001",
  63179=>"101110000",
  63180=>"010010011",
  63181=>"000011110",
  63182=>"010111010",
  63183=>"011101110",
  63184=>"010110010",
  63185=>"100010101",
  63186=>"001110101",
  63187=>"000101101",
  63188=>"001000110",
  63189=>"100101001",
  63190=>"100011101",
  63191=>"110011000",
  63192=>"111111011",
  63193=>"000110101",
  63194=>"101011101",
  63195=>"001010110",
  63196=>"101001010",
  63197=>"111101010",
  63198=>"101100011",
  63199=>"111111100",
  63200=>"010011100",
  63201=>"101100010",
  63202=>"010011010",
  63203=>"000010001",
  63204=>"001010000",
  63205=>"111101001",
  63206=>"110000011",
  63207=>"011001101",
  63208=>"110000100",
  63209=>"101101100",
  63210=>"111111111",
  63211=>"110011110",
  63212=>"010100110",
  63213=>"010011011",
  63214=>"111100101",
  63215=>"110101000",
  63216=>"011100000",
  63217=>"000101011",
  63218=>"010010100",
  63219=>"111011001",
  63220=>"110011111",
  63221=>"011000011",
  63222=>"011111100",
  63223=>"010001000",
  63224=>"010101000",
  63225=>"111110110",
  63226=>"001000001",
  63227=>"100010010",
  63228=>"101111101",
  63229=>"100110110",
  63230=>"111000011",
  63231=>"111111001",
  63232=>"011101100",
  63233=>"010111010",
  63234=>"000011110",
  63235=>"010100110",
  63236=>"111011000",
  63237=>"100011001",
  63238=>"010001101",
  63239=>"110010011",
  63240=>"000101101",
  63241=>"101011101",
  63242=>"011001010",
  63243=>"000100110",
  63244=>"111001111",
  63245=>"111011100",
  63246=>"110010000",
  63247=>"010101001",
  63248=>"001110110",
  63249=>"110111111",
  63250=>"001001000",
  63251=>"000011100",
  63252=>"100110110",
  63253=>"001000010",
  63254=>"101101010",
  63255=>"101001111",
  63256=>"011001000",
  63257=>"000100000",
  63258=>"001001011",
  63259=>"011101011",
  63260=>"000110111",
  63261=>"001001110",
  63262=>"110111110",
  63263=>"000001101",
  63264=>"110000001",
  63265=>"101110010",
  63266=>"000000101",
  63267=>"101001111",
  63268=>"010110010",
  63269=>"111110001",
  63270=>"010100010",
  63271=>"001110111",
  63272=>"010010001",
  63273=>"011101111",
  63274=>"110001110",
  63275=>"010000100",
  63276=>"100101011",
  63277=>"000100000",
  63278=>"000110100",
  63279=>"010001000",
  63280=>"010011011",
  63281=>"110000101",
  63282=>"100000111",
  63283=>"100111111",
  63284=>"001010101",
  63285=>"110100010",
  63286=>"011101000",
  63287=>"000110010",
  63288=>"000101001",
  63289=>"100000101",
  63290=>"001110111",
  63291=>"101010011",
  63292=>"011100000",
  63293=>"111000011",
  63294=>"100001100",
  63295=>"011111110",
  63296=>"100010100",
  63297=>"011000011",
  63298=>"111011001",
  63299=>"101011111",
  63300=>"010101101",
  63301=>"111010011",
  63302=>"000110010",
  63303=>"101111101",
  63304=>"010011100",
  63305=>"010110100",
  63306=>"010011000",
  63307=>"100000010",
  63308=>"011110011",
  63309=>"100111010",
  63310=>"111100010",
  63311=>"111011011",
  63312=>"100001111",
  63313=>"010101000",
  63314=>"100011011",
  63315=>"111001111",
  63316=>"001111000",
  63317=>"110010100",
  63318=>"100111100",
  63319=>"110001101",
  63320=>"000100111",
  63321=>"010101000",
  63322=>"111001000",
  63323=>"000111100",
  63324=>"000111000",
  63325=>"000101111",
  63326=>"111110000",
  63327=>"001000101",
  63328=>"000011010",
  63329=>"001101100",
  63330=>"101010101",
  63331=>"001010000",
  63332=>"011011111",
  63333=>"001100100",
  63334=>"100100110",
  63335=>"110101101",
  63336=>"100011101",
  63337=>"110111000",
  63338=>"111111100",
  63339=>"101010011",
  63340=>"000110011",
  63341=>"010001100",
  63342=>"011100001",
  63343=>"100000100",
  63344=>"100100111",
  63345=>"001100011",
  63346=>"000000110",
  63347=>"000101000",
  63348=>"001111000",
  63349=>"110111101",
  63350=>"000111011",
  63351=>"010010011",
  63352=>"000011011",
  63353=>"100110000",
  63354=>"111011101",
  63355=>"000000000",
  63356=>"111111101",
  63357=>"000000010",
  63358=>"000100001",
  63359=>"110010111",
  63360=>"110011000",
  63361=>"001010100",
  63362=>"010010011",
  63363=>"010010111",
  63364=>"001100000",
  63365=>"101011111",
  63366=>"110101100",
  63367=>"110100011",
  63368=>"100111110",
  63369=>"111001000",
  63370=>"010110110",
  63371=>"011000001",
  63372=>"010000001",
  63373=>"011001111",
  63374=>"110000101",
  63375=>"111111000",
  63376=>"111001011",
  63377=>"111010110",
  63378=>"011110100",
  63379=>"011001011",
  63380=>"011010100",
  63381=>"011111010",
  63382=>"111100111",
  63383=>"001001011",
  63384=>"001100011",
  63385=>"100110011",
  63386=>"000011110",
  63387=>"111101111",
  63388=>"001000110",
  63389=>"101010111",
  63390=>"011101000",
  63391=>"111000000",
  63392=>"100110001",
  63393=>"100110110",
  63394=>"000010000",
  63395=>"011111101",
  63396=>"100101100",
  63397=>"011011101",
  63398=>"100010011",
  63399=>"011001111",
  63400=>"011101111",
  63401=>"110111001",
  63402=>"100111110",
  63403=>"000101110",
  63404=>"010000100",
  63405=>"110111100",
  63406=>"100100101",
  63407=>"100100011",
  63408=>"001001100",
  63409=>"001110111",
  63410=>"011001100",
  63411=>"000011001",
  63412=>"101011001",
  63413=>"000101110",
  63414=>"100111010",
  63415=>"111111001",
  63416=>"000100000",
  63417=>"110010011",
  63418=>"111010010",
  63419=>"010011011",
  63420=>"010111110",
  63421=>"001111011",
  63422=>"100000001",
  63423=>"111100111",
  63424=>"111111010",
  63425=>"010111110",
  63426=>"101100011",
  63427=>"110100000",
  63428=>"011111010",
  63429=>"100000010",
  63430=>"100000101",
  63431=>"010011101",
  63432=>"010101111",
  63433=>"000111000",
  63434=>"000001000",
  63435=>"010100101",
  63436=>"010100010",
  63437=>"001001111",
  63438=>"010111000",
  63439=>"100010111",
  63440=>"001101011",
  63441=>"111100110",
  63442=>"101011010",
  63443=>"100100111",
  63444=>"001000111",
  63445=>"000000100",
  63446=>"111000111",
  63447=>"110111111",
  63448=>"010010100",
  63449=>"011010101",
  63450=>"011110011",
  63451=>"111101011",
  63452=>"111111101",
  63453=>"101000111",
  63454=>"011011011",
  63455=>"000110111",
  63456=>"101010100",
  63457=>"001011101",
  63458=>"110010100",
  63459=>"011100100",
  63460=>"101001011",
  63461=>"101100101",
  63462=>"000100101",
  63463=>"101100001",
  63464=>"010101001",
  63465=>"100100100",
  63466=>"011101100",
  63467=>"111110101",
  63468=>"011001001",
  63469=>"101000101",
  63470=>"010101101",
  63471=>"001011010",
  63472=>"000100001",
  63473=>"111100101",
  63474=>"110000011",
  63475=>"010011001",
  63476=>"001010100",
  63477=>"100100000",
  63478=>"001000001",
  63479=>"110000100",
  63480=>"110011101",
  63481=>"101011011",
  63482=>"100101001",
  63483=>"101101010",
  63484=>"001000111",
  63485=>"010001011",
  63486=>"001100110",
  63487=>"001000000",
  63488=>"010100111",
  63489=>"000101101",
  63490=>"101001010",
  63491=>"001000101",
  63492=>"010110010",
  63493=>"001111110",
  63494=>"111101001",
  63495=>"101001001",
  63496=>"111101000",
  63497=>"010100110",
  63498=>"011011011",
  63499=>"101101110",
  63500=>"100001000",
  63501=>"001110011",
  63502=>"010001001",
  63503=>"011011111",
  63504=>"001100001",
  63505=>"100100011",
  63506=>"111101010",
  63507=>"000110001",
  63508=>"001000010",
  63509=>"110110100",
  63510=>"001101010",
  63511=>"010001100",
  63512=>"011111100",
  63513=>"010101111",
  63514=>"010000101",
  63515=>"101100101",
  63516=>"101001001",
  63517=>"111101001",
  63518=>"110010101",
  63519=>"000010011",
  63520=>"101001111",
  63521=>"000011010",
  63522=>"011000001",
  63523=>"101001000",
  63524=>"100110110",
  63525=>"100010000",
  63526=>"011000110",
  63527=>"101000010",
  63528=>"110100100",
  63529=>"000010011",
  63530=>"010111111",
  63531=>"010001000",
  63532=>"001000011",
  63533=>"111101000",
  63534=>"110110101",
  63535=>"110110001",
  63536=>"100100111",
  63537=>"000101010",
  63538=>"001101001",
  63539=>"011001100",
  63540=>"110110100",
  63541=>"000011110",
  63542=>"111000000",
  63543=>"100011001",
  63544=>"011100100",
  63545=>"001101001",
  63546=>"100001011",
  63547=>"111001010",
  63548=>"011100110",
  63549=>"001000100",
  63550=>"000011000",
  63551=>"100111101",
  63552=>"111001111",
  63553=>"101010010",
  63554=>"010010001",
  63555=>"001001100",
  63556=>"111100100",
  63557=>"110110110",
  63558=>"110110010",
  63559=>"010001000",
  63560=>"111100101",
  63561=>"011011011",
  63562=>"010100111",
  63563=>"111001001",
  63564=>"000001111",
  63565=>"110100000",
  63566=>"111011100",
  63567=>"000001010",
  63568=>"011001000",
  63569=>"000100101",
  63570=>"001010111",
  63571=>"100010100",
  63572=>"111100110",
  63573=>"000100110",
  63574=>"100000100",
  63575=>"000100010",
  63576=>"111111010",
  63577=>"011000010",
  63578=>"111000110",
  63579=>"000011011",
  63580=>"000000000",
  63581=>"110101111",
  63582=>"010000111",
  63583=>"101001101",
  63584=>"100011110",
  63585=>"011110101",
  63586=>"110101000",
  63587=>"101101101",
  63588=>"001100011",
  63589=>"111001101",
  63590=>"100101011",
  63591=>"000010000",
  63592=>"000011000",
  63593=>"010011000",
  63594=>"011010011",
  63595=>"000101011",
  63596=>"010000000",
  63597=>"011010010",
  63598=>"000011011",
  63599=>"010100010",
  63600=>"111100001",
  63601=>"101011111",
  63602=>"000011000",
  63603=>"001001011",
  63604=>"000001000",
  63605=>"010101100",
  63606=>"110011101",
  63607=>"111101110",
  63608=>"001100100",
  63609=>"011010011",
  63610=>"010010101",
  63611=>"100101011",
  63612=>"001101111",
  63613=>"101000110",
  63614=>"000000001",
  63615=>"111010011",
  63616=>"000010100",
  63617=>"001000111",
  63618=>"010001111",
  63619=>"100100100",
  63620=>"001110010",
  63621=>"100110111",
  63622=>"001101111",
  63623=>"001010001",
  63624=>"000001110",
  63625=>"101001010",
  63626=>"111010000",
  63627=>"011110000",
  63628=>"111111001",
  63629=>"001000000",
  63630=>"111010011",
  63631=>"110011000",
  63632=>"011100110",
  63633=>"011110000",
  63634=>"101011010",
  63635=>"101000101",
  63636=>"111000110",
  63637=>"000010010",
  63638=>"111000110",
  63639=>"001001101",
  63640=>"101101111",
  63641=>"000000001",
  63642=>"000100011",
  63643=>"100110011",
  63644=>"111101101",
  63645=>"111110110",
  63646=>"010010010",
  63647=>"001001111",
  63648=>"010011001",
  63649=>"000100100",
  63650=>"011001000",
  63651=>"110101001",
  63652=>"000110001",
  63653=>"111111101",
  63654=>"101101101",
  63655=>"100000001",
  63656=>"101011011",
  63657=>"001010000",
  63658=>"100011101",
  63659=>"011100101",
  63660=>"110100001",
  63661=>"100001111",
  63662=>"001101100",
  63663=>"101111111",
  63664=>"011000010",
  63665=>"001100111",
  63666=>"000010100",
  63667=>"101001000",
  63668=>"000111100",
  63669=>"000101011",
  63670=>"111000110",
  63671=>"110000011",
  63672=>"110011111",
  63673=>"010110111",
  63674=>"111001101",
  63675=>"011011110",
  63676=>"001101000",
  63677=>"100000000",
  63678=>"111101110",
  63679=>"011000111",
  63680=>"001000000",
  63681=>"111000000",
  63682=>"101001111",
  63683=>"101110100",
  63684=>"111100011",
  63685=>"101111101",
  63686=>"011010110",
  63687=>"100011110",
  63688=>"000010010",
  63689=>"100100000",
  63690=>"101111111",
  63691=>"010010011",
  63692=>"111001010",
  63693=>"101110100",
  63694=>"010101111",
  63695=>"101100000",
  63696=>"001100111",
  63697=>"101111100",
  63698=>"101010010",
  63699=>"001011001",
  63700=>"000100011",
  63701=>"110000010",
  63702=>"110110001",
  63703=>"101001001",
  63704=>"011010001",
  63705=>"000110111",
  63706=>"011110111",
  63707=>"001101010",
  63708=>"110101101",
  63709=>"011100101",
  63710=>"011101100",
  63711=>"010101001",
  63712=>"001000101",
  63713=>"000000101",
  63714=>"101011010",
  63715=>"010101001",
  63716=>"101000101",
  63717=>"001011001",
  63718=>"100011100",
  63719=>"001111111",
  63720=>"010010010",
  63721=>"010011010",
  63722=>"001011011",
  63723=>"100000101",
  63724=>"111101000",
  63725=>"100000101",
  63726=>"110011100",
  63727=>"111110000",
  63728=>"011110111",
  63729=>"000000001",
  63730=>"001111010",
  63731=>"101000101",
  63732=>"001100110",
  63733=>"100001000",
  63734=>"001010010",
  63735=>"010111000",
  63736=>"101100010",
  63737=>"101101010",
  63738=>"000101000",
  63739=>"000001011",
  63740=>"001101010",
  63741=>"101001001",
  63742=>"110001101",
  63743=>"101000000",
  63744=>"010000011",
  63745=>"100000000",
  63746=>"101110001",
  63747=>"010111000",
  63748=>"010000000",
  63749=>"000010001",
  63750=>"010010110",
  63751=>"000000100",
  63752=>"110110010",
  63753=>"011010111",
  63754=>"101111000",
  63755=>"111100110",
  63756=>"011000011",
  63757=>"101001011",
  63758=>"001110000",
  63759=>"100000111",
  63760=>"010000011",
  63761=>"011111101",
  63762=>"011010000",
  63763=>"111011001",
  63764=>"101000110",
  63765=>"111010001",
  63766=>"000101111",
  63767=>"001001110",
  63768=>"111000100",
  63769=>"000011000",
  63770=>"010111111",
  63771=>"100101110",
  63772=>"011010111",
  63773=>"101100100",
  63774=>"011010001",
  63775=>"010110111",
  63776=>"110111100",
  63777=>"101010110",
  63778=>"010000100",
  63779=>"000000101",
  63780=>"110010111",
  63781=>"010010111",
  63782=>"100110001",
  63783=>"101011010",
  63784=>"111110100",
  63785=>"011111111",
  63786=>"111001010",
  63787=>"011010110",
  63788=>"010010110",
  63789=>"110111110",
  63790=>"101101000",
  63791=>"000001111",
  63792=>"111111101",
  63793=>"001001111",
  63794=>"110101011",
  63795=>"100100000",
  63796=>"011101011",
  63797=>"101101111",
  63798=>"010010111",
  63799=>"110010100",
  63800=>"011010110",
  63801=>"000010011",
  63802=>"101000001",
  63803=>"111111000",
  63804=>"101010011",
  63805=>"011000010",
  63806=>"000101101",
  63807=>"010100001",
  63808=>"111010100",
  63809=>"001000000",
  63810=>"000000101",
  63811=>"110101001",
  63812=>"101111110",
  63813=>"000111101",
  63814=>"110001101",
  63815=>"110011011",
  63816=>"001011110",
  63817=>"001010001",
  63818=>"000110111",
  63819=>"100101010",
  63820=>"001110010",
  63821=>"000101100",
  63822=>"000110000",
  63823=>"101000011",
  63824=>"001010100",
  63825=>"001101000",
  63826=>"010101111",
  63827=>"011001101",
  63828=>"100011100",
  63829=>"001110010",
  63830=>"111011011",
  63831=>"100000111",
  63832=>"010001010",
  63833=>"100111111",
  63834=>"010101100",
  63835=>"111100100",
  63836=>"001111111",
  63837=>"010011011",
  63838=>"110110100",
  63839=>"011100011",
  63840=>"101000000",
  63841=>"010001000",
  63842=>"010101011",
  63843=>"010001100",
  63844=>"010101101",
  63845=>"100010110",
  63846=>"111001101",
  63847=>"101010100",
  63848=>"100111111",
  63849=>"110010000",
  63850=>"111001101",
  63851=>"101110001",
  63852=>"111110111",
  63853=>"100101110",
  63854=>"000010100",
  63855=>"110110101",
  63856=>"001010010",
  63857=>"001010111",
  63858=>"011000101",
  63859=>"100100100",
  63860=>"110010100",
  63861=>"100111000",
  63862=>"101100010",
  63863=>"011111110",
  63864=>"000100001",
  63865=>"111011000",
  63866=>"001111110",
  63867=>"111110010",
  63868=>"011011000",
  63869=>"000000111",
  63870=>"101100110",
  63871=>"101101000",
  63872=>"001110011",
  63873=>"010000000",
  63874=>"010110001",
  63875=>"000111000",
  63876=>"110101110",
  63877=>"000010000",
  63878=>"111011010",
  63879=>"010110110",
  63880=>"000000110",
  63881=>"101101001",
  63882=>"000000101",
  63883=>"010101110",
  63884=>"011110110",
  63885=>"001001010",
  63886=>"100010001",
  63887=>"010000010",
  63888=>"111000101",
  63889=>"100001111",
  63890=>"001111001",
  63891=>"101100101",
  63892=>"101001101",
  63893=>"001101110",
  63894=>"000011001",
  63895=>"100010000",
  63896=>"111111111",
  63897=>"111111000",
  63898=>"001011011",
  63899=>"001101011",
  63900=>"100001101",
  63901=>"111110111",
  63902=>"111100110",
  63903=>"010001110",
  63904=>"101100111",
  63905=>"111100111",
  63906=>"100000010",
  63907=>"110011000",
  63908=>"100011111",
  63909=>"001101110",
  63910=>"011111110",
  63911=>"101011001",
  63912=>"111110111",
  63913=>"010110000",
  63914=>"001110110",
  63915=>"000110010",
  63916=>"001010001",
  63917=>"001110001",
  63918=>"101110100",
  63919=>"111110010",
  63920=>"101111011",
  63921=>"001010001",
  63922=>"000111111",
  63923=>"101011100",
  63924=>"110001110",
  63925=>"101011110",
  63926=>"000100100",
  63927=>"011111001",
  63928=>"101101001",
  63929=>"011100100",
  63930=>"010100010",
  63931=>"111110010",
  63932=>"101000010",
  63933=>"011101011",
  63934=>"111111001",
  63935=>"000100011",
  63936=>"101110111",
  63937=>"000010001",
  63938=>"010101100",
  63939=>"001101010",
  63940=>"100110101",
  63941=>"100110011",
  63942=>"001001101",
  63943=>"101000011",
  63944=>"100101100",
  63945=>"001100011",
  63946=>"101100101",
  63947=>"111100110",
  63948=>"110111111",
  63949=>"110011101",
  63950=>"100011011",
  63951=>"011000100",
  63952=>"011000000",
  63953=>"011011001",
  63954=>"011110101",
  63955=>"111110111",
  63956=>"100010000",
  63957=>"010011100",
  63958=>"001100010",
  63959=>"011100000",
  63960=>"010010011",
  63961=>"110010111",
  63962=>"101100100",
  63963=>"001000110",
  63964=>"100011111",
  63965=>"001111011",
  63966=>"001101010",
  63967=>"001111001",
  63968=>"010101010",
  63969=>"100111011",
  63970=>"000011011",
  63971=>"011110100",
  63972=>"110010001",
  63973=>"111011000",
  63974=>"101000110",
  63975=>"011000101",
  63976=>"010101010",
  63977=>"000111111",
  63978=>"101101110",
  63979=>"110110110",
  63980=>"000101010",
  63981=>"101100101",
  63982=>"010010100",
  63983=>"001110000",
  63984=>"110111110",
  63985=>"100010101",
  63986=>"000000000",
  63987=>"001111111",
  63988=>"100101011",
  63989=>"010011101",
  63990=>"000010000",
  63991=>"101000100",
  63992=>"011000010",
  63993=>"100100000",
  63994=>"000101000",
  63995=>"001010000",
  63996=>"100100000",
  63997=>"111011001",
  63998=>"110100010",
  63999=>"010000000",
  64000=>"011010110",
  64001=>"100010100",
  64002=>"001011000",
  64003=>"001000000",
  64004=>"001011100",
  64005=>"110010100",
  64006=>"010110000",
  64007=>"101110101",
  64008=>"000111001",
  64009=>"010001011",
  64010=>"001110110",
  64011=>"111111111",
  64012=>"010010000",
  64013=>"010100110",
  64014=>"100000100",
  64015=>"011110100",
  64016=>"001100101",
  64017=>"011011111",
  64018=>"000100011",
  64019=>"110000111",
  64020=>"001100011",
  64021=>"011111011",
  64022=>"010010010",
  64023=>"101000011",
  64024=>"010010110",
  64025=>"100000111",
  64026=>"100111101",
  64027=>"101011111",
  64028=>"010010011",
  64029=>"101101101",
  64030=>"010001110",
  64031=>"010111100",
  64032=>"000010101",
  64033=>"001111011",
  64034=>"111010000",
  64035=>"100000010",
  64036=>"100010010",
  64037=>"011000000",
  64038=>"111101000",
  64039=>"100000000",
  64040=>"101110101",
  64041=>"010000000",
  64042=>"111000000",
  64043=>"111110010",
  64044=>"101111001",
  64045=>"000011000",
  64046=>"101001000",
  64047=>"101111110",
  64048=>"010000010",
  64049=>"001000001",
  64050=>"110100101",
  64051=>"000000010",
  64052=>"110110100",
  64053=>"101010111",
  64054=>"110110011",
  64055=>"110101011",
  64056=>"010111100",
  64057=>"010011100",
  64058=>"111001000",
  64059=>"000001100",
  64060=>"011111110",
  64061=>"000011001",
  64062=>"011000000",
  64063=>"011110001",
  64064=>"101011111",
  64065=>"010000000",
  64066=>"011111001",
  64067=>"010010111",
  64068=>"000100100",
  64069=>"110010010",
  64070=>"110100101",
  64071=>"010100001",
  64072=>"010010110",
  64073=>"111010001",
  64074=>"101101000",
  64075=>"100101110",
  64076=>"001001100",
  64077=>"001111110",
  64078=>"010001100",
  64079=>"011110100",
  64080=>"011101111",
  64081=>"011001110",
  64082=>"100111001",
  64083=>"001111101",
  64084=>"001010011",
  64085=>"110101110",
  64086=>"111001110",
  64087=>"000011110",
  64088=>"010100111",
  64089=>"010100010",
  64090=>"100100101",
  64091=>"000110001",
  64092=>"001111001",
  64093=>"010100000",
  64094=>"111001110",
  64095=>"000000001",
  64096=>"100101010",
  64097=>"110100000",
  64098=>"100010001",
  64099=>"100101011",
  64100=>"001011110",
  64101=>"110111111",
  64102=>"001000100",
  64103=>"101000010",
  64104=>"101110110",
  64105=>"010010001",
  64106=>"011100011",
  64107=>"110100101",
  64108=>"110001001",
  64109=>"111011011",
  64110=>"000101110",
  64111=>"111100001",
  64112=>"000101100",
  64113=>"001000000",
  64114=>"100101011",
  64115=>"100001011",
  64116=>"011111111",
  64117=>"101001101",
  64118=>"111001001",
  64119=>"111000110",
  64120=>"100001111",
  64121=>"111100000",
  64122=>"001100001",
  64123=>"010100011",
  64124=>"110001101",
  64125=>"100011111",
  64126=>"100001010",
  64127=>"111000001",
  64128=>"000000001",
  64129=>"100000100",
  64130=>"010111110",
  64131=>"111110111",
  64132=>"111010010",
  64133=>"110000001",
  64134=>"001010011",
  64135=>"100010000",
  64136=>"010110111",
  64137=>"111110001",
  64138=>"111001111",
  64139=>"110000111",
  64140=>"110010000",
  64141=>"001001101",
  64142=>"110110110",
  64143=>"000001111",
  64144=>"001000010",
  64145=>"111111000",
  64146=>"101001000",
  64147=>"011111111",
  64148=>"010101100",
  64149=>"011101010",
  64150=>"000010001",
  64151=>"010100110",
  64152=>"100001001",
  64153=>"010011000",
  64154=>"010010111",
  64155=>"111010000",
  64156=>"000100111",
  64157=>"010001101",
  64158=>"001110001",
  64159=>"101110111",
  64160=>"000000010",
  64161=>"001011101",
  64162=>"111100000",
  64163=>"111100100",
  64164=>"100001010",
  64165=>"001100101",
  64166=>"001011011",
  64167=>"000000001",
  64168=>"011011010",
  64169=>"001001011",
  64170=>"100111111",
  64171=>"010011100",
  64172=>"101110000",
  64173=>"000000011",
  64174=>"110000110",
  64175=>"010101101",
  64176=>"111000101",
  64177=>"111001110",
  64178=>"001010101",
  64179=>"001001100",
  64180=>"111010110",
  64181=>"010110010",
  64182=>"011010110",
  64183=>"110000001",
  64184=>"101011100",
  64185=>"000011011",
  64186=>"011010111",
  64187=>"000000100",
  64188=>"010011000",
  64189=>"001001010",
  64190=>"111100100",
  64191=>"110100101",
  64192=>"100100111",
  64193=>"011101111",
  64194=>"001101111",
  64195=>"010000001",
  64196=>"111110001",
  64197=>"111101101",
  64198=>"000000100",
  64199=>"000100001",
  64200=>"000000010",
  64201=>"010111000",
  64202=>"101010100",
  64203=>"011100100",
  64204=>"110011111",
  64205=>"001011110",
  64206=>"101001101",
  64207=>"001011111",
  64208=>"011111110",
  64209=>"000001001",
  64210=>"101000010",
  64211=>"000100001",
  64212=>"011111111",
  64213=>"000100100",
  64214=>"111111110",
  64215=>"010011100",
  64216=>"111001101",
  64217=>"100101000",
  64218=>"000001010",
  64219=>"011101111",
  64220=>"010100100",
  64221=>"100010011",
  64222=>"111111010",
  64223=>"001001000",
  64224=>"000111110",
  64225=>"010011000",
  64226=>"010010011",
  64227=>"110100110",
  64228=>"111001111",
  64229=>"010100101",
  64230=>"011000101",
  64231=>"100111110",
  64232=>"101011100",
  64233=>"001000111",
  64234=>"011111111",
  64235=>"100001001",
  64236=>"010010111",
  64237=>"111011110",
  64238=>"101001101",
  64239=>"100000101",
  64240=>"011100101",
  64241=>"100011001",
  64242=>"100110000",
  64243=>"010010110",
  64244=>"101101101",
  64245=>"000000010",
  64246=>"000110010",
  64247=>"110001101",
  64248=>"110001111",
  64249=>"111000011",
  64250=>"101110000",
  64251=>"101110101",
  64252=>"000100000",
  64253=>"110100000",
  64254=>"000111010",
  64255=>"101111011",
  64256=>"010011001",
  64257=>"101011101",
  64258=>"010011000",
  64259=>"001100011",
  64260=>"100000010",
  64261=>"100100010",
  64262=>"101101000",
  64263=>"100111101",
  64264=>"001011010",
  64265=>"110100000",
  64266=>"011101111",
  64267=>"001011101",
  64268=>"000110100",
  64269=>"000011000",
  64270=>"000101110",
  64271=>"010000111",
  64272=>"110011001",
  64273=>"110100111",
  64274=>"010100000",
  64275=>"111001100",
  64276=>"111001111",
  64277=>"100010000",
  64278=>"000000011",
  64279=>"100000111",
  64280=>"001000111",
  64281=>"110011011",
  64282=>"111001001",
  64283=>"110000100",
  64284=>"100111010",
  64285=>"100111000",
  64286=>"010101011",
  64287=>"110010001",
  64288=>"100000001",
  64289=>"010111110",
  64290=>"011000000",
  64291=>"011111110",
  64292=>"000001010",
  64293=>"001010011",
  64294=>"110011111",
  64295=>"001101111",
  64296=>"100101111",
  64297=>"010100010",
  64298=>"011100011",
  64299=>"110000101",
  64300=>"100001001",
  64301=>"101110110",
  64302=>"011111101",
  64303=>"110010101",
  64304=>"011101111",
  64305=>"111111000",
  64306=>"110110100",
  64307=>"011110010",
  64308=>"010001110",
  64309=>"010110010",
  64310=>"110110011",
  64311=>"011100100",
  64312=>"110100011",
  64313=>"000101001",
  64314=>"001001001",
  64315=>"111101011",
  64316=>"001110000",
  64317=>"111111010",
  64318=>"010001101",
  64319=>"000101100",
  64320=>"101001100",
  64321=>"010101000",
  64322=>"000011101",
  64323=>"001010100",
  64324=>"111001001",
  64325=>"001011101",
  64326=>"010110100",
  64327=>"100010100",
  64328=>"111010101",
  64329=>"101001001",
  64330=>"011011111",
  64331=>"111000100",
  64332=>"101111110",
  64333=>"110110100",
  64334=>"101011001",
  64335=>"000100111",
  64336=>"110101101",
  64337=>"010000001",
  64338=>"100110110",
  64339=>"110001110",
  64340=>"110110100",
  64341=>"101100110",
  64342=>"000001111",
  64343=>"111110000",
  64344=>"010111111",
  64345=>"100101110",
  64346=>"100011111",
  64347=>"010010101",
  64348=>"111001110",
  64349=>"110011011",
  64350=>"010111111",
  64351=>"001000110",
  64352=>"110111010",
  64353=>"111000010",
  64354=>"010111101",
  64355=>"110000001",
  64356=>"110000100",
  64357=>"010111011",
  64358=>"101101001",
  64359=>"000100001",
  64360=>"101001000",
  64361=>"010110001",
  64362=>"011110111",
  64363=>"001111110",
  64364=>"001101000",
  64365=>"111010000",
  64366=>"101011010",
  64367=>"111001110",
  64368=>"100111000",
  64369=>"101110110",
  64370=>"110011101",
  64371=>"111101001",
  64372=>"111000001",
  64373=>"101111100",
  64374=>"100111111",
  64375=>"010010110",
  64376=>"100110000",
  64377=>"001101111",
  64378=>"001011010",
  64379=>"101000001",
  64380=>"100011111",
  64381=>"001011000",
  64382=>"100101100",
  64383=>"110111111",
  64384=>"100111011",
  64385=>"100101111",
  64386=>"010111101",
  64387=>"000111101",
  64388=>"101101000",
  64389=>"110101111",
  64390=>"111011111",
  64391=>"001010110",
  64392=>"011110110",
  64393=>"111000010",
  64394=>"110111111",
  64395=>"100000110",
  64396=>"111000011",
  64397=>"111000011",
  64398=>"111000110",
  64399=>"000001010",
  64400=>"010001100",
  64401=>"111111000",
  64402=>"010001101",
  64403=>"111110110",
  64404=>"111101110",
  64405=>"010000110",
  64406=>"110101011",
  64407=>"010100010",
  64408=>"010010101",
  64409=>"000010001",
  64410=>"110111010",
  64411=>"100101010",
  64412=>"000100000",
  64413=>"001001001",
  64414=>"000110111",
  64415=>"001101001",
  64416=>"111001000",
  64417=>"100011001",
  64418=>"111111110",
  64419=>"110011011",
  64420=>"110010000",
  64421=>"000110101",
  64422=>"001010111",
  64423=>"001011100",
  64424=>"100010001",
  64425=>"001001111",
  64426=>"001111101",
  64427=>"111000001",
  64428=>"110010011",
  64429=>"011101001",
  64430=>"001100111",
  64431=>"101011010",
  64432=>"100000010",
  64433=>"000111100",
  64434=>"111001001",
  64435=>"011101111",
  64436=>"011011010",
  64437=>"000000010",
  64438=>"001100010",
  64439=>"110110100",
  64440=>"111000110",
  64441=>"111110110",
  64442=>"110010100",
  64443=>"100110010",
  64444=>"101001000",
  64445=>"010000111",
  64446=>"100100010",
  64447=>"001100100",
  64448=>"100100000",
  64449=>"010000000",
  64450=>"111111111",
  64451=>"101011111",
  64452=>"110000001",
  64453=>"010001011",
  64454=>"011111110",
  64455=>"110111011",
  64456=>"111010000",
  64457=>"100101000",
  64458=>"110010001",
  64459=>"101110011",
  64460=>"010011110",
  64461=>"100100111",
  64462=>"011110111",
  64463=>"110010110",
  64464=>"111100110",
  64465=>"011111110",
  64466=>"001101011",
  64467=>"110101010",
  64468=>"011011010",
  64469=>"010011000",
  64470=>"011100010",
  64471=>"110101111",
  64472=>"111110001",
  64473=>"110111110",
  64474=>"011101100",
  64475=>"100110000",
  64476=>"111101100",
  64477=>"101110111",
  64478=>"000001010",
  64479=>"100010100",
  64480=>"011110001",
  64481=>"111101100",
  64482=>"011110011",
  64483=>"011111000",
  64484=>"000011101",
  64485=>"100111101",
  64486=>"101100111",
  64487=>"100100000",
  64488=>"001100011",
  64489=>"110110011",
  64490=>"001111011",
  64491=>"000110111",
  64492=>"011010000",
  64493=>"000101001",
  64494=>"011010011",
  64495=>"011110111",
  64496=>"111001100",
  64497=>"011010010",
  64498=>"101001101",
  64499=>"110110010",
  64500=>"001000011",
  64501=>"010001011",
  64502=>"110011100",
  64503=>"101010100",
  64504=>"101111000",
  64505=>"101101110",
  64506=>"110101100",
  64507=>"101011011",
  64508=>"110101100",
  64509=>"101110000",
  64510=>"011111011",
  64511=>"010010010",
  64512=>"011001001",
  64513=>"000100001",
  64514=>"000100010",
  64515=>"101101011",
  64516=>"010011110",
  64517=>"110000101",
  64518=>"011011000",
  64519=>"110100100",
  64520=>"011010100",
  64521=>"111101000",
  64522=>"011011101",
  64523=>"100101010",
  64524=>"100000010",
  64525=>"100011110",
  64526=>"000000001",
  64527=>"011111110",
  64528=>"010100000",
  64529=>"101010100",
  64530=>"010110011",
  64531=>"000110111",
  64532=>"101000011",
  64533=>"100101000",
  64534=>"010100011",
  64535=>"000110101",
  64536=>"100110101",
  64537=>"101001001",
  64538=>"011111111",
  64539=>"111000101",
  64540=>"110001000",
  64541=>"011110010",
  64542=>"010001111",
  64543=>"001011011",
  64544=>"010011011",
  64545=>"101111101",
  64546=>"000010010",
  64547=>"101001011",
  64548=>"000100110",
  64549=>"101110001",
  64550=>"001101110",
  64551=>"000111100",
  64552=>"111100001",
  64553=>"000110111",
  64554=>"011101010",
  64555=>"110100011",
  64556=>"010001010",
  64557=>"100110001",
  64558=>"011001111",
  64559=>"101011111",
  64560=>"001110011",
  64561=>"110111000",
  64562=>"111100111",
  64563=>"100011000",
  64564=>"000001111",
  64565=>"111100101",
  64566=>"110001110",
  64567=>"011000010",
  64568=>"001100011",
  64569=>"111001111",
  64570=>"110000111",
  64571=>"111110010",
  64572=>"110011001",
  64573=>"100110111",
  64574=>"011111010",
  64575=>"101011000",
  64576=>"001101010",
  64577=>"000010001",
  64578=>"110011100",
  64579=>"110001111",
  64580=>"000100011",
  64581=>"110010011",
  64582=>"111110111",
  64583=>"001101001",
  64584=>"000010000",
  64585=>"011000001",
  64586=>"100000000",
  64587=>"110101101",
  64588=>"010000011",
  64589=>"001010101",
  64590=>"100001011",
  64591=>"100011010",
  64592=>"111100010",
  64593=>"010111111",
  64594=>"100011001",
  64595=>"011011010",
  64596=>"001011100",
  64597=>"100010101",
  64598=>"110101000",
  64599=>"100110111",
  64600=>"010100110",
  64601=>"101101111",
  64602=>"010011001",
  64603=>"010001011",
  64604=>"110101110",
  64605=>"001101101",
  64606=>"011001111",
  64607=>"010000111",
  64608=>"001110000",
  64609=>"000111110",
  64610=>"000010000",
  64611=>"010001010",
  64612=>"000111100",
  64613=>"101111011",
  64614=>"010001011",
  64615=>"110101010",
  64616=>"010100011",
  64617=>"010010001",
  64618=>"000100100",
  64619=>"110011111",
  64620=>"111111011",
  64621=>"001100111",
  64622=>"110001011",
  64623=>"110110000",
  64624=>"000110100",
  64625=>"010110111",
  64626=>"100100011",
  64627=>"000010111",
  64628=>"100000011",
  64629=>"111110110",
  64630=>"111100111",
  64631=>"110101111",
  64632=>"111100000",
  64633=>"010111110",
  64634=>"101100011",
  64635=>"100011000",
  64636=>"110000001",
  64637=>"111011110",
  64638=>"111110100",
  64639=>"011001010",
  64640=>"100001011",
  64641=>"010110011",
  64642=>"000011100",
  64643=>"110110100",
  64644=>"111011100",
  64645=>"110100011",
  64646=>"100010000",
  64647=>"101110110",
  64648=>"111100111",
  64649=>"001010000",
  64650=>"111001000",
  64651=>"010101010",
  64652=>"110010010",
  64653=>"000111100",
  64654=>"010111010",
  64655=>"011000010",
  64656=>"001011101",
  64657=>"100111111",
  64658=>"010000111",
  64659=>"010001011",
  64660=>"000101000",
  64661=>"111100111",
  64662=>"000100011",
  64663=>"111110011",
  64664=>"111001110",
  64665=>"110010111",
  64666=>"010110101",
  64667=>"110100100",
  64668=>"000010000",
  64669=>"101101011",
  64670=>"000000101",
  64671=>"110100011",
  64672=>"001100010",
  64673=>"010101000",
  64674=>"110000100",
  64675=>"011100110",
  64676=>"101011010",
  64677=>"010001010",
  64678=>"011101101",
  64679=>"101101101",
  64680=>"111110101",
  64681=>"010100000",
  64682=>"110000000",
  64683=>"011110010",
  64684=>"100000110",
  64685=>"100010001",
  64686=>"111011110",
  64687=>"010010011",
  64688=>"101001101",
  64689=>"111000000",
  64690=>"101001001",
  64691=>"010010110",
  64692=>"111001011",
  64693=>"110100100",
  64694=>"111001100",
  64695=>"101010011",
  64696=>"010000101",
  64697=>"100000110",
  64698=>"011011011",
  64699=>"100011110",
  64700=>"100001001",
  64701=>"010100001",
  64702=>"010000100",
  64703=>"101100001",
  64704=>"011101011",
  64705=>"001101010",
  64706=>"011100011",
  64707=>"101000000",
  64708=>"100110000",
  64709=>"000011000",
  64710=>"000100101",
  64711=>"101000000",
  64712=>"001100011",
  64713=>"010011011",
  64714=>"000011100",
  64715=>"100111001",
  64716=>"010010011",
  64717=>"101111010",
  64718=>"110111010",
  64719=>"101000100",
  64720=>"011010101",
  64721=>"000100001",
  64722=>"111001010",
  64723=>"001001001",
  64724=>"101011101",
  64725=>"110001011",
  64726=>"100000011",
  64727=>"111000011",
  64728=>"101010101",
  64729=>"000001101",
  64730=>"000110101",
  64731=>"100000010",
  64732=>"000111111",
  64733=>"110101110",
  64734=>"011101000",
  64735=>"010111110",
  64736=>"110001101",
  64737=>"011110010",
  64738=>"011000010",
  64739=>"010000000",
  64740=>"001011111",
  64741=>"110000011",
  64742=>"000000001",
  64743=>"000001000",
  64744=>"101001100",
  64745=>"001110011",
  64746=>"001011000",
  64747=>"101001001",
  64748=>"101000010",
  64749=>"001010111",
  64750=>"110111000",
  64751=>"101000011",
  64752=>"001011010",
  64753=>"011001000",
  64754=>"101011010",
  64755=>"110001111",
  64756=>"010000011",
  64757=>"101011000",
  64758=>"010000110",
  64759=>"101000111",
  64760=>"111111011",
  64761=>"000110101",
  64762=>"101011010",
  64763=>"001111100",
  64764=>"111110001",
  64765=>"110010110",
  64766=>"011110001",
  64767=>"000111111",
  64768=>"111101110",
  64769=>"100100110",
  64770=>"111111001",
  64771=>"100010000",
  64772=>"111011010",
  64773=>"000101110",
  64774=>"101011001",
  64775=>"001101011",
  64776=>"000011100",
  64777=>"000110011",
  64778=>"001110100",
  64779=>"111100011",
  64780=>"100100100",
  64781=>"010100101",
  64782=>"010111001",
  64783=>"000001101",
  64784=>"001001001",
  64785=>"101001010",
  64786=>"001011111",
  64787=>"101000010",
  64788=>"100111101",
  64789=>"100010011",
  64790=>"101001010",
  64791=>"000111110",
  64792=>"010000001",
  64793=>"011000111",
  64794=>"111001010",
  64795=>"000101000",
  64796=>"001010111",
  64797=>"010100000",
  64798=>"011101101",
  64799=>"001111111",
  64800=>"000100001",
  64801=>"010101111",
  64802=>"001110011",
  64803=>"000101100",
  64804=>"101001011",
  64805=>"010010100",
  64806=>"001110000",
  64807=>"101111000",
  64808=>"011010100",
  64809=>"010001111",
  64810=>"101111011",
  64811=>"100101111",
  64812=>"011011010",
  64813=>"110110000",
  64814=>"000101100",
  64815=>"111100110",
  64816=>"100111101",
  64817=>"110100011",
  64818=>"111111101",
  64819=>"010001100",
  64820=>"111011101",
  64821=>"011110111",
  64822=>"101011100",
  64823=>"101111111",
  64824=>"100000101",
  64825=>"110100010",
  64826=>"000100000",
  64827=>"011101010",
  64828=>"010010001",
  64829=>"110110010",
  64830=>"010111000",
  64831=>"111111000",
  64832=>"110001001",
  64833=>"100000001",
  64834=>"001111111",
  64835=>"011000001",
  64836=>"011101011",
  64837=>"010001110",
  64838=>"000110110",
  64839=>"011000111",
  64840=>"100100000",
  64841=>"110010011",
  64842=>"010100000",
  64843=>"101011010",
  64844=>"001110110",
  64845=>"110101110",
  64846=>"110111100",
  64847=>"100000011",
  64848=>"100000010",
  64849=>"011010011",
  64850=>"101001000",
  64851=>"011010111",
  64852=>"110110101",
  64853=>"000111011",
  64854=>"000010011",
  64855=>"010100000",
  64856=>"010101000",
  64857=>"101111110",
  64858=>"110100001",
  64859=>"100101000",
  64860=>"100001010",
  64861=>"000100001",
  64862=>"101011111",
  64863=>"011110010",
  64864=>"100000011",
  64865=>"111000111",
  64866=>"100010010",
  64867=>"000100111",
  64868=>"000010001",
  64869=>"000011101",
  64870=>"100110111",
  64871=>"000110100",
  64872=>"100010100",
  64873=>"000001101",
  64874=>"110101111",
  64875=>"000011101",
  64876=>"110000000",
  64877=>"110110010",
  64878=>"111101111",
  64879=>"001100001",
  64880=>"111101110",
  64881=>"100101010",
  64882=>"010100111",
  64883=>"011001001",
  64884=>"111111001",
  64885=>"101001001",
  64886=>"111000001",
  64887=>"010100111",
  64888=>"110111101",
  64889=>"101111001",
  64890=>"011011001",
  64891=>"101000110",
  64892=>"000001111",
  64893=>"111000011",
  64894=>"100011101",
  64895=>"010000000",
  64896=>"000111100",
  64897=>"101111001",
  64898=>"111011111",
  64899=>"010110110",
  64900=>"110111101",
  64901=>"001000010",
  64902=>"100111010",
  64903=>"001101010",
  64904=>"000001011",
  64905=>"110111110",
  64906=>"011101001",
  64907=>"001000111",
  64908=>"101110111",
  64909=>"001100000",
  64910=>"011111110",
  64911=>"011001110",
  64912=>"111100101",
  64913=>"000000100",
  64914=>"100010110",
  64915=>"100000000",
  64916=>"010001010",
  64917=>"111001111",
  64918=>"110001111",
  64919=>"011101010",
  64920=>"111000000",
  64921=>"001010001",
  64922=>"110110110",
  64923=>"011011011",
  64924=>"101110111",
  64925=>"001110100",
  64926=>"000000011",
  64927=>"111101001",
  64928=>"011001000",
  64929=>"110010001",
  64930=>"000010101",
  64931=>"001001011",
  64932=>"000000000",
  64933=>"110110100",
  64934=>"110100111",
  64935=>"100111011",
  64936=>"100111101",
  64937=>"001100111",
  64938=>"111011010",
  64939=>"000010000",
  64940=>"100111000",
  64941=>"101001111",
  64942=>"110010100",
  64943=>"101100111",
  64944=>"000110111",
  64945=>"010110000",
  64946=>"110010100",
  64947=>"110100110",
  64948=>"001101100",
  64949=>"110110111",
  64950=>"010110001",
  64951=>"100111101",
  64952=>"010110011",
  64953=>"011010111",
  64954=>"010000100",
  64955=>"010010111",
  64956=>"001011111",
  64957=>"100110001",
  64958=>"111110111",
  64959=>"100111010",
  64960=>"010110000",
  64961=>"111100000",
  64962=>"111010110",
  64963=>"111111110",
  64964=>"001101101",
  64965=>"011001111",
  64966=>"010000000",
  64967=>"101011000",
  64968=>"110110110",
  64969=>"110000101",
  64970=>"000000001",
  64971=>"011001101",
  64972=>"010101011",
  64973=>"111010000",
  64974=>"001000011",
  64975=>"011110011",
  64976=>"111000101",
  64977=>"001000010",
  64978=>"000001101",
  64979=>"000101111",
  64980=>"000000011",
  64981=>"011101100",
  64982=>"100010011",
  64983=>"100110101",
  64984=>"001001111",
  64985=>"111100000",
  64986=>"110010000",
  64987=>"110010101",
  64988=>"001001011",
  64989=>"000010011",
  64990=>"101101011",
  64991=>"111100110",
  64992=>"000010001",
  64993=>"011011010",
  64994=>"110101010",
  64995=>"000000010",
  64996=>"111100011",
  64997=>"110001010",
  64998=>"000101010",
  64999=>"001011100",
  65000=>"101000001",
  65001=>"010011001",
  65002=>"100111100",
  65003=>"010111001",
  65004=>"111001000",
  65005=>"111000101",
  65006=>"000111011",
  65007=>"111101101",
  65008=>"010111000",
  65009=>"010100110",
  65010=>"101100111",
  65011=>"011011001",
  65012=>"001111101",
  65013=>"001001011",
  65014=>"001110110",
  65015=>"101000101",
  65016=>"011000100",
  65017=>"100011010",
  65018=>"010101110",
  65019=>"100010010",
  65020=>"001101011",
  65021=>"111010011",
  65022=>"101000010",
  65023=>"011100000",
  65024=>"001110010",
  65025=>"001101101",
  65026=>"010010110",
  65027=>"011011011",
  65028=>"110101001",
  65029=>"110111111",
  65030=>"110010101",
  65031=>"110111001",
  65032=>"111111101",
  65033=>"110010100",
  65034=>"101111001",
  65035=>"110111101",
  65036=>"001111111",
  65037=>"101001011",
  65038=>"100111110",
  65039=>"111111010",
  65040=>"001101100",
  65041=>"001101111",
  65042=>"111101110",
  65043=>"000000000",
  65044=>"000011010",
  65045=>"100111000",
  65046=>"000001011",
  65047=>"101000111",
  65048=>"010111101",
  65049=>"111011101",
  65050=>"011111010",
  65051=>"101010101",
  65052=>"100100011",
  65053=>"000001101",
  65054=>"111101111",
  65055=>"101100000",
  65056=>"010010111",
  65057=>"001000110",
  65058=>"001110000",
  65059=>"001000010",
  65060=>"111100000",
  65061=>"110101010",
  65062=>"101000000",
  65063=>"101101101",
  65064=>"110101001",
  65065=>"111111001",
  65066=>"110101100",
  65067=>"010000100",
  65068=>"000110110",
  65069=>"000011110",
  65070=>"010111000",
  65071=>"000001101",
  65072=>"010001010",
  65073=>"001001001",
  65074=>"100100001",
  65075=>"011101011",
  65076=>"111011100",
  65077=>"111101100",
  65078=>"011111101",
  65079=>"100000111",
  65080=>"110011100",
  65081=>"100011010",
  65082=>"101001110",
  65083=>"111110111",
  65084=>"110111100",
  65085=>"101001000",
  65086=>"000001010",
  65087=>"010000000",
  65088=>"010011111",
  65089=>"000111111",
  65090=>"010100011",
  65091=>"101101010",
  65092=>"001111001",
  65093=>"110000101",
  65094=>"100000111",
  65095=>"000101000",
  65096=>"101101010",
  65097=>"100001011",
  65098=>"101011100",
  65099=>"010110111",
  65100=>"011000100",
  65101=>"001000010",
  65102=>"101110100",
  65103=>"001100100",
  65104=>"110010010",
  65105=>"110111011",
  65106=>"111101011",
  65107=>"001100010",
  65108=>"110000101",
  65109=>"111100001",
  65110=>"100110011",
  65111=>"010100111",
  65112=>"110111000",
  65113=>"000100110",
  65114=>"110001100",
  65115=>"000110111",
  65116=>"101000010",
  65117=>"101001111",
  65118=>"111010010",
  65119=>"011101100",
  65120=>"110011001",
  65121=>"001000000",
  65122=>"100101101",
  65123=>"011111111",
  65124=>"010010011",
  65125=>"001101111",
  65126=>"010100101",
  65127=>"110010110",
  65128=>"111110010",
  65129=>"001011111",
  65130=>"010010101",
  65131=>"010000000",
  65132=>"000011001",
  65133=>"011001010",
  65134=>"010110001",
  65135=>"111111000",
  65136=>"110110000",
  65137=>"101110001",
  65138=>"000111111",
  65139=>"011011101",
  65140=>"001000011",
  65141=>"101100110",
  65142=>"000100111",
  65143=>"110011001",
  65144=>"001011000",
  65145=>"100001000",
  65146=>"011011011",
  65147=>"101110100",
  65148=>"101101001",
  65149=>"110111110",
  65150=>"111111111",
  65151=>"111100000",
  65152=>"001000011",
  65153=>"000010110",
  65154=>"100010111",
  65155=>"000100001",
  65156=>"001100011",
  65157=>"110001001",
  65158=>"100101110",
  65159=>"010100101",
  65160=>"001000101",
  65161=>"111001101",
  65162=>"011100000",
  65163=>"011000110",
  65164=>"001000101",
  65165=>"100111000",
  65166=>"100010110",
  65167=>"110001011",
  65168=>"101010000",
  65169=>"011101011",
  65170=>"011111111",
  65171=>"110001010",
  65172=>"000110011",
  65173=>"010101000",
  65174=>"001111010",
  65175=>"101000000",
  65176=>"001111010",
  65177=>"000100000",
  65178=>"001010010",
  65179=>"001110101",
  65180=>"111111001",
  65181=>"111001101",
  65182=>"101110010",
  65183=>"101000011",
  65184=>"010000010",
  65185=>"000011111",
  65186=>"100011101",
  65187=>"011011001",
  65188=>"001001101",
  65189=>"101000111",
  65190=>"010111010",
  65191=>"101111010",
  65192=>"110101010",
  65193=>"101010111",
  65194=>"110011101",
  65195=>"001000011",
  65196=>"100100010",
  65197=>"111001100",
  65198=>"011001111",
  65199=>"010101000",
  65200=>"110111110",
  65201=>"010110000",
  65202=>"011011110",
  65203=>"111100000",
  65204=>"101110010",
  65205=>"000100000",
  65206=>"001010001",
  65207=>"110110111",
  65208=>"010111101",
  65209=>"011001111",
  65210=>"010101000",
  65211=>"010101011",
  65212=>"110111111",
  65213=>"010001100",
  65214=>"001001101",
  65215=>"110111101",
  65216=>"111000101",
  65217=>"111001100",
  65218=>"010110001",
  65219=>"011100001",
  65220=>"111011011",
  65221=>"010000111",
  65222=>"000100011",
  65223=>"101001001",
  65224=>"111010000",
  65225=>"100101111",
  65226=>"101111100",
  65227=>"001110110",
  65228=>"110011011",
  65229=>"110111000",
  65230=>"010010111",
  65231=>"011010111",
  65232=>"001101011",
  65233=>"010011011",
  65234=>"100110111",
  65235=>"101111101",
  65236=>"010100001",
  65237=>"101010111",
  65238=>"111110011",
  65239=>"000010110",
  65240=>"101101011",
  65241=>"110010100",
  65242=>"100110010",
  65243=>"100101110",
  65244=>"110101000",
  65245=>"000000000",
  65246=>"111001001",
  65247=>"111110100",
  65248=>"111100001",
  65249=>"100100110",
  65250=>"011110110",
  65251=>"100001000",
  65252=>"000001101",
  65253=>"100010111",
  65254=>"011001101",
  65255=>"000011100",
  65256=>"011010111",
  65257=>"100001100",
  65258=>"000111110",
  65259=>"000100110",
  65260=>"111101011",
  65261=>"111111000",
  65262=>"111110001",
  65263=>"110101111",
  65264=>"011011111",
  65265=>"100111011",
  65266=>"000111010",
  65267=>"110110001",
  65268=>"011001011",
  65269=>"000110110",
  65270=>"010010000",
  65271=>"010010110",
  65272=>"101001111",
  65273=>"110001001",
  65274=>"100011111",
  65275=>"110000100",
  65276=>"110011010",
  65277=>"110001011",
  65278=>"000111000",
  65279=>"001110011",
  65280=>"100110000",
  65281=>"011100011",
  65282=>"010001111",
  65283=>"001010110",
  65284=>"101001011",
  65285=>"010010100",
  65286=>"000010110",
  65287=>"011111001",
  65288=>"011111001",
  65289=>"001011000",
  65290=>"100100010",
  65291=>"000000000",
  65292=>"100111010",
  65293=>"001111110",
  65294=>"000100011",
  65295=>"011000111",
  65296=>"010010100",
  65297=>"100001000",
  65298=>"101100011",
  65299=>"100000101",
  65300=>"010100000",
  65301=>"100110101",
  65302=>"010110011",
  65303=>"000110111",
  65304=>"011010010",
  65305=>"001101000",
  65306=>"111011010",
  65307=>"001000010",
  65308=>"010110011",
  65309=>"110101101",
  65310=>"100101100",
  65311=>"000111101",
  65312=>"011111011",
  65313=>"100101001",
  65314=>"010100110",
  65315=>"101100000",
  65316=>"000011110",
  65317=>"000000010",
  65318=>"110011111",
  65319=>"011111001",
  65320=>"011011100",
  65321=>"110110011",
  65322=>"111110000",
  65323=>"110011101",
  65324=>"110100011",
  65325=>"011111011",
  65326=>"111100000",
  65327=>"011100000",
  65328=>"000101101",
  65329=>"111001000",
  65330=>"111000110",
  65331=>"101001000",
  65332=>"111010000",
  65333=>"101111111",
  65334=>"111011111",
  65335=>"100010111",
  65336=>"111011000",
  65337=>"100000101",
  65338=>"000000000",
  65339=>"101011000",
  65340=>"101110010",
  65341=>"111101101",
  65342=>"011101001",
  65343=>"111100011",
  65344=>"101000101",
  65345=>"011101111",
  65346=>"001010000",
  65347=>"010011001",
  65348=>"110011010",
  65349=>"001011011",
  65350=>"100100001",
  65351=>"001000000",
  65352=>"000010010",
  65353=>"111010001",
  65354=>"011000110",
  65355=>"010101000",
  65356=>"110100001",
  65357=>"000010110",
  65358=>"011101001",
  65359=>"010000000",
  65360=>"000001000",
  65361=>"000100111",
  65362=>"001001010",
  65363=>"011100000",
  65364=>"110100001",
  65365=>"110101000",
  65366=>"011001000",
  65367=>"001001111",
  65368=>"111111110",
  65369=>"111111110",
  65370=>"000100011",
  65371=>"110110011",
  65372=>"000001110",
  65373=>"110100111",
  65374=>"010101011",
  65375=>"001000101",
  65376=>"100011001",
  65377=>"101000101",
  65378=>"000110011",
  65379=>"000100000",
  65380=>"010010001",
  65381=>"101000010",
  65382=>"101110010",
  65383=>"111100000",
  65384=>"011001000",
  65385=>"111010001",
  65386=>"011100101",
  65387=>"101010110",
  65388=>"111101111",
  65389=>"011100000",
  65390=>"101001111",
  65391=>"000100100",
  65392=>"001101011",
  65393=>"001110100",
  65394=>"101000110",
  65395=>"000010111",
  65396=>"010001111",
  65397=>"011001000",
  65398=>"000101001",
  65399=>"101100011",
  65400=>"101010010",
  65401=>"110010010",
  65402=>"011101100",
  65403=>"110000111",
  65404=>"000001101",
  65405=>"001101011",
  65406=>"100011010",
  65407=>"011011001",
  65408=>"001001111",
  65409=>"010101000",
  65410=>"010010000",
  65411=>"110010101",
  65412=>"110001110",
  65413=>"101000000",
  65414=>"100001011",
  65415=>"001101110",
  65416=>"101011010",
  65417=>"111100001",
  65418=>"010011001",
  65419=>"100101111",
  65420=>"110101011",
  65421=>"100011011",
  65422=>"010010011",
  65423=>"010101001",
  65424=>"011000000",
  65425=>"010100001",
  65426=>"101000001",
  65427=>"111100100",
  65428=>"001111111",
  65429=>"110100111",
  65430=>"110110110",
  65431=>"010111000",
  65432=>"111101111",
  65433=>"111110100",
  65434=>"100001111",
  65435=>"001101110",
  65436=>"010111001",
  65437=>"100000001",
  65438=>"111000000",
  65439=>"010001100",
  65440=>"011001111",
  65441=>"111011111",
  65442=>"101001100",
  65443=>"000110010",
  65444=>"001110111",
  65445=>"011010001",
  65446=>"111001010",
  65447=>"101100001",
  65448=>"111111111",
  65449=>"001000000",
  65450=>"000011011",
  65451=>"100011100",
  65452=>"011101101",
  65453=>"111010001",
  65454=>"110101100",
  65455=>"101010011",
  65456=>"100101110",
  65457=>"111011010",
  65458=>"011111111",
  65459=>"011100000",
  65460=>"110000011",
  65461=>"001000111",
  65462=>"101100001",
  65463=>"000001000",
  65464=>"001000110",
  65465=>"001000111",
  65466=>"011011011",
  65467=>"110011011",
  65468=>"010011011",
  65469=>"110110000",
  65470=>"010011111",
  65471=>"110110101",
  65472=>"111110111",
  65473=>"000110001",
  65474=>"100000100",
  65475=>"100101111",
  65476=>"010101010",
  65477=>"010011100",
  65478=>"110011011",
  65479=>"111110110",
  65480=>"000010111",
  65481=>"110110101",
  65482=>"011100011",
  65483=>"001111111",
  65484=>"100110111",
  65485=>"100111001",
  65486=>"110101101",
  65487=>"110011011",
  65488=>"010111101",
  65489=>"110001110",
  65490=>"110010110",
  65491=>"011000111",
  65492=>"010111010",
  65493=>"010110111",
  65494=>"001010011",
  65495=>"100011010",
  65496=>"010011100",
  65497=>"000101010",
  65498=>"110111011",
  65499=>"100100010",
  65500=>"010110111",
  65501=>"000110111",
  65502=>"011001000",
  65503=>"100100110",
  65504=>"011111001",
  65505=>"100110010",
  65506=>"101010100",
  65507=>"100101011",
  65508=>"000010110",
  65509=>"001010111",
  65510=>"100011110",
  65511=>"000000011",
  65512=>"101111100",
  65513=>"101110001",
  65514=>"010101100",
  65515=>"101100010",
  65516=>"010010110",
  65517=>"110101011",
  65518=>"000000011",
  65519=>"000000001",
  65520=>"101111011",
  65521=>"010001001",
  65522=>"101011110",
  65523=>"101111111",
  65524=>"110111000",
  65525=>"100101000",
  65526=>"011011001",
  65527=>"111010111",
  65528=>"110101100",
  65529=>"110110101",
  65530=>"110010011",
  65531=>"101010000",
  65532=>"101011101",
  65533=>"111010011",
  65534=>"110001100",
  65535=>"011001100");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;