LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L6_1_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(7 DOWNTO 0));
END L6_1_BNROM;

ARCHITECTURE RTL OF L6_1_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"1111000011010101"&"0001110000110010",
  1=>"1111100010010011"&"0001010110100011",
  2=>"1111110100011110"&"0001001011011000",
  3=>"1111101111110001"&"0001111000010001",
  4=>"1111011001111010"&"0001111110011111",
  5=>"1110101010110000"&"0010000001111101",
  6=>"1111110101011011"&"0000111010001001",
  7=>"1111110010000011"&"0001011101011010",
  8=>"1111110010111011"&"0001100000101001",
  9=>"1111011011101100"&"0001111001100010",
  10=>"1111110001111011"&"0001011010000100",
  11=>"1111011010100111"&"0001111001011110",
  12=>"1111101000011001"&"0001010011101101",
  13=>"1111001111001110"&"0001101100000110",
  14=>"1111010001111100"&"0010001000011010",
  15=>"1111111110101111"&"0001000101010001",
  16=>"1111010100001110"&"0010000000000000",
  17=>"1111101100111100"&"0001011101100100",
  18=>"1111110110000000"&"0001010101110011",
  19=>"1111100111110100"&"0001011011010100",
  20=>"1111111111010011"&"0001100010100001",
  21=>"1111110011100110"&"0001001011111011",
  22=>"1111011000001011"&"0001100011111001",
  23=>"1111100001110011"&"0001101001100010",
  24=>"1111100111100101"&"0001111100110001",
  25=>"1111010111001101"&"0001110010100101",
  26=>"1111100000110000"&"0001010111111011",
  27=>"1111010000010010"&"0010000110010100",
  28=>"0000000011010100"&"0001000011000100",
  29=>"1111100011110111"&"0010001000000000",
  30=>"1111101011000100"&"0001110010100000",
  31=>"1111010000101111"&"0001111110100100",
  32=>"1110111100100110"&"0001111111100110",
  33=>"1111001010110100"&"0010010101101101",
  34=>"1111110010111011"&"0001101011000001",
  35=>"1111000000000010"&"0010010110010101",
  36=>"1111100011010001"&"0001101001110010",
  37=>"1111010011101101"&"0001110101010000",
  38=>"1111001110000100"&"0001101100000111",
  39=>"1111000111001101"&"0001110011101011",
  40=>"1111001100101101"&"0010001010000100",
  41=>"1111010010010011"&"0001000110010001",
  42=>"0000000110110010"&"0001010010011001",
  43=>"1111010000111011"&"0001111100001100",
  44=>"1111110010000001"&"0001011111000100",
  45=>"1111110111100010"&"0001101101100100",
  46=>"1111010110000111"&"0001100110101100",
  47=>"1111001111100100"&"0001110011101010",
  48=>"1111011110101001"&"0001111100101100",
  49=>"1111110001010111"&"0000111010111001",
  50=>"1111100000111001"&"0001011011011011",
  51=>"1111001011001101"&"0001110101010000",
  52=>"1111101011010100"&"0001010010011100",
  53=>"1111101000001010"&"0001011101000010",
  54=>"1110111101110001"&"0001101100110101",
  55=>"1111001001101000"&"0010001000000010",
  56=>"1111101101010001"&"0001100011110011",
  57=>"1111011011110101"&"0001101101101010",
  58=>"0000000001100000"&"0000101101110001",
  59=>"1111001111000110"&"0001101000110010",
  60=>"1111110011001001"&"0001001111001000",
  61=>"1111001010100111"&"0001011111010010",
  62=>"1111100000100100"&"0001111101001011",
  63=>"0000000000110100"&"0001000100100011",
  64=>"1110100011010011"&"0010010000111101",
  65=>"1111101011000011"&"0001011100001101",
  66=>"1111100111001010"&"0001101001101101",
  67=>"1111011100011111"&"0001111101111011",
  68=>"1111100110101011"&"0001100110011110",
  69=>"1111101010001110"&"0001001111010111",
  70=>"1111010000111100"&"0001100011001110",
  71=>"1111000010010101"&"0001011000111111",
  72=>"1111100000111010"&"0001101110001011",
  73=>"0000000111011001"&"0001001011101100",
  74=>"1111100011110011"&"0001101001100010",
  75=>"1110110101010101"&"0010011011010011",
  76=>"1111110100111110"&"0001100111100101",
  77=>"1111100011111010"&"0001101010111011",
  78=>"1111011100110000"&"0001100101110111",
  79=>"1111101110110111"&"0001010010110101",
  80=>"1111101000100001"&"0001010000101001",
  81=>"1111100001110000"&"0001111101010010",
  82=>"1110110001100111"&"0001111010001101",
  83=>"1111010000001010"&"0001111000000011",
  84=>"1111110110101110"&"0000111010000101",
  85=>"1111000101100001"&"0001100101000111",
  86=>"1110101001010010"&"0010000110100101",
  87=>"1111110100001111"&"0001001100011010",
  88=>"1111100011011010"&"0001110000100011",
  89=>"1111101011001110"&"0001010000001111",
  90=>"1111101011101010"&"0001110111111100",
  91=>"1111010101001101"&"0001101110100011",
  92=>"1111111110011010"&"0001000000101010",
  93=>"1111100100111100"&"0001001001111100",
  94=>"1111010011101001"&"0010010011001110",
  95=>"1111001010101111"&"0010000011010010",
  96=>"1111111010110000"&"0001100000011001",
  97=>"1111100101010010"&"0001011000000100",
  98=>"1111001001011101"&"0001111000100001",
  99=>"1111100101100010"&"0001000010001111",
  100=>"1111001011011000"&"0001110100101001",
  101=>"1111001000010010"&"0010000001011101",
  102=>"1111011100000000"&"0001100011100000",
  103=>"1111100011101110"&"0001100111101011",
  104=>"1111101010010101"&"0001010100111110",
  105=>"0000000000010111"&"0001011101010110",
  106=>"1111101001001001"&"0001011000010100",
  107=>"1111010110111011"&"0001010010001101",
  108=>"1111010011110000"&"0010000100111100",
  109=>"1111011001001101"&"0001101001111101",
  110=>"1111110101010110"&"0001001110111111",
  111=>"1111011000011000"&"0001011100101000",
  112=>"1111100101010010"&"0001011101011100",
  113=>"1111010010101111"&"0001101110111010",
  114=>"1111110010110010"&"0001010111000000",
  115=>"1111000010110000"&"0010000001101111",
  116=>"1111100101110111"&"0001010010101110",
  117=>"1111100110101001"&"0001100111001001",
  118=>"1111110010010100"&"0001001110001001",
  119=>"1111100011011100"&"0001000011000101",
  120=>"1111100010110110"&"0001100101010110",
  121=>"1111001001100100"&"0010010011101111",
  122=>"1110111110010011"&"0001110100011011",
  123=>"1111110001111011"&"0001000111111011",
  124=>"1111011100110110"&"0001100001110101",
  125=>"1110110010011101"&"0001101000111110",
  126=>"1111001010000111"&"0001101100000010",
  127=>"1111101001001111"&"0000111110101011",
  128=>"1111110101011100"&"0001000110000010",
  129=>"1110111011000101"&"0010000111100011",
  130=>"1111011100011110"&"0001100101101110",
  131=>"1111011111101100"&"0001100111011110",
  132=>"1111101000110001"&"0001100101100110",
  133=>"1110110101011111"&"0001111010110111",
  134=>"1111010110101111"&"0010011101111011",
  135=>"1111100110100001"&"0001010001010100",
  136=>"1111101000100111"&"0001011110000111",
  137=>"1111100110000100"&"0001011101111110",
  138=>"1111110001101111"&"0001001000010001",
  139=>"1111001001110101"&"0001110001010010",
  140=>"1111010100010011"&"0010000011000001",
  141=>"1111110110000101"&"0001011101101101",
  142=>"1110111111011101"&"0010011000101000",
  143=>"1111010010001000"&"0001100001000111",
  144=>"1111111111011100"&"0000110111111010",
  145=>"1111110110001110"&"0001000010110110",
  146=>"1111001011000000"&"0001100001111101",
  147=>"1111000000100000"&"0010000101100100",
  148=>"1111010010101011"&"0001100100010000",
  149=>"1111010111001011"&"0001011101100000",
  150=>"1111101000100001"&"0001000010100001",
  151=>"1111010101110001"&"0001100011011101",
  152=>"1110101011000001"&"0001101111100101",
  153=>"1110111101100111"&"0010100110010000",
  154=>"1111100010000000"&"0001101001111111",
  155=>"1111110101110011"&"0001010111011011",
  156=>"1111010001101011"&"0001111010011000",
  157=>"1110101110000001"&"0010001000000111",
  158=>"1111011000000001"&"0001111000101111",
  159=>"1111101010110100"&"0001011010010100",
  160=>"1111000011011011"&"0001110100010011",
  161=>"1111011100000000"&"0010000000100000",
  162=>"1111111111011110"&"0001000000111010",
  163=>"1111011111111010"&"0001101000011101",
  164=>"1111010001001111"&"0001101011110011",
  165=>"1111001010010011"&"0010001000010101",
  166=>"0000000001001010"&"0001000011001010",
  167=>"1111101110001000"&"0001010110110011",
  168=>"1101100110111011"&"0001110110100010",
  169=>"1111100110110001"&"0000111010111011",
  170=>"1111010000000100"&"0001001110010001",
  171=>"0000000010010110"&"0001001011111001",
  172=>"1111100111101011"&"0001100101111100",
  173=>"1111001110110010"&"0001110111001100",
  174=>"1111011011001010"&"0001111100100110",
  175=>"1111001101010011"&"0001101111111100",
  176=>"1111010011010110"&"0001000101101111",
  177=>"1111100011010111"&"0001110101101111",
  178=>"0000011110011000"&"0001000101010010",
  179=>"1111010110100111"&"0001101011001101",
  180=>"1110111000100001"&"0010000001111110",
  181=>"1111100000010110"&"0001100011110011",
  182=>"1111101111111111"&"0000111011111110",
  183=>"1111010110101110"&"0001110010011001",
  184=>"1110100110001100"&"0010101001000000",
  185=>"1111110000110000"&"0001001100001001",
  186=>"1110111101000111"&"0001100111100000",
  187=>"1111001011001010"&"0001110110110001",
  188=>"1111101011100011"&"0001100000001101",
  189=>"1111101100000100"&"0001101001111100",
  190=>"1110101110110110"&"0010100000000111",
  191=>"1111100110010110"&"0001011100001111",
  192=>"1111101011011100"&"0001100000100101",
  193=>"1111100111100111"&"0001111110001111",
  194=>"1111100000101011"&"0001011011010000",
  195=>"1111010011001000"&"0001011000101011",
  196=>"1111111010100000"&"0001010000010000",
  197=>"1111101111100000"&"0000111001100010",
  198=>"1110111000100110"&"0010010011101001",
  199=>"1111011100000000"&"0001101101011100",
  200=>"1111000001010101"&"0001110100110100",
  201=>"1111011010111101"&"0001011101011111",
  202=>"1110100000100001"&"0010010101011100",
  203=>"1111100000000100"&"0001011010000010",
  204=>"1111010110010100"&"0010000011001001",
  205=>"1111011010101100"&"0001100111001001",
  206=>"1111011110010100"&"0001100000010110",
  207=>"1110111011110011"&"0001011101111101",
  208=>"1111010010000101"&"0001011110110110",
  209=>"1111001111011110"&"0001100110111100",
  210=>"1111100000010011"&"0001011100110110",
  211=>"1111011110000000"&"0001010000010101",
  212=>"1111110000011001"&"0001011100001110",
  213=>"1111100100100000"&"0010001000010000",
  214=>"1111100110000110"&"0001000011111111",
  215=>"1110101001010100"&"0010011101001110",
  216=>"1111011110010100"&"0001101100001000",
  217=>"1110010101000100"&"0010101000101001",
  218=>"1111011110111001"&"0001010100100110",
  219=>"1111011010100001"&"0001101010000000",
  220=>"1111010010111100"&"0001110010101110",
  221=>"1110101100011100"&"0001111111001100",
  222=>"0000001100000011"&"0000111101101001",
  223=>"1110111101111100"&"0001110010110010",
  224=>"1111111100110000"&"0000111011110011",
  225=>"1111101001001110"&"0001010111010001",
  226=>"1111001110110110"&"0001110010110100",
  227=>"1111011101111000"&"0001100001010001",
  228=>"1111001000101110"&"0001111001011101",
  229=>"1111011001110011"&"0001111100000001",
  230=>"1111010010010101"&"0010000011100111",
  231=>"1111001000000101"&"0010000101100110",
  232=>"1111011101010000"&"0001101110011111",
  233=>"1111101001001110"&"0001011101100000",
  234=>"1111011010001101"&"0010000100111001",
  235=>"1111001010000011"&"0001111101111011",
  236=>"1111111101001010"&"0000111111100011",
  237=>"1111100111111010"&"0001010000011011",
  238=>"1111110101101101"&"0001100001011000",
  239=>"1111101000011101"&"0001010001111000",
  240=>"1111010001001010"&"0010001110101010",
  241=>"1111001100010100"&"0001110011100000",
  242=>"1111010101011110"&"0001101010011101",
  243=>"1111001101001100"&"0001100100001000",
  244=>"1111011001010001"&"0001101101010110",
  245=>"1110101110010111"&"0010010110110101",
  246=>"1111110010010111"&"0001100011001110",
  247=>"1111100101111001"&"0001100000011111",
  248=>"1111011111100001"&"0001010011111010",
  249=>"1111100101001000"&"0001001010000111",
  250=>"1111011010000000"&"0001000001010000",
  251=>"1111011100000000"&"0001011100100100",
  252=>"1111011100111110"&"0001101100111110",
  253=>"1110110100101011"&"0010000001001001",
  254=>"1111100110111010"&"0001011010000000",
  255=>"1110110100000011"&"0010011001111100");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;