LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_10_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_10_WROM;

ARCHITECTURE RTL OF L8_10_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"000010110",
  1=>"010101110",
  2=>"010000110",
  3=>"100111110",
  4=>"011011101",
  5=>"001111010",
  6=>"011110101",
  7=>"011110000",
  8=>"011001100",
  9=>"100110011",
  10=>"111000110",
  11=>"101101000",
  12=>"001110110",
  13=>"001100010",
  14=>"000110010",
  15=>"011001011",
  16=>"000001000",
  17=>"000011001",
  18=>"110110100",
  19=>"101000110",
  20=>"010001100",
  21=>"111000100",
  22=>"111101110",
  23=>"100010001",
  24=>"000110100",
  25=>"100000101",
  26=>"100001000",
  27=>"011011111",
  28=>"101100001",
  29=>"000110010",
  30=>"011100010",
  31=>"001110010",
  32=>"010010011",
  33=>"001101011",
  34=>"101001010",
  35=>"011000100",
  36=>"001011110",
  37=>"001001100",
  38=>"101011100",
  39=>"000001011",
  40=>"000011011",
  41=>"110001001",
  42=>"101100000",
  43=>"011110001",
  44=>"000000000",
  45=>"000111010",
  46=>"100001001",
  47=>"001101101",
  48=>"011010100",
  49=>"111110011",
  50=>"111110010",
  51=>"001110110",
  52=>"101011010",
  53=>"011111101",
  54=>"011110011",
  55=>"111111111",
  56=>"111011110",
  57=>"011001110",
  58=>"110101000",
  59=>"100101011",
  60=>"100001001",
  61=>"100001010",
  62=>"000100111",
  63=>"000000101",
  64=>"010000010",
  65=>"000010100",
  66=>"110000000",
  67=>"001101100",
  68=>"010010011",
  69=>"111011111",
  70=>"101001000",
  71=>"111110000",
  72=>"110011010",
  73=>"100000101",
  74=>"101111111",
  75=>"010001011",
  76=>"011001001",
  77=>"110010011",
  78=>"111111111",
  79=>"101100110",
  80=>"110100101",
  81=>"100100110",
  82=>"001000100",
  83=>"100000000",
  84=>"010011011",
  85=>"011000011",
  86=>"001000100",
  87=>"101101101",
  88=>"001010110",
  89=>"001100011",
  90=>"110110010",
  91=>"010100001",
  92=>"101111000",
  93=>"101101110",
  94=>"000000101",
  95=>"010101000",
  96=>"011000001",
  97=>"001000100",
  98=>"000000001",
  99=>"111000111",
  100=>"001001100",
  101=>"001001100",
  102=>"110111010",
  103=>"011001000",
  104=>"000001100",
  105=>"101101110",
  106=>"110100110",
  107=>"000000011",
  108=>"100110010",
  109=>"001001100",
  110=>"100100001",
  111=>"000011011",
  112=>"000101110",
  113=>"001101100",
  114=>"100010101",
  115=>"000011000",
  116=>"001010000",
  117=>"110100010",
  118=>"000000101",
  119=>"110111100",
  120=>"110001000",
  121=>"011111000",
  122=>"001001010",
  123=>"010011110",
  124=>"100100110",
  125=>"110101101",
  126=>"010010000",
  127=>"001111111",
  128=>"101111011",
  129=>"001011101",
  130=>"101101001",
  131=>"000010110",
  132=>"001100100",
  133=>"001111111",
  134=>"110111111",
  135=>"010011010",
  136=>"101110010",
  137=>"000100010",
  138=>"100000011",
  139=>"101010111",
  140=>"101100101",
  141=>"001000101",
  142=>"101111011",
  143=>"010000101",
  144=>"000001110",
  145=>"000101111",
  146=>"100000101",
  147=>"000000111",
  148=>"010111011",
  149=>"100010001",
  150=>"110001100",
  151=>"011110001",
  152=>"100101001",
  153=>"111011111",
  154=>"010111001",
  155=>"110101000",
  156=>"000010001",
  157=>"101100100",
  158=>"010010000",
  159=>"100111011",
  160=>"000001000",
  161=>"111100001",
  162=>"110001000",
  163=>"111000111",
  164=>"111001000",
  165=>"000010000",
  166=>"100001101",
  167=>"001000100",
  168=>"000101010",
  169=>"010110010",
  170=>"110101001",
  171=>"001010000",
  172=>"100010010",
  173=>"110111000",
  174=>"110110011",
  175=>"110110100",
  176=>"001010001",
  177=>"000001010",
  178=>"100010001",
  179=>"100100100",
  180=>"100110110",
  181=>"110010000",
  182=>"000000001",
  183=>"110111110",
  184=>"001101100",
  185=>"001011100",
  186=>"001000011",
  187=>"110011011",
  188=>"111110100",
  189=>"110001001",
  190=>"100001101",
  191=>"000100111",
  192=>"111011011",
  193=>"111100110",
  194=>"001010001",
  195=>"101001001",
  196=>"010100110",
  197=>"110001000",
  198=>"000000101",
  199=>"001111011",
  200=>"001100111",
  201=>"011100001",
  202=>"111010001",
  203=>"100101010",
  204=>"111000001",
  205=>"001110000",
  206=>"110010101",
  207=>"111110110",
  208=>"011101101",
  209=>"011001010",
  210=>"110110000",
  211=>"001101001",
  212=>"111000011",
  213=>"001011100",
  214=>"101111100",
  215=>"111100011",
  216=>"100100111",
  217=>"000010010",
  218=>"010101000",
  219=>"010100001",
  220=>"010011001",
  221=>"111101010",
  222=>"110000001",
  223=>"100111011",
  224=>"010100010",
  225=>"010011000",
  226=>"101100101",
  227=>"100001100",
  228=>"110011011",
  229=>"001010011",
  230=>"011000011",
  231=>"000100101",
  232=>"101111011",
  233=>"100111010",
  234=>"101000111",
  235=>"101100101",
  236=>"001001111",
  237=>"101010110",
  238=>"001101110",
  239=>"000111001",
  240=>"001001101",
  241=>"110000000",
  242=>"000011110",
  243=>"011001001",
  244=>"111011110",
  245=>"110011001",
  246=>"110000111",
  247=>"100001001",
  248=>"011000011",
  249=>"000110001",
  250=>"100111100",
  251=>"010010101",
  252=>"100110110",
  253=>"010100101",
  254=>"110001111",
  255=>"101010111",
  256=>"110110100",
  257=>"000010000",
  258=>"011111011",
  259=>"001010010",
  260=>"000110110",
  261=>"100000011",
  262=>"011110000",
  263=>"101000111",
  264=>"011011111",
  265=>"001000111",
  266=>"101001110",
  267=>"000101110",
  268=>"110110010",
  269=>"110111010",
  270=>"111010010",
  271=>"110011000",
  272=>"111000010",
  273=>"001110100",
  274=>"110001011",
  275=>"011110011",
  276=>"111111110",
  277=>"011100110",
  278=>"111011100",
  279=>"010001011",
  280=>"101110000",
  281=>"010001001",
  282=>"100010100",
  283=>"000000101",
  284=>"010111100",
  285=>"101000100",
  286=>"110101101",
  287=>"000001011",
  288=>"110101111",
  289=>"100111011",
  290=>"110101101",
  291=>"111100010",
  292=>"111101101",
  293=>"110001100",
  294=>"010010111",
  295=>"100000100",
  296=>"001110011",
  297=>"011101111",
  298=>"000100101",
  299=>"100010100",
  300=>"011010001",
  301=>"100111010",
  302=>"011101100",
  303=>"001001000",
  304=>"101001000",
  305=>"101001010",
  306=>"111111110",
  307=>"000001000",
  308=>"000011001",
  309=>"001000010",
  310=>"100011111",
  311=>"100000101",
  312=>"001000110",
  313=>"000010001",
  314=>"111000000",
  315=>"011000001",
  316=>"010100111",
  317=>"000000000",
  318=>"011001011",
  319=>"101011110",
  320=>"011101001",
  321=>"000010001",
  322=>"110101110",
  323=>"111110000",
  324=>"011000000",
  325=>"100001010",
  326=>"110001001",
  327=>"110010000",
  328=>"011001101",
  329=>"111110001",
  330=>"101110000",
  331=>"001110011",
  332=>"101111110",
  333=>"010111000",
  334=>"100011100",
  335=>"101000000",
  336=>"011011100",
  337=>"111110111",
  338=>"010010001",
  339=>"001010011",
  340=>"010100101",
  341=>"111111100",
  342=>"001010101",
  343=>"011011001",
  344=>"101100110",
  345=>"010101000",
  346=>"110011100",
  347=>"000000110",
  348=>"011010100",
  349=>"010000000",
  350=>"100001110",
  351=>"010111000",
  352=>"111001101",
  353=>"010110110",
  354=>"010110111",
  355=>"001101101",
  356=>"110011100",
  357=>"011001100",
  358=>"100110111",
  359=>"010001001",
  360=>"101001110",
  361=>"000000010",
  362=>"010011011",
  363=>"010110011",
  364=>"110101000",
  365=>"101010001",
  366=>"100000000",
  367=>"111001100",
  368=>"010001010",
  369=>"101110001",
  370=>"111100111",
  371=>"000010111",
  372=>"000001110",
  373=>"001110101",
  374=>"010110000",
  375=>"110000100",
  376=>"100111001",
  377=>"010110010",
  378=>"100111110",
  379=>"011111110",
  380=>"010001000",
  381=>"010110101",
  382=>"111010111",
  383=>"001001101",
  384=>"010101110",
  385=>"110010110",
  386=>"001001010",
  387=>"100000110",
  388=>"000101111",
  389=>"010000101",
  390=>"100100010",
  391=>"100010001",
  392=>"000000111",
  393=>"011100100",
  394=>"111010011",
  395=>"100101111",
  396=>"011111101",
  397=>"100010101",
  398=>"101101101",
  399=>"111111010",
  400=>"101111111",
  401=>"001000101",
  402=>"101011001",
  403=>"100010000",
  404=>"100000011",
  405=>"010000000",
  406=>"111101111",
  407=>"011110001",
  408=>"001111100",
  409=>"001111100",
  410=>"000011010",
  411=>"010011011",
  412=>"111110011",
  413=>"000001001",
  414=>"000101111",
  415=>"110111011",
  416=>"111111001",
  417=>"110110101",
  418=>"100110001",
  419=>"000100000",
  420=>"110001000",
  421=>"011011001",
  422=>"000001000",
  423=>"100111010",
  424=>"101111110",
  425=>"000010101",
  426=>"010010111",
  427=>"010111000",
  428=>"010110000",
  429=>"010010110",
  430=>"111000100",
  431=>"100100110",
  432=>"010000101",
  433=>"111100011",
  434=>"011000100",
  435=>"101001110",
  436=>"100100100",
  437=>"110011110",
  438=>"001001010",
  439=>"000010000",
  440=>"101100001",
  441=>"101000111",
  442=>"110000000",
  443=>"110101011",
  444=>"101010000",
  445=>"100010100",
  446=>"000000000",
  447=>"110010000",
  448=>"101011101",
  449=>"111011101",
  450=>"101001010",
  451=>"100111001",
  452=>"111111010",
  453=>"011111110",
  454=>"000110010",
  455=>"000001001",
  456=>"100010111",
  457=>"101011001",
  458=>"010001001",
  459=>"010101011",
  460=>"010111110",
  461=>"110000010",
  462=>"001100101",
  463=>"100000101",
  464=>"101111111",
  465=>"100001000",
  466=>"010100011",
  467=>"110000100",
  468=>"001001000",
  469=>"010010011",
  470=>"001011001",
  471=>"100110111",
  472=>"010111011",
  473=>"011001001",
  474=>"111010101",
  475=>"111000101",
  476=>"101010110",
  477=>"111001010",
  478=>"011011100",
  479=>"110011010",
  480=>"100101000",
  481=>"101011100",
  482=>"101111110",
  483=>"011000000",
  484=>"011100111",
  485=>"110000111",
  486=>"010101010",
  487=>"000001000",
  488=>"011001001",
  489=>"101100110",
  490=>"100110001",
  491=>"001011000",
  492=>"110000111",
  493=>"010101100",
  494=>"010110110",
  495=>"010100110",
  496=>"011001110",
  497=>"111010101",
  498=>"101001000",
  499=>"111101100",
  500=>"000100000",
  501=>"001101000",
  502=>"111110111",
  503=>"011000110",
  504=>"011001111",
  505=>"110000000",
  506=>"101101010",
  507=>"101001111",
  508=>"111100101",
  509=>"010110100",
  510=>"101100111",
  511=>"011000000",
  512=>"100000001",
  513=>"110111110",
  514=>"000011110",
  515=>"001001000",
  516=>"100111110",
  517=>"000110101",
  518=>"101000100",
  519=>"010101000",
  520=>"010101101",
  521=>"101011100",
  522=>"110000101",
  523=>"010101000",
  524=>"110000010",
  525=>"010000111",
  526=>"100101110",
  527=>"111110001",
  528=>"110010100",
  529=>"010011010",
  530=>"011001100",
  531=>"001110001",
  532=>"011101101",
  533=>"010011000",
  534=>"100001111",
  535=>"001101001",
  536=>"111000000",
  537=>"010011111",
  538=>"011011100",
  539=>"010000010",
  540=>"111111000",
  541=>"111000000",
  542=>"000001010",
  543=>"011101100",
  544=>"000000011",
  545=>"101001000",
  546=>"000011010",
  547=>"100001010",
  548=>"111011011",
  549=>"000001111",
  550=>"010110111",
  551=>"110110100",
  552=>"101100110",
  553=>"100000000",
  554=>"100011111",
  555=>"101000100",
  556=>"010110111",
  557=>"111001010",
  558=>"000001100",
  559=>"000001100",
  560=>"111011110",
  561=>"101010010",
  562=>"000001000",
  563=>"000100111",
  564=>"001100001",
  565=>"010101101",
  566=>"001110000",
  567=>"010001010",
  568=>"010100010",
  569=>"000111101",
  570=>"001100111",
  571=>"110011110",
  572=>"100100001",
  573=>"011100001",
  574=>"110001001",
  575=>"100101000",
  576=>"100010000",
  577=>"011010000",
  578=>"001000110",
  579=>"000001111",
  580=>"101001100",
  581=>"010111101",
  582=>"111000011",
  583=>"010101111",
  584=>"010011111",
  585=>"011011110",
  586=>"001111011",
  587=>"100101110",
  588=>"001011111",
  589=>"010011001",
  590=>"110110001",
  591=>"000101000",
  592=>"000010100",
  593=>"001001000",
  594=>"100100011",
  595=>"000111010",
  596=>"001110110",
  597=>"010001101",
  598=>"011011011",
  599=>"100010110",
  600=>"111001111",
  601=>"011111000",
  602=>"100000111",
  603=>"000010100",
  604=>"100000000",
  605=>"000101010",
  606=>"001010110",
  607=>"110101000",
  608=>"110101000",
  609=>"100001010",
  610=>"010000100",
  611=>"010001000",
  612=>"000001100",
  613=>"100011000",
  614=>"010101110",
  615=>"111111001",
  616=>"110111010",
  617=>"111000110",
  618=>"010111011",
  619=>"111101101",
  620=>"001100010",
  621=>"100000001",
  622=>"000101010",
  623=>"111101000",
  624=>"101100001",
  625=>"001110001",
  626=>"001010101",
  627=>"111000010",
  628=>"000101100",
  629=>"100000000",
  630=>"101001001",
  631=>"000000011",
  632=>"000000111",
  633=>"101110100",
  634=>"000101011",
  635=>"001000011",
  636=>"101111011",
  637=>"001000100",
  638=>"110110001",
  639=>"101101010",
  640=>"000010001",
  641=>"001110100",
  642=>"010011100",
  643=>"010000101",
  644=>"100010001",
  645=>"000110010",
  646=>"011010011",
  647=>"101100101",
  648=>"110101010",
  649=>"000101011",
  650=>"111010110",
  651=>"011010000",
  652=>"000010001",
  653=>"000001001",
  654=>"100100001",
  655=>"110010000",
  656=>"111100010",
  657=>"011001001",
  658=>"010001101",
  659=>"010110110",
  660=>"110011111",
  661=>"101111101",
  662=>"110111100",
  663=>"001101101",
  664=>"101101111",
  665=>"000100110",
  666=>"111011011",
  667=>"100111111",
  668=>"100001100",
  669=>"010011011",
  670=>"110101111",
  671=>"110010010",
  672=>"010010001",
  673=>"001000111",
  674=>"010100011",
  675=>"000111011",
  676=>"001000110",
  677=>"110111110",
  678=>"100001101",
  679=>"000011101",
  680=>"110111100",
  681=>"010101000",
  682=>"010000010",
  683=>"000111111",
  684=>"111001000",
  685=>"101101100",
  686=>"010010110",
  687=>"101000111",
  688=>"011110100",
  689=>"000100111",
  690=>"000011110",
  691=>"011100010",
  692=>"000110011",
  693=>"100101100",
  694=>"100111101",
  695=>"011100011",
  696=>"001011100",
  697=>"100010011",
  698=>"010001111",
  699=>"011100111",
  700=>"011100111",
  701=>"010000000",
  702=>"011000111",
  703=>"111111110",
  704=>"101111011",
  705=>"101011100",
  706=>"000011010",
  707=>"101100111",
  708=>"000000011",
  709=>"000010011",
  710=>"110000100",
  711=>"100000010",
  712=>"010000101",
  713=>"111010011",
  714=>"111101110",
  715=>"010000100",
  716=>"011001100",
  717=>"101111011",
  718=>"001111101",
  719=>"100001100",
  720=>"101110001",
  721=>"011110111",
  722=>"000000001",
  723=>"000000100",
  724=>"111111111",
  725=>"000000011",
  726=>"001010111",
  727=>"110000101",
  728=>"000111010",
  729=>"010000010",
  730=>"011111001",
  731=>"001000100",
  732=>"101011100",
  733=>"001001110",
  734=>"001011010",
  735=>"010011011",
  736=>"000000000",
  737=>"100011010",
  738=>"111101011",
  739=>"010000011",
  740=>"010011000",
  741=>"111001111",
  742=>"100100000",
  743=>"000001101",
  744=>"010011011",
  745=>"010000001",
  746=>"110100100",
  747=>"100000110",
  748=>"001111001",
  749=>"110011111",
  750=>"110100111",
  751=>"110111010",
  752=>"011011010",
  753=>"011000001",
  754=>"101000110",
  755=>"001111110",
  756=>"100111111",
  757=>"001100110",
  758=>"101010001",
  759=>"111101101",
  760=>"110001001",
  761=>"111111111",
  762=>"110011000",
  763=>"100000100",
  764=>"110110011",
  765=>"110000101",
  766=>"110111001",
  767=>"001010100",
  768=>"100001000",
  769=>"111000001",
  770=>"101101010",
  771=>"111010100",
  772=>"101110010",
  773=>"010010111",
  774=>"101001110",
  775=>"110001100",
  776=>"111000001",
  777=>"101010000",
  778=>"100111001",
  779=>"110011110",
  780=>"000011001",
  781=>"001101111",
  782=>"001001101",
  783=>"000001111",
  784=>"111000010",
  785=>"100111111",
  786=>"101010001",
  787=>"110010010",
  788=>"101100011",
  789=>"110001010",
  790=>"010010011",
  791=>"001111011",
  792=>"011101001",
  793=>"010010101",
  794=>"001011011",
  795=>"010000101",
  796=>"000000111",
  797=>"111001001",
  798=>"010010011",
  799=>"111110110",
  800=>"000111000",
  801=>"000001101",
  802=>"000101111",
  803=>"011001101",
  804=>"010011100",
  805=>"110011111",
  806=>"101001111",
  807=>"001010000",
  808=>"010011001",
  809=>"010101101",
  810=>"101111011",
  811=>"111100000",
  812=>"010110010",
  813=>"001001010",
  814=>"010101010",
  815=>"010110010",
  816=>"010101100",
  817=>"101000000",
  818=>"100101001",
  819=>"101001100",
  820=>"110111000",
  821=>"011100001",
  822=>"011011000",
  823=>"110001010",
  824=>"001100010",
  825=>"001101001",
  826=>"001000101",
  827=>"110110001",
  828=>"001111100",
  829=>"110101111",
  830=>"001100001",
  831=>"001110001",
  832=>"110010100",
  833=>"001101101",
  834=>"101100011",
  835=>"110011011",
  836=>"001101001",
  837=>"010111101",
  838=>"111101101",
  839=>"110010111",
  840=>"010001010",
  841=>"001101100",
  842=>"101010010",
  843=>"100000100",
  844=>"110010011",
  845=>"010000101",
  846=>"101001110",
  847=>"101001011",
  848=>"100000000",
  849=>"000001001",
  850=>"111010111",
  851=>"000001100",
  852=>"111101000",
  853=>"101111100",
  854=>"000111001",
  855=>"011010111",
  856=>"111111111",
  857=>"001011111",
  858=>"101001100",
  859=>"010000001",
  860=>"011100100",
  861=>"101001101",
  862=>"000011011",
  863=>"001001011",
  864=>"100111001",
  865=>"100111110",
  866=>"101011110",
  867=>"111001101",
  868=>"001001001",
  869=>"110000110",
  870=>"001011100",
  871=>"100111011",
  872=>"001001100",
  873=>"011000010",
  874=>"100001011",
  875=>"101111111",
  876=>"000111001",
  877=>"000001111",
  878=>"010010000",
  879=>"101000101",
  880=>"000011000",
  881=>"011000101",
  882=>"110110101",
  883=>"111100101",
  884=>"111101000",
  885=>"110111111",
  886=>"011111101",
  887=>"101110100",
  888=>"111101111",
  889=>"110010110",
  890=>"111010101",
  891=>"010101101",
  892=>"001110001",
  893=>"101000011",
  894=>"010100001",
  895=>"110110010",
  896=>"100101000",
  897=>"101111000",
  898=>"100101101",
  899=>"111010000",
  900=>"010000000",
  901=>"111110001",
  902=>"001100101",
  903=>"101111011",
  904=>"111011010",
  905=>"011111001",
  906=>"101010111",
  907=>"001111000",
  908=>"001110110",
  909=>"101000110",
  910=>"100101001",
  911=>"111101010",
  912=>"111100110",
  913=>"001000001",
  914=>"101001100",
  915=>"110011110",
  916=>"101001011",
  917=>"111111100",
  918=>"000111110",
  919=>"101100111",
  920=>"110000101",
  921=>"111111011",
  922=>"000010010",
  923=>"100011000",
  924=>"010011000",
  925=>"011101001",
  926=>"000010001",
  927=>"000001001",
  928=>"001111000",
  929=>"001010111",
  930=>"101100110",
  931=>"100000010",
  932=>"001111010",
  933=>"001001000",
  934=>"010110111",
  935=>"110011100",
  936=>"001111110",
  937=>"110000011",
  938=>"000101001",
  939=>"011000100",
  940=>"100111000",
  941=>"001011011",
  942=>"011111111",
  943=>"011111111",
  944=>"110110000",
  945=>"011110110",
  946=>"110001111",
  947=>"111101101",
  948=>"001011111",
  949=>"000000000",
  950=>"011110101",
  951=>"101100101",
  952=>"000101011",
  953=>"011101010",
  954=>"111011010",
  955=>"011001010",
  956=>"011101001",
  957=>"011111011",
  958=>"010101000",
  959=>"111011110",
  960=>"101110001",
  961=>"001101110",
  962=>"110111011",
  963=>"011101011",
  964=>"111000011",
  965=>"010000100",
  966=>"010010100",
  967=>"110000110",
  968=>"010111110",
  969=>"100101010",
  970=>"000000100",
  971=>"101001101",
  972=>"111111111",
  973=>"110111000",
  974=>"001001000",
  975=>"100010101",
  976=>"100000011",
  977=>"100100000",
  978=>"111111110",
  979=>"011110011",
  980=>"000000001",
  981=>"110001011",
  982=>"100010001",
  983=>"010000010",
  984=>"001110100",
  985=>"101000101",
  986=>"010000101",
  987=>"010111010",
  988=>"010011001",
  989=>"011011011",
  990=>"100000111",
  991=>"001100100",
  992=>"110011111",
  993=>"001010100",
  994=>"100100010",
  995=>"111100100",
  996=>"100010000",
  997=>"000110011",
  998=>"011010111",
  999=>"101001011",
  1000=>"010101000",
  1001=>"111011100",
  1002=>"101010010",
  1003=>"101111000",
  1004=>"101110001",
  1005=>"110011110",
  1006=>"111111111",
  1007=>"011100110",
  1008=>"101100101",
  1009=>"100110110",
  1010=>"101000010",
  1011=>"000101001",
  1012=>"001111111",
  1013=>"101110010",
  1014=>"110000111",
  1015=>"011101001",
  1016=>"000100101",
  1017=>"101001011",
  1018=>"111111110",
  1019=>"110101000",
  1020=>"010011100",
  1021=>"010001001",
  1022=>"000011010",
  1023=>"110101101",
  1024=>"101010001",
  1025=>"001110100",
  1026=>"110100110",
  1027=>"111111011",
  1028=>"100001000",
  1029=>"111010000",
  1030=>"110000111",
  1031=>"111001010",
  1032=>"010110111",
  1033=>"010001110",
  1034=>"000000000",
  1035=>"000010101",
  1036=>"100100111",
  1037=>"000111101",
  1038=>"010101110",
  1039=>"101001010",
  1040=>"111000010",
  1041=>"110110100",
  1042=>"100010100",
  1043=>"110101100",
  1044=>"001000100",
  1045=>"100010000",
  1046=>"110110010",
  1047=>"001010001",
  1048=>"111100000",
  1049=>"010100111",
  1050=>"100001100",
  1051=>"110000010",
  1052=>"011101010",
  1053=>"010011011",
  1054=>"010001111",
  1055=>"110010011",
  1056=>"110011100",
  1057=>"000001010",
  1058=>"000101000",
  1059=>"111000111",
  1060=>"000111010",
  1061=>"101000001",
  1062=>"111010010",
  1063=>"100011000",
  1064=>"000001110",
  1065=>"000100011",
  1066=>"001111110",
  1067=>"001111100",
  1068=>"111100011",
  1069=>"001000000",
  1070=>"101110001",
  1071=>"000011001",
  1072=>"101010111",
  1073=>"001110101",
  1074=>"100110100",
  1075=>"101111100",
  1076=>"100010010",
  1077=>"001001000",
  1078=>"001101111",
  1079=>"110010100",
  1080=>"100011000",
  1081=>"001011111",
  1082=>"100000111",
  1083=>"101000000",
  1084=>"110011101",
  1085=>"000011101",
  1086=>"010011011",
  1087=>"000011101",
  1088=>"010110100",
  1089=>"000001111",
  1090=>"010011000",
  1091=>"110010000",
  1092=>"100111010",
  1093=>"011111011",
  1094=>"000110011",
  1095=>"100101101",
  1096=>"000000001",
  1097=>"101011111",
  1098=>"101110000",
  1099=>"110001100",
  1100=>"110111010",
  1101=>"010010111",
  1102=>"110111011",
  1103=>"010010001",
  1104=>"001010010",
  1105=>"101110110",
  1106=>"100100001",
  1107=>"010111000",
  1108=>"111110110",
  1109=>"111101111",
  1110=>"110101111",
  1111=>"100110111",
  1112=>"010011110",
  1113=>"001011111",
  1114=>"111001101",
  1115=>"110010010",
  1116=>"010001011",
  1117=>"100111101",
  1118=>"110010101",
  1119=>"001001110",
  1120=>"111000001",
  1121=>"000011000",
  1122=>"001001000",
  1123=>"111100101",
  1124=>"100010010",
  1125=>"000101011",
  1126=>"011000000",
  1127=>"101110101",
  1128=>"011101000",
  1129=>"101010001",
  1130=>"110111001",
  1131=>"001011100",
  1132=>"100111100",
  1133=>"111111000",
  1134=>"100011010",
  1135=>"110110001",
  1136=>"100011010",
  1137=>"111111111",
  1138=>"010010010",
  1139=>"111111111",
  1140=>"010110000",
  1141=>"111011101",
  1142=>"011000000",
  1143=>"110110011",
  1144=>"000111111",
  1145=>"111010101",
  1146=>"011010000",
  1147=>"000110001",
  1148=>"111101111",
  1149=>"001101100",
  1150=>"010001000",
  1151=>"101101100",
  1152=>"011110111",
  1153=>"000010110",
  1154=>"011001011",
  1155=>"111111101",
  1156=>"110011101",
  1157=>"110010101",
  1158=>"111100101",
  1159=>"000011011",
  1160=>"100101111",
  1161=>"111000011",
  1162=>"010000000",
  1163=>"001011000",
  1164=>"011100110",
  1165=>"110100110",
  1166=>"111011101",
  1167=>"111110000",
  1168=>"111111010",
  1169=>"001000110",
  1170=>"100001011",
  1171=>"101111101",
  1172=>"010001010",
  1173=>"111100000",
  1174=>"111011010",
  1175=>"101110110",
  1176=>"001010010",
  1177=>"011110100",
  1178=>"100010101",
  1179=>"001000010",
  1180=>"111001010",
  1181=>"010000101",
  1182=>"001001010",
  1183=>"000011001",
  1184=>"100010101",
  1185=>"001101100",
  1186=>"001110001",
  1187=>"110100000",
  1188=>"010110111",
  1189=>"110101100",
  1190=>"101110101",
  1191=>"000011001",
  1192=>"110000101",
  1193=>"001101111",
  1194=>"100011111",
  1195=>"101101110",
  1196=>"100111001",
  1197=>"001000011",
  1198=>"001101110",
  1199=>"101100111",
  1200=>"000000000",
  1201=>"101001111",
  1202=>"100110101",
  1203=>"100011111",
  1204=>"010101100",
  1205=>"011000001",
  1206=>"110000000",
  1207=>"111111011",
  1208=>"101011110",
  1209=>"000100011",
  1210=>"111101111",
  1211=>"010110110",
  1212=>"110000101",
  1213=>"111100100",
  1214=>"000000011",
  1215=>"010101000",
  1216=>"101110111",
  1217=>"000110011",
  1218=>"001010011",
  1219=>"010010010",
  1220=>"111000110",
  1221=>"100100001",
  1222=>"010010000",
  1223=>"100100110",
  1224=>"001000110",
  1225=>"111101000",
  1226=>"000100010",
  1227=>"011010001",
  1228=>"010111110",
  1229=>"110001101",
  1230=>"000010000",
  1231=>"000101001",
  1232=>"010010000",
  1233=>"111110000",
  1234=>"000011110",
  1235=>"101000000",
  1236=>"010110101",
  1237=>"000111001",
  1238=>"101111010",
  1239=>"101110011",
  1240=>"000011001",
  1241=>"001101111",
  1242=>"010001101",
  1243=>"000011111",
  1244=>"100101000",
  1245=>"011101000",
  1246=>"100010111",
  1247=>"101101110",
  1248=>"000110010",
  1249=>"111010100",
  1250=>"100000011",
  1251=>"100011101",
  1252=>"001101000",
  1253=>"111010000",
  1254=>"101011100",
  1255=>"011111000",
  1256=>"110011110",
  1257=>"010000100",
  1258=>"110000110",
  1259=>"100110011",
  1260=>"010111100",
  1261=>"010010110",
  1262=>"100110000",
  1263=>"100010011",
  1264=>"010011100",
  1265=>"110110000",
  1266=>"111001001",
  1267=>"011000011",
  1268=>"010111110",
  1269=>"001111011",
  1270=>"100110000",
  1271=>"111110100",
  1272=>"010110100",
  1273=>"100100101",
  1274=>"110011111",
  1275=>"100011011",
  1276=>"010111110",
  1277=>"111110110",
  1278=>"111011011",
  1279=>"011000011",
  1280=>"001001101",
  1281=>"000011100",
  1282=>"111011000",
  1283=>"100011011",
  1284=>"000111110",
  1285=>"101100100",
  1286=>"111101110",
  1287=>"000011011",
  1288=>"110101101",
  1289=>"010000001",
  1290=>"101101100",
  1291=>"010011000",
  1292=>"100100011",
  1293=>"001000100",
  1294=>"101011001",
  1295=>"001000110",
  1296=>"101111110",
  1297=>"111111110",
  1298=>"100111101",
  1299=>"110111101",
  1300=>"111100001",
  1301=>"011101111",
  1302=>"001010110",
  1303=>"011101010",
  1304=>"101111101",
  1305=>"001101011",
  1306=>"101010110",
  1307=>"000011100",
  1308=>"100110001",
  1309=>"011111010",
  1310=>"110101010",
  1311=>"110010001",
  1312=>"010010110",
  1313=>"001001001",
  1314=>"101010011",
  1315=>"100101011",
  1316=>"001011011",
  1317=>"001001101",
  1318=>"001000010",
  1319=>"011000010",
  1320=>"111010000",
  1321=>"010111110",
  1322=>"001001010",
  1323=>"111111111",
  1324=>"110010110",
  1325=>"010010000",
  1326=>"010010100",
  1327=>"010111101",
  1328=>"010010001",
  1329=>"000000011",
  1330=>"111101111",
  1331=>"111100000",
  1332=>"000011010",
  1333=>"001011010",
  1334=>"110110110",
  1335=>"101101011",
  1336=>"101111011",
  1337=>"010011010",
  1338=>"100100000",
  1339=>"100010010",
  1340=>"111001101",
  1341=>"110111101",
  1342=>"101001011",
  1343=>"011110000",
  1344=>"001111000",
  1345=>"111111111",
  1346=>"011001100",
  1347=>"011000001",
  1348=>"101101011",
  1349=>"100110000",
  1350=>"011111000",
  1351=>"101010010",
  1352=>"010011100",
  1353=>"111001010",
  1354=>"101011101",
  1355=>"100001000",
  1356=>"011111101",
  1357=>"000000010",
  1358=>"110010010",
  1359=>"010111011",
  1360=>"001111000",
  1361=>"100101001",
  1362=>"110101111",
  1363=>"000011110",
  1364=>"010111111",
  1365=>"100000010",
  1366=>"010101010",
  1367=>"101001110",
  1368=>"011100100",
  1369=>"010010110",
  1370=>"001100100",
  1371=>"110111010",
  1372=>"010110000",
  1373=>"010000010",
  1374=>"110000110",
  1375=>"111101100",
  1376=>"111010000",
  1377=>"010111001",
  1378=>"010110011",
  1379=>"000010100",
  1380=>"100000001",
  1381=>"110110001",
  1382=>"000001011",
  1383=>"011111110",
  1384=>"011011011",
  1385=>"011000101",
  1386=>"011000100",
  1387=>"111011111",
  1388=>"100001010",
  1389=>"000010010",
  1390=>"101100100",
  1391=>"110100011",
  1392=>"010010101",
  1393=>"101000001",
  1394=>"100101111",
  1395=>"000100110",
  1396=>"000001001",
  1397=>"011100110",
  1398=>"001000100",
  1399=>"101010000",
  1400=>"001001000",
  1401=>"011001000",
  1402=>"001101001",
  1403=>"111111101",
  1404=>"100001100",
  1405=>"100001110",
  1406=>"100010010",
  1407=>"100100110",
  1408=>"101111010",
  1409=>"011000101",
  1410=>"111100001",
  1411=>"010100101",
  1412=>"101100111",
  1413=>"100101000",
  1414=>"101010011",
  1415=>"100110010",
  1416=>"111010000",
  1417=>"110100010",
  1418=>"111110101",
  1419=>"001010001",
  1420=>"001010101",
  1421=>"000000011",
  1422=>"011010100",
  1423=>"100001010",
  1424=>"101000010",
  1425=>"000001011",
  1426=>"001100011",
  1427=>"101010111",
  1428=>"100010001",
  1429=>"100011000",
  1430=>"001001100",
  1431=>"101011101",
  1432=>"001010110",
  1433=>"011010001",
  1434=>"000110000",
  1435=>"000110110",
  1436=>"001011111",
  1437=>"010110100",
  1438=>"011011111",
  1439=>"000011110",
  1440=>"111101111",
  1441=>"111010101",
  1442=>"111000000",
  1443=>"100001110",
  1444=>"111001101",
  1445=>"100011010",
  1446=>"100000101",
  1447=>"111111111",
  1448=>"000110001",
  1449=>"001011001",
  1450=>"001111100",
  1451=>"010100100",
  1452=>"000101101",
  1453=>"010110110",
  1454=>"111011011",
  1455=>"000000000",
  1456=>"111101001",
  1457=>"111111011",
  1458=>"100111110",
  1459=>"110000001",
  1460=>"101011110",
  1461=>"110010000",
  1462=>"111111110",
  1463=>"101001001",
  1464=>"100110001",
  1465=>"100101100",
  1466=>"010000100",
  1467=>"001010110",
  1468=>"110110101",
  1469=>"011111000",
  1470=>"010000100",
  1471=>"011011010",
  1472=>"111010000",
  1473=>"100100100",
  1474=>"001001100",
  1475=>"110111010",
  1476=>"001111011",
  1477=>"011111100",
  1478=>"110010001",
  1479=>"110001111",
  1480=>"100101011",
  1481=>"001101100",
  1482=>"001100011",
  1483=>"100101111",
  1484=>"001000110",
  1485=>"010100011",
  1486=>"100000010",
  1487=>"000110101",
  1488=>"101111111",
  1489=>"101011101",
  1490=>"010111111",
  1491=>"000100000",
  1492=>"011101101",
  1493=>"010101101",
  1494=>"111100101",
  1495=>"110011101",
  1496=>"110010010",
  1497=>"100010000",
  1498=>"011111110",
  1499=>"001001110",
  1500=>"101111011",
  1501=>"101001010",
  1502=>"110101111",
  1503=>"010011110",
  1504=>"110000000",
  1505=>"100011001",
  1506=>"000000100",
  1507=>"001010100",
  1508=>"001001110",
  1509=>"101110011",
  1510=>"101100010",
  1511=>"110111111",
  1512=>"011101110",
  1513=>"100011000",
  1514=>"110001101",
  1515=>"000001100",
  1516=>"001001000",
  1517=>"011000011",
  1518=>"000011101",
  1519=>"100110101",
  1520=>"110001100",
  1521=>"010001110",
  1522=>"011101001",
  1523=>"110000000",
  1524=>"001111100",
  1525=>"010111010",
  1526=>"110110010",
  1527=>"001100000",
  1528=>"010011000",
  1529=>"100011001",
  1530=>"000100101",
  1531=>"101000010",
  1532=>"010010010",
  1533=>"001111100",
  1534=>"010110000",
  1535=>"100001111",
  1536=>"100010100",
  1537=>"100000110",
  1538=>"100000101",
  1539=>"010011110",
  1540=>"010000011",
  1541=>"111110100",
  1542=>"001001000",
  1543=>"100101011",
  1544=>"101010010",
  1545=>"100101011",
  1546=>"110011000",
  1547=>"111111001",
  1548=>"111111111",
  1549=>"111111111",
  1550=>"101111000",
  1551=>"001000110",
  1552=>"001001000",
  1553=>"000001010",
  1554=>"010001111",
  1555=>"001010110",
  1556=>"000100010",
  1557=>"101101000",
  1558=>"111111110",
  1559=>"110100001",
  1560=>"110101101",
  1561=>"000001000",
  1562=>"010110000",
  1563=>"101010011",
  1564=>"110101110",
  1565=>"000010110",
  1566=>"001111110",
  1567=>"000001011",
  1568=>"000001100",
  1569=>"011100000",
  1570=>"010100000",
  1571=>"111110011",
  1572=>"011100010",
  1573=>"101101111",
  1574=>"010011010",
  1575=>"111010011",
  1576=>"010000111",
  1577=>"011011001",
  1578=>"111001111",
  1579=>"000111110",
  1580=>"000011111",
  1581=>"000001000",
  1582=>"000100101",
  1583=>"010100001",
  1584=>"111101110",
  1585=>"010011110",
  1586=>"110110001",
  1587=>"001101011",
  1588=>"000010100",
  1589=>"101100111",
  1590=>"101010000",
  1591=>"111000011",
  1592=>"010100010",
  1593=>"111100110",
  1594=>"111100001",
  1595=>"100001010",
  1596=>"111111001",
  1597=>"101100001",
  1598=>"001111000",
  1599=>"010001010",
  1600=>"100110010",
  1601=>"100011111",
  1602=>"110111101",
  1603=>"010110000",
  1604=>"110110010",
  1605=>"010100100",
  1606=>"100001111",
  1607=>"001011000",
  1608=>"001001100",
  1609=>"000010001",
  1610=>"010100110",
  1611=>"101001100",
  1612=>"100100101",
  1613=>"011101001",
  1614=>"110110100",
  1615=>"001000000",
  1616=>"110001001",
  1617=>"001111001",
  1618=>"011101110",
  1619=>"000110101",
  1620=>"011111100",
  1621=>"001110111",
  1622=>"000000100",
  1623=>"010100011",
  1624=>"100110010",
  1625=>"101111011",
  1626=>"110010101",
  1627=>"101110110",
  1628=>"011000101",
  1629=>"101000100",
  1630=>"111000011",
  1631=>"010110011",
  1632=>"111000000",
  1633=>"110111001",
  1634=>"100011100",
  1635=>"110000110",
  1636=>"011000000",
  1637=>"000000110",
  1638=>"100001101",
  1639=>"101001000",
  1640=>"110101110",
  1641=>"001000010",
  1642=>"111110100",
  1643=>"001011001",
  1644=>"101100111",
  1645=>"011111010",
  1646=>"111111111",
  1647=>"001001100",
  1648=>"110101011",
  1649=>"101010101",
  1650=>"110101001",
  1651=>"001001011",
  1652=>"011011110",
  1653=>"100101111",
  1654=>"010111101",
  1655=>"010100111",
  1656=>"010011111",
  1657=>"000010000",
  1658=>"011101001",
  1659=>"110011101",
  1660=>"001100011",
  1661=>"000000100",
  1662=>"010001101",
  1663=>"110010111",
  1664=>"010010001",
  1665=>"001101101",
  1666=>"100111111",
  1667=>"100101010",
  1668=>"001011000",
  1669=>"111010101",
  1670=>"000110010",
  1671=>"011101101",
  1672=>"011100111",
  1673=>"100010110",
  1674=>"011011001",
  1675=>"010001100",
  1676=>"011010001",
  1677=>"110100101",
  1678=>"000010011",
  1679=>"010010100",
  1680=>"000110010",
  1681=>"011110000",
  1682=>"000101011",
  1683=>"011010110",
  1684=>"111010110",
  1685=>"111000101",
  1686=>"101010011",
  1687=>"000100110",
  1688=>"011101010",
  1689=>"000111001",
  1690=>"000011100",
  1691=>"011010111",
  1692=>"110111000",
  1693=>"011101100",
  1694=>"001000000",
  1695=>"000001110",
  1696=>"011110011",
  1697=>"011110001",
  1698=>"100111110",
  1699=>"111101101",
  1700=>"000111101",
  1701=>"111001100",
  1702=>"010100100",
  1703=>"010110100",
  1704=>"111111110",
  1705=>"010000000",
  1706=>"000000110",
  1707=>"111011110",
  1708=>"010101111",
  1709=>"111010101",
  1710=>"111101101",
  1711=>"010100010",
  1712=>"011011111",
  1713=>"110100011",
  1714=>"101001001",
  1715=>"011110111",
  1716=>"001101111",
  1717=>"010111100",
  1718=>"101011001",
  1719=>"010010100",
  1720=>"000101001",
  1721=>"110000010",
  1722=>"010001000",
  1723=>"111111111",
  1724=>"101011110",
  1725=>"110101100",
  1726=>"110011101",
  1727=>"101111101",
  1728=>"011000001",
  1729=>"001001101",
  1730=>"010110010",
  1731=>"001100011",
  1732=>"101000100",
  1733=>"110000001",
  1734=>"111111000",
  1735=>"000110100",
  1736=>"110011011",
  1737=>"000100011",
  1738=>"000000111",
  1739=>"010010011",
  1740=>"001101001",
  1741=>"011101110",
  1742=>"000001010",
  1743=>"011110010",
  1744=>"011000100",
  1745=>"101100101",
  1746=>"111111000",
  1747=>"110110010",
  1748=>"100100100",
  1749=>"001010101",
  1750=>"011111100",
  1751=>"110011111",
  1752=>"001111011",
  1753=>"110000011",
  1754=>"110000001",
  1755=>"100101110",
  1756=>"100111101",
  1757=>"000101110",
  1758=>"011001001",
  1759=>"111100110",
  1760=>"100000001",
  1761=>"010001100",
  1762=>"000011010",
  1763=>"010010000",
  1764=>"011111101",
  1765=>"111110100",
  1766=>"101111100",
  1767=>"000110101",
  1768=>"001111100",
  1769=>"001011011",
  1770=>"111110010",
  1771=>"001011000",
  1772=>"000101000",
  1773=>"011101011",
  1774=>"101111000",
  1775=>"111011000",
  1776=>"000100010",
  1777=>"000011110",
  1778=>"110111100",
  1779=>"111111000",
  1780=>"010110000",
  1781=>"110000100",
  1782=>"100010001",
  1783=>"000110110",
  1784=>"100000110",
  1785=>"000110111",
  1786=>"111110111",
  1787=>"101000101",
  1788=>"100011010",
  1789=>"011100100",
  1790=>"001100101",
  1791=>"011100010",
  1792=>"111110110",
  1793=>"001110111",
  1794=>"101011010",
  1795=>"001110110",
  1796=>"000001010",
  1797=>"101010111",
  1798=>"100111111",
  1799=>"001000010",
  1800=>"000000010",
  1801=>"110001000",
  1802=>"110000001",
  1803=>"010100010",
  1804=>"111100011",
  1805=>"100100000",
  1806=>"111000010",
  1807=>"101111110",
  1808=>"011100110",
  1809=>"011000100",
  1810=>"000010000",
  1811=>"001001010",
  1812=>"011011100",
  1813=>"110010000",
  1814=>"111111110",
  1815=>"110110101",
  1816=>"010111011",
  1817=>"101000111",
  1818=>"011100001",
  1819=>"011011011",
  1820=>"111111110",
  1821=>"111111110",
  1822=>"000110011",
  1823=>"010111000",
  1824=>"110011001",
  1825=>"000101011",
  1826=>"000011110",
  1827=>"001111101",
  1828=>"100010100",
  1829=>"111111101",
  1830=>"110010001",
  1831=>"100000010",
  1832=>"100111010",
  1833=>"001110101",
  1834=>"100011000",
  1835=>"101010010",
  1836=>"101001001",
  1837=>"001001111",
  1838=>"011110100",
  1839=>"111001110",
  1840=>"100100011",
  1841=>"000010000",
  1842=>"010001010",
  1843=>"110100011",
  1844=>"100010111",
  1845=>"011000011",
  1846=>"101000000",
  1847=>"000001010",
  1848=>"011011111",
  1849=>"010010011",
  1850=>"110010101",
  1851=>"011010011",
  1852=>"010100000",
  1853=>"101100100",
  1854=>"011111101",
  1855=>"101111111",
  1856=>"111100101",
  1857=>"000001101",
  1858=>"111110110",
  1859=>"000000101",
  1860=>"010000011",
  1861=>"111101101",
  1862=>"010000101",
  1863=>"001100011",
  1864=>"110011101",
  1865=>"111111111",
  1866=>"011011110",
  1867=>"011000001",
  1868=>"101100000",
  1869=>"100101011",
  1870=>"010010010",
  1871=>"101011100",
  1872=>"010010001",
  1873=>"000011001",
  1874=>"001101100",
  1875=>"101100000",
  1876=>"111000101",
  1877=>"101110011",
  1878=>"111000011",
  1879=>"101111001",
  1880=>"001010000",
  1881=>"001100111",
  1882=>"011001110",
  1883=>"111010100",
  1884=>"000011111",
  1885=>"001000100",
  1886=>"000010000",
  1887=>"000000000",
  1888=>"100111010",
  1889=>"011001001",
  1890=>"010100110",
  1891=>"010001100",
  1892=>"110111100",
  1893=>"011011101",
  1894=>"010101010",
  1895=>"101000000",
  1896=>"000111011",
  1897=>"110100111",
  1898=>"100001111",
  1899=>"001010010",
  1900=>"001000111",
  1901=>"010111011",
  1902=>"101101001",
  1903=>"111010100",
  1904=>"000101000",
  1905=>"001110111",
  1906=>"010011110",
  1907=>"110000010",
  1908=>"101101101",
  1909=>"110110101",
  1910=>"011111101",
  1911=>"000001001",
  1912=>"011101011",
  1913=>"001011011",
  1914=>"111001101",
  1915=>"000001101",
  1916=>"110111000",
  1917=>"001010001",
  1918=>"100100101",
  1919=>"001100001",
  1920=>"100000000",
  1921=>"011001001",
  1922=>"110011011",
  1923=>"010100110",
  1924=>"010001100",
  1925=>"111111100",
  1926=>"111100011",
  1927=>"110011010",
  1928=>"010000010",
  1929=>"100110010",
  1930=>"010101011",
  1931=>"111011101",
  1932=>"100111001",
  1933=>"000110110",
  1934=>"110110010",
  1935=>"100101000",
  1936=>"101110000",
  1937=>"101100110",
  1938=>"111100110",
  1939=>"000000010",
  1940=>"110101100",
  1941=>"011100110",
  1942=>"100110110",
  1943=>"000010111",
  1944=>"011111101",
  1945=>"010011000",
  1946=>"110100100",
  1947=>"101000000",
  1948=>"111001110",
  1949=>"111101011",
  1950=>"101101110",
  1951=>"010111100",
  1952=>"001010111",
  1953=>"010100001",
  1954=>"010010111",
  1955=>"011010011",
  1956=>"101011001",
  1957=>"110011101",
  1958=>"100110100",
  1959=>"101110011",
  1960=>"110110101",
  1961=>"000001110",
  1962=>"100111001",
  1963=>"010000110",
  1964=>"100111101",
  1965=>"010100000",
  1966=>"111100000",
  1967=>"010011101",
  1968=>"101011000",
  1969=>"101000010",
  1970=>"001101010",
  1971=>"111001110",
  1972=>"011111101",
  1973=>"101011100",
  1974=>"010101101",
  1975=>"001101011",
  1976=>"011101111",
  1977=>"000111001",
  1978=>"100100100",
  1979=>"110001001",
  1980=>"010111111",
  1981=>"000010001",
  1982=>"110100100",
  1983=>"000001100",
  1984=>"111000010",
  1985=>"111000100",
  1986=>"111110001",
  1987=>"011001001",
  1988=>"010000011",
  1989=>"000100100",
  1990=>"101000011",
  1991=>"110100000",
  1992=>"110101010",
  1993=>"100001110",
  1994=>"101010110",
  1995=>"111000000",
  1996=>"000100100",
  1997=>"111111101",
  1998=>"011101110",
  1999=>"001101001",
  2000=>"000111010",
  2001=>"110111111",
  2002=>"100100000",
  2003=>"111101001",
  2004=>"101110111",
  2005=>"111001010",
  2006=>"111011001",
  2007=>"100110000",
  2008=>"000101010",
  2009=>"001110000",
  2010=>"100101110",
  2011=>"001000101",
  2012=>"110111000",
  2013=>"111111000",
  2014=>"001100101",
  2015=>"111110000",
  2016=>"111010111",
  2017=>"100010001",
  2018=>"111011000",
  2019=>"001101001",
  2020=>"000001000",
  2021=>"100000001",
  2022=>"010101011",
  2023=>"011100000",
  2024=>"100011000",
  2025=>"110110000",
  2026=>"010011000",
  2027=>"110101111",
  2028=>"100101111",
  2029=>"110000011",
  2030=>"000010101",
  2031=>"110001001",
  2032=>"010010101",
  2033=>"101111001",
  2034=>"010000101",
  2035=>"010111101",
  2036=>"111000001",
  2037=>"000100111",
  2038=>"110011001",
  2039=>"001101111",
  2040=>"111010010",
  2041=>"100011010",
  2042=>"111001100",
  2043=>"011000000",
  2044=>"000111000",
  2045=>"010100001",
  2046=>"111110010",
  2047=>"101000010",
  2048=>"100010100",
  2049=>"011101111",
  2050=>"001111000",
  2051=>"110111011",
  2052=>"101001100",
  2053=>"101001011",
  2054=>"101010111",
  2055=>"011110101",
  2056=>"000101111",
  2057=>"111001011",
  2058=>"100110001",
  2059=>"000110000",
  2060=>"101010011",
  2061=>"101011100",
  2062=>"000100100",
  2063=>"000101110",
  2064=>"010011100",
  2065=>"100000011",
  2066=>"110101100",
  2067=>"011101000",
  2068=>"100001101",
  2069=>"111011011",
  2070=>"010000010",
  2071=>"111100000",
  2072=>"100011001",
  2073=>"111000000",
  2074=>"100101100",
  2075=>"100101011",
  2076=>"010111001",
  2077=>"010101101",
  2078=>"101110011",
  2079=>"100100100",
  2080=>"100110101",
  2081=>"001001001",
  2082=>"101001110",
  2083=>"000000100",
  2084=>"010100100",
  2085=>"110110100",
  2086=>"110100111",
  2087=>"010111011",
  2088=>"100000001",
  2089=>"101111010",
  2090=>"100011011",
  2091=>"010010010",
  2092=>"110100000",
  2093=>"000001001",
  2094=>"011101011",
  2095=>"100110001",
  2096=>"010011111",
  2097=>"100110011",
  2098=>"011001001",
  2099=>"100111101",
  2100=>"010011010",
  2101=>"001101100",
  2102=>"100111100",
  2103=>"110100000",
  2104=>"101000000",
  2105=>"100101010",
  2106=>"010110100",
  2107=>"000100101",
  2108=>"111111000",
  2109=>"110011100",
  2110=>"001011001",
  2111=>"000011000",
  2112=>"011000000",
  2113=>"011010000",
  2114=>"001101000",
  2115=>"111011011",
  2116=>"111000110",
  2117=>"010010110",
  2118=>"111011100",
  2119=>"101011101",
  2120=>"110000100",
  2121=>"000110010",
  2122=>"110111111",
  2123=>"001001101",
  2124=>"110000000",
  2125=>"000000100",
  2126=>"001000100",
  2127=>"110100110",
  2128=>"010111001",
  2129=>"001111011",
  2130=>"011100111",
  2131=>"100001111",
  2132=>"111010001",
  2133=>"011111110",
  2134=>"011111110",
  2135=>"100010001",
  2136=>"001100000",
  2137=>"011010011",
  2138=>"110001011",
  2139=>"001110010",
  2140=>"011000000",
  2141=>"000001110",
  2142=>"011011000",
  2143=>"110101011",
  2144=>"000101100",
  2145=>"110101101",
  2146=>"010001000",
  2147=>"011100001",
  2148=>"001110100",
  2149=>"101010010",
  2150=>"000001000",
  2151=>"110010110",
  2152=>"011100011",
  2153=>"101111110",
  2154=>"010011111",
  2155=>"011011000",
  2156=>"001010001",
  2157=>"010000011",
  2158=>"001010101",
  2159=>"000111000",
  2160=>"101001000",
  2161=>"001000110",
  2162=>"110101011",
  2163=>"001111111",
  2164=>"001000001",
  2165=>"100111011",
  2166=>"111001101",
  2167=>"110000011",
  2168=>"011101001",
  2169=>"001011101",
  2170=>"000000000",
  2171=>"101011001",
  2172=>"011010110",
  2173=>"000010100",
  2174=>"010101000",
  2175=>"011100101",
  2176=>"110000000",
  2177=>"011000101",
  2178=>"010100101",
  2179=>"111110111",
  2180=>"001110010",
  2181=>"101101001",
  2182=>"110000010",
  2183=>"110011010",
  2184=>"000001110",
  2185=>"000011100",
  2186=>"000111011",
  2187=>"100001101",
  2188=>"000111110",
  2189=>"011101111",
  2190=>"000001111",
  2191=>"000101110",
  2192=>"010101111",
  2193=>"001011100",
  2194=>"111110110",
  2195=>"001111111",
  2196=>"111110010",
  2197=>"000001111",
  2198=>"100111100",
  2199=>"001011100",
  2200=>"111111111",
  2201=>"110000001",
  2202=>"010001001",
  2203=>"111001000",
  2204=>"001010101",
  2205=>"001101000",
  2206=>"100000000",
  2207=>"111100101",
  2208=>"001000101",
  2209=>"111110111",
  2210=>"000101010",
  2211=>"111000001",
  2212=>"101010001",
  2213=>"101101011",
  2214=>"001011101",
  2215=>"100010001",
  2216=>"111000011",
  2217=>"001111101",
  2218=>"101111000",
  2219=>"011000010",
  2220=>"000101000",
  2221=>"000010110",
  2222=>"101010101",
  2223=>"000010100",
  2224=>"010000111",
  2225=>"001000100",
  2226=>"011101011",
  2227=>"100011100",
  2228=>"001000100",
  2229=>"000100000",
  2230=>"001110110",
  2231=>"000000000",
  2232=>"011100011",
  2233=>"111111111",
  2234=>"001000010",
  2235=>"011100101",
  2236=>"100110010",
  2237=>"101111110",
  2238=>"001001110",
  2239=>"000011000",
  2240=>"001100101",
  2241=>"011011101",
  2242=>"101111111",
  2243=>"110100001",
  2244=>"001111111",
  2245=>"111101110",
  2246=>"000110001",
  2247=>"111000000",
  2248=>"101011001",
  2249=>"111100100",
  2250=>"001011011",
  2251=>"110100111",
  2252=>"011110001",
  2253=>"101101110",
  2254=>"001011011",
  2255=>"100100001",
  2256=>"010010011",
  2257=>"000011001",
  2258=>"110101100",
  2259=>"100110010",
  2260=>"101110000",
  2261=>"110110001",
  2262=>"111111000",
  2263=>"110111100",
  2264=>"100101000",
  2265=>"001111011",
  2266=>"010111100",
  2267=>"111110001",
  2268=>"101100001",
  2269=>"011101110",
  2270=>"110100110",
  2271=>"110010011",
  2272=>"010011110",
  2273=>"001011100",
  2274=>"110000010",
  2275=>"011110110",
  2276=>"100110100",
  2277=>"100110001",
  2278=>"100111001",
  2279=>"100000001",
  2280=>"110000000",
  2281=>"111000011",
  2282=>"000100000",
  2283=>"001001101",
  2284=>"111000000",
  2285=>"010110110",
  2286=>"001101010",
  2287=>"100100010",
  2288=>"001110110",
  2289=>"100010001",
  2290=>"100101111",
  2291=>"000001111",
  2292=>"000001100",
  2293=>"100000000",
  2294=>"101101010",
  2295=>"001110101",
  2296=>"011111101",
  2297=>"001110001",
  2298=>"110011010",
  2299=>"000011100",
  2300=>"110110110",
  2301=>"111011010",
  2302=>"110000000",
  2303=>"000100010",
  2304=>"111001110",
  2305=>"100000000",
  2306=>"111000010",
  2307=>"000001010",
  2308=>"101111001",
  2309=>"000101001",
  2310=>"101010000",
  2311=>"000101000",
  2312=>"000000011",
  2313=>"101110100",
  2314=>"100101011",
  2315=>"101000000",
  2316=>"010010000",
  2317=>"101110110",
  2318=>"101111110",
  2319=>"100010011",
  2320=>"110100010",
  2321=>"001001001",
  2322=>"010010111",
  2323=>"000110101",
  2324=>"010011000",
  2325=>"100000011",
  2326=>"011011110",
  2327=>"001110000",
  2328=>"100001010",
  2329=>"010001000",
  2330=>"110101111",
  2331=>"111010110",
  2332=>"001101111",
  2333=>"001001001",
  2334=>"011011011",
  2335=>"000011001",
  2336=>"100001010",
  2337=>"000001011",
  2338=>"110010101",
  2339=>"110111000",
  2340=>"011000101",
  2341=>"100000111",
  2342=>"111111111",
  2343=>"001010111",
  2344=>"101010111",
  2345=>"101100010",
  2346=>"011100111",
  2347=>"001100011",
  2348=>"111110000",
  2349=>"000001010",
  2350=>"011010110",
  2351=>"100101011",
  2352=>"000101101",
  2353=>"101100100",
  2354=>"000101011",
  2355=>"011111100",
  2356=>"101111110",
  2357=>"011000101",
  2358=>"111011010",
  2359=>"110000010",
  2360=>"000000000",
  2361=>"000110011",
  2362=>"000100100",
  2363=>"111100110",
  2364=>"111110010",
  2365=>"011001111",
  2366=>"110001100",
  2367=>"001111111",
  2368=>"011000101",
  2369=>"101111101",
  2370=>"000000000",
  2371=>"111100110",
  2372=>"011111001",
  2373=>"100110110",
  2374=>"000010110",
  2375=>"010011010",
  2376=>"011011000",
  2377=>"000000110",
  2378=>"010011100",
  2379=>"001111111",
  2380=>"010101100",
  2381=>"110111111",
  2382=>"011101110",
  2383=>"000011110",
  2384=>"101110011",
  2385=>"010101111",
  2386=>"001010100",
  2387=>"011100100",
  2388=>"011110010",
  2389=>"101111000",
  2390=>"110110001",
  2391=>"110001100",
  2392=>"001100011",
  2393=>"101110000",
  2394=>"001001001",
  2395=>"000100110",
  2396=>"110000000",
  2397=>"001111101",
  2398=>"001000001",
  2399=>"110011000",
  2400=>"000001111",
  2401=>"001010101",
  2402=>"110001101",
  2403=>"001010101",
  2404=>"101010001",
  2405=>"010001011",
  2406=>"001110101",
  2407=>"010110011",
  2408=>"010001100",
  2409=>"000110010",
  2410=>"100101111",
  2411=>"001101010",
  2412=>"001000000",
  2413=>"111001000",
  2414=>"000000101",
  2415=>"111111000",
  2416=>"111100001",
  2417=>"000001000",
  2418=>"101000100",
  2419=>"110011110",
  2420=>"111010100",
  2421=>"011111011",
  2422=>"011110010",
  2423=>"001000110",
  2424=>"101010001",
  2425=>"101010000",
  2426=>"010001101",
  2427=>"000101011",
  2428=>"111100010",
  2429=>"111011001",
  2430=>"010001111",
  2431=>"001110101",
  2432=>"000101011",
  2433=>"101000001",
  2434=>"101011010",
  2435=>"111010100",
  2436=>"000001110",
  2437=>"001001011",
  2438=>"110001011",
  2439=>"011000010",
  2440=>"110011001",
  2441=>"100000111",
  2442=>"111111000",
  2443=>"000000101",
  2444=>"010001101",
  2445=>"110011000",
  2446=>"100011100",
  2447=>"100111011",
  2448=>"101000111",
  2449=>"010110011",
  2450=>"010010001",
  2451=>"110111111",
  2452=>"101110111",
  2453=>"111101100",
  2454=>"011101010",
  2455=>"101100111",
  2456=>"010001001",
  2457=>"100011000",
  2458=>"101110000",
  2459=>"000001000",
  2460=>"010101101",
  2461=>"100100110",
  2462=>"001111110",
  2463=>"001101101",
  2464=>"000001011",
  2465=>"000001001",
  2466=>"001001010",
  2467=>"010111001",
  2468=>"000010101",
  2469=>"100000010",
  2470=>"100000001",
  2471=>"010110110",
  2472=>"011100001",
  2473=>"011110011",
  2474=>"000000010",
  2475=>"010110011",
  2476=>"110101100",
  2477=>"110010111",
  2478=>"101111111",
  2479=>"000000011",
  2480=>"001110011",
  2481=>"011000100",
  2482=>"011100010",
  2483=>"011001101",
  2484=>"101110101",
  2485=>"011001000",
  2486=>"010011111",
  2487=>"111110011",
  2488=>"011011000",
  2489=>"100101001",
  2490=>"101111110",
  2491=>"110101011",
  2492=>"111111001",
  2493=>"011010100",
  2494=>"110100000",
  2495=>"111001010",
  2496=>"101000000",
  2497=>"101110011",
  2498=>"011110100",
  2499=>"100110101",
  2500=>"011001111",
  2501=>"001011110",
  2502=>"010101010",
  2503=>"000100000",
  2504=>"110011010",
  2505=>"011100011",
  2506=>"000110000",
  2507=>"101000110",
  2508=>"011001001",
  2509=>"101011110",
  2510=>"000000111",
  2511=>"110110100",
  2512=>"101011011",
  2513=>"000011000",
  2514=>"011100100",
  2515=>"100011110",
  2516=>"000001111",
  2517=>"001000001",
  2518=>"100110101",
  2519=>"000111111",
  2520=>"011111000",
  2521=>"110100110",
  2522=>"101011101",
  2523=>"010101001",
  2524=>"111000010",
  2525=>"110000110",
  2526=>"000010110",
  2527=>"000001100",
  2528=>"110101100",
  2529=>"001010110",
  2530=>"100010010",
  2531=>"000111100",
  2532=>"100101010",
  2533=>"101000000",
  2534=>"010101010",
  2535=>"011001000",
  2536=>"111100111",
  2537=>"011001010",
  2538=>"000001010",
  2539=>"011101110",
  2540=>"101011011",
  2541=>"011000010",
  2542=>"000111001",
  2543=>"010111101",
  2544=>"011011010",
  2545=>"001000101",
  2546=>"001101010",
  2547=>"011110011",
  2548=>"011110100",
  2549=>"111011011",
  2550=>"101000101",
  2551=>"110100111",
  2552=>"110011111",
  2553=>"000000100",
  2554=>"100001111",
  2555=>"011000001",
  2556=>"011111011",
  2557=>"100000110",
  2558=>"010111111",
  2559=>"111010111",
  2560=>"101000111",
  2561=>"010111110",
  2562=>"000010110",
  2563=>"011000110",
  2564=>"110000000",
  2565=>"011000111",
  2566=>"101110111",
  2567=>"100100001",
  2568=>"010010001",
  2569=>"010010011",
  2570=>"110111001",
  2571=>"010001100",
  2572=>"011001111",
  2573=>"010011110",
  2574=>"011001101",
  2575=>"001100001",
  2576=>"001101001",
  2577=>"000100011",
  2578=>"010100010",
  2579=>"110010010",
  2580=>"001101000",
  2581=>"100000000",
  2582=>"010001111",
  2583=>"110011010",
  2584=>"100011110",
  2585=>"111011100",
  2586=>"001011101",
  2587=>"000100011",
  2588=>"001000011",
  2589=>"100000110",
  2590=>"100011100",
  2591=>"000010101",
  2592=>"110100101",
  2593=>"110011100",
  2594=>"011100100",
  2595=>"000111110",
  2596=>"001110010",
  2597=>"100010111",
  2598=>"111011001",
  2599=>"010001000",
  2600=>"001100101",
  2601=>"011111111",
  2602=>"111001000",
  2603=>"110100100",
  2604=>"000110001",
  2605=>"011101101",
  2606=>"100111101",
  2607=>"000111000",
  2608=>"000010110",
  2609=>"001101110",
  2610=>"101110111",
  2611=>"110111100",
  2612=>"100001101",
  2613=>"101010100",
  2614=>"010001011",
  2615=>"001100001",
  2616=>"010000100",
  2617=>"100100000",
  2618=>"001010010",
  2619=>"101010101",
  2620=>"101110011",
  2621=>"000101000",
  2622=>"010111111",
  2623=>"100010110",
  2624=>"011000010",
  2625=>"101011100",
  2626=>"000011001",
  2627=>"010001011",
  2628=>"010010000",
  2629=>"100100110",
  2630=>"000010000",
  2631=>"010100011",
  2632=>"100101010",
  2633=>"001000110",
  2634=>"111000000",
  2635=>"000010010",
  2636=>"010001010",
  2637=>"000111110",
  2638=>"010000000",
  2639=>"110110000",
  2640=>"111100111",
  2641=>"111110101",
  2642=>"111110011",
  2643=>"011000001",
  2644=>"100000010",
  2645=>"110100100",
  2646=>"000010100",
  2647=>"011110000",
  2648=>"110111101",
  2649=>"011010000",
  2650=>"010100001",
  2651=>"011110101",
  2652=>"000000111",
  2653=>"001000101",
  2654=>"011100111",
  2655=>"011011010",
  2656=>"000100111",
  2657=>"000000000",
  2658=>"110011001",
  2659=>"100111101",
  2660=>"001100000",
  2661=>"011011011",
  2662=>"011000011",
  2663=>"110110011",
  2664=>"100010000",
  2665=>"110111011",
  2666=>"111001111",
  2667=>"100100000",
  2668=>"100000100",
  2669=>"010010001",
  2670=>"111001000",
  2671=>"011010110",
  2672=>"001010000",
  2673=>"000011000",
  2674=>"011101111",
  2675=>"111110110",
  2676=>"100110011",
  2677=>"001110101",
  2678=>"011101110",
  2679=>"100100111",
  2680=>"001101110",
  2681=>"001110100",
  2682=>"001010110",
  2683=>"010010111",
  2684=>"100100001",
  2685=>"010000010",
  2686=>"111110110",
  2687=>"110001000",
  2688=>"011100111",
  2689=>"100111101",
  2690=>"000111000",
  2691=>"100011101",
  2692=>"100000111",
  2693=>"110000010",
  2694=>"111110101",
  2695=>"101011111",
  2696=>"111101101",
  2697=>"100010100",
  2698=>"100011000",
  2699=>"111110100",
  2700=>"001101000",
  2701=>"111111011",
  2702=>"110111000",
  2703=>"100101001",
  2704=>"111111110",
  2705=>"011011001",
  2706=>"010000001",
  2707=>"000111111",
  2708=>"110100101",
  2709=>"110010011",
  2710=>"110111111",
  2711=>"110010100",
  2712=>"101111001",
  2713=>"111100101",
  2714=>"011001110",
  2715=>"111101111",
  2716=>"111001111",
  2717=>"101101010",
  2718=>"111101001",
  2719=>"011111111",
  2720=>"000010101",
  2721=>"111010000",
  2722=>"010010111",
  2723=>"000111010",
  2724=>"010001111",
  2725=>"000010101",
  2726=>"011000101",
  2727=>"011011000",
  2728=>"000001110",
  2729=>"100100010",
  2730=>"101001111",
  2731=>"100110110",
  2732=>"001100001",
  2733=>"011101000",
  2734=>"100111110",
  2735=>"100011001",
  2736=>"101100000",
  2737=>"111001000",
  2738=>"101011000",
  2739=>"010000101",
  2740=>"010011110",
  2741=>"001101101",
  2742=>"010111001",
  2743=>"101100101",
  2744=>"110101110",
  2745=>"110110111",
  2746=>"100000100",
  2747=>"110110111",
  2748=>"100111001",
  2749=>"011000000",
  2750=>"000000100",
  2751=>"011101010",
  2752=>"111101101",
  2753=>"110101111",
  2754=>"110101010",
  2755=>"011111110",
  2756=>"000010000",
  2757=>"100110010",
  2758=>"100010110",
  2759=>"100101010",
  2760=>"010010001",
  2761=>"111011010",
  2762=>"110110001",
  2763=>"001000000",
  2764=>"010011011",
  2765=>"100001010",
  2766=>"100101010",
  2767=>"000010001",
  2768=>"100001000",
  2769=>"110100001",
  2770=>"000010110",
  2771=>"010000100",
  2772=>"111001000",
  2773=>"010110000",
  2774=>"001111000",
  2775=>"101001101",
  2776=>"100101100",
  2777=>"011101011",
  2778=>"011010010",
  2779=>"100100110",
  2780=>"000100111",
  2781=>"010010001",
  2782=>"000011101",
  2783=>"010010110",
  2784=>"101000010",
  2785=>"010001001",
  2786=>"100001111",
  2787=>"110001100",
  2788=>"110111000",
  2789=>"001111100",
  2790=>"111110011",
  2791=>"111000010",
  2792=>"000001111",
  2793=>"111111111",
  2794=>"001100100",
  2795=>"011110000",
  2796=>"101011010",
  2797=>"100011001",
  2798=>"101000101",
  2799=>"111100011",
  2800=>"011100010",
  2801=>"110011001",
  2802=>"110001011",
  2803=>"000010111",
  2804=>"010010101",
  2805=>"001001011",
  2806=>"110100001",
  2807=>"000100110",
  2808=>"101110000",
  2809=>"101101011",
  2810=>"011100100",
  2811=>"010110010",
  2812=>"000111000",
  2813=>"010111110",
  2814=>"110010110",
  2815=>"000011100",
  2816=>"000110110",
  2817=>"110111011",
  2818=>"000011011",
  2819=>"110001011",
  2820=>"000101100",
  2821=>"100011100",
  2822=>"000011001",
  2823=>"111010100",
  2824=>"100011111",
  2825=>"101010111",
  2826=>"000011100",
  2827=>"111111110",
  2828=>"101000001",
  2829=>"111011011",
  2830=>"101001100",
  2831=>"110100111",
  2832=>"100110011",
  2833=>"000000000",
  2834=>"100001001",
  2835=>"101001110",
  2836=>"100010000",
  2837=>"101001101",
  2838=>"000011111",
  2839=>"011101111",
  2840=>"101000100",
  2841=>"011000011",
  2842=>"101110001",
  2843=>"110111010",
  2844=>"101000111",
  2845=>"110000010",
  2846=>"100000000",
  2847=>"010101000",
  2848=>"100101111",
  2849=>"110011101",
  2850=>"100000111",
  2851=>"000110010",
  2852=>"000110111",
  2853=>"001000000",
  2854=>"000001001",
  2855=>"110111100",
  2856=>"100101110",
  2857=>"101110011",
  2858=>"100101110",
  2859=>"101101010",
  2860=>"100100110",
  2861=>"001000000",
  2862=>"001110010",
  2863=>"111100001",
  2864=>"101101010",
  2865=>"111111011",
  2866=>"011000000",
  2867=>"101111001",
  2868=>"100010110",
  2869=>"001100010",
  2870=>"010011000",
  2871=>"010101000",
  2872=>"010100011",
  2873=>"100100001",
  2874=>"010011001",
  2875=>"110101110",
  2876=>"001100001",
  2877=>"110011011",
  2878=>"110001110",
  2879=>"010100101",
  2880=>"100001010",
  2881=>"010100010",
  2882=>"000011010",
  2883=>"100000011",
  2884=>"010010111",
  2885=>"100100011",
  2886=>"011010010",
  2887=>"001101000",
  2888=>"101010111",
  2889=>"110000001",
  2890=>"010100000",
  2891=>"010110010",
  2892=>"110010000",
  2893=>"000101100",
  2894=>"011111100",
  2895=>"010001001",
  2896=>"111111010",
  2897=>"110011000",
  2898=>"000110100",
  2899=>"101011011",
  2900=>"111100110",
  2901=>"011111111",
  2902=>"111101010",
  2903=>"010001001",
  2904=>"101011011",
  2905=>"100111111",
  2906=>"101000011",
  2907=>"100101001",
  2908=>"000111111",
  2909=>"111111110",
  2910=>"111101001",
  2911=>"000000001",
  2912=>"111000000",
  2913=>"101100101",
  2914=>"001000010",
  2915=>"110110011",
  2916=>"011010001",
  2917=>"001110100",
  2918=>"010011100",
  2919=>"111011110",
  2920=>"001100000",
  2921=>"100110111",
  2922=>"110011111",
  2923=>"000010010",
  2924=>"001010011",
  2925=>"111011000",
  2926=>"111111100",
  2927=>"001001001",
  2928=>"011010100",
  2929=>"100101011",
  2930=>"100100001",
  2931=>"110001101",
  2932=>"001001100",
  2933=>"111100101",
  2934=>"110100110",
  2935=>"111111111",
  2936=>"001010000",
  2937=>"011110010",
  2938=>"001010010",
  2939=>"001101010",
  2940=>"110110001",
  2941=>"011110110",
  2942=>"111001010",
  2943=>"101110010",
  2944=>"001011101",
  2945=>"011011101",
  2946=>"001101011",
  2947=>"110000101",
  2948=>"100001011",
  2949=>"101100010",
  2950=>"001101001",
  2951=>"001011010",
  2952=>"001010010",
  2953=>"000101101",
  2954=>"000100010",
  2955=>"000110010",
  2956=>"001101101",
  2957=>"110010110",
  2958=>"110010010",
  2959=>"000110101",
  2960=>"010110010",
  2961=>"000101110",
  2962=>"111000011",
  2963=>"111101010",
  2964=>"100111000",
  2965=>"010110010",
  2966=>"110001000",
  2967=>"011100101",
  2968=>"101110011",
  2969=>"001011001",
  2970=>"010101110",
  2971=>"010101011",
  2972=>"111111010",
  2973=>"011111011",
  2974=>"100101000",
  2975=>"011110000",
  2976=>"110000000",
  2977=>"110000001",
  2978=>"110000001",
  2979=>"101101000",
  2980=>"101011000",
  2981=>"111111011",
  2982=>"001111111",
  2983=>"010000010",
  2984=>"111110000",
  2985=>"110011100",
  2986=>"100000111",
  2987=>"100010110",
  2988=>"001010101",
  2989=>"110001110",
  2990=>"110110110",
  2991=>"110100000",
  2992=>"010110101",
  2993=>"001110100",
  2994=>"001001011",
  2995=>"100111010",
  2996=>"111100000",
  2997=>"011011000",
  2998=>"100100111",
  2999=>"101111100",
  3000=>"010110110",
  3001=>"111111100",
  3002=>"001011111",
  3003=>"101101100",
  3004=>"111101000",
  3005=>"001000011",
  3006=>"011101110",
  3007=>"010000000",
  3008=>"011001001",
  3009=>"011010111",
  3010=>"000101010",
  3011=>"101000111",
  3012=>"010000000",
  3013=>"101110111",
  3014=>"011010000",
  3015=>"011111111",
  3016=>"111100101",
  3017=>"010010001",
  3018=>"001111101",
  3019=>"111111110",
  3020=>"111111010",
  3021=>"000001000",
  3022=>"001011100",
  3023=>"101101000",
  3024=>"111100011",
  3025=>"111001000",
  3026=>"110000011",
  3027=>"101010100",
  3028=>"000101011",
  3029=>"000111100",
  3030=>"000100100",
  3031=>"011100111",
  3032=>"101111101",
  3033=>"000110010",
  3034=>"101111111",
  3035=>"110111100",
  3036=>"100111110",
  3037=>"111100101",
  3038=>"101000010",
  3039=>"011011000",
  3040=>"000011000",
  3041=>"000000000",
  3042=>"011111011",
  3043=>"000001000",
  3044=>"000001001",
  3045=>"111100000",
  3046=>"010111000",
  3047=>"110111001",
  3048=>"111011000",
  3049=>"110001110",
  3050=>"010111011",
  3051=>"100111111",
  3052=>"100111100",
  3053=>"011001111",
  3054=>"011011110",
  3055=>"100010000",
  3056=>"000001001",
  3057=>"010100000",
  3058=>"011111101",
  3059=>"000000011",
  3060=>"000010010",
  3061=>"001001010",
  3062=>"001100010",
  3063=>"101110111",
  3064=>"110011011",
  3065=>"011011010",
  3066=>"000010000",
  3067=>"010010010",
  3068=>"111011100",
  3069=>"100000010",
  3070=>"011001101",
  3071=>"011100110",
  3072=>"100100001",
  3073=>"000110110",
  3074=>"001011110",
  3075=>"001010011",
  3076=>"110100011",
  3077=>"011111010",
  3078=>"001000010",
  3079=>"001001000",
  3080=>"100101000",
  3081=>"100000111",
  3082=>"001001100",
  3083=>"110110101",
  3084=>"001001010",
  3085=>"101100000",
  3086=>"001000001",
  3087=>"100111010",
  3088=>"011110001",
  3089=>"110011001",
  3090=>"000100111",
  3091=>"001111110",
  3092=>"100010101",
  3093=>"101110101",
  3094=>"101111010",
  3095=>"001000100",
  3096=>"100111000",
  3097=>"011000001",
  3098=>"011010001",
  3099=>"001001110",
  3100=>"001110110",
  3101=>"100011011",
  3102=>"011100010",
  3103=>"100010111",
  3104=>"001011000",
  3105=>"011011110",
  3106=>"011010000",
  3107=>"101100001",
  3108=>"110111111",
  3109=>"110100100",
  3110=>"010110100",
  3111=>"111110010",
  3112=>"100100010",
  3113=>"011101111",
  3114=>"101010110",
  3115=>"010001101",
  3116=>"011011001",
  3117=>"000011101",
  3118=>"010001111",
  3119=>"001010000",
  3120=>"011101111",
  3121=>"001101011",
  3122=>"001110110",
  3123=>"010011111",
  3124=>"100001001",
  3125=>"100111010",
  3126=>"001100010",
  3127=>"111111010",
  3128=>"111100001",
  3129=>"111000101",
  3130=>"101001100",
  3131=>"000000001",
  3132=>"010011010",
  3133=>"110011111",
  3134=>"011100110",
  3135=>"100101100",
  3136=>"110100011",
  3137=>"001000001",
  3138=>"001001110",
  3139=>"010101000",
  3140=>"001000011",
  3141=>"110000000",
  3142=>"000111110",
  3143=>"010001001",
  3144=>"111000110",
  3145=>"101000010",
  3146=>"001011101",
  3147=>"110000110",
  3148=>"000100111",
  3149=>"001010011",
  3150=>"110100011",
  3151=>"010011000",
  3152=>"100000011",
  3153=>"011111111",
  3154=>"100100010",
  3155=>"001011000",
  3156=>"101101100",
  3157=>"011001100",
  3158=>"101111111",
  3159=>"001000010",
  3160=>"101010111",
  3161=>"000001110",
  3162=>"111111001",
  3163=>"000100101",
  3164=>"011110000",
  3165=>"000110101",
  3166=>"000000101",
  3167=>"111000010",
  3168=>"011011101",
  3169=>"101111111",
  3170=>"011001111",
  3171=>"000100000",
  3172=>"011000001",
  3173=>"001110101",
  3174=>"111101010",
  3175=>"110010001",
  3176=>"000010001",
  3177=>"001011101",
  3178=>"000011000",
  3179=>"101010111",
  3180=>"110100101",
  3181=>"001010101",
  3182=>"011000100",
  3183=>"001111011",
  3184=>"001000010",
  3185=>"001011110",
  3186=>"100011111",
  3187=>"011101101",
  3188=>"100000010",
  3189=>"010011001",
  3190=>"111010101",
  3191=>"100111010",
  3192=>"001101110",
  3193=>"110110100",
  3194=>"000001001",
  3195=>"011001010",
  3196=>"111001001",
  3197=>"101111000",
  3198=>"101000010",
  3199=>"100110100",
  3200=>"101010001",
  3201=>"010011100",
  3202=>"100000010",
  3203=>"000001011",
  3204=>"000000010",
  3205=>"101001010",
  3206=>"100000011",
  3207=>"011111110",
  3208=>"110110101",
  3209=>"000000011",
  3210=>"101010011",
  3211=>"011001011",
  3212=>"111000111",
  3213=>"110110000",
  3214=>"001001011",
  3215=>"001111011",
  3216=>"000000010",
  3217=>"100011111",
  3218=>"011011010",
  3219=>"110110011",
  3220=>"001101101",
  3221=>"010001101",
  3222=>"010010001",
  3223=>"011101001",
  3224=>"100101101",
  3225=>"100010001",
  3226=>"110010100",
  3227=>"101001011",
  3228=>"100110110",
  3229=>"101100000",
  3230=>"001000000",
  3231=>"100001111",
  3232=>"111110000",
  3233=>"100101111",
  3234=>"100000101",
  3235=>"111010100",
  3236=>"101111111",
  3237=>"010011011",
  3238=>"111100010",
  3239=>"000111001",
  3240=>"111100001",
  3241=>"001000011",
  3242=>"010000010",
  3243=>"000010111",
  3244=>"111100001",
  3245=>"000100101",
  3246=>"101111010",
  3247=>"001101001",
  3248=>"100000001",
  3249=>"111010101",
  3250=>"100011010",
  3251=>"100110011",
  3252=>"100111101",
  3253=>"100010110",
  3254=>"100100110",
  3255=>"000111011",
  3256=>"001000011",
  3257=>"111111101",
  3258=>"011100101",
  3259=>"000000111",
  3260=>"011110101",
  3261=>"001001001",
  3262=>"101010111",
  3263=>"100000101",
  3264=>"000110000",
  3265=>"010011000",
  3266=>"101100011",
  3267=>"000010011",
  3268=>"101111010",
  3269=>"001111111",
  3270=>"110001011",
  3271=>"110000000",
  3272=>"110001000",
  3273=>"101100011",
  3274=>"101111101",
  3275=>"010011100",
  3276=>"101000111",
  3277=>"111000101",
  3278=>"000100011",
  3279=>"101001111",
  3280=>"011001110",
  3281=>"100110001",
  3282=>"000100100",
  3283=>"100111010",
  3284=>"011000101",
  3285=>"100101000",
  3286=>"111001000",
  3287=>"100011011",
  3288=>"100000111",
  3289=>"000010101",
  3290=>"101000000",
  3291=>"111100101",
  3292=>"011011011",
  3293=>"010001011",
  3294=>"111110100",
  3295=>"011110011",
  3296=>"000010011",
  3297=>"000010011",
  3298=>"100010000",
  3299=>"001000111",
  3300=>"011110011",
  3301=>"001000001",
  3302=>"100010110",
  3303=>"011011110",
  3304=>"110100011",
  3305=>"011110010",
  3306=>"011011010",
  3307=>"110000000",
  3308=>"111000000",
  3309=>"100100111",
  3310=>"011010010",
  3311=>"101100100",
  3312=>"101111010",
  3313=>"001001111",
  3314=>"011100000",
  3315=>"111100001",
  3316=>"101001100",
  3317=>"101110000",
  3318=>"001011001",
  3319=>"001000101",
  3320=>"001100110",
  3321=>"011101011",
  3322=>"101110111",
  3323=>"101000000",
  3324=>"110110010",
  3325=>"110010001",
  3326=>"011000111",
  3327=>"011100100",
  3328=>"101001011",
  3329=>"011111110",
  3330=>"110110001",
  3331=>"000101101",
  3332=>"011011110",
  3333=>"101110001",
  3334=>"011111011",
  3335=>"100111011",
  3336=>"110100100",
  3337=>"101000011",
  3338=>"110110010",
  3339=>"111010111",
  3340=>"000001010",
  3341=>"010110001",
  3342=>"100000010",
  3343=>"101110000",
  3344=>"100110001",
  3345=>"010101010",
  3346=>"001101101",
  3347=>"101010011",
  3348=>"010010010",
  3349=>"000011101",
  3350=>"011100101",
  3351=>"001010110",
  3352=>"100011111",
  3353=>"010011001",
  3354=>"000111110",
  3355=>"000111101",
  3356=>"010011100",
  3357=>"001000001",
  3358=>"010101111",
  3359=>"011101000",
  3360=>"011011100",
  3361=>"100110001",
  3362=>"000100100",
  3363=>"101111110",
  3364=>"011110100",
  3365=>"010110111",
  3366=>"111001101",
  3367=>"111100011",
  3368=>"110100000",
  3369=>"000001011",
  3370=>"110101110",
  3371=>"001001111",
  3372=>"101110101",
  3373=>"100100100",
  3374=>"000011011",
  3375=>"101001001",
  3376=>"001010100",
  3377=>"101000000",
  3378=>"000101111",
  3379=>"000110101",
  3380=>"110010110",
  3381=>"000000100",
  3382=>"111110110",
  3383=>"100100100",
  3384=>"011000010",
  3385=>"100001011",
  3386=>"100111111",
  3387=>"110111100",
  3388=>"110011101",
  3389=>"001011011",
  3390=>"100100110",
  3391=>"110100011",
  3392=>"101110001",
  3393=>"001000110",
  3394=>"101111010",
  3395=>"111110000",
  3396=>"001111010",
  3397=>"011010011",
  3398=>"010000011",
  3399=>"000010001",
  3400=>"011000010",
  3401=>"001001110",
  3402=>"110111011",
  3403=>"000000001",
  3404=>"100001111",
  3405=>"101001000",
  3406=>"110100011",
  3407=>"000100101",
  3408=>"111111010",
  3409=>"100001000",
  3410=>"111110110",
  3411=>"110001111",
  3412=>"111101011",
  3413=>"010011011",
  3414=>"000001010",
  3415=>"001100111",
  3416=>"111110101",
  3417=>"100110110",
  3418=>"101100001",
  3419=>"100001111",
  3420=>"010100111",
  3421=>"111100111",
  3422=>"110101101",
  3423=>"000000101",
  3424=>"011100000",
  3425=>"111110101",
  3426=>"011101011",
  3427=>"011000000",
  3428=>"110101011",
  3429=>"001000000",
  3430=>"010010001",
  3431=>"110110101",
  3432=>"111010001",
  3433=>"100010010",
  3434=>"011000100",
  3435=>"001111100",
  3436=>"110101010",
  3437=>"100110010",
  3438=>"010010010",
  3439=>"111101000",
  3440=>"011100011",
  3441=>"011110000",
  3442=>"110000001",
  3443=>"110011011",
  3444=>"011000011",
  3445=>"000111100",
  3446=>"000001111",
  3447=>"010010100",
  3448=>"010000000",
  3449=>"010101100",
  3450=>"011110000",
  3451=>"011000110",
  3452=>"111100111",
  3453=>"101111101",
  3454=>"000010000",
  3455=>"001100010",
  3456=>"001101100",
  3457=>"011100000",
  3458=>"110001100",
  3459=>"001010011",
  3460=>"001011011",
  3461=>"100011101",
  3462=>"111110001",
  3463=>"110111010",
  3464=>"100010010",
  3465=>"100111111",
  3466=>"101110110",
  3467=>"000000101",
  3468=>"000001010",
  3469=>"000001100",
  3470=>"001001100",
  3471=>"111011100",
  3472=>"101010011",
  3473=>"010010101",
  3474=>"001110001",
  3475=>"001010011",
  3476=>"100010011",
  3477=>"001110110",
  3478=>"010100001",
  3479=>"111001111",
  3480=>"100111010",
  3481=>"010010000",
  3482=>"010001000",
  3483=>"100001101",
  3484=>"011100101",
  3485=>"000011111",
  3486=>"110111001",
  3487=>"001100000",
  3488=>"101101101",
  3489=>"100101101",
  3490=>"100000001",
  3491=>"111111100",
  3492=>"011111100",
  3493=>"100010001",
  3494=>"100011111",
  3495=>"101011110",
  3496=>"001001101",
  3497=>"011110010",
  3498=>"111110111",
  3499=>"001110110",
  3500=>"000010111",
  3501=>"011010001",
  3502=>"111111111",
  3503=>"100101000",
  3504=>"000011101",
  3505=>"001001111",
  3506=>"100011101",
  3507=>"000011100",
  3508=>"000001000",
  3509=>"101010100",
  3510=>"010111011",
  3511=>"101111010",
  3512=>"001011001",
  3513=>"001101000",
  3514=>"011000001",
  3515=>"001100110",
  3516=>"001000000",
  3517=>"001000000",
  3518=>"111001101",
  3519=>"010111110",
  3520=>"000101110",
  3521=>"010100000",
  3522=>"000100011",
  3523=>"101011111",
  3524=>"000000100",
  3525=>"101001100",
  3526=>"001110000",
  3527=>"100001100",
  3528=>"111011110",
  3529=>"000001001",
  3530=>"100000001",
  3531=>"011101010",
  3532=>"001110001",
  3533=>"010110111",
  3534=>"001100101",
  3535=>"000101001",
  3536=>"101001000",
  3537=>"110000000",
  3538=>"110100011",
  3539=>"000111000",
  3540=>"101011111",
  3541=>"100110100",
  3542=>"011101101",
  3543=>"111110011",
  3544=>"101011111",
  3545=>"111110010",
  3546=>"011100101",
  3547=>"101001011",
  3548=>"010100001",
  3549=>"001110110",
  3550=>"100101110",
  3551=>"001111011",
  3552=>"111000000",
  3553=>"010111010",
  3554=>"001000000",
  3555=>"111111000",
  3556=>"101010100",
  3557=>"111110111",
  3558=>"000000111",
  3559=>"101001001",
  3560=>"011101000",
  3561=>"111110010",
  3562=>"011000100",
  3563=>"101010011",
  3564=>"001100010",
  3565=>"100100101",
  3566=>"101000100",
  3567=>"111001000",
  3568=>"111010100",
  3569=>"001101101",
  3570=>"000010000",
  3571=>"011011000",
  3572=>"001000111",
  3573=>"110000110",
  3574=>"001101001",
  3575=>"000000010",
  3576=>"110001000",
  3577=>"000000010",
  3578=>"001101011",
  3579=>"010010110",
  3580=>"000001111",
  3581=>"111001110",
  3582=>"110000100",
  3583=>"011011100",
  3584=>"000000000",
  3585=>"000010010",
  3586=>"011011000",
  3587=>"001010101",
  3588=>"000000101",
  3589=>"011010000",
  3590=>"101001101",
  3591=>"101000011",
  3592=>"101000010",
  3593=>"110111110",
  3594=>"000011001",
  3595=>"111001111",
  3596=>"010010111",
  3597=>"101101010",
  3598=>"100111111",
  3599=>"111111100",
  3600=>"111101000",
  3601=>"001010100",
  3602=>"100010100",
  3603=>"010010111",
  3604=>"101111101",
  3605=>"100011001",
  3606=>"001000111",
  3607=>"100011000",
  3608=>"100101011",
  3609=>"101000100",
  3610=>"010001010",
  3611=>"110010100",
  3612=>"110010110",
  3613=>"011111000",
  3614=>"101001000",
  3615=>"110101110",
  3616=>"101011111",
  3617=>"011010000",
  3618=>"011111101",
  3619=>"110100100",
  3620=>"101010001",
  3621=>"001101100",
  3622=>"000111110",
  3623=>"101110001",
  3624=>"101000001",
  3625=>"111000001",
  3626=>"000001011",
  3627=>"001111100",
  3628=>"110010010",
  3629=>"001001111",
  3630=>"011110010",
  3631=>"011001010",
  3632=>"010100000",
  3633=>"011010110",
  3634=>"010000001",
  3635=>"100010000",
  3636=>"010010011",
  3637=>"010010100",
  3638=>"011001101",
  3639=>"010011101",
  3640=>"001110000",
  3641=>"010100101",
  3642=>"010011100",
  3643=>"100000100",
  3644=>"000010110",
  3645=>"001111111",
  3646=>"111110001",
  3647=>"111011001",
  3648=>"010100110",
  3649=>"010101001",
  3650=>"011101000",
  3651=>"011001011",
  3652=>"111110001",
  3653=>"111111001",
  3654=>"001000000",
  3655=>"001010111",
  3656=>"011000111",
  3657=>"011100111",
  3658=>"100011110",
  3659=>"111100001",
  3660=>"101000101",
  3661=>"110001100",
  3662=>"100100110",
  3663=>"000011111",
  3664=>"011101010",
  3665=>"001000100",
  3666=>"110000110",
  3667=>"111110101",
  3668=>"110111101",
  3669=>"111111111",
  3670=>"000001011",
  3671=>"110011111",
  3672=>"101011010",
  3673=>"011111111",
  3674=>"101010101",
  3675=>"000001001",
  3676=>"110111000",
  3677=>"000000110",
  3678=>"001100001",
  3679=>"100101111",
  3680=>"100001110",
  3681=>"001110001",
  3682=>"000101011",
  3683=>"011101000",
  3684=>"001001001",
  3685=>"110001010",
  3686=>"011111010",
  3687=>"001111010",
  3688=>"001001111",
  3689=>"011011011",
  3690=>"100100101",
  3691=>"000111010",
  3692=>"000000100",
  3693=>"001001101",
  3694=>"110101001",
  3695=>"110110010",
  3696=>"111101000",
  3697=>"000100010",
  3698=>"000111111",
  3699=>"001011001",
  3700=>"100110000",
  3701=>"111111111",
  3702=>"100010000",
  3703=>"101101110",
  3704=>"001101010",
  3705=>"010001100",
  3706=>"010100101",
  3707=>"101001100",
  3708=>"011111111",
  3709=>"001110010",
  3710=>"100110001",
  3711=>"110101101",
  3712=>"110011111",
  3713=>"010010100",
  3714=>"001110111",
  3715=>"110011010",
  3716=>"011100101",
  3717=>"001100010",
  3718=>"111001011",
  3719=>"000111011",
  3720=>"000011011",
  3721=>"010000011",
  3722=>"011111111",
  3723=>"100001110",
  3724=>"000110010",
  3725=>"101001100",
  3726=>"100110111",
  3727=>"111011011",
  3728=>"000111000",
  3729=>"000000010",
  3730=>"010001101",
  3731=>"101010100",
  3732=>"010100001",
  3733=>"111010101",
  3734=>"010111010",
  3735=>"111111101",
  3736=>"100101001",
  3737=>"101010001",
  3738=>"011100111",
  3739=>"101010100",
  3740=>"001111000",
  3741=>"110111001",
  3742=>"101111111",
  3743=>"011011111",
  3744=>"011111100",
  3745=>"111111011",
  3746=>"011110011",
  3747=>"010100111",
  3748=>"111110100",
  3749=>"110011100",
  3750=>"110110110",
  3751=>"011100101",
  3752=>"111001010",
  3753=>"110001101",
  3754=>"110010110",
  3755=>"000100111",
  3756=>"000000101",
  3757=>"110010110",
  3758=>"010011111",
  3759=>"010011000",
  3760=>"001010100",
  3761=>"100101101",
  3762=>"001100000",
  3763=>"110101100",
  3764=>"111111111",
  3765=>"110111011",
  3766=>"111111101",
  3767=>"101000111",
  3768=>"001000111",
  3769=>"001010001",
  3770=>"101001111",
  3771=>"100010010",
  3772=>"111011111",
  3773=>"111010011",
  3774=>"000100001",
  3775=>"011010000",
  3776=>"010100101",
  3777=>"001111101",
  3778=>"100101111",
  3779=>"011000111",
  3780=>"101110001",
  3781=>"000110001",
  3782=>"101101011",
  3783=>"110101001",
  3784=>"101101101",
  3785=>"000001111",
  3786=>"010001111",
  3787=>"100001011",
  3788=>"100110001",
  3789=>"110110000",
  3790=>"110111111",
  3791=>"000001011",
  3792=>"111110110",
  3793=>"110100001",
  3794=>"111101000",
  3795=>"101011001",
  3796=>"010001100",
  3797=>"000001001",
  3798=>"000000110",
  3799=>"111110101",
  3800=>"011000000",
  3801=>"001010010",
  3802=>"001101010",
  3803=>"000100000",
  3804=>"010011010",
  3805=>"111100010",
  3806=>"000010001",
  3807=>"010001111",
  3808=>"101011100",
  3809=>"000010111",
  3810=>"111001001",
  3811=>"001000001",
  3812=>"100001011",
  3813=>"010110100",
  3814=>"011000011",
  3815=>"010111100",
  3816=>"000100000",
  3817=>"011100111",
  3818=>"100000100",
  3819=>"000100011",
  3820=>"000010100",
  3821=>"000111000",
  3822=>"101101110",
  3823=>"101100101",
  3824=>"001000110",
  3825=>"100110010",
  3826=>"100010111",
  3827=>"110110010",
  3828=>"110100000",
  3829=>"001101100",
  3830=>"000111000",
  3831=>"010001010",
  3832=>"100101110",
  3833=>"111011110",
  3834=>"110010000",
  3835=>"010010111",
  3836=>"001010101",
  3837=>"100111101",
  3838=>"111001011",
  3839=>"000001001",
  3840=>"000010010",
  3841=>"110111010",
  3842=>"001111001",
  3843=>"100011010",
  3844=>"001100100",
  3845=>"111111101",
  3846=>"111001100",
  3847=>"110100101",
  3848=>"011010110",
  3849=>"100001000",
  3850=>"100010111",
  3851=>"011111111",
  3852=>"110001000",
  3853=>"100100010",
  3854=>"100101110",
  3855=>"001001000",
  3856=>"100010001",
  3857=>"111011100",
  3858=>"001110100",
  3859=>"101101000",
  3860=>"111101011",
  3861=>"101001101",
  3862=>"011000100",
  3863=>"000100010",
  3864=>"011010111",
  3865=>"110011101",
  3866=>"000101001",
  3867=>"011101111",
  3868=>"111110110",
  3869=>"000110111",
  3870=>"101000000",
  3871=>"010111001",
  3872=>"010111110",
  3873=>"010100010",
  3874=>"100001101",
  3875=>"101111011",
  3876=>"000100100",
  3877=>"010110110",
  3878=>"110101100",
  3879=>"001010011",
  3880=>"011110010",
  3881=>"010111011",
  3882=>"101011000",
  3883=>"100111111",
  3884=>"010010011",
  3885=>"111111100",
  3886=>"010000010",
  3887=>"001011110",
  3888=>"110111011",
  3889=>"000011001",
  3890=>"111100101",
  3891=>"000010010",
  3892=>"101000010",
  3893=>"000101100",
  3894=>"110101011",
  3895=>"000100101",
  3896=>"010010011",
  3897=>"101101011",
  3898=>"000001111",
  3899=>"100010010",
  3900=>"101000001",
  3901=>"111111000",
  3902=>"001110001",
  3903=>"000001011",
  3904=>"100100011",
  3905=>"010010010",
  3906=>"100011110",
  3907=>"100000111",
  3908=>"000000000",
  3909=>"010000001",
  3910=>"101110000",
  3911=>"010101010",
  3912=>"101100100",
  3913=>"001011001",
  3914=>"001011110",
  3915=>"010110000",
  3916=>"000010110",
  3917=>"111100110",
  3918=>"101011100",
  3919=>"110111000",
  3920=>"101000111",
  3921=>"001010111",
  3922=>"000001101",
  3923=>"111000000",
  3924=>"101100101",
  3925=>"100100100",
  3926=>"001011101",
  3927=>"010001001",
  3928=>"000010010",
  3929=>"100110010",
  3930=>"110011100",
  3931=>"111101101",
  3932=>"011010101",
  3933=>"101000010",
  3934=>"000000110",
  3935=>"001110101",
  3936=>"101101001",
  3937=>"110110001",
  3938=>"000101101",
  3939=>"110010100",
  3940=>"111100100",
  3941=>"110101011",
  3942=>"000100111",
  3943=>"110001110",
  3944=>"111100010",
  3945=>"110111100",
  3946=>"101100111",
  3947=>"101011111",
  3948=>"000111101",
  3949=>"101001001",
  3950=>"100000100",
  3951=>"100100111",
  3952=>"000110100",
  3953=>"010001111",
  3954=>"100001011",
  3955=>"011110101",
  3956=>"000111100",
  3957=>"010000111",
  3958=>"010000100",
  3959=>"000010001",
  3960=>"000111001",
  3961=>"010101100",
  3962=>"100111011",
  3963=>"000000110",
  3964=>"000101100",
  3965=>"101011111",
  3966=>"010100100",
  3967=>"010000001",
  3968=>"000010100",
  3969=>"001010000",
  3970=>"001100011",
  3971=>"010010111",
  3972=>"101000101",
  3973=>"100011101",
  3974=>"000000001",
  3975=>"111011101",
  3976=>"111110011",
  3977=>"100100000",
  3978=>"010010010",
  3979=>"100000011",
  3980=>"010110000",
  3981=>"100010111",
  3982=>"000111100",
  3983=>"101111100",
  3984=>"111110010",
  3985=>"001000110",
  3986=>"110110100",
  3987=>"111011100",
  3988=>"010011001",
  3989=>"010000101",
  3990=>"010000100",
  3991=>"011010010",
  3992=>"110001110",
  3993=>"101101010",
  3994=>"001010111",
  3995=>"000010000",
  3996=>"001001000",
  3997=>"010010001",
  3998=>"010010100",
  3999=>"100000001",
  4000=>"011001000",
  4001=>"011101000",
  4002=>"011011100",
  4003=>"000011100",
  4004=>"001101011",
  4005=>"001101011",
  4006=>"011000001",
  4007=>"010110111",
  4008=>"100101110",
  4009=>"001101001",
  4010=>"111111100",
  4011=>"010101100",
  4012=>"011010010",
  4013=>"001110101",
  4014=>"010101010",
  4015=>"100101111",
  4016=>"000000101",
  4017=>"000111111",
  4018=>"010110111",
  4019=>"011010010",
  4020=>"111010010",
  4021=>"011001110",
  4022=>"010011110",
  4023=>"100010111",
  4024=>"001010100",
  4025=>"000110111",
  4026=>"111111000",
  4027=>"000001100",
  4028=>"001110000",
  4029=>"101001001",
  4030=>"111011010",
  4031=>"111010000",
  4032=>"100110000",
  4033=>"001100101",
  4034=>"010001101",
  4035=>"111001111",
  4036=>"000011101",
  4037=>"001111001",
  4038=>"010100000",
  4039=>"100011111",
  4040=>"111111111",
  4041=>"100000100",
  4042=>"110000111",
  4043=>"011101011",
  4044=>"001111000",
  4045=>"100001011",
  4046=>"110101010",
  4047=>"001111011",
  4048=>"000010010",
  4049=>"101000111",
  4050=>"011010011",
  4051=>"100000100",
  4052=>"100011110",
  4053=>"011001101",
  4054=>"100100110",
  4055=>"011100110",
  4056=>"010000000",
  4057=>"111010001",
  4058=>"101111111",
  4059=>"000101011",
  4060=>"100110111",
  4061=>"000110010",
  4062=>"101001110",
  4063=>"001001111",
  4064=>"111111111",
  4065=>"000001111",
  4066=>"011101000",
  4067=>"001011111",
  4068=>"001010001",
  4069=>"001011001",
  4070=>"001001001",
  4071=>"110101000",
  4072=>"101010111",
  4073=>"001101111",
  4074=>"111011110",
  4075=>"010001010",
  4076=>"110110101",
  4077=>"011101100",
  4078=>"001001110",
  4079=>"100101100",
  4080=>"000101100",
  4081=>"100001010",
  4082=>"010000111",
  4083=>"011011110",
  4084=>"100100011",
  4085=>"110111001",
  4086=>"000110110",
  4087=>"000000011",
  4088=>"000110010",
  4089=>"110101100",
  4090=>"011000010",
  4091=>"110101100",
  4092=>"000011000",
  4093=>"100000010",
  4094=>"100011110",
  4095=>"100000010",
  4096=>"001000111",
  4097=>"101011001",
  4098=>"010011010",
  4099=>"110100010",
  4100=>"100011001",
  4101=>"001000010",
  4102=>"011001111",
  4103=>"101001101",
  4104=>"011000101",
  4105=>"000010000",
  4106=>"001011111",
  4107=>"001010010",
  4108=>"111000111",
  4109=>"010010100",
  4110=>"110101000",
  4111=>"110010101",
  4112=>"110100110",
  4113=>"010101100",
  4114=>"011011110",
  4115=>"110000010",
  4116=>"011000011",
  4117=>"010001001",
  4118=>"110111010",
  4119=>"000110100",
  4120=>"110011101",
  4121=>"000111011",
  4122=>"010010110",
  4123=>"100011000",
  4124=>"111001101",
  4125=>"011111000",
  4126=>"010010010",
  4127=>"000110000",
  4128=>"011100110",
  4129=>"110100011",
  4130=>"101100000",
  4131=>"000101011",
  4132=>"101111010",
  4133=>"110011011",
  4134=>"010000110",
  4135=>"101101011",
  4136=>"010000000",
  4137=>"110101110",
  4138=>"011100000",
  4139=>"110011100",
  4140=>"001100000",
  4141=>"011011001",
  4142=>"001010000",
  4143=>"110101000",
  4144=>"101100101",
  4145=>"011011000",
  4146=>"011000101",
  4147=>"001001100",
  4148=>"001111010",
  4149=>"111000111",
  4150=>"010101100",
  4151=>"100101110",
  4152=>"010010001",
  4153=>"000011110",
  4154=>"100110100",
  4155=>"110100100",
  4156=>"101001111",
  4157=>"100110001",
  4158=>"100110100",
  4159=>"101000000",
  4160=>"001111111",
  4161=>"010000001",
  4162=>"000110010",
  4163=>"011010110",
  4164=>"111111110",
  4165=>"000010000",
  4166=>"000111110",
  4167=>"111110010",
  4168=>"011011011",
  4169=>"111100101",
  4170=>"011101011",
  4171=>"100101111",
  4172=>"100010100",
  4173=>"111101010",
  4174=>"011110000",
  4175=>"001101101",
  4176=>"001101111",
  4177=>"000010011",
  4178=>"110111101",
  4179=>"001001100",
  4180=>"011100001",
  4181=>"010110001",
  4182=>"110100101",
  4183=>"101111111",
  4184=>"110011100",
  4185=>"110011100",
  4186=>"011111001",
  4187=>"010001010",
  4188=>"011111000",
  4189=>"111000110",
  4190=>"111010010",
  4191=>"000001010",
  4192=>"100000100",
  4193=>"101011101",
  4194=>"111011000",
  4195=>"000000100",
  4196=>"101001001",
  4197=>"011100011",
  4198=>"001000010",
  4199=>"101001101",
  4200=>"101000100",
  4201=>"111110101",
  4202=>"110010110",
  4203=>"011100001",
  4204=>"101111010",
  4205=>"001000011",
  4206=>"100000100",
  4207=>"000101111",
  4208=>"000101101",
  4209=>"100001100",
  4210=>"100111100",
  4211=>"100000000",
  4212=>"001100100",
  4213=>"001101100",
  4214=>"111001001",
  4215=>"001011101",
  4216=>"001011100",
  4217=>"000100100",
  4218=>"001111110",
  4219=>"010011010",
  4220=>"010000110",
  4221=>"111111111",
  4222=>"000001111",
  4223=>"001000100",
  4224=>"000111110",
  4225=>"001100011",
  4226=>"000110011",
  4227=>"100110101",
  4228=>"101101100",
  4229=>"110011110",
  4230=>"000111011",
  4231=>"000010111",
  4232=>"111011011",
  4233=>"000000101",
  4234=>"110011011",
  4235=>"111101100",
  4236=>"011010001",
  4237=>"110100110",
  4238=>"111010010",
  4239=>"011000000",
  4240=>"111011010",
  4241=>"111110010",
  4242=>"111111100",
  4243=>"000010010",
  4244=>"010010100",
  4245=>"110100100",
  4246=>"010111011",
  4247=>"011011110",
  4248=>"110110111",
  4249=>"001000110",
  4250=>"011011111",
  4251=>"110111000",
  4252=>"001100000",
  4253=>"010101001",
  4254=>"111001101",
  4255=>"001100000",
  4256=>"101000000",
  4257=>"011110111",
  4258=>"101010000",
  4259=>"101101100",
  4260=>"001101000",
  4261=>"100111000",
  4262=>"000111111",
  4263=>"001100010",
  4264=>"101011000",
  4265=>"111000111",
  4266=>"010111111",
  4267=>"101001001",
  4268=>"110010000",
  4269=>"000101011",
  4270=>"101101010",
  4271=>"010010100",
  4272=>"100011000",
  4273=>"011110001",
  4274=>"011001110",
  4275=>"100000001",
  4276=>"001000001",
  4277=>"001101001",
  4278=>"100100111",
  4279=>"011100111",
  4280=>"001000001",
  4281=>"001001111",
  4282=>"100010110",
  4283=>"000111011",
  4284=>"110010110",
  4285=>"100001101",
  4286=>"000001110",
  4287=>"100010000",
  4288=>"110101101",
  4289=>"101100111",
  4290=>"110010000",
  4291=>"110111001",
  4292=>"000000011",
  4293=>"010111111",
  4294=>"000010001",
  4295=>"110000111",
  4296=>"010111000",
  4297=>"101101110",
  4298=>"101111100",
  4299=>"011110110",
  4300=>"111111000",
  4301=>"000101010",
  4302=>"011010100",
  4303=>"000011110",
  4304=>"011101011",
  4305=>"101010110",
  4306=>"001001111",
  4307=>"000111000",
  4308=>"011100011",
  4309=>"101010101",
  4310=>"100010100",
  4311=>"001111110",
  4312=>"101011001",
  4313=>"111000011",
  4314=>"101010101",
  4315=>"110101010",
  4316=>"000010001",
  4317=>"011111011",
  4318=>"101110011",
  4319=>"101111011",
  4320=>"111010111",
  4321=>"100111000",
  4322=>"000000111",
  4323=>"000010100",
  4324=>"010100001",
  4325=>"000101111",
  4326=>"011000111",
  4327=>"010111110",
  4328=>"110000101",
  4329=>"001010110",
  4330=>"000001010",
  4331=>"101001000",
  4332=>"110001000",
  4333=>"001101100",
  4334=>"010111111",
  4335=>"100110111",
  4336=>"111100110",
  4337=>"011010111",
  4338=>"100011011",
  4339=>"000101111",
  4340=>"101010010",
  4341=>"111000110",
  4342=>"111010000",
  4343=>"111110010",
  4344=>"001100010",
  4345=>"111101000",
  4346=>"101111100",
  4347=>"010000011",
  4348=>"001100101",
  4349=>"110011101",
  4350=>"000101001",
  4351=>"111010010",
  4352=>"111100111",
  4353=>"000010000",
  4354=>"111100010",
  4355=>"010011110",
  4356=>"001000011",
  4357=>"010111101",
  4358=>"100000110",
  4359=>"011111100",
  4360=>"100001101",
  4361=>"011010111",
  4362=>"010100000",
  4363=>"010100111",
  4364=>"100010010",
  4365=>"010110000",
  4366=>"001001010",
  4367=>"110001100",
  4368=>"010011101",
  4369=>"001110111",
  4370=>"001110111",
  4371=>"100101010",
  4372=>"111110011",
  4373=>"101101111",
  4374=>"111001000",
  4375=>"000101011",
  4376=>"000010010",
  4377=>"110111001",
  4378=>"011000010",
  4379=>"001011000",
  4380=>"101101001",
  4381=>"001001010",
  4382=>"001000010",
  4383=>"100000001",
  4384=>"101000000",
  4385=>"100110110",
  4386=>"000010101",
  4387=>"001001110",
  4388=>"010111110",
  4389=>"000010000",
  4390=>"110001101",
  4391=>"100100011",
  4392=>"110011000",
  4393=>"111111001",
  4394=>"100010100",
  4395=>"100000101",
  4396=>"010101001",
  4397=>"101011001",
  4398=>"110010100",
  4399=>"101000001",
  4400=>"110000100",
  4401=>"110000101",
  4402=>"110010101",
  4403=>"011000110",
  4404=>"101001001",
  4405=>"110010111",
  4406=>"111010001",
  4407=>"010100000",
  4408=>"001111001",
  4409=>"010001110",
  4410=>"001110111",
  4411=>"000100000",
  4412=>"111110000",
  4413=>"110010011",
  4414=>"001001100",
  4415=>"010101001",
  4416=>"101101111",
  4417=>"010001101",
  4418=>"000011100",
  4419=>"000011011",
  4420=>"011110111",
  4421=>"000010111",
  4422=>"011101111",
  4423=>"000001110",
  4424=>"000110000",
  4425=>"010001110",
  4426=>"111001110",
  4427=>"111100001",
  4428=>"101111010",
  4429=>"110111101",
  4430=>"000110110",
  4431=>"110011011",
  4432=>"000100101",
  4433=>"110000111",
  4434=>"101001000",
  4435=>"011110101",
  4436=>"001001010",
  4437=>"111100001",
  4438=>"001110001",
  4439=>"110011111",
  4440=>"000111101",
  4441=>"110001000",
  4442=>"111110111",
  4443=>"110000010",
  4444=>"111100111",
  4445=>"010000101",
  4446=>"100110101",
  4447=>"111101000",
  4448=>"100111011",
  4449=>"001100000",
  4450=>"101100001",
  4451=>"000001101",
  4452=>"001000001",
  4453=>"111101111",
  4454=>"111110111",
  4455=>"101010100",
  4456=>"001010101",
  4457=>"111000000",
  4458=>"111100010",
  4459=>"010110011",
  4460=>"110110010",
  4461=>"111001011",
  4462=>"001000000",
  4463=>"110110100",
  4464=>"110010110",
  4465=>"010000111",
  4466=>"101011000",
  4467=>"011010101",
  4468=>"111000001",
  4469=>"101001100",
  4470=>"111110010",
  4471=>"110110001",
  4472=>"100110000",
  4473=>"000011111",
  4474=>"000110011",
  4475=>"011010010",
  4476=>"101001111",
  4477=>"000110000",
  4478=>"101101100",
  4479=>"010000100",
  4480=>"111010011",
  4481=>"010001001",
  4482=>"110011000",
  4483=>"001110011",
  4484=>"110101011",
  4485=>"010110110",
  4486=>"111101010",
  4487=>"110110100",
  4488=>"000000111",
  4489=>"111001100",
  4490=>"110011100",
  4491=>"111010011",
  4492=>"110100000",
  4493=>"001010000",
  4494=>"101101100",
  4495=>"100101001",
  4496=>"000110110",
  4497=>"100001001",
  4498=>"110001001",
  4499=>"010011010",
  4500=>"100000111",
  4501=>"011010010",
  4502=>"001100101",
  4503=>"111100010",
  4504=>"000110001",
  4505=>"100000001",
  4506=>"110111010",
  4507=>"110010000",
  4508=>"010101000",
  4509=>"111011001",
  4510=>"111000000",
  4511=>"101110001",
  4512=>"001111010",
  4513=>"011101101",
  4514=>"001000100",
  4515=>"000100011",
  4516=>"000101111",
  4517=>"101110111",
  4518=>"011010001",
  4519=>"110010001",
  4520=>"000001110",
  4521=>"000101110",
  4522=>"100010110",
  4523=>"001100010",
  4524=>"100000001",
  4525=>"011111110",
  4526=>"011000111",
  4527=>"100010001",
  4528=>"011010100",
  4529=>"010011001",
  4530=>"111011011",
  4531=>"111001010",
  4532=>"100010000",
  4533=>"010100101",
  4534=>"001010100",
  4535=>"111110001",
  4536=>"000101001",
  4537=>"100000010",
  4538=>"011100111",
  4539=>"111000101",
  4540=>"010001010",
  4541=>"101000111",
  4542=>"000000101",
  4543=>"100101000",
  4544=>"110100111",
  4545=>"101011101",
  4546=>"011111011",
  4547=>"000000100",
  4548=>"111000011",
  4549=>"110111011",
  4550=>"110110000",
  4551=>"011010011",
  4552=>"101001100",
  4553=>"100110011",
  4554=>"010111111",
  4555=>"100110101",
  4556=>"001111101",
  4557=>"100110110",
  4558=>"111111011",
  4559=>"101001001",
  4560=>"000001111",
  4561=>"111100010",
  4562=>"001001010",
  4563=>"000011111",
  4564=>"101000000",
  4565=>"100111001",
  4566=>"011000001",
  4567=>"100101010",
  4568=>"100110110",
  4569=>"000000100",
  4570=>"111011110",
  4571=>"110100100",
  4572=>"000010100",
  4573=>"111001110",
  4574=>"011110101",
  4575=>"000000110",
  4576=>"110101110",
  4577=>"000111101",
  4578=>"011010011",
  4579=>"001110011",
  4580=>"110000010",
  4581=>"110110010",
  4582=>"010000000",
  4583=>"000000000",
  4584=>"100101100",
  4585=>"000000100",
  4586=>"010000000",
  4587=>"101111110",
  4588=>"010110100",
  4589=>"111110000",
  4590=>"010111001",
  4591=>"110100011",
  4592=>"011111000",
  4593=>"011100010",
  4594=>"100110010",
  4595=>"000111110",
  4596=>"101000111",
  4597=>"000011111",
  4598=>"010010001",
  4599=>"101111110",
  4600=>"010100010",
  4601=>"001100011",
  4602=>"100111111",
  4603=>"101111001",
  4604=>"000110010",
  4605=>"100110010",
  4606=>"001101100",
  4607=>"101010111",
  4608=>"100001111",
  4609=>"100111101",
  4610=>"011110001",
  4611=>"111111011",
  4612=>"101000110",
  4613=>"111010010",
  4614=>"011000101",
  4615=>"001000010",
  4616=>"000010000",
  4617=>"000111000",
  4618=>"100111001",
  4619=>"000001111",
  4620=>"011110010",
  4621=>"100010000",
  4622=>"000110000",
  4623=>"110110011",
  4624=>"111111011",
  4625=>"101000010",
  4626=>"100100110",
  4627=>"111100001",
  4628=>"011111011",
  4629=>"101111101",
  4630=>"010010100",
  4631=>"001001110",
  4632=>"001010010",
  4633=>"110100010",
  4634=>"101001100",
  4635=>"111101111",
  4636=>"100100001",
  4637=>"100110100",
  4638=>"011001000",
  4639=>"101001000",
  4640=>"011000110",
  4641=>"100010001",
  4642=>"010000101",
  4643=>"001011110",
  4644=>"000010000",
  4645=>"001100011",
  4646=>"111111000",
  4647=>"000000100",
  4648=>"010011111",
  4649=>"011111101",
  4650=>"110110101",
  4651=>"010011111",
  4652=>"011010100",
  4653=>"000010010",
  4654=>"110111100",
  4655=>"110000101",
  4656=>"010000110",
  4657=>"111111110",
  4658=>"101101011",
  4659=>"001010010",
  4660=>"110011111",
  4661=>"000111011",
  4662=>"100011010",
  4663=>"000001001",
  4664=>"101100100",
  4665=>"110000111",
  4666=>"011001100",
  4667=>"100100101",
  4668=>"010001110",
  4669=>"100111010",
  4670=>"000011110",
  4671=>"100110101",
  4672=>"110111110",
  4673=>"111110001",
  4674=>"110011111",
  4675=>"001111011",
  4676=>"111111111",
  4677=>"110111010",
  4678=>"100101101",
  4679=>"001111110",
  4680=>"001001011",
  4681=>"101001101",
  4682=>"111000111",
  4683=>"001101110",
  4684=>"000010110",
  4685=>"010010010",
  4686=>"110011010",
  4687=>"001001110",
  4688=>"000010000",
  4689=>"110001001",
  4690=>"100000010",
  4691=>"101010001",
  4692=>"111000000",
  4693=>"010100010",
  4694=>"101110010",
  4695=>"100011010",
  4696=>"101001101",
  4697=>"101001111",
  4698=>"001101111",
  4699=>"000001011",
  4700=>"101100100",
  4701=>"000101011",
  4702=>"000111010",
  4703=>"111110110",
  4704=>"101101000",
  4705=>"110001000",
  4706=>"001001010",
  4707=>"101101100",
  4708=>"101001011",
  4709=>"011110000",
  4710=>"100010111",
  4711=>"101111010",
  4712=>"101100101",
  4713=>"101001010",
  4714=>"100011111",
  4715=>"110011100",
  4716=>"000001100",
  4717=>"001110100",
  4718=>"000000101",
  4719=>"100001000",
  4720=>"101111111",
  4721=>"100010100",
  4722=>"110001111",
  4723=>"011100001",
  4724=>"010110110",
  4725=>"000011100",
  4726=>"101001000",
  4727=>"000100101",
  4728=>"010011101",
  4729=>"000111111",
  4730=>"111100100",
  4731=>"110100000",
  4732=>"000000100",
  4733=>"011001101",
  4734=>"001011110",
  4735=>"110001000",
  4736=>"110110111",
  4737=>"011011001",
  4738=>"101100000",
  4739=>"001001101",
  4740=>"110100101",
  4741=>"100000101",
  4742=>"011110011",
  4743=>"101001111",
  4744=>"110011101",
  4745=>"011000110",
  4746=>"001100101",
  4747=>"010001011",
  4748=>"111011111",
  4749=>"111101101",
  4750=>"010100100",
  4751=>"100001011",
  4752=>"111111111",
  4753=>"011011001",
  4754=>"111000110",
  4755=>"111111011",
  4756=>"111100100",
  4757=>"011111110",
  4758=>"011100110",
  4759=>"010010111",
  4760=>"100100101",
  4761=>"101100011",
  4762=>"100111010",
  4763=>"100110111",
  4764=>"000110111",
  4765=>"001101010",
  4766=>"001100110",
  4767=>"011111101",
  4768=>"001100010",
  4769=>"001000000",
  4770=>"001000010",
  4771=>"011111111",
  4772=>"110110101",
  4773=>"000000010",
  4774=>"110001101",
  4775=>"010000000",
  4776=>"111000000",
  4777=>"001101011",
  4778=>"011100001",
  4779=>"110001100",
  4780=>"001011011",
  4781=>"110001001",
  4782=>"100111001",
  4783=>"100001111",
  4784=>"011100001",
  4785=>"101001011",
  4786=>"011110000",
  4787=>"001001000",
  4788=>"100001011",
  4789=>"001111100",
  4790=>"111001000",
  4791=>"110001010",
  4792=>"011000110",
  4793=>"101001101",
  4794=>"000000100",
  4795=>"100100100",
  4796=>"000111011",
  4797=>"110111001",
  4798=>"001101101",
  4799=>"100001000",
  4800=>"100001101",
  4801=>"000001101",
  4802=>"111001110",
  4803=>"110111010",
  4804=>"110111110",
  4805=>"000110111",
  4806=>"111011111",
  4807=>"001100000",
  4808=>"010010111",
  4809=>"001100000",
  4810=>"101110110",
  4811=>"001110100",
  4812=>"101000000",
  4813=>"111101001",
  4814=>"010100101",
  4815=>"111101010",
  4816=>"110011000",
  4817=>"100110100",
  4818=>"011100111",
  4819=>"100010001",
  4820=>"100000011",
  4821=>"110010110",
  4822=>"000101100",
  4823=>"011101100",
  4824=>"001010101",
  4825=>"101101000",
  4826=>"010011110",
  4827=>"111111001",
  4828=>"100100010",
  4829=>"111111011",
  4830=>"001000011",
  4831=>"001010010",
  4832=>"000100001",
  4833=>"110111101",
  4834=>"000111011",
  4835=>"000111011",
  4836=>"110101000",
  4837=>"011001111",
  4838=>"101011010",
  4839=>"111011000",
  4840=>"000100001",
  4841=>"010100101",
  4842=>"000000111",
  4843=>"011011101",
  4844=>"100010000",
  4845=>"011010111",
  4846=>"110100000",
  4847=>"010010011",
  4848=>"111111111",
  4849=>"001001101",
  4850=>"110100011",
  4851=>"010000011",
  4852=>"111010011",
  4853=>"001000101",
  4854=>"100000101",
  4855=>"011110011",
  4856=>"110011101",
  4857=>"000101000",
  4858=>"000100101",
  4859=>"010000110",
  4860=>"110111111",
  4861=>"110100110",
  4862=>"011100101",
  4863=>"001010100",
  4864=>"001000010",
  4865=>"010000110",
  4866=>"111110000",
  4867=>"110100001",
  4868=>"111101001",
  4869=>"011010011",
  4870=>"100111011",
  4871=>"110100110",
  4872=>"101101011",
  4873=>"010010100",
  4874=>"011001101",
  4875=>"110100100",
  4876=>"000110001",
  4877=>"100101110",
  4878=>"000010011",
  4879=>"100010110",
  4880=>"111001000",
  4881=>"011001101",
  4882=>"100001001",
  4883=>"010001100",
  4884=>"010010111",
  4885=>"101010101",
  4886=>"100011110",
  4887=>"000000010",
  4888=>"110001011",
  4889=>"101000111",
  4890=>"100101010",
  4891=>"001001111",
  4892=>"001010001",
  4893=>"001010111",
  4894=>"010101100",
  4895=>"001001101",
  4896=>"000001110",
  4897=>"100101110",
  4898=>"111100000",
  4899=>"110011110",
  4900=>"011100010",
  4901=>"110111101",
  4902=>"100110000",
  4903=>"111100101",
  4904=>"100000000",
  4905=>"010001101",
  4906=>"000001110",
  4907=>"001101001",
  4908=>"011111011",
  4909=>"100101101",
  4910=>"100101010",
  4911=>"110101000",
  4912=>"101110100",
  4913=>"000101000",
  4914=>"000000100",
  4915=>"001111100",
  4916=>"111100000",
  4917=>"000010011",
  4918=>"011110110",
  4919=>"000110011",
  4920=>"011011010",
  4921=>"100110011",
  4922=>"001011110",
  4923=>"111000010",
  4924=>"100111111",
  4925=>"000101011",
  4926=>"000000011",
  4927=>"110110001",
  4928=>"110010111",
  4929=>"100001010",
  4930=>"011010010",
  4931=>"110010110",
  4932=>"101101010",
  4933=>"011001101",
  4934=>"010001110",
  4935=>"100000101",
  4936=>"100101110",
  4937=>"110011110",
  4938=>"000101101",
  4939=>"000110011",
  4940=>"011010010",
  4941=>"011111110",
  4942=>"000011000",
  4943=>"110110011",
  4944=>"000111011",
  4945=>"111101100",
  4946=>"111010000",
  4947=>"011000000",
  4948=>"010101010",
  4949=>"111001000",
  4950=>"111101110",
  4951=>"011010110",
  4952=>"100101000",
  4953=>"010010011",
  4954=>"001101011",
  4955=>"110010111",
  4956=>"001001100",
  4957=>"110001110",
  4958=>"000100001",
  4959=>"010010111",
  4960=>"110100110",
  4961=>"100011011",
  4962=>"001010010",
  4963=>"100011111",
  4964=>"101100000",
  4965=>"110000001",
  4966=>"100101101",
  4967=>"110111001",
  4968=>"011000110",
  4969=>"101111110",
  4970=>"110100001",
  4971=>"101111001",
  4972=>"011001101",
  4973=>"011110101",
  4974=>"011000001",
  4975=>"001101100",
  4976=>"100000110",
  4977=>"011110100",
  4978=>"100000001",
  4979=>"111011111",
  4980=>"111110010",
  4981=>"010100010",
  4982=>"000000001",
  4983=>"010010110",
  4984=>"110000010",
  4985=>"000110011",
  4986=>"111101000",
  4987=>"000110010",
  4988=>"000101000",
  4989=>"110101110",
  4990=>"011001101",
  4991=>"011111000",
  4992=>"010011011",
  4993=>"011111001",
  4994=>"001100000",
  4995=>"011010000",
  4996=>"001110100",
  4997=>"000110011",
  4998=>"110111010",
  4999=>"100101101",
  5000=>"110111110",
  5001=>"011100000",
  5002=>"010000111",
  5003=>"011111110",
  5004=>"010110011",
  5005=>"010011110",
  5006=>"000100110",
  5007=>"010111011",
  5008=>"000000110",
  5009=>"001110101",
  5010=>"000111001",
  5011=>"000101011",
  5012=>"100101000",
  5013=>"101101110",
  5014=>"000100110",
  5015=>"001111110",
  5016=>"100000101",
  5017=>"111000111",
  5018=>"000111000",
  5019=>"101000011",
  5020=>"101001100",
  5021=>"000011100",
  5022=>"101010111",
  5023=>"111010001",
  5024=>"010011100",
  5025=>"110110000",
  5026=>"100111010",
  5027=>"110010100",
  5028=>"010000100",
  5029=>"011111011",
  5030=>"110000010",
  5031=>"100111010",
  5032=>"110010111",
  5033=>"110010111",
  5034=>"110101001",
  5035=>"100010101",
  5036=>"100100111",
  5037=>"001100000",
  5038=>"100000100",
  5039=>"011100001",
  5040=>"000100111",
  5041=>"011100011",
  5042=>"110011110",
  5043=>"000000100",
  5044=>"110101100",
  5045=>"100010000",
  5046=>"101001111",
  5047=>"101111011",
  5048=>"101000111",
  5049=>"110110111",
  5050=>"000111010",
  5051=>"010110101",
  5052=>"100100111",
  5053=>"001100011",
  5054=>"011011000",
  5055=>"010010100",
  5056=>"100111111",
  5057=>"000010011",
  5058=>"100010001",
  5059=>"110110101",
  5060=>"011000110",
  5061=>"001110100",
  5062=>"110100111",
  5063=>"110000010",
  5064=>"001101000",
  5065=>"111110100",
  5066=>"110110110",
  5067=>"100011100",
  5068=>"111110100",
  5069=>"101000011",
  5070=>"001101000",
  5071=>"101111010",
  5072=>"001011110",
  5073=>"001110100",
  5074=>"111000001",
  5075=>"100010000",
  5076=>"000100100",
  5077=>"011110111",
  5078=>"011010001",
  5079=>"101101000",
  5080=>"110101000",
  5081=>"011001101",
  5082=>"111100111",
  5083=>"101111101",
  5084=>"110100111",
  5085=>"101000000",
  5086=>"010110100",
  5087=>"110000100",
  5088=>"101000111",
  5089=>"101010001",
  5090=>"111111000",
  5091=>"000110000",
  5092=>"110010101",
  5093=>"010001100",
  5094=>"111101011",
  5095=>"001001000",
  5096=>"100000101",
  5097=>"001110010",
  5098=>"000001111",
  5099=>"110010111",
  5100=>"111000110",
  5101=>"001110011",
  5102=>"010100111",
  5103=>"000100110",
  5104=>"000111100",
  5105=>"000111010",
  5106=>"001000000",
  5107=>"010101101",
  5108=>"010010011",
  5109=>"010000000",
  5110=>"010110111",
  5111=>"101000010",
  5112=>"101101111",
  5113=>"010001111",
  5114=>"110000110",
  5115=>"101110111",
  5116=>"010000110",
  5117=>"100001000",
  5118=>"101101111",
  5119=>"110010001",
  5120=>"100011100",
  5121=>"101101011",
  5122=>"011100010",
  5123=>"111001110",
  5124=>"011000110",
  5125=>"000101000",
  5126=>"100000111",
  5127=>"011100000",
  5128=>"100100100",
  5129=>"010011110",
  5130=>"000100111",
  5131=>"101111100",
  5132=>"110000011",
  5133=>"000010011",
  5134=>"000111110",
  5135=>"110110010",
  5136=>"101000110",
  5137=>"101100110",
  5138=>"011000000",
  5139=>"110100111",
  5140=>"001000000",
  5141=>"000001011",
  5142=>"101111011",
  5143=>"000101101",
  5144=>"110010001",
  5145=>"111101100",
  5146=>"001111001",
  5147=>"110101101",
  5148=>"010101011",
  5149=>"000000000",
  5150=>"001000010",
  5151=>"011010001",
  5152=>"110111101",
  5153=>"110111001",
  5154=>"011100101",
  5155=>"100100111",
  5156=>"110110111",
  5157=>"010111111",
  5158=>"101100011",
  5159=>"010001100",
  5160=>"101100100",
  5161=>"000010111",
  5162=>"111000000",
  5163=>"101101010",
  5164=>"110011001",
  5165=>"110000111",
  5166=>"010011001",
  5167=>"100101001",
  5168=>"010111000",
  5169=>"101100100",
  5170=>"000001100",
  5171=>"001001001",
  5172=>"011011001",
  5173=>"010011110",
  5174=>"001110101",
  5175=>"111011100",
  5176=>"000000001",
  5177=>"011001101",
  5178=>"001100111",
  5179=>"011000100",
  5180=>"110110101",
  5181=>"001001010",
  5182=>"101111101",
  5183=>"110110010",
  5184=>"110000001",
  5185=>"111000001",
  5186=>"110111111",
  5187=>"110110010",
  5188=>"111110101",
  5189=>"011010000",
  5190=>"100101111",
  5191=>"100000100",
  5192=>"010101100",
  5193=>"000101000",
  5194=>"000111011",
  5195=>"010011010",
  5196=>"000010101",
  5197=>"010100001",
  5198=>"110110100",
  5199=>"101110110",
  5200=>"111111100",
  5201=>"100001001",
  5202=>"011010101",
  5203=>"101110110",
  5204=>"010001110",
  5205=>"110010001",
  5206=>"010011001",
  5207=>"000101100",
  5208=>"100111001",
  5209=>"000010111",
  5210=>"011101010",
  5211=>"101100110",
  5212=>"100101110",
  5213=>"111101000",
  5214=>"001100001",
  5215=>"000010111",
  5216=>"010010001",
  5217=>"011010011",
  5218=>"001101001",
  5219=>"111101110",
  5220=>"010111101",
  5221=>"111011010",
  5222=>"110101001",
  5223=>"110110010",
  5224=>"000101000",
  5225=>"111011000",
  5226=>"010000011",
  5227=>"001101101",
  5228=>"110100111",
  5229=>"011100110",
  5230=>"100110001",
  5231=>"000000011",
  5232=>"000111100",
  5233=>"100100111",
  5234=>"000110001",
  5235=>"110101001",
  5236=>"110011101",
  5237=>"111101110",
  5238=>"101101001",
  5239=>"101101110",
  5240=>"001011111",
  5241=>"101101110",
  5242=>"001010101",
  5243=>"001011111",
  5244=>"101111010",
  5245=>"111011001",
  5246=>"101011010",
  5247=>"010110100",
  5248=>"000001011",
  5249=>"011101011",
  5250=>"011000111",
  5251=>"101010111",
  5252=>"010001100",
  5253=>"101011101",
  5254=>"001100111",
  5255=>"001111111",
  5256=>"111100111",
  5257=>"101000001",
  5258=>"101001101",
  5259=>"110011100",
  5260=>"010111101",
  5261=>"001010101",
  5262=>"101011110",
  5263=>"010110111",
  5264=>"001110110",
  5265=>"010100111",
  5266=>"001010101",
  5267=>"001010010",
  5268=>"001101101",
  5269=>"010010100",
  5270=>"001001100",
  5271=>"001010001",
  5272=>"111100110",
  5273=>"000001101",
  5274=>"101100001",
  5275=>"101011100",
  5276=>"001110000",
  5277=>"111001100",
  5278=>"111001011",
  5279=>"000001110",
  5280=>"100010010",
  5281=>"000010101",
  5282=>"100110111",
  5283=>"111011100",
  5284=>"000011110",
  5285=>"111000001",
  5286=>"111010010",
  5287=>"100011110",
  5288=>"011101010",
  5289=>"100010101",
  5290=>"000001000",
  5291=>"100001111",
  5292=>"100111010",
  5293=>"011100110",
  5294=>"001100000",
  5295=>"100110010",
  5296=>"110011011",
  5297=>"010110110",
  5298=>"101001011",
  5299=>"110010000",
  5300=>"100000000",
  5301=>"010001000",
  5302=>"011111011",
  5303=>"001001000",
  5304=>"110101000",
  5305=>"001001000",
  5306=>"100000010",
  5307=>"001011001",
  5308=>"010010001",
  5309=>"101011011",
  5310=>"001101001",
  5311=>"110110000",
  5312=>"110001000",
  5313=>"110000011",
  5314=>"010100001",
  5315=>"000011101",
  5316=>"010011001",
  5317=>"111010111",
  5318=>"111011100",
  5319=>"001010010",
  5320=>"101110101",
  5321=>"111000010",
  5322=>"010001001",
  5323=>"100111100",
  5324=>"111100010",
  5325=>"100101100",
  5326=>"110001000",
  5327=>"101010011",
  5328=>"011101001",
  5329=>"000010101",
  5330=>"101100011",
  5331=>"111101000",
  5332=>"110010100",
  5333=>"111100001",
  5334=>"010010001",
  5335=>"111100001",
  5336=>"000101101",
  5337=>"110000111",
  5338=>"110010010",
  5339=>"001001001",
  5340=>"010000010",
  5341=>"111000011",
  5342=>"111100111",
  5343=>"111010111",
  5344=>"101011110",
  5345=>"001011000",
  5346=>"010100000",
  5347=>"110110110",
  5348=>"111101110",
  5349=>"000110110",
  5350=>"101111010",
  5351=>"110011100",
  5352=>"101010110",
  5353=>"011101101",
  5354=>"000001110",
  5355=>"101100000",
  5356=>"001101000",
  5357=>"010101010",
  5358=>"001111101",
  5359=>"110100100",
  5360=>"111111011",
  5361=>"010011000",
  5362=>"011100101",
  5363=>"101111011",
  5364=>"110101011",
  5365=>"001001010",
  5366=>"111111100",
  5367=>"000001001",
  5368=>"100001011",
  5369=>"011100010",
  5370=>"110101101",
  5371=>"001000111",
  5372=>"101001110",
  5373=>"001001010",
  5374=>"100110001",
  5375=>"010001100",
  5376=>"100100100",
  5377=>"111100011",
  5378=>"001111001",
  5379=>"110110111",
  5380=>"111000010",
  5381=>"010010110",
  5382=>"110100111",
  5383=>"010100010",
  5384=>"001101100",
  5385=>"100001011",
  5386=>"011000111",
  5387=>"101111100",
  5388=>"010010000",
  5389=>"100110000",
  5390=>"010000000",
  5391=>"000010100",
  5392=>"100011001",
  5393=>"101010011",
  5394=>"100001111",
  5395=>"101001101",
  5396=>"011110011",
  5397=>"110111111",
  5398=>"000001101",
  5399=>"010000011",
  5400=>"100000100",
  5401=>"000010110",
  5402=>"011011011",
  5403=>"011001011",
  5404=>"100011011",
  5405=>"111110111",
  5406=>"000110010",
  5407=>"000000110",
  5408=>"010111011",
  5409=>"001101010",
  5410=>"000101110",
  5411=>"001001100",
  5412=>"111011111",
  5413=>"011101010",
  5414=>"101110000",
  5415=>"011000101",
  5416=>"111001101",
  5417=>"100001010",
  5418=>"011110111",
  5419=>"111000001",
  5420=>"101101001",
  5421=>"001110100",
  5422=>"000101111",
  5423=>"100100000",
  5424=>"001010011",
  5425=>"101100111",
  5426=>"100001111",
  5427=>"000001010",
  5428=>"011101011",
  5429=>"010001110",
  5430=>"001001010",
  5431=>"101000101",
  5432=>"001011001",
  5433=>"011010110",
  5434=>"110100011",
  5435=>"011110110",
  5436=>"001000100",
  5437=>"100010111",
  5438=>"000110111",
  5439=>"101111111",
  5440=>"000010100",
  5441=>"110111010",
  5442=>"010000001",
  5443=>"110110100",
  5444=>"010010111",
  5445=>"111000001",
  5446=>"111000101",
  5447=>"000011101",
  5448=>"110001010",
  5449=>"111000111",
  5450=>"000000011",
  5451=>"000101011",
  5452=>"000011100",
  5453=>"111100101",
  5454=>"000111100",
  5455=>"101010011",
  5456=>"111101101",
  5457=>"110111010",
  5458=>"111010011",
  5459=>"000111111",
  5460=>"001001010",
  5461=>"110011110",
  5462=>"100001111",
  5463=>"010011001",
  5464=>"000100010",
  5465=>"100100110",
  5466=>"000001011",
  5467=>"101100011",
  5468=>"010110100",
  5469=>"111100101",
  5470=>"010010001",
  5471=>"000110000",
  5472=>"110000001",
  5473=>"000110001",
  5474=>"100000100",
  5475=>"011000101",
  5476=>"001000001",
  5477=>"100110111",
  5478=>"010001111",
  5479=>"000111111",
  5480=>"100100110",
  5481=>"001011101",
  5482=>"000000100",
  5483=>"110110001",
  5484=>"111010100",
  5485=>"110000101",
  5486=>"111100010",
  5487=>"110001000",
  5488=>"000011110",
  5489=>"100000001",
  5490=>"101010001",
  5491=>"101101110",
  5492=>"001100000",
  5493=>"010001100",
  5494=>"100000111",
  5495=>"000011011",
  5496=>"000111010",
  5497=>"110001111",
  5498=>"000101011",
  5499=>"110101111",
  5500=>"000100011",
  5501=>"000111011",
  5502=>"010010011",
  5503=>"000111111",
  5504=>"101111111",
  5505=>"001101011",
  5506=>"110101000",
  5507=>"011010100",
  5508=>"101011000",
  5509=>"111101101",
  5510=>"001010010",
  5511=>"100010100",
  5512=>"101000100",
  5513=>"111010001",
  5514=>"110101001",
  5515=>"101001100",
  5516=>"001110011",
  5517=>"100011100",
  5518=>"011001000",
  5519=>"000011110",
  5520=>"110100011",
  5521=>"100111001",
  5522=>"000100001",
  5523=>"100000001",
  5524=>"101111111",
  5525=>"001001010",
  5526=>"110011111",
  5527=>"101111001",
  5528=>"001110110",
  5529=>"000010101",
  5530=>"101011111",
  5531=>"100100001",
  5532=>"100011011",
  5533=>"011011111",
  5534=>"111011000",
  5535=>"010010110",
  5536=>"101000100",
  5537=>"100110001",
  5538=>"010000101",
  5539=>"111100111",
  5540=>"001001000",
  5541=>"111000110",
  5542=>"110110111",
  5543=>"100001110",
  5544=>"101010100",
  5545=>"001001110",
  5546=>"000100001",
  5547=>"001011011",
  5548=>"111110100",
  5549=>"011110110",
  5550=>"001000100",
  5551=>"110010001",
  5552=>"000001101",
  5553=>"001101010",
  5554=>"101000000",
  5555=>"011001000",
  5556=>"111001100",
  5557=>"111110010",
  5558=>"111101011",
  5559=>"011111011",
  5560=>"110001001",
  5561=>"001100111",
  5562=>"001010101",
  5563=>"001001000",
  5564=>"110111000",
  5565=>"100001000",
  5566=>"001011011",
  5567=>"111000101",
  5568=>"100010001",
  5569=>"010111100",
  5570=>"111011010",
  5571=>"110000000",
  5572=>"101000100",
  5573=>"011000000",
  5574=>"111110011",
  5575=>"101100100",
  5576=>"000111001",
  5577=>"111010110",
  5578=>"011100000",
  5579=>"111000010",
  5580=>"110101011",
  5581=>"111110110",
  5582=>"100010010",
  5583=>"101101010",
  5584=>"001110010",
  5585=>"110000011",
  5586=>"101010100",
  5587=>"100110100",
  5588=>"010001010",
  5589=>"001011010",
  5590=>"011110100",
  5591=>"000000001",
  5592=>"011001011",
  5593=>"011000110",
  5594=>"000000010",
  5595=>"001100100",
  5596=>"101101001",
  5597=>"110111011",
  5598=>"111001100",
  5599=>"011110101",
  5600=>"111010110",
  5601=>"010001110",
  5602=>"110110011",
  5603=>"010000111",
  5604=>"110110011",
  5605=>"010011001",
  5606=>"111101100",
  5607=>"001100000",
  5608=>"000001010",
  5609=>"001010000",
  5610=>"111101010",
  5611=>"000011011",
  5612=>"110000011",
  5613=>"111011101",
  5614=>"101101100",
  5615=>"101001010",
  5616=>"111010011",
  5617=>"100010000",
  5618=>"100011001",
  5619=>"111010101",
  5620=>"001000011",
  5621=>"010100000",
  5622=>"000101001",
  5623=>"101100100",
  5624=>"101101110",
  5625=>"011001001",
  5626=>"111110110",
  5627=>"001000010",
  5628=>"100010111",
  5629=>"000110111",
  5630=>"101011101",
  5631=>"101010000",
  5632=>"110011111",
  5633=>"110101011",
  5634=>"001101001",
  5635=>"001001100",
  5636=>"000111000",
  5637=>"011100000",
  5638=>"011110110",
  5639=>"001111010",
  5640=>"110001110",
  5641=>"111011110",
  5642=>"111110011",
  5643=>"100011101",
  5644=>"110110011",
  5645=>"100100100",
  5646=>"111111011",
  5647=>"101001011",
  5648=>"011010111",
  5649=>"111011100",
  5650=>"100101101",
  5651=>"100000110",
  5652=>"001100101",
  5653=>"010101100",
  5654=>"010101100",
  5655=>"000101010",
  5656=>"101100111",
  5657=>"001110101",
  5658=>"110000000",
  5659=>"010011001",
  5660=>"101110110",
  5661=>"010100100",
  5662=>"111011010",
  5663=>"001000110",
  5664=>"100100000",
  5665=>"011010111",
  5666=>"001100011",
  5667=>"000000001",
  5668=>"101100010",
  5669=>"111001011",
  5670=>"010101101",
  5671=>"111111000",
  5672=>"111101011",
  5673=>"010000110",
  5674=>"001100111",
  5675=>"110111101",
  5676=>"011000001",
  5677=>"000101001",
  5678=>"000010010",
  5679=>"000010110",
  5680=>"011111010",
  5681=>"100110100",
  5682=>"011000100",
  5683=>"011110110",
  5684=>"110100011",
  5685=>"100101111",
  5686=>"100101010",
  5687=>"101000000",
  5688=>"101000010",
  5689=>"011000011",
  5690=>"001101011",
  5691=>"110111111",
  5692=>"000110101",
  5693=>"010100111",
  5694=>"000010001",
  5695=>"001111101",
  5696=>"100100000",
  5697=>"111101011",
  5698=>"000100110",
  5699=>"010011000",
  5700=>"010100001",
  5701=>"000100101",
  5702=>"011001100",
  5703=>"011001111",
  5704=>"111011110",
  5705=>"001000101",
  5706=>"110001100",
  5707=>"000000110",
  5708=>"100110001",
  5709=>"000000000",
  5710=>"001000100",
  5711=>"010111111",
  5712=>"011100000",
  5713=>"000000011",
  5714=>"100011000",
  5715=>"100111011",
  5716=>"011010011",
  5717=>"000011011",
  5718=>"110000000",
  5719=>"000110100",
  5720=>"111111000",
  5721=>"010100111",
  5722=>"001000101",
  5723=>"110101000",
  5724=>"010101100",
  5725=>"110100101",
  5726=>"101101110",
  5727=>"001110110",
  5728=>"111111101",
  5729=>"001110110",
  5730=>"100110111",
  5731=>"101000111",
  5732=>"000100100",
  5733=>"101011011",
  5734=>"100001101",
  5735=>"000000001",
  5736=>"100100001",
  5737=>"000111011",
  5738=>"010000001",
  5739=>"110100100",
  5740=>"101111110",
  5741=>"110000010",
  5742=>"100010100",
  5743=>"001100001",
  5744=>"101011101",
  5745=>"110000110",
  5746=>"111011101",
  5747=>"101101111",
  5748=>"000101101",
  5749=>"111110110",
  5750=>"001000111",
  5751=>"100110101",
  5752=>"001001000",
  5753=>"010001001",
  5754=>"011100101",
  5755=>"000100010",
  5756=>"010101111",
  5757=>"010000010",
  5758=>"111011010",
  5759=>"100000011",
  5760=>"010000110",
  5761=>"110000110",
  5762=>"101110110",
  5763=>"100001111",
  5764=>"100010000",
  5765=>"010000000",
  5766=>"101100000",
  5767=>"001010100",
  5768=>"110011000",
  5769=>"111000010",
  5770=>"101001111",
  5771=>"000011001",
  5772=>"011001111",
  5773=>"111001100",
  5774=>"101001000",
  5775=>"001100101",
  5776=>"001000100",
  5777=>"001001101",
  5778=>"110010111",
  5779=>"010000101",
  5780=>"010100001",
  5781=>"011001001",
  5782=>"110000111",
  5783=>"101000111",
  5784=>"100111011",
  5785=>"011111011",
  5786=>"000100011",
  5787=>"101001010",
  5788=>"110010011",
  5789=>"110111111",
  5790=>"010100010",
  5791=>"110111111",
  5792=>"111010110",
  5793=>"001001000",
  5794=>"101011000",
  5795=>"010000111",
  5796=>"000010011",
  5797=>"100001011",
  5798=>"101001010",
  5799=>"001010010",
  5800=>"110110110",
  5801=>"110010011",
  5802=>"100101100",
  5803=>"111001010",
  5804=>"010000101",
  5805=>"011111100",
  5806=>"101110101",
  5807=>"011110011",
  5808=>"000100101",
  5809=>"101111111",
  5810=>"010001101",
  5811=>"100101000",
  5812=>"011101001",
  5813=>"000001001",
  5814=>"000100010",
  5815=>"011110011",
  5816=>"011101010",
  5817=>"111111111",
  5818=>"011000010",
  5819=>"100000001",
  5820=>"000001011",
  5821=>"010110100",
  5822=>"111100011",
  5823=>"110010000",
  5824=>"010110111",
  5825=>"100111110",
  5826=>"011110110",
  5827=>"000100011",
  5828=>"010000000",
  5829=>"010100011",
  5830=>"111111001",
  5831=>"001000110",
  5832=>"111110100",
  5833=>"010100011",
  5834=>"000011111",
  5835=>"110001101",
  5836=>"011101011",
  5837=>"001000111",
  5838=>"001101101",
  5839=>"000100101",
  5840=>"001011010",
  5841=>"011101111",
  5842=>"010100011",
  5843=>"101010001",
  5844=>"100000100",
  5845=>"010001010",
  5846=>"000011010",
  5847=>"010010011",
  5848=>"100010010",
  5849=>"010000010",
  5850=>"111000101",
  5851=>"011011110",
  5852=>"111111101",
  5853=>"011000100",
  5854=>"000100011",
  5855=>"011111111",
  5856=>"000001110",
  5857=>"101101001",
  5858=>"010010111",
  5859=>"010101101",
  5860=>"010001011",
  5861=>"000010010",
  5862=>"111001111",
  5863=>"101001111",
  5864=>"101101100",
  5865=>"110100011",
  5866=>"101101010",
  5867=>"001011000",
  5868=>"111000101",
  5869=>"011101001",
  5870=>"000011011",
  5871=>"111011000",
  5872=>"101010101",
  5873=>"111000110",
  5874=>"111001001",
  5875=>"110011110",
  5876=>"011111001",
  5877=>"100111100",
  5878=>"101101100",
  5879=>"001000000",
  5880=>"111011111",
  5881=>"111111101",
  5882=>"100111111",
  5883=>"000010110",
  5884=>"111001100",
  5885=>"111101000",
  5886=>"101001000",
  5887=>"100111101",
  5888=>"100011110",
  5889=>"110001111",
  5890=>"001000000",
  5891=>"000110010",
  5892=>"010011110",
  5893=>"001110111",
  5894=>"001001101",
  5895=>"001100110",
  5896=>"010111110",
  5897=>"110100101",
  5898=>"001000101",
  5899=>"011010000",
  5900=>"110011000",
  5901=>"110001000",
  5902=>"000100001",
  5903=>"110110110",
  5904=>"101100010",
  5905=>"110000000",
  5906=>"111100010",
  5907=>"011001001",
  5908=>"100100000",
  5909=>"110101101",
  5910=>"001000010",
  5911=>"011101001",
  5912=>"000001101",
  5913=>"111011000",
  5914=>"001110101",
  5915=>"101010111",
  5916=>"110101101",
  5917=>"000111011",
  5918=>"101110000",
  5919=>"100000001",
  5920=>"010100010",
  5921=>"010010000",
  5922=>"011101001",
  5923=>"011010010",
  5924=>"010010011",
  5925=>"001010101",
  5926=>"111001111",
  5927=>"000100101",
  5928=>"010101000",
  5929=>"111001011",
  5930=>"110010100",
  5931=>"100110000",
  5932=>"011010010",
  5933=>"110110010",
  5934=>"101001000",
  5935=>"001000111",
  5936=>"001100111",
  5937=>"101011100",
  5938=>"100000111",
  5939=>"011011101",
  5940=>"011011100",
  5941=>"110111110",
  5942=>"010010000",
  5943=>"001000010",
  5944=>"100010111",
  5945=>"010101101",
  5946=>"010010101",
  5947=>"110001001",
  5948=>"111011001",
  5949=>"011011101",
  5950=>"111101011",
  5951=>"100010111",
  5952=>"111001001",
  5953=>"111010001",
  5954=>"101111000",
  5955=>"011001101",
  5956=>"000000101",
  5957=>"011000000",
  5958=>"000010110",
  5959=>"101010100",
  5960=>"101000001",
  5961=>"010000101",
  5962=>"101110100",
  5963=>"000010100",
  5964=>"011111111",
  5965=>"001000110",
  5966=>"100001010",
  5967=>"001110000",
  5968=>"000100111",
  5969=>"110001110",
  5970=>"010001010",
  5971=>"011001101",
  5972=>"010011011",
  5973=>"000011000",
  5974=>"001000111",
  5975=>"101001000",
  5976=>"010111000",
  5977=>"110011001",
  5978=>"011001010",
  5979=>"101011011",
  5980=>"101001000",
  5981=>"100110001",
  5982=>"001111110",
  5983=>"001010011",
  5984=>"100001101",
  5985=>"111001001",
  5986=>"001111101",
  5987=>"100111100",
  5988=>"111011001",
  5989=>"010110000",
  5990=>"011101010",
  5991=>"011100111",
  5992=>"010011011",
  5993=>"101110011",
  5994=>"101100011",
  5995=>"110100111",
  5996=>"111000001",
  5997=>"101111010",
  5998=>"110011100",
  5999=>"100111000",
  6000=>"100110000",
  6001=>"011111110",
  6002=>"111111100",
  6003=>"110001000",
  6004=>"111110001",
  6005=>"011111011",
  6006=>"110011110",
  6007=>"010111111",
  6008=>"001001100",
  6009=>"000101011",
  6010=>"100010101",
  6011=>"100000011",
  6012=>"000000000",
  6013=>"001111100",
  6014=>"010111010",
  6015=>"101111101",
  6016=>"110010010",
  6017=>"110110111",
  6018=>"011000001",
  6019=>"011010000",
  6020=>"001000101",
  6021=>"111100011",
  6022=>"110010010",
  6023=>"100101001",
  6024=>"101101011",
  6025=>"110110010",
  6026=>"000011111",
  6027=>"101001111",
  6028=>"111101000",
  6029=>"100110000",
  6030=>"111001001",
  6031=>"011110000",
  6032=>"010101001",
  6033=>"000110001",
  6034=>"101111011",
  6035=>"111110001",
  6036=>"100011101",
  6037=>"000111000",
  6038=>"011011010",
  6039=>"010110001",
  6040=>"111100011",
  6041=>"100001011",
  6042=>"000101001",
  6043=>"000100111",
  6044=>"010010001",
  6045=>"001101110",
  6046=>"000101011",
  6047=>"101010000",
  6048=>"100000000",
  6049=>"110101000",
  6050=>"101100000",
  6051=>"010001010",
  6052=>"110000101",
  6053=>"001010001",
  6054=>"111110100",
  6055=>"010011100",
  6056=>"110001010",
  6057=>"011000100",
  6058=>"101011011",
  6059=>"101100011",
  6060=>"110100111",
  6061=>"000110101",
  6062=>"001100101",
  6063=>"100011110",
  6064=>"011110100",
  6065=>"000110001",
  6066=>"111011011",
  6067=>"001000000",
  6068=>"101000011",
  6069=>"100011001",
  6070=>"100111010",
  6071=>"111101111",
  6072=>"100001001",
  6073=>"101010101",
  6074=>"010110100",
  6075=>"000100010",
  6076=>"001110101",
  6077=>"001010001",
  6078=>"100011001",
  6079=>"100110110",
  6080=>"000100111",
  6081=>"001001001",
  6082=>"110001011",
  6083=>"110110110",
  6084=>"110110010",
  6085=>"001001111",
  6086=>"011110000",
  6087=>"011110010",
  6088=>"110000010",
  6089=>"100011110",
  6090=>"110000101",
  6091=>"010100111",
  6092=>"000110101",
  6093=>"011001010",
  6094=>"111001010",
  6095=>"001101101",
  6096=>"111101100",
  6097=>"000001111",
  6098=>"110001000",
  6099=>"000110100",
  6100=>"100101110",
  6101=>"111011110",
  6102=>"000000100",
  6103=>"111011100",
  6104=>"000011111",
  6105=>"111111101",
  6106=>"011011110",
  6107=>"101001011",
  6108=>"111100000",
  6109=>"110001000",
  6110=>"111011110",
  6111=>"111011111",
  6112=>"101100000",
  6113=>"110100010",
  6114=>"001111101",
  6115=>"110110100",
  6116=>"111000011",
  6117=>"000100000",
  6118=>"011011000",
  6119=>"111000011",
  6120=>"100110111",
  6121=>"001111110",
  6122=>"000000001",
  6123=>"010110001",
  6124=>"111001010",
  6125=>"100111001",
  6126=>"000110001",
  6127=>"111111101",
  6128=>"101000111",
  6129=>"000000001",
  6130=>"100111101",
  6131=>"001010100",
  6132=>"010110010",
  6133=>"001000110",
  6134=>"000111111",
  6135=>"111010010",
  6136=>"010101011",
  6137=>"101110111",
  6138=>"101000010",
  6139=>"111101001",
  6140=>"100010010",
  6141=>"111001110",
  6142=>"011001111",
  6143=>"001010110",
  6144=>"011000100",
  6145=>"111111111",
  6146=>"011001101",
  6147=>"010111001",
  6148=>"101011011",
  6149=>"111010010",
  6150=>"111100010",
  6151=>"001011011",
  6152=>"110010100",
  6153=>"100001110",
  6154=>"011011000",
  6155=>"100110001",
  6156=>"001001000",
  6157=>"001000110",
  6158=>"100111010",
  6159=>"010111001",
  6160=>"011111100",
  6161=>"111001101",
  6162=>"101000100",
  6163=>"110001011",
  6164=>"001001000",
  6165=>"010011001",
  6166=>"110111111",
  6167=>"010011111",
  6168=>"001101001",
  6169=>"110000101",
  6170=>"011000001",
  6171=>"011101100",
  6172=>"001110000",
  6173=>"011000101",
  6174=>"111011000",
  6175=>"001001100",
  6176=>"011001100",
  6177=>"010000101",
  6178=>"000101111",
  6179=>"000101001",
  6180=>"000010111",
  6181=>"101110110",
  6182=>"101001110",
  6183=>"000010001",
  6184=>"110011000",
  6185=>"000100110",
  6186=>"101110101",
  6187=>"011100001",
  6188=>"100010000",
  6189=>"000011011",
  6190=>"011111111",
  6191=>"010001001",
  6192=>"000111101",
  6193=>"100011000",
  6194=>"101000111",
  6195=>"110011101",
  6196=>"000101100",
  6197=>"001100110",
  6198=>"001100100",
  6199=>"101000110",
  6200=>"011101100",
  6201=>"111010100",
  6202=>"000100110",
  6203=>"111000111",
  6204=>"101100100",
  6205=>"001110010",
  6206=>"100000101",
  6207=>"110011100",
  6208=>"011011101",
  6209=>"010111110",
  6210=>"101010111",
  6211=>"111111000",
  6212=>"001101010",
  6213=>"000000110",
  6214=>"001111101",
  6215=>"111110110",
  6216=>"110111111",
  6217=>"000011011",
  6218=>"100111111",
  6219=>"011101110",
  6220=>"010010011",
  6221=>"000111111",
  6222=>"111000010",
  6223=>"110011101",
  6224=>"111011111",
  6225=>"111111011",
  6226=>"110010010",
  6227=>"010001110",
  6228=>"100111010",
  6229=>"111111111",
  6230=>"110100000",
  6231=>"101010001",
  6232=>"010001000",
  6233=>"101001101",
  6234=>"100110100",
  6235=>"011111011",
  6236=>"101010001",
  6237=>"011011001",
  6238=>"101010010",
  6239=>"111101111",
  6240=>"001001110",
  6241=>"111100111",
  6242=>"111111101",
  6243=>"011101100",
  6244=>"101110001",
  6245=>"100001000",
  6246=>"111111101",
  6247=>"000100111",
  6248=>"100000001",
  6249=>"010111010",
  6250=>"111100110",
  6251=>"100111011",
  6252=>"100111101",
  6253=>"110111000",
  6254=>"000000011",
  6255=>"101101111",
  6256=>"011100001",
  6257=>"010010101",
  6258=>"100101111",
  6259=>"111000000",
  6260=>"111111011",
  6261=>"000110000",
  6262=>"001110010",
  6263=>"110111100",
  6264=>"011001111",
  6265=>"100000100",
  6266=>"010101000",
  6267=>"011100000",
  6268=>"000001001",
  6269=>"000101111",
  6270=>"001000100",
  6271=>"011100000",
  6272=>"101101100",
  6273=>"010010111",
  6274=>"000100000",
  6275=>"100001011",
  6276=>"011001000",
  6277=>"111100101",
  6278=>"011110011",
  6279=>"000110110",
  6280=>"100010001",
  6281=>"101001010",
  6282=>"010111011",
  6283=>"101111001",
  6284=>"101010000",
  6285=>"100010000",
  6286=>"011101111",
  6287=>"001000010",
  6288=>"100101111",
  6289=>"111111111",
  6290=>"001001000",
  6291=>"110100011",
  6292=>"000101011",
  6293=>"011000111",
  6294=>"101011111",
  6295=>"001101110",
  6296=>"101101000",
  6297=>"100100110",
  6298=>"100001111",
  6299=>"111101111",
  6300=>"010100101",
  6301=>"010100100",
  6302=>"101010100",
  6303=>"011001000",
  6304=>"111000011",
  6305=>"110100101",
  6306=>"000000010",
  6307=>"010110000",
  6308=>"100101011",
  6309=>"111111100",
  6310=>"111111110",
  6311=>"010111001",
  6312=>"111110000",
  6313=>"111100000",
  6314=>"111000001",
  6315=>"000001111",
  6316=>"000111010",
  6317=>"001000101",
  6318=>"111101100",
  6319=>"101010001",
  6320=>"001111010",
  6321=>"111000100",
  6322=>"100111110",
  6323=>"100100111",
  6324=>"101010111",
  6325=>"011011111",
  6326=>"101101110",
  6327=>"000010000",
  6328=>"000001001",
  6329=>"010110000",
  6330=>"000011100",
  6331=>"001111111",
  6332=>"010010010",
  6333=>"011111001",
  6334=>"111000111",
  6335=>"101010010",
  6336=>"110101011",
  6337=>"111011111",
  6338=>"001111100",
  6339=>"000001000",
  6340=>"010100101",
  6341=>"100101011",
  6342=>"111111111",
  6343=>"010100100",
  6344=>"101110011",
  6345=>"110010001",
  6346=>"010000110",
  6347=>"011110110",
  6348=>"101110100",
  6349=>"100100010",
  6350=>"110011010",
  6351=>"000000010",
  6352=>"011110000",
  6353=>"100011100",
  6354=>"001011101",
  6355=>"101010011",
  6356=>"001100100",
  6357=>"110101110",
  6358=>"101101001",
  6359=>"111011001",
  6360=>"100011110",
  6361=>"001100011",
  6362=>"000010100",
  6363=>"111001110",
  6364=>"100111001",
  6365=>"011000010",
  6366=>"000010001",
  6367=>"010110111",
  6368=>"000010010",
  6369=>"010000110",
  6370=>"001101000",
  6371=>"110100010",
  6372=>"011111101",
  6373=>"001100001",
  6374=>"011010001",
  6375=>"110111001",
  6376=>"011111100",
  6377=>"111000111",
  6378=>"000011000",
  6379=>"011110111",
  6380=>"011100011",
  6381=>"110110110",
  6382=>"000000000",
  6383=>"000001100",
  6384=>"011100011",
  6385=>"111101010",
  6386=>"000011110",
  6387=>"010011100",
  6388=>"100111111",
  6389=>"000110000",
  6390=>"111111100",
  6391=>"100011011",
  6392=>"010001111",
  6393=>"010100010",
  6394=>"100100000",
  6395=>"110111100",
  6396=>"111100000",
  6397=>"010010101",
  6398=>"110001001",
  6399=>"111111001",
  6400=>"110110001",
  6401=>"111111110",
  6402=>"100110010",
  6403=>"001000110",
  6404=>"100111010",
  6405=>"111101011",
  6406=>"111111110",
  6407=>"111101001",
  6408=>"100011100",
  6409=>"110101001",
  6410=>"010010110",
  6411=>"011010100",
  6412=>"111010001",
  6413=>"101101010",
  6414=>"011011000",
  6415=>"100110111",
  6416=>"101010011",
  6417=>"100011001",
  6418=>"101011011",
  6419=>"010000010",
  6420=>"001000010",
  6421=>"110111010",
  6422=>"110001110",
  6423=>"111100001",
  6424=>"110110101",
  6425=>"011100111",
  6426=>"111100010",
  6427=>"101111010",
  6428=>"011010111",
  6429=>"111100001",
  6430=>"010100101",
  6431=>"101000100",
  6432=>"101000110",
  6433=>"000100101",
  6434=>"100010000",
  6435=>"000000000",
  6436=>"010011101",
  6437=>"000010000",
  6438=>"001110000",
  6439=>"101000110",
  6440=>"010010110",
  6441=>"101101001",
  6442=>"111101110",
  6443=>"001010101",
  6444=>"101001110",
  6445=>"101010010",
  6446=>"011011111",
  6447=>"000000001",
  6448=>"110000111",
  6449=>"110110101",
  6450=>"010101000",
  6451=>"000100111",
  6452=>"101110110",
  6453=>"010010110",
  6454=>"111100010",
  6455=>"011011100",
  6456=>"110011011",
  6457=>"010110000",
  6458=>"100001110",
  6459=>"110100100",
  6460=>"010000011",
  6461=>"101011010",
  6462=>"010111100",
  6463=>"111000111",
  6464=>"000101000",
  6465=>"001111001",
  6466=>"101000101",
  6467=>"001111011",
  6468=>"100101100",
  6469=>"000101001",
  6470=>"000001100",
  6471=>"000010110",
  6472=>"000011111",
  6473=>"000000101",
  6474=>"101110001",
  6475=>"110111011",
  6476=>"100111000",
  6477=>"110010011",
  6478=>"011001100",
  6479=>"101010110",
  6480=>"110110111",
  6481=>"010001010",
  6482=>"111111110",
  6483=>"101111001",
  6484=>"000100001",
  6485=>"001011111",
  6486=>"101000000",
  6487=>"100110011",
  6488=>"111010100",
  6489=>"111110001",
  6490=>"001110001",
  6491=>"101000000",
  6492=>"101100110",
  6493=>"110101111",
  6494=>"011100010",
  6495=>"111101101",
  6496=>"111000010",
  6497=>"111001100",
  6498=>"001011110",
  6499=>"100101100",
  6500=>"011101000",
  6501=>"000010110",
  6502=>"111110010",
  6503=>"110101100",
  6504=>"101100100",
  6505=>"001011111",
  6506=>"010111010",
  6507=>"011110100",
  6508=>"101100111",
  6509=>"111000011",
  6510=>"000011001",
  6511=>"010110001",
  6512=>"000010110",
  6513=>"010010101",
  6514=>"100111110",
  6515=>"001111001",
  6516=>"010000100",
  6517=>"100010100",
  6518=>"101001111",
  6519=>"111011001",
  6520=>"100110111",
  6521=>"000100111",
  6522=>"000001111",
  6523=>"100010000",
  6524=>"001000100",
  6525=>"011110110",
  6526=>"011000001",
  6527=>"111111000",
  6528=>"010010100",
  6529=>"010001000",
  6530=>"110001101",
  6531=>"011001000",
  6532=>"001000101",
  6533=>"011100111",
  6534=>"101000010",
  6535=>"101001111",
  6536=>"100010000",
  6537=>"101001011",
  6538=>"110010110",
  6539=>"111001001",
  6540=>"001110100",
  6541=>"100100001",
  6542=>"010000000",
  6543=>"011111111",
  6544=>"100111011",
  6545=>"110001110",
  6546=>"111010110",
  6547=>"101110111",
  6548=>"111111111",
  6549=>"100000110",
  6550=>"001001010",
  6551=>"110010001",
  6552=>"101110011",
  6553=>"000001011",
  6554=>"100000111",
  6555=>"000010100",
  6556=>"010111101",
  6557=>"001101000",
  6558=>"010000000",
  6559=>"011010010",
  6560=>"101110001",
  6561=>"101011010",
  6562=>"101101111",
  6563=>"000111110",
  6564=>"110011110",
  6565=>"010110101",
  6566=>"000000000",
  6567=>"000001000",
  6568=>"111001010",
  6569=>"111011111",
  6570=>"000111111",
  6571=>"000100000",
  6572=>"010010100",
  6573=>"000001100",
  6574=>"010101001",
  6575=>"010010000",
  6576=>"100010001",
  6577=>"011111110",
  6578=>"011000100",
  6579=>"001001100",
  6580=>"111110110",
  6581=>"000000110",
  6582=>"000001100",
  6583=>"111110010",
  6584=>"101110010",
  6585=>"001000111",
  6586=>"000100001",
  6587=>"110000011",
  6588=>"110001111",
  6589=>"001111111",
  6590=>"001100000",
  6591=>"110000000",
  6592=>"000001000",
  6593=>"101101001",
  6594=>"010000010",
  6595=>"010010101",
  6596=>"110100111",
  6597=>"011010010",
  6598=>"100110110",
  6599=>"110001101",
  6600=>"110011001",
  6601=>"000110011",
  6602=>"011111101",
  6603=>"010010100",
  6604=>"100011111",
  6605=>"010000011",
  6606=>"101010111",
  6607=>"111000011",
  6608=>"100110011",
  6609=>"011101011",
  6610=>"111100000",
  6611=>"011010100",
  6612=>"111010101",
  6613=>"110111000",
  6614=>"011100000",
  6615=>"101010011",
  6616=>"010100000",
  6617=>"110111001",
  6618=>"100011100",
  6619=>"000101010",
  6620=>"100101000",
  6621=>"101100100",
  6622=>"101100011",
  6623=>"010001000",
  6624=>"000010001",
  6625=>"000010110",
  6626=>"100101111",
  6627=>"111101000",
  6628=>"101010110",
  6629=>"110110111",
  6630=>"011101000",
  6631=>"001111100",
  6632=>"010000100",
  6633=>"011100111",
  6634=>"101111101",
  6635=>"001101010",
  6636=>"110111111",
  6637=>"101010011",
  6638=>"100010000",
  6639=>"110110111",
  6640=>"101101011",
  6641=>"111011010",
  6642=>"010000101",
  6643=>"110111001",
  6644=>"011000101",
  6645=>"010000101",
  6646=>"101111010",
  6647=>"101100011",
  6648=>"110111011",
  6649=>"010011001",
  6650=>"111000001",
  6651=>"011010011",
  6652=>"011110011",
  6653=>"010011100",
  6654=>"000101111",
  6655=>"110110110",
  6656=>"000100101",
  6657=>"101001100",
  6658=>"010110111",
  6659=>"101001000",
  6660=>"100010000",
  6661=>"011001111",
  6662=>"111111110",
  6663=>"111101111",
  6664=>"001001111",
  6665=>"011010011",
  6666=>"101110100",
  6667=>"110010110",
  6668=>"010000101",
  6669=>"010100100",
  6670=>"111000000",
  6671=>"011101001",
  6672=>"010111010",
  6673=>"100001000",
  6674=>"001100001",
  6675=>"001101101",
  6676=>"100001010",
  6677=>"010000101",
  6678=>"001000111",
  6679=>"111010110",
  6680=>"111101011",
  6681=>"111000000",
  6682=>"101110001",
  6683=>"010110110",
  6684=>"000001001",
  6685=>"110000100",
  6686=>"110111111",
  6687=>"000111111",
  6688=>"010001110",
  6689=>"100101011",
  6690=>"100001010",
  6691=>"011111100",
  6692=>"110011111",
  6693=>"010011000",
  6694=>"010111011",
  6695=>"001011101",
  6696=>"100100100",
  6697=>"110110110",
  6698=>"011110100",
  6699=>"000100001",
  6700=>"100110000",
  6701=>"101110101",
  6702=>"011000101",
  6703=>"000000111",
  6704=>"101111011",
  6705=>"110110100",
  6706=>"000101100",
  6707=>"001011111",
  6708=>"100011001",
  6709=>"000100011",
  6710=>"010000000",
  6711=>"011111010",
  6712=>"001011011",
  6713=>"111101111",
  6714=>"110100111",
  6715=>"000101111",
  6716=>"110110110",
  6717=>"000001100",
  6718=>"111000101",
  6719=>"010111000",
  6720=>"010000010",
  6721=>"100100101",
  6722=>"111000001",
  6723=>"001001110",
  6724=>"110101110",
  6725=>"000000110",
  6726=>"111101111",
  6727=>"101110001",
  6728=>"000001011",
  6729=>"111000110",
  6730=>"011100110",
  6731=>"100001001",
  6732=>"110101100",
  6733=>"010011011",
  6734=>"001111000",
  6735=>"100101011",
  6736=>"110101001",
  6737=>"101110100",
  6738=>"000000110",
  6739=>"111110100",
  6740=>"011100100",
  6741=>"111100110",
  6742=>"000101000",
  6743=>"101000010",
  6744=>"110110100",
  6745=>"100000001",
  6746=>"010100111",
  6747=>"000000010",
  6748=>"101101110",
  6749=>"010101110",
  6750=>"101011111",
  6751=>"101010100",
  6752=>"101111000",
  6753=>"000101110",
  6754=>"001100001",
  6755=>"000110111",
  6756=>"111101110",
  6757=>"000101001",
  6758=>"110100111",
  6759=>"011100110",
  6760=>"010101000",
  6761=>"011101101",
  6762=>"011101011",
  6763=>"111100011",
  6764=>"000100101",
  6765=>"000001010",
  6766=>"111010100",
  6767=>"111010101",
  6768=>"000010001",
  6769=>"001001010",
  6770=>"101010111",
  6771=>"110100101",
  6772=>"011100100",
  6773=>"000001001",
  6774=>"000100100",
  6775=>"011110110",
  6776=>"101100010",
  6777=>"010011100",
  6778=>"110001101",
  6779=>"000110101",
  6780=>"110011101",
  6781=>"010010010",
  6782=>"010010110",
  6783=>"001110011",
  6784=>"000000001",
  6785=>"011000000",
  6786=>"111101111",
  6787=>"100101111",
  6788=>"000100100",
  6789=>"110010110",
  6790=>"100000110",
  6791=>"011010110",
  6792=>"101101010",
  6793=>"010000110",
  6794=>"111111111",
  6795=>"000001010",
  6796=>"101011001",
  6797=>"100000110",
  6798=>"111100101",
  6799=>"100110101",
  6800=>"001100111",
  6801=>"000011011",
  6802=>"110000000",
  6803=>"110011011",
  6804=>"000010101",
  6805=>"110001110",
  6806=>"110010010",
  6807=>"001010110",
  6808=>"110100111",
  6809=>"100110101",
  6810=>"001001101",
  6811=>"001010000",
  6812=>"101011011",
  6813=>"001000111",
  6814=>"000010010",
  6815=>"101111111",
  6816=>"010000001",
  6817=>"110001010",
  6818=>"110000110",
  6819=>"101011111",
  6820=>"100000101",
  6821=>"010111011",
  6822=>"001010001",
  6823=>"000000010",
  6824=>"011000100",
  6825=>"001010001",
  6826=>"011001000",
  6827=>"110011100",
  6828=>"010001010",
  6829=>"111000001",
  6830=>"110000110",
  6831=>"110101110",
  6832=>"100010100",
  6833=>"000001110",
  6834=>"100101101",
  6835=>"101111010",
  6836=>"001110010",
  6837=>"001110110",
  6838=>"001011110",
  6839=>"010001111",
  6840=>"110011001",
  6841=>"010100001",
  6842=>"000011111",
  6843=>"110001110",
  6844=>"011010000",
  6845=>"111011101",
  6846=>"010001000",
  6847=>"011100000",
  6848=>"010100111",
  6849=>"001111011",
  6850=>"100010001",
  6851=>"111101000",
  6852=>"010100110",
  6853=>"010011010",
  6854=>"101010001",
  6855=>"101101101",
  6856=>"011000100",
  6857=>"110100011",
  6858=>"111000000",
  6859=>"001101011",
  6860=>"100111110",
  6861=>"000111010",
  6862=>"001101100",
  6863=>"011001001",
  6864=>"001101100",
  6865=>"111011111",
  6866=>"111110001",
  6867=>"000010001",
  6868=>"101000000",
  6869=>"100011011",
  6870=>"101010000",
  6871=>"000101111",
  6872=>"010000110",
  6873=>"100010000",
  6874=>"110001000",
  6875=>"000000111",
  6876=>"111100111",
  6877=>"110001100",
  6878=>"100111011",
  6879=>"111001010",
  6880=>"100001001",
  6881=>"010000110",
  6882=>"110101110",
  6883=>"100010101",
  6884=>"001011000",
  6885=>"111100101",
  6886=>"001110101",
  6887=>"010100000",
  6888=>"000001100",
  6889=>"001011111",
  6890=>"101111101",
  6891=>"011110111",
  6892=>"001110111",
  6893=>"100101100",
  6894=>"000010101",
  6895=>"011010101",
  6896=>"000101010",
  6897=>"110001100",
  6898=>"101001101",
  6899=>"100000111",
  6900=>"110110010",
  6901=>"100011000",
  6902=>"101111111",
  6903=>"000010111",
  6904=>"101011001",
  6905=>"011100000",
  6906=>"110101011",
  6907=>"000001101",
  6908=>"111000010",
  6909=>"000000100",
  6910=>"110001101",
  6911=>"000110000",
  6912=>"000111011",
  6913=>"111000011",
  6914=>"111110101",
  6915=>"110000010",
  6916=>"100111110",
  6917=>"101000010",
  6918=>"111011000",
  6919=>"000101110",
  6920=>"100000111",
  6921=>"011000000",
  6922=>"010100011",
  6923=>"110100101",
  6924=>"100010100",
  6925=>"011001011",
  6926=>"101010101",
  6927=>"111010101",
  6928=>"100101000",
  6929=>"111011100",
  6930=>"001111111",
  6931=>"001011011",
  6932=>"001011001",
  6933=>"001100101",
  6934=>"111001101",
  6935=>"101011111",
  6936=>"101001010",
  6937=>"010010110",
  6938=>"011010111",
  6939=>"111101011",
  6940=>"001111111",
  6941=>"010100010",
  6942=>"111010101",
  6943=>"000011000",
  6944=>"111010011",
  6945=>"110100101",
  6946=>"100011000",
  6947=>"000100100",
  6948=>"011111011",
  6949=>"011000111",
  6950=>"010101011",
  6951=>"111111101",
  6952=>"000010000",
  6953=>"011111000",
  6954=>"001010101",
  6955=>"100001100",
  6956=>"000010001",
  6957=>"010001000",
  6958=>"001011000",
  6959=>"101000011",
  6960=>"101001110",
  6961=>"010010001",
  6962=>"000100000",
  6963=>"111101010",
  6964=>"111001001",
  6965=>"001010011",
  6966=>"001101010",
  6967=>"000101000",
  6968=>"010110000",
  6969=>"101011001",
  6970=>"111011001",
  6971=>"110111101",
  6972=>"011110111",
  6973=>"010011011",
  6974=>"101110011",
  6975=>"110100111",
  6976=>"001111010",
  6977=>"110010000",
  6978=>"001010100",
  6979=>"100100001",
  6980=>"101111010",
  6981=>"111100001",
  6982=>"011111110",
  6983=>"000010110",
  6984=>"010101001",
  6985=>"100001010",
  6986=>"010010010",
  6987=>"111101011",
  6988=>"000101011",
  6989=>"111010010",
  6990=>"101000000",
  6991=>"100101101",
  6992=>"100101001",
  6993=>"011011011",
  6994=>"101110000",
  6995=>"100010101",
  6996=>"001011111",
  6997=>"010011011",
  6998=>"001001111",
  6999=>"101011000",
  7000=>"010000001",
  7001=>"101000011",
  7002=>"000100000",
  7003=>"011010000",
  7004=>"010011110",
  7005=>"011101111",
  7006=>"000000101",
  7007=>"010011110",
  7008=>"001001000",
  7009=>"111101011",
  7010=>"010110011",
  7011=>"100010001",
  7012=>"101101111",
  7013=>"010000100",
  7014=>"000111110",
  7015=>"000111111",
  7016=>"000000011",
  7017=>"000000000",
  7018=>"000000100",
  7019=>"010100110",
  7020=>"111000101",
  7021=>"010101011",
  7022=>"100011110",
  7023=>"101010101",
  7024=>"011011010",
  7025=>"011010001",
  7026=>"011111011",
  7027=>"111011011",
  7028=>"010010000",
  7029=>"100111000",
  7030=>"001100000",
  7031=>"000101001",
  7032=>"001010001",
  7033=>"001000000",
  7034=>"111001010",
  7035=>"010000010",
  7036=>"010101100",
  7037=>"111011111",
  7038=>"010011111",
  7039=>"011101101",
  7040=>"111111010",
  7041=>"001111011",
  7042=>"111110000",
  7043=>"101110110",
  7044=>"001100101",
  7045=>"101000110",
  7046=>"001001111",
  7047=>"000010000",
  7048=>"000111000",
  7049=>"100100011",
  7050=>"100000001",
  7051=>"111011111",
  7052=>"100110110",
  7053=>"101000001",
  7054=>"010010011",
  7055=>"111101101",
  7056=>"111011001",
  7057=>"110000111",
  7058=>"000000011",
  7059=>"001111000",
  7060=>"000111111",
  7061=>"001100010",
  7062=>"011111111",
  7063=>"001000011",
  7064=>"011010110",
  7065=>"101111111",
  7066=>"101101100",
  7067=>"011011111",
  7068=>"110100101",
  7069=>"110110100",
  7070=>"001010100",
  7071=>"010001100",
  7072=>"100110011",
  7073=>"100111101",
  7074=>"001010011",
  7075=>"001001001",
  7076=>"111111010",
  7077=>"110111011",
  7078=>"100101100",
  7079=>"001010111",
  7080=>"001100000",
  7081=>"010110001",
  7082=>"010000110",
  7083=>"111000001",
  7084=>"001100100",
  7085=>"000101100",
  7086=>"001010100",
  7087=>"001101100",
  7088=>"010010110",
  7089=>"111110101",
  7090=>"101001000",
  7091=>"000010100",
  7092=>"111010000",
  7093=>"010010011",
  7094=>"001101010",
  7095=>"000000101",
  7096=>"000000111",
  7097=>"111001010",
  7098=>"011110000",
  7099=>"111001000",
  7100=>"111011101",
  7101=>"010100101",
  7102=>"101001101",
  7103=>"100110111",
  7104=>"010000110",
  7105=>"111100111",
  7106=>"110000101",
  7107=>"101010101",
  7108=>"001110111",
  7109=>"111000101",
  7110=>"100100110",
  7111=>"011110000",
  7112=>"010101001",
  7113=>"010010010",
  7114=>"100101001",
  7115=>"101001100",
  7116=>"111000100",
  7117=>"011010011",
  7118=>"100011000",
  7119=>"011100000",
  7120=>"001101110",
  7121=>"011011101",
  7122=>"100011100",
  7123=>"100010001",
  7124=>"110100111",
  7125=>"001100000",
  7126=>"110111010",
  7127=>"101010100",
  7128=>"100101111",
  7129=>"111101111",
  7130=>"110011100",
  7131=>"011110001",
  7132=>"111111011",
  7133=>"010010111",
  7134=>"010110111",
  7135=>"110011110",
  7136=>"001101010",
  7137=>"110101101",
  7138=>"111110101",
  7139=>"101000000",
  7140=>"110010001",
  7141=>"000010100",
  7142=>"010100111",
  7143=>"110011111",
  7144=>"011110111",
  7145=>"011011110",
  7146=>"101001100",
  7147=>"011101101",
  7148=>"100111001",
  7149=>"010011001",
  7150=>"110011110",
  7151=>"000001010",
  7152=>"001100011",
  7153=>"101010100",
  7154=>"000001001",
  7155=>"011101100",
  7156=>"000110100",
  7157=>"100010101",
  7158=>"100110011",
  7159=>"001010001",
  7160=>"000101100",
  7161=>"011100000",
  7162=>"100001010",
  7163=>"001010010",
  7164=>"000100001",
  7165=>"010111010",
  7166=>"000100100",
  7167=>"111110011",
  7168=>"011100010",
  7169=>"011111110",
  7170=>"101011101",
  7171=>"000011000",
  7172=>"001001111",
  7173=>"100000111",
  7174=>"110011000",
  7175=>"010010111",
  7176=>"011010011",
  7177=>"110101111",
  7178=>"001111100",
  7179=>"111001100",
  7180=>"111100101",
  7181=>"100100011",
  7182=>"101001011",
  7183=>"110101011",
  7184=>"011111101",
  7185=>"000101110",
  7186=>"011001001",
  7187=>"011001010",
  7188=>"111111011",
  7189=>"000001011",
  7190=>"100100100",
  7191=>"010111001",
  7192=>"100011010",
  7193=>"101111101",
  7194=>"100011011",
  7195=>"001110001",
  7196=>"101001101",
  7197=>"000010001",
  7198=>"000101100",
  7199=>"100001001",
  7200=>"001101101",
  7201=>"101110010",
  7202=>"100001000",
  7203=>"001101111",
  7204=>"101100110",
  7205=>"011110010",
  7206=>"001000001",
  7207=>"010111111",
  7208=>"100110011",
  7209=>"101111001",
  7210=>"001011011",
  7211=>"101010001",
  7212=>"111101000",
  7213=>"101111001",
  7214=>"010100001",
  7215=>"110111000",
  7216=>"110111010",
  7217=>"100101111",
  7218=>"101110100",
  7219=>"110110000",
  7220=>"110111000",
  7221=>"111110000",
  7222=>"000000101",
  7223=>"101110110",
  7224=>"100100101",
  7225=>"010011000",
  7226=>"101000011",
  7227=>"000000101",
  7228=>"100101011",
  7229=>"010101011",
  7230=>"010000011",
  7231=>"101000111",
  7232=>"100110101",
  7233=>"000011011",
  7234=>"000100110",
  7235=>"000100001",
  7236=>"001110011",
  7237=>"101110110",
  7238=>"011110011",
  7239=>"010010000",
  7240=>"100111101",
  7241=>"111011011",
  7242=>"010000001",
  7243=>"111001000",
  7244=>"000110001",
  7245=>"101110011",
  7246=>"011010010",
  7247=>"000010010",
  7248=>"110110010",
  7249=>"010000000",
  7250=>"100101111",
  7251=>"010000101",
  7252=>"000010100",
  7253=>"101110100",
  7254=>"000111000",
  7255=>"001101111",
  7256=>"011001011",
  7257=>"101100100",
  7258=>"110010111",
  7259=>"100000010",
  7260=>"000110110",
  7261=>"010001011",
  7262=>"111111101",
  7263=>"101000101",
  7264=>"101000001",
  7265=>"011001010",
  7266=>"000100100",
  7267=>"100100011",
  7268=>"101110010",
  7269=>"101011111",
  7270=>"100010010",
  7271=>"111010101",
  7272=>"101001001",
  7273=>"110111110",
  7274=>"100011010",
  7275=>"000001100",
  7276=>"101011000",
  7277=>"110010000",
  7278=>"001110000",
  7279=>"100001011",
  7280=>"100011001",
  7281=>"101101111",
  7282=>"111111001",
  7283=>"101011001",
  7284=>"011100000",
  7285=>"011101100",
  7286=>"110000000",
  7287=>"100100100",
  7288=>"111110111",
  7289=>"011001011",
  7290=>"101000101",
  7291=>"111000100",
  7292=>"000101101",
  7293=>"001010101",
  7294=>"011001010",
  7295=>"110100110",
  7296=>"011011111",
  7297=>"111101100",
  7298=>"100010010",
  7299=>"010111111",
  7300=>"111001011",
  7301=>"100111010",
  7302=>"010010001",
  7303=>"100111100",
  7304=>"101010011",
  7305=>"110010101",
  7306=>"001100011",
  7307=>"110100100",
  7308=>"111010100",
  7309=>"110111111",
  7310=>"111110111",
  7311=>"101100000",
  7312=>"100000011",
  7313=>"001000011",
  7314=>"000100100",
  7315=>"010010110",
  7316=>"100111001",
  7317=>"001010111",
  7318=>"001100100",
  7319=>"010111101",
  7320=>"111000011",
  7321=>"010110101",
  7322=>"101001010",
  7323=>"101001010",
  7324=>"010101100",
  7325=>"011111110",
  7326=>"011110011",
  7327=>"010001110",
  7328=>"000101101",
  7329=>"100100100",
  7330=>"010110010",
  7331=>"001010111",
  7332=>"100010111",
  7333=>"001010011",
  7334=>"010011011",
  7335=>"000010010",
  7336=>"000111010",
  7337=>"001100110",
  7338=>"011000001",
  7339=>"101100100",
  7340=>"001111000",
  7341=>"101000110",
  7342=>"011001100",
  7343=>"000001000",
  7344=>"011011010",
  7345=>"000010111",
  7346=>"010110001",
  7347=>"100111010",
  7348=>"110101101",
  7349=>"001010010",
  7350=>"110001100",
  7351=>"000100001",
  7352=>"110100000",
  7353=>"011011100",
  7354=>"010101101",
  7355=>"000110100",
  7356=>"101101100",
  7357=>"011000111",
  7358=>"011110001",
  7359=>"001011011",
  7360=>"100110001",
  7361=>"010110111",
  7362=>"110001111",
  7363=>"110001100",
  7364=>"101110110",
  7365=>"110100110",
  7366=>"111011000",
  7367=>"010111001",
  7368=>"100001010",
  7369=>"111100110",
  7370=>"001011100",
  7371=>"011110010",
  7372=>"101011110",
  7373=>"001001110",
  7374=>"000110000",
  7375=>"010111110",
  7376=>"010000000",
  7377=>"001100000",
  7378=>"011000100",
  7379=>"010001101",
  7380=>"111101111",
  7381=>"101110001",
  7382=>"111001000",
  7383=>"000011000",
  7384=>"101000100",
  7385=>"100100011",
  7386=>"000000111",
  7387=>"110111110",
  7388=>"000000100",
  7389=>"111011100",
  7390=>"111111110",
  7391=>"001100111",
  7392=>"111000101",
  7393=>"010110001",
  7394=>"010010101",
  7395=>"011110010",
  7396=>"100111100",
  7397=>"101100000",
  7398=>"100011100",
  7399=>"011000101",
  7400=>"110010110",
  7401=>"011000111",
  7402=>"001111100",
  7403=>"000011100",
  7404=>"010100000",
  7405=>"111001010",
  7406=>"100011100",
  7407=>"010110100",
  7408=>"100010010",
  7409=>"111111111",
  7410=>"101100100",
  7411=>"001011100",
  7412=>"100101110",
  7413=>"100110001",
  7414=>"100100100",
  7415=>"110011001",
  7416=>"001001000",
  7417=>"111101100",
  7418=>"001001100",
  7419=>"000111000",
  7420=>"001100011",
  7421=>"010011101",
  7422=>"000111010",
  7423=>"010001001",
  7424=>"111000100",
  7425=>"101000000",
  7426=>"001101111",
  7427=>"111111000",
  7428=>"101011000",
  7429=>"010000111",
  7430=>"010000111",
  7431=>"101011101",
  7432=>"001001001",
  7433=>"101110101",
  7434=>"010111111",
  7435=>"000001010",
  7436=>"010011101",
  7437=>"100011111",
  7438=>"001101011",
  7439=>"101101000",
  7440=>"100111110",
  7441=>"001001011",
  7442=>"000100010",
  7443=>"110010001",
  7444=>"011100011",
  7445=>"110100010",
  7446=>"100010111",
  7447=>"100110001",
  7448=>"000100000",
  7449=>"000101011",
  7450=>"000011010",
  7451=>"110001101",
  7452=>"110110101",
  7453=>"001101111",
  7454=>"100010010",
  7455=>"000000010",
  7456=>"110110001",
  7457=>"110010110",
  7458=>"101010110",
  7459=>"001111011",
  7460=>"010110011",
  7461=>"111100011",
  7462=>"100000110",
  7463=>"101000001",
  7464=>"101000011",
  7465=>"000111101",
  7466=>"000000011",
  7467=>"100011001",
  7468=>"001011001",
  7469=>"000000000",
  7470=>"000001110",
  7471=>"011001101",
  7472=>"101000001",
  7473=>"010010011",
  7474=>"111001101",
  7475=>"011001000",
  7476=>"010001000",
  7477=>"110011010",
  7478=>"110010101",
  7479=>"100001010",
  7480=>"011110110",
  7481=>"111100110",
  7482=>"000000001",
  7483=>"010010011",
  7484=>"111100101",
  7485=>"100000111",
  7486=>"101110000",
  7487=>"110011100",
  7488=>"010110111",
  7489=>"000101110",
  7490=>"001000011",
  7491=>"000010101",
  7492=>"101001000",
  7493=>"010110001",
  7494=>"010110000",
  7495=>"000001100",
  7496=>"100100110",
  7497=>"100010010",
  7498=>"010001110",
  7499=>"000101101",
  7500=>"100100011",
  7501=>"101101110",
  7502=>"001010101",
  7503=>"100111111",
  7504=>"001111101",
  7505=>"010001010",
  7506=>"000001101",
  7507=>"101111101",
  7508=>"111101110",
  7509=>"101010000",
  7510=>"000000110",
  7511=>"110111001",
  7512=>"011000110",
  7513=>"011111100",
  7514=>"010011000",
  7515=>"100010010",
  7516=>"111100010",
  7517=>"110100011",
  7518=>"110001100",
  7519=>"010011111",
  7520=>"011101101",
  7521=>"100101111",
  7522=>"000000100",
  7523=>"100101000",
  7524=>"101101110",
  7525=>"011100110",
  7526=>"011011101",
  7527=>"101101011",
  7528=>"001111001",
  7529=>"001000011",
  7530=>"101110011",
  7531=>"111101010",
  7532=>"101100001",
  7533=>"100001101",
  7534=>"000101010",
  7535=>"001101000",
  7536=>"101011000",
  7537=>"100100011",
  7538=>"100001110",
  7539=>"100010100",
  7540=>"111111000",
  7541=>"001000100",
  7542=>"100111001",
  7543=>"011000101",
  7544=>"100110111",
  7545=>"111000100",
  7546=>"000111010",
  7547=>"111101111",
  7548=>"101110101",
  7549=>"111101011",
  7550=>"111100110",
  7551=>"101001111",
  7552=>"101111011",
  7553=>"010111001",
  7554=>"101111001",
  7555=>"011110001",
  7556=>"001101010",
  7557=>"100111100",
  7558=>"010010101",
  7559=>"110101110",
  7560=>"010010110",
  7561=>"101101100",
  7562=>"001001001",
  7563=>"111101110",
  7564=>"000001110",
  7565=>"111010011",
  7566=>"001111111",
  7567=>"110011111",
  7568=>"111000100",
  7569=>"001111010",
  7570=>"100001100",
  7571=>"100100100",
  7572=>"101000111",
  7573=>"111111101",
  7574=>"001010010",
  7575=>"101101001",
  7576=>"101111000",
  7577=>"001101101",
  7578=>"110100000",
  7579=>"001101000",
  7580=>"100001100",
  7581=>"010110010",
  7582=>"101000101",
  7583=>"100001101",
  7584=>"001101000",
  7585=>"110100001",
  7586=>"000111100",
  7587=>"001100000",
  7588=>"010101101",
  7589=>"001000101",
  7590=>"100010011",
  7591=>"101010000",
  7592=>"111011100",
  7593=>"000000000",
  7594=>"110100101",
  7595=>"000000111",
  7596=>"100110101",
  7597=>"010111101",
  7598=>"101100100",
  7599=>"101110001",
  7600=>"100110011",
  7601=>"000111101",
  7602=>"111110111",
  7603=>"110100001",
  7604=>"011011010",
  7605=>"100100111",
  7606=>"111110111",
  7607=>"011101000",
  7608=>"011000100",
  7609=>"000011111",
  7610=>"000011010",
  7611=>"001010001",
  7612=>"001101111",
  7613=>"000000001",
  7614=>"001010111",
  7615=>"001100111",
  7616=>"000001101",
  7617=>"111110100",
  7618=>"101111000",
  7619=>"111010001",
  7620=>"010000000",
  7621=>"110101110",
  7622=>"100111111",
  7623=>"001111000",
  7624=>"101100100",
  7625=>"010011110",
  7626=>"110000001",
  7627=>"010001001",
  7628=>"001111001",
  7629=>"010100010",
  7630=>"100101010",
  7631=>"110101101",
  7632=>"001010011",
  7633=>"111111101",
  7634=>"100010101",
  7635=>"100110000",
  7636=>"100110001",
  7637=>"111001001",
  7638=>"100101110",
  7639=>"011011110",
  7640=>"111111010",
  7641=>"010111001",
  7642=>"110110101",
  7643=>"110010101",
  7644=>"001110101",
  7645=>"011101110",
  7646=>"100110111",
  7647=>"110110001",
  7648=>"111001011",
  7649=>"100110000",
  7650=>"000000000",
  7651=>"110000010",
  7652=>"110100001",
  7653=>"100100010",
  7654=>"011000111",
  7655=>"000010010",
  7656=>"111001000",
  7657=>"111101011",
  7658=>"001001010",
  7659=>"000110111",
  7660=>"101010101",
  7661=>"000010001",
  7662=>"100111011",
  7663=>"000100100",
  7664=>"111000001",
  7665=>"110001111",
  7666=>"000000110",
  7667=>"001001111",
  7668=>"010101010",
  7669=>"101000110",
  7670=>"000100111",
  7671=>"110011110",
  7672=>"111100111",
  7673=>"110111100",
  7674=>"001001010",
  7675=>"100010011",
  7676=>"100010111",
  7677=>"111101001",
  7678=>"100001101",
  7679=>"100111100",
  7680=>"010101001",
  7681=>"010110011",
  7682=>"001100001",
  7683=>"100000000",
  7684=>"011011110",
  7685=>"110010010",
  7686=>"110111011",
  7687=>"000101100",
  7688=>"011100110",
  7689=>"001111110",
  7690=>"010001011",
  7691=>"100010000",
  7692=>"000000000",
  7693=>"111011011",
  7694=>"000000001",
  7695=>"101001100",
  7696=>"100011001",
  7697=>"100111010",
  7698=>"111001111",
  7699=>"001001001",
  7700=>"001100000",
  7701=>"000000100",
  7702=>"010100001",
  7703=>"001111100",
  7704=>"000111011",
  7705=>"111010010",
  7706=>"111010011",
  7707=>"111110110",
  7708=>"110111111",
  7709=>"010001011",
  7710=>"111001011",
  7711=>"111101101",
  7712=>"000100011",
  7713=>"101110010",
  7714=>"000111110",
  7715=>"000110011",
  7716=>"010010101",
  7717=>"101000001",
  7718=>"011001111",
  7719=>"000110000",
  7720=>"110101000",
  7721=>"011010100",
  7722=>"111101011",
  7723=>"101110001",
  7724=>"000011101",
  7725=>"001111001",
  7726=>"101011111",
  7727=>"111110100",
  7728=>"011001110",
  7729=>"111111111",
  7730=>"110011101",
  7731=>"011111001",
  7732=>"111011110",
  7733=>"100100100",
  7734=>"100111101",
  7735=>"001011110",
  7736=>"011110100",
  7737=>"000010001",
  7738=>"011100101",
  7739=>"011100110",
  7740=>"100000010",
  7741=>"001001011",
  7742=>"000010000",
  7743=>"010101011",
  7744=>"000111101",
  7745=>"011000011",
  7746=>"011101001",
  7747=>"110101010",
  7748=>"111110000",
  7749=>"000111100",
  7750=>"111010100",
  7751=>"100111011",
  7752=>"000110111",
  7753=>"110001110",
  7754=>"000110110",
  7755=>"011110010",
  7756=>"011000111",
  7757=>"001010001",
  7758=>"110011111",
  7759=>"110101100",
  7760=>"111111111",
  7761=>"101000110",
  7762=>"101001001",
  7763=>"110101100",
  7764=>"100011100",
  7765=>"110000100",
  7766=>"011100001",
  7767=>"100010111",
  7768=>"110000001",
  7769=>"101000110",
  7770=>"011001010",
  7771=>"010001010",
  7772=>"001111111",
  7773=>"001010100",
  7774=>"101101110",
  7775=>"100110001",
  7776=>"011110100",
  7777=>"010001010",
  7778=>"110001010",
  7779=>"110110010",
  7780=>"000100010",
  7781=>"110010100",
  7782=>"001000110",
  7783=>"000110111",
  7784=>"010001110",
  7785=>"100111000",
  7786=>"000000111",
  7787=>"111010001",
  7788=>"001100110",
  7789=>"110011000",
  7790=>"001011101",
  7791=>"101101011",
  7792=>"111111010",
  7793=>"101101111",
  7794=>"111011100",
  7795=>"101101111",
  7796=>"010110111",
  7797=>"101000101",
  7798=>"100011011",
  7799=>"111000101",
  7800=>"001010110",
  7801=>"010010010",
  7802=>"110001000",
  7803=>"000000101",
  7804=>"101001000",
  7805=>"010001000",
  7806=>"001110110",
  7807=>"011111110",
  7808=>"000100110",
  7809=>"111111100",
  7810=>"110011111",
  7811=>"100100100",
  7812=>"111000100",
  7813=>"010000011",
  7814=>"001100001",
  7815=>"011001000",
  7816=>"010001110",
  7817=>"000101001",
  7818=>"110101101",
  7819=>"000010000",
  7820=>"010000110",
  7821=>"101001111",
  7822=>"001010011",
  7823=>"101000001",
  7824=>"010100100",
  7825=>"100001010",
  7826=>"000010011",
  7827=>"000001100",
  7828=>"101110110",
  7829=>"001001111",
  7830=>"011101100",
  7831=>"110101110",
  7832=>"101001010",
  7833=>"010101001",
  7834=>"101010001",
  7835=>"101011110",
  7836=>"101001010",
  7837=>"100110011",
  7838=>"000101001",
  7839=>"000000000",
  7840=>"110100000",
  7841=>"010010001",
  7842=>"100111011",
  7843=>"111000101",
  7844=>"101000010",
  7845=>"111011010",
  7846=>"001110101",
  7847=>"000010010",
  7848=>"101111101",
  7849=>"000000000",
  7850=>"000101010",
  7851=>"111101100",
  7852=>"101011000",
  7853=>"000000101",
  7854=>"100000101",
  7855=>"000100011",
  7856=>"110111000",
  7857=>"101011100",
  7858=>"010010001",
  7859=>"100100101",
  7860=>"100110001",
  7861=>"000001011",
  7862=>"000010101",
  7863=>"011001011",
  7864=>"101101100",
  7865=>"111001011",
  7866=>"100001011",
  7867=>"111111011",
  7868=>"110011111",
  7869=>"100011000",
  7870=>"101101110",
  7871=>"000001001",
  7872=>"010000000",
  7873=>"011111100",
  7874=>"011111001",
  7875=>"100111110",
  7876=>"001000010",
  7877=>"100110100",
  7878=>"100101111",
  7879=>"100110001",
  7880=>"001101001",
  7881=>"111110110",
  7882=>"101110011",
  7883=>"100101001",
  7884=>"011101111",
  7885=>"100100111",
  7886=>"001011001",
  7887=>"100001100",
  7888=>"011000001",
  7889=>"000001100",
  7890=>"000001110",
  7891=>"000010000",
  7892=>"101011101",
  7893=>"011000110",
  7894=>"000110000",
  7895=>"111111010",
  7896=>"001101111",
  7897=>"000111100",
  7898=>"011100001",
  7899=>"101010111",
  7900=>"111000101",
  7901=>"000110000",
  7902=>"110101111",
  7903=>"010101111",
  7904=>"100111010",
  7905=>"100101010",
  7906=>"010110010",
  7907=>"011100000",
  7908=>"101000100",
  7909=>"000111001",
  7910=>"010010100",
  7911=>"011000110",
  7912=>"101010001",
  7913=>"000101111",
  7914=>"010111110",
  7915=>"010100011",
  7916=>"010011011",
  7917=>"000101000",
  7918=>"000111100",
  7919=>"111101011",
  7920=>"100001100",
  7921=>"110010101",
  7922=>"010111110",
  7923=>"110110101",
  7924=>"100101111",
  7925=>"001011011",
  7926=>"001101110",
  7927=>"100010000",
  7928=>"101000111",
  7929=>"100001101",
  7930=>"000001111",
  7931=>"000010001",
  7932=>"010010001",
  7933=>"001111100",
  7934=>"110011001",
  7935=>"000000100",
  7936=>"010001000",
  7937=>"101110101",
  7938=>"001011101",
  7939=>"011100011",
  7940=>"110001100",
  7941=>"010101001",
  7942=>"111001010",
  7943=>"111111101",
  7944=>"111011111",
  7945=>"110011000",
  7946=>"111101111",
  7947=>"011101101",
  7948=>"010011001",
  7949=>"111110110",
  7950=>"000101100",
  7951=>"101111110",
  7952=>"100111001",
  7953=>"010111010",
  7954=>"001011100",
  7955=>"000011101",
  7956=>"101010110",
  7957=>"110111001",
  7958=>"001100011",
  7959=>"100010000",
  7960=>"111000000",
  7961=>"010111111",
  7962=>"000100110",
  7963=>"000000001",
  7964=>"010111001",
  7965=>"100111111",
  7966=>"000011101",
  7967=>"101111100",
  7968=>"111001101",
  7969=>"011110001",
  7970=>"111110111",
  7971=>"001010001",
  7972=>"110100010",
  7973=>"000000111",
  7974=>"100001010",
  7975=>"111110110",
  7976=>"110101101",
  7977=>"001101010",
  7978=>"110011100",
  7979=>"011011101",
  7980=>"001101000",
  7981=>"000000010",
  7982=>"001111110",
  7983=>"000000101",
  7984=>"000001111",
  7985=>"100111110",
  7986=>"000011100",
  7987=>"000010011",
  7988=>"111110101",
  7989=>"010111101",
  7990=>"011000100",
  7991=>"001101000",
  7992=>"000001000",
  7993=>"011000010",
  7994=>"101110101",
  7995=>"111100101",
  7996=>"111011000",
  7997=>"011110001",
  7998=>"001111101",
  7999=>"111111100",
  8000=>"101110101",
  8001=>"000111110",
  8002=>"101001011",
  8003=>"110001110",
  8004=>"010011010",
  8005=>"110000101",
  8006=>"010000100",
  8007=>"110111011",
  8008=>"001100100",
  8009=>"001100111",
  8010=>"101111111",
  8011=>"100101001",
  8012=>"000111001",
  8013=>"110001110",
  8014=>"010110001",
  8015=>"011011011",
  8016=>"100110010",
  8017=>"110100011",
  8018=>"100001101",
  8019=>"110010100",
  8020=>"100010110",
  8021=>"111001000",
  8022=>"100011100",
  8023=>"110001111",
  8024=>"110010010",
  8025=>"001000111",
  8026=>"100110000",
  8027=>"101011111",
  8028=>"110101101",
  8029=>"101100100",
  8030=>"000000110",
  8031=>"100000101",
  8032=>"011001010",
  8033=>"010101100",
  8034=>"101110010",
  8035=>"101001011",
  8036=>"001000101",
  8037=>"111100101",
  8038=>"001110001",
  8039=>"000001011",
  8040=>"010001000",
  8041=>"011011101",
  8042=>"110000001",
  8043=>"101011010",
  8044=>"110001001",
  8045=>"111111110",
  8046=>"001110011",
  8047=>"010010011",
  8048=>"011110111",
  8049=>"111011011",
  8050=>"011111010",
  8051=>"100010110",
  8052=>"001010010",
  8053=>"011100000",
  8054=>"001100101",
  8055=>"000000011",
  8056=>"110111111",
  8057=>"011111100",
  8058=>"100100111",
  8059=>"010101000",
  8060=>"101001110",
  8061=>"101101000",
  8062=>"101011001",
  8063=>"110001111",
  8064=>"010111000",
  8065=>"111101101",
  8066=>"010001010",
  8067=>"001000101",
  8068=>"100111011",
  8069=>"101000000",
  8070=>"100010001",
  8071=>"110111001",
  8072=>"100110110",
  8073=>"011101000",
  8074=>"001001110",
  8075=>"100110011",
  8076=>"011110010",
  8077=>"110010001",
  8078=>"110000101",
  8079=>"000001000",
  8080=>"001111111",
  8081=>"011111011",
  8082=>"001010000",
  8083=>"101001011",
  8084=>"100110000",
  8085=>"101110111",
  8086=>"000011100",
  8087=>"111000010",
  8088=>"100101110",
  8089=>"110110110",
  8090=>"100111110",
  8091=>"000010010",
  8092=>"101000001",
  8093=>"010001001",
  8094=>"111111001",
  8095=>"001100000",
  8096=>"101000101",
  8097=>"101101001",
  8098=>"100111011",
  8099=>"111100000",
  8100=>"000000000",
  8101=>"111011100",
  8102=>"111001000",
  8103=>"011000000",
  8104=>"001100000",
  8105=>"000010000",
  8106=>"000011110",
  8107=>"010001111",
  8108=>"000001111",
  8109=>"001011010",
  8110=>"010110110",
  8111=>"010010000",
  8112=>"100000110",
  8113=>"101001011",
  8114=>"111000010",
  8115=>"011110101",
  8116=>"110110110",
  8117=>"000010110",
  8118=>"000100101",
  8119=>"000111100",
  8120=>"010100010",
  8121=>"001000110",
  8122=>"011011000",
  8123=>"000000011",
  8124=>"101101111",
  8125=>"111010100",
  8126=>"001001111",
  8127=>"001101010",
  8128=>"110111111",
  8129=>"101101010",
  8130=>"111110110",
  8131=>"010101111",
  8132=>"100010001",
  8133=>"011010000",
  8134=>"111101000",
  8135=>"110100010",
  8136=>"000000011",
  8137=>"100100101",
  8138=>"101100111",
  8139=>"000011001",
  8140=>"110000001",
  8141=>"010000101",
  8142=>"011111000",
  8143=>"100111010",
  8144=>"011100101",
  8145=>"000011111",
  8146=>"011010111",
  8147=>"001110000",
  8148=>"011000100",
  8149=>"111111000",
  8150=>"010011000",
  8151=>"000001011",
  8152=>"111101111",
  8153=>"101111100",
  8154=>"101010001",
  8155=>"000000000",
  8156=>"111100001",
  8157=>"001100000",
  8158=>"110010011",
  8159=>"000001110",
  8160=>"101100010",
  8161=>"100011101",
  8162=>"011111011",
  8163=>"110001000",
  8164=>"000000110",
  8165=>"111000110",
  8166=>"011011000",
  8167=>"000001011",
  8168=>"101011111",
  8169=>"011001001",
  8170=>"111100011",
  8171=>"110111010",
  8172=>"010110110",
  8173=>"001111111",
  8174=>"010110000",
  8175=>"111101000",
  8176=>"010100000",
  8177=>"001001110",
  8178=>"011001001",
  8179=>"110000011",
  8180=>"101101001",
  8181=>"111010101",
  8182=>"100101101",
  8183=>"101010100",
  8184=>"101001111",
  8185=>"000100011",
  8186=>"111100111",
  8187=>"110001110",
  8188=>"000010010",
  8189=>"111010011",
  8190=>"001011011",
  8191=>"111110011",
  8192=>"001000000",
  8193=>"010110110",
  8194=>"000010111",
  8195=>"101110100",
  8196=>"010111111",
  8197=>"001011111",
  8198=>"011101110",
  8199=>"101000010",
  8200=>"111010000",
  8201=>"001100100",
  8202=>"010100001",
  8203=>"101100111",
  8204=>"010010010",
  8205=>"000110110",
  8206=>"011111100",
  8207=>"101111011",
  8208=>"001110001",
  8209=>"000000101",
  8210=>"110111100",
  8211=>"000010101",
  8212=>"100100110",
  8213=>"010100001",
  8214=>"101111110",
  8215=>"000001011",
  8216=>"100110010",
  8217=>"010100101",
  8218=>"000001101",
  8219=>"011000001",
  8220=>"000110111",
  8221=>"010110011",
  8222=>"001010101",
  8223=>"101100000",
  8224=>"111011011",
  8225=>"100000101",
  8226=>"001101010",
  8227=>"100110100",
  8228=>"111010011",
  8229=>"000010111",
  8230=>"101001010",
  8231=>"111000001",
  8232=>"000111111",
  8233=>"011111111",
  8234=>"001101101",
  8235=>"001100011",
  8236=>"011010111",
  8237=>"001110010",
  8238=>"100101100",
  8239=>"111111010",
  8240=>"100111000",
  8241=>"111111000",
  8242=>"011010001",
  8243=>"010001001",
  8244=>"010100001",
  8245=>"101001100",
  8246=>"101100000",
  8247=>"010011010",
  8248=>"110011010",
  8249=>"100000110",
  8250=>"001100110",
  8251=>"001010010",
  8252=>"011010111",
  8253=>"110001100",
  8254=>"101101100",
  8255=>"000010001",
  8256=>"010010010",
  8257=>"001101001",
  8258=>"010100100",
  8259=>"110101000",
  8260=>"010100110",
  8261=>"110000110",
  8262=>"111011001",
  8263=>"011100100",
  8264=>"010100000",
  8265=>"101001100",
  8266=>"010010100",
  8267=>"000110000",
  8268=>"011000010",
  8269=>"111110101",
  8270=>"100111001",
  8271=>"001101000",
  8272=>"111000100",
  8273=>"110100001",
  8274=>"101010001",
  8275=>"010010011",
  8276=>"011010001",
  8277=>"101011011",
  8278=>"001001110",
  8279=>"110001000",
  8280=>"010001100",
  8281=>"100011001",
  8282=>"101011101",
  8283=>"000011111",
  8284=>"110101000",
  8285=>"101100111",
  8286=>"000100110",
  8287=>"100001101",
  8288=>"110011000",
  8289=>"011001000",
  8290=>"111100101",
  8291=>"110100111",
  8292=>"110111010",
  8293=>"010110001",
  8294=>"101011111",
  8295=>"100011000",
  8296=>"010000111",
  8297=>"100110010",
  8298=>"101011101",
  8299=>"000110010",
  8300=>"011001010",
  8301=>"010100000",
  8302=>"010101010",
  8303=>"010000000",
  8304=>"101001001",
  8305=>"000000111",
  8306=>"010100011",
  8307=>"011110111",
  8308=>"100101000",
  8309=>"010000100",
  8310=>"001111110",
  8311=>"100111101",
  8312=>"100011001",
  8313=>"010011000",
  8314=>"000111011",
  8315=>"111100100",
  8316=>"100110111",
  8317=>"000101110",
  8318=>"010011000",
  8319=>"001101011",
  8320=>"000010001",
  8321=>"001010110",
  8322=>"111100000",
  8323=>"101010010",
  8324=>"110110000",
  8325=>"101000101",
  8326=>"011000001",
  8327=>"110110000",
  8328=>"100001100",
  8329=>"000001011",
  8330=>"011110001",
  8331=>"010011100",
  8332=>"101101100",
  8333=>"111011010",
  8334=>"011010000",
  8335=>"100110010",
  8336=>"010001111",
  8337=>"110000101",
  8338=>"000010011",
  8339=>"011010011",
  8340=>"111010111",
  8341=>"001011001",
  8342=>"000001001",
  8343=>"111101010",
  8344=>"101010110",
  8345=>"100011100",
  8346=>"100111010",
  8347=>"111100111",
  8348=>"010001110",
  8349=>"100111011",
  8350=>"110110111",
  8351=>"100111010",
  8352=>"101111000",
  8353=>"110010110",
  8354=>"101010000",
  8355=>"010001101",
  8356=>"100001111",
  8357=>"100110100",
  8358=>"101110011",
  8359=>"111000000",
  8360=>"011011001",
  8361=>"111110111",
  8362=>"000001001",
  8363=>"000111011",
  8364=>"011111110",
  8365=>"001100011",
  8366=>"100110001",
  8367=>"001110101",
  8368=>"000100101",
  8369=>"001101000",
  8370=>"000001110",
  8371=>"011100001",
  8372=>"111001111",
  8373=>"010000111",
  8374=>"010010010",
  8375=>"010100000",
  8376=>"010000001",
  8377=>"010010000",
  8378=>"001111010",
  8379=>"101101111",
  8380=>"001111011",
  8381=>"111110001",
  8382=>"011011111",
  8383=>"110010111",
  8384=>"000110101",
  8385=>"110111110",
  8386=>"001110001",
  8387=>"111101000",
  8388=>"110100111",
  8389=>"001010100",
  8390=>"011010101",
  8391=>"001011100",
  8392=>"001000111",
  8393=>"010010111",
  8394=>"111110100",
  8395=>"001101010",
  8396=>"101100010",
  8397=>"000001101",
  8398=>"011000000",
  8399=>"110000001",
  8400=>"100111110",
  8401=>"110011111",
  8402=>"110010101",
  8403=>"101110011",
  8404=>"100001000",
  8405=>"110110000",
  8406=>"010011101",
  8407=>"010111011",
  8408=>"111011000",
  8409=>"111101000",
  8410=>"101000111",
  8411=>"010011111",
  8412=>"100011011",
  8413=>"011110100",
  8414=>"000110011",
  8415=>"011101011",
  8416=>"111001010",
  8417=>"101101000",
  8418=>"001010111",
  8419=>"110111001",
  8420=>"011101100",
  8421=>"000111111",
  8422=>"100001000",
  8423=>"010011100",
  8424=>"010100000",
  8425=>"110111100",
  8426=>"010111101",
  8427=>"001111110",
  8428=>"111110100",
  8429=>"111110110",
  8430=>"100111001",
  8431=>"000100011",
  8432=>"111001101",
  8433=>"100110110",
  8434=>"111001101",
  8435=>"101101110",
  8436=>"000110110",
  8437=>"101000111",
  8438=>"101100011",
  8439=>"001000000",
  8440=>"011010111",
  8441=>"000110100",
  8442=>"010110101",
  8443=>"001111110",
  8444=>"110010010",
  8445=>"101000000",
  8446=>"110101010",
  8447=>"000001000",
  8448=>"110001100",
  8449=>"010100110",
  8450=>"000000110",
  8451=>"000101000",
  8452=>"010101010",
  8453=>"010010000",
  8454=>"101100000",
  8455=>"010010110",
  8456=>"111111000",
  8457=>"101101000",
  8458=>"111110000",
  8459=>"011101100",
  8460=>"000011001",
  8461=>"001111010",
  8462=>"011100101",
  8463=>"010000110",
  8464=>"101000011",
  8465=>"110000110",
  8466=>"011011001",
  8467=>"100010100",
  8468=>"000101000",
  8469=>"101001111",
  8470=>"000110010",
  8471=>"010111011",
  8472=>"100110101",
  8473=>"101001000",
  8474=>"100111010",
  8475=>"110110100",
  8476=>"000000100",
  8477=>"111001001",
  8478=>"100001100",
  8479=>"100111011",
  8480=>"111011110",
  8481=>"111010100",
  8482=>"011110111",
  8483=>"011100101",
  8484=>"100011100",
  8485=>"111110011",
  8486=>"110000110",
  8487=>"111001110",
  8488=>"100010111",
  8489=>"001100010",
  8490=>"000100011",
  8491=>"101001101",
  8492=>"101101100",
  8493=>"100000000",
  8494=>"110101011",
  8495=>"010100100",
  8496=>"000101011",
  8497=>"000001000",
  8498=>"000101100",
  8499=>"000101000",
  8500=>"101010010",
  8501=>"100101010",
  8502=>"111001110",
  8503=>"010111010",
  8504=>"101100100",
  8505=>"000100000",
  8506=>"011001111",
  8507=>"000010110",
  8508=>"011001111",
  8509=>"100110110",
  8510=>"100011011",
  8511=>"000111001",
  8512=>"011010011",
  8513=>"010101110",
  8514=>"010000000",
  8515=>"011011010",
  8516=>"011100011",
  8517=>"011001111",
  8518=>"001010000",
  8519=>"101011011",
  8520=>"001100101",
  8521=>"100001010",
  8522=>"111011100",
  8523=>"100010010",
  8524=>"011001011",
  8525=>"000101011",
  8526=>"101010010",
  8527=>"110101000",
  8528=>"110100011",
  8529=>"001110100",
  8530=>"111100111",
  8531=>"110011000",
  8532=>"100110010",
  8533=>"000101001",
  8534=>"101001000",
  8535=>"000001111",
  8536=>"101110100",
  8537=>"101101110",
  8538=>"001011101",
  8539=>"110000011",
  8540=>"010111000",
  8541=>"011001100",
  8542=>"000100000",
  8543=>"000010001",
  8544=>"000010010",
  8545=>"111010110",
  8546=>"111000001",
  8547=>"001010100",
  8548=>"101000110",
  8549=>"100101100",
  8550=>"100010100",
  8551=>"100101100",
  8552=>"001111111",
  8553=>"000101010",
  8554=>"000100100",
  8555=>"101101101",
  8556=>"010001000",
  8557=>"111010100",
  8558=>"100001111",
  8559=>"101011101",
  8560=>"101100110",
  8561=>"001000100",
  8562=>"000011000",
  8563=>"110001001",
  8564=>"100000101",
  8565=>"100011010",
  8566=>"010110101",
  8567=>"111001001",
  8568=>"100010011",
  8569=>"101010100",
  8570=>"101011010",
  8571=>"010110000",
  8572=>"110100001",
  8573=>"111110011",
  8574=>"000000001",
  8575=>"100111110",
  8576=>"010100101",
  8577=>"101000010",
  8578=>"110111111",
  8579=>"100101000",
  8580=>"010001010",
  8581=>"001011100",
  8582=>"001111000",
  8583=>"100010001",
  8584=>"000100111",
  8585=>"100011110",
  8586=>"001100001",
  8587=>"001100010",
  8588=>"001000100",
  8589=>"011100001",
  8590=>"000000001",
  8591=>"001010010",
  8592=>"010110110",
  8593=>"011100010",
  8594=>"100101010",
  8595=>"101101100",
  8596=>"001001000",
  8597=>"000100110",
  8598=>"000010010",
  8599=>"110010001",
  8600=>"001110111",
  8601=>"101011101",
  8602=>"001001010",
  8603=>"110011000",
  8604=>"011000111",
  8605=>"100101001",
  8606=>"110100010",
  8607=>"101011011",
  8608=>"001000010",
  8609=>"111101100",
  8610=>"100100001",
  8611=>"101111111",
  8612=>"101000111",
  8613=>"100100100",
  8614=>"111110001",
  8615=>"111111111",
  8616=>"111101110",
  8617=>"010110000",
  8618=>"011011100",
  8619=>"010001111",
  8620=>"111101010",
  8621=>"000101100",
  8622=>"100111000",
  8623=>"100100010",
  8624=>"001011110",
  8625=>"111000101",
  8626=>"100111001",
  8627=>"011011000",
  8628=>"000101001",
  8629=>"111111111",
  8630=>"010101011",
  8631=>"011100110",
  8632=>"000110101",
  8633=>"110000000",
  8634=>"001011001",
  8635=>"000001100",
  8636=>"111100110",
  8637=>"001010010",
  8638=>"111001000",
  8639=>"110100010",
  8640=>"110001000",
  8641=>"010000000",
  8642=>"001010011",
  8643=>"101001111",
  8644=>"100011100",
  8645=>"011111010",
  8646=>"100100111",
  8647=>"000100001",
  8648=>"000101010",
  8649=>"110010000",
  8650=>"011110110",
  8651=>"000100110",
  8652=>"100110111",
  8653=>"010100011",
  8654=>"111111110",
  8655=>"010100100",
  8656=>"101101000",
  8657=>"001011100",
  8658=>"100111000",
  8659=>"000010011",
  8660=>"010000001",
  8661=>"110010011",
  8662=>"110100000",
  8663=>"111111001",
  8664=>"101111111",
  8665=>"100111111",
  8666=>"001010010",
  8667=>"000000010",
  8668=>"101000100",
  8669=>"001001101",
  8670=>"110011010",
  8671=>"100101101",
  8672=>"101101110",
  8673=>"101000111",
  8674=>"111001000",
  8675=>"100110011",
  8676=>"011001110",
  8677=>"011000000",
  8678=>"010000110",
  8679=>"000111000",
  8680=>"000101000",
  8681=>"101111011",
  8682=>"101101110",
  8683=>"101111001",
  8684=>"010001000",
  8685=>"101111011",
  8686=>"011110111",
  8687=>"011010111",
  8688=>"100100110",
  8689=>"000001100",
  8690=>"101000010",
  8691=>"110111110",
  8692=>"100000111",
  8693=>"100100111",
  8694=>"010011101",
  8695=>"110011000",
  8696=>"111001011",
  8697=>"111100000",
  8698=>"000110001",
  8699=>"111100000",
  8700=>"000010110",
  8701=>"001000110",
  8702=>"100111011",
  8703=>"100000010",
  8704=>"110000000",
  8705=>"000110100",
  8706=>"101101111",
  8707=>"000010100",
  8708=>"001011110",
  8709=>"101100111",
  8710=>"100010100",
  8711=>"100101001",
  8712=>"000011001",
  8713=>"100011100",
  8714=>"110100001",
  8715=>"010010001",
  8716=>"000101000",
  8717=>"110010111",
  8718=>"011100100",
  8719=>"110111111",
  8720=>"110010111",
  8721=>"111111001",
  8722=>"111001111",
  8723=>"010000000",
  8724=>"101100011",
  8725=>"100001000",
  8726=>"110101100",
  8727=>"011001101",
  8728=>"110001001",
  8729=>"000110100",
  8730=>"110110011",
  8731=>"011000110",
  8732=>"011000110",
  8733=>"110101101",
  8734=>"111011011",
  8735=>"001111101",
  8736=>"111000011",
  8737=>"001101110",
  8738=>"010000110",
  8739=>"000001101",
  8740=>"010111110",
  8741=>"001111100",
  8742=>"000010111",
  8743=>"000001101",
  8744=>"010101111",
  8745=>"100111100",
  8746=>"111000111",
  8747=>"101001111",
  8748=>"100111111",
  8749=>"101111100",
  8750=>"001111101",
  8751=>"000001110",
  8752=>"110001001",
  8753=>"111111111",
  8754=>"111110000",
  8755=>"111000011",
  8756=>"001011110",
  8757=>"110010010",
  8758=>"010110110",
  8759=>"010000111",
  8760=>"101010110",
  8761=>"000110001",
  8762=>"010010110",
  8763=>"011110000",
  8764=>"011010000",
  8765=>"101010100",
  8766=>"110000011",
  8767=>"011001010",
  8768=>"101011101",
  8769=>"011111010",
  8770=>"000011000",
  8771=>"101010000",
  8772=>"100000001",
  8773=>"101000011",
  8774=>"011010000",
  8775=>"000000111",
  8776=>"111110111",
  8777=>"110000001",
  8778=>"100101011",
  8779=>"100000010",
  8780=>"011111001",
  8781=>"010000001",
  8782=>"010110100",
  8783=>"110100101",
  8784=>"100111110",
  8785=>"000101101",
  8786=>"011110111",
  8787=>"011101001",
  8788=>"110011010",
  8789=>"111011000",
  8790=>"110011110",
  8791=>"010110010",
  8792=>"001000110",
  8793=>"011110100",
  8794=>"010000101",
  8795=>"101010100",
  8796=>"011111101",
  8797=>"110100011",
  8798=>"100100110",
  8799=>"110110111",
  8800=>"101001101",
  8801=>"010000000",
  8802=>"110000000",
  8803=>"101011011",
  8804=>"111001101",
  8805=>"110110111",
  8806=>"101011011",
  8807=>"100100110",
  8808=>"001000010",
  8809=>"101001001",
  8810=>"100101001",
  8811=>"001110100",
  8812=>"110000100",
  8813=>"100101100",
  8814=>"100111000",
  8815=>"011100101",
  8816=>"100101000",
  8817=>"000011000",
  8818=>"110000011",
  8819=>"000001100",
  8820=>"010101011",
  8821=>"110101110",
  8822=>"011000010",
  8823=>"001110000",
  8824=>"101010011",
  8825=>"011011111",
  8826=>"000110001",
  8827=>"000000000",
  8828=>"000001011",
  8829=>"010101110",
  8830=>"110111101",
  8831=>"101011000",
  8832=>"111011101",
  8833=>"100110011",
  8834=>"110100000",
  8835=>"110001011",
  8836=>"100110010",
  8837=>"010111101",
  8838=>"010011110",
  8839=>"111110100",
  8840=>"001111110",
  8841=>"000011100",
  8842=>"010011001",
  8843=>"001000011",
  8844=>"010011101",
  8845=>"001011101",
  8846=>"110010100",
  8847=>"010011111",
  8848=>"101010000",
  8849=>"011100111",
  8850=>"010110011",
  8851=>"001110101",
  8852=>"000111110",
  8853=>"111110010",
  8854=>"011010110",
  8855=>"010101110",
  8856=>"100001010",
  8857=>"110101001",
  8858=>"101100000",
  8859=>"110011001",
  8860=>"101010001",
  8861=>"011101100",
  8862=>"000011101",
  8863=>"001111101",
  8864=>"010111110",
  8865=>"101101110",
  8866=>"101111001",
  8867=>"000101000",
  8868=>"111010101",
  8869=>"100011100",
  8870=>"100110111",
  8871=>"011000010",
  8872=>"111011001",
  8873=>"010001000",
  8874=>"110011100",
  8875=>"110100100",
  8876=>"111000011",
  8877=>"010101101",
  8878=>"111001000",
  8879=>"110000110",
  8880=>"000011010",
  8881=>"111000111",
  8882=>"011001010",
  8883=>"000001111",
  8884=>"010100101",
  8885=>"010110101",
  8886=>"100110101",
  8887=>"110010111",
  8888=>"001010110",
  8889=>"111000011",
  8890=>"000000100",
  8891=>"110101101",
  8892=>"110001101",
  8893=>"011000011",
  8894=>"110010110",
  8895=>"011100001",
  8896=>"101101111",
  8897=>"101111000",
  8898=>"111011110",
  8899=>"010111110",
  8900=>"010101101",
  8901=>"011110110",
  8902=>"110110011",
  8903=>"111110011",
  8904=>"101000000",
  8905=>"001111111",
  8906=>"110111001",
  8907=>"000101010",
  8908=>"011001010",
  8909=>"100000111",
  8910=>"110011110",
  8911=>"000101000",
  8912=>"011000100",
  8913=>"101110000",
  8914=>"110000001",
  8915=>"010011100",
  8916=>"101011111",
  8917=>"011111110",
  8918=>"101100100",
  8919=>"101100001",
  8920=>"001111100",
  8921=>"110110101",
  8922=>"110001001",
  8923=>"010010110",
  8924=>"100100100",
  8925=>"011010000",
  8926=>"100001111",
  8927=>"110001111",
  8928=>"101110010",
  8929=>"000110001",
  8930=>"100100110",
  8931=>"111010000",
  8932=>"110100101",
  8933=>"000101110",
  8934=>"111111110",
  8935=>"001011010",
  8936=>"110111110",
  8937=>"001011010",
  8938=>"100001011",
  8939=>"100011101",
  8940=>"010000010",
  8941=>"011010110",
  8942=>"000100001",
  8943=>"010100000",
  8944=>"111011001",
  8945=>"001111101",
  8946=>"111111111",
  8947=>"010010011",
  8948=>"010110001",
  8949=>"100001011",
  8950=>"110010101",
  8951=>"101100110",
  8952=>"001111011",
  8953=>"010100011",
  8954=>"010000101",
  8955=>"001101000",
  8956=>"000001110",
  8957=>"000010011",
  8958=>"011001111",
  8959=>"011000000",
  8960=>"110010011",
  8961=>"001000111",
  8962=>"100110000",
  8963=>"001110110",
  8964=>"101111011",
  8965=>"110000010",
  8966=>"100011110",
  8967=>"000100111",
  8968=>"001010011",
  8969=>"101111001",
  8970=>"110111001",
  8971=>"000010000",
  8972=>"001000100",
  8973=>"000011011",
  8974=>"110101111",
  8975=>"011000000",
  8976=>"000101111",
  8977=>"101111001",
  8978=>"100000010",
  8979=>"001011100",
  8980=>"100010010",
  8981=>"010011000",
  8982=>"000100001",
  8983=>"010000010",
  8984=>"111110111",
  8985=>"100101111",
  8986=>"001000011",
  8987=>"110110010",
  8988=>"110100101",
  8989=>"011101000",
  8990=>"100010100",
  8991=>"111011100",
  8992=>"010100010",
  8993=>"001011111",
  8994=>"000000010",
  8995=>"010010010",
  8996=>"000000000",
  8997=>"101100011",
  8998=>"101000110",
  8999=>"011111101",
  9000=>"000010011",
  9001=>"011001110",
  9002=>"101100101",
  9003=>"011010000",
  9004=>"101000001",
  9005=>"100101000",
  9006=>"110110100",
  9007=>"000101111",
  9008=>"010100100",
  9009=>"110010100",
  9010=>"100111010",
  9011=>"101101010",
  9012=>"011111011",
  9013=>"001001000",
  9014=>"001000110",
  9015=>"011001010",
  9016=>"111010100",
  9017=>"101101101",
  9018=>"101111011",
  9019=>"101010010",
  9020=>"111101000",
  9021=>"000101100",
  9022=>"000000100",
  9023=>"010111000",
  9024=>"000000100",
  9025=>"110111111",
  9026=>"010000100",
  9027=>"001111111",
  9028=>"001011111",
  9029=>"010000010",
  9030=>"100011100",
  9031=>"111110100",
  9032=>"010101011",
  9033=>"000100000",
  9034=>"000000010",
  9035=>"101011011",
  9036=>"001011011",
  9037=>"110000000",
  9038=>"110011111",
  9039=>"010000101",
  9040=>"110110110",
  9041=>"101010000",
  9042=>"101001111",
  9043=>"111100010",
  9044=>"000101011",
  9045=>"111111000",
  9046=>"010111101",
  9047=>"011010101",
  9048=>"111100111",
  9049=>"001101100",
  9050=>"001000111",
  9051=>"001100111",
  9052=>"101101110",
  9053=>"011111011",
  9054=>"011110111",
  9055=>"100000101",
  9056=>"111000110",
  9057=>"110101011",
  9058=>"010110001",
  9059=>"001001100",
  9060=>"001001001",
  9061=>"001001100",
  9062=>"100010001",
  9063=>"001001010",
  9064=>"001001000",
  9065=>"101111001",
  9066=>"111001000",
  9067=>"011100000",
  9068=>"011100001",
  9069=>"010101111",
  9070=>"010110100",
  9071=>"111010000",
  9072=>"011010001",
  9073=>"000010000",
  9074=>"101101001",
  9075=>"011100001",
  9076=>"110010101",
  9077=>"010100010",
  9078=>"100111111",
  9079=>"100111101",
  9080=>"001111001",
  9081=>"100001000",
  9082=>"101100111",
  9083=>"110110111",
  9084=>"000000000",
  9085=>"011001001",
  9086=>"100010001",
  9087=>"110011110",
  9088=>"101110111",
  9089=>"000010100",
  9090=>"110000111",
  9091=>"101111001",
  9092=>"011101100",
  9093=>"011000010",
  9094=>"010000111",
  9095=>"100100000",
  9096=>"001111110",
  9097=>"111000011",
  9098=>"011001000",
  9099=>"011111010",
  9100=>"100101100",
  9101=>"011110111",
  9102=>"000101101",
  9103=>"111100110",
  9104=>"110110110",
  9105=>"000010000",
  9106=>"000110000",
  9107=>"100101011",
  9108=>"010011101",
  9109=>"001111011",
  9110=>"010101001",
  9111=>"000110010",
  9112=>"000111000",
  9113=>"111001001",
  9114=>"100010111",
  9115=>"111111011",
  9116=>"100111011",
  9117=>"101110101",
  9118=>"011111111",
  9119=>"110000101",
  9120=>"001001010",
  9121=>"010010010",
  9122=>"100011010",
  9123=>"110011001",
  9124=>"001010110",
  9125=>"001111010",
  9126=>"000011000",
  9127=>"000101110",
  9128=>"100110100",
  9129=>"000110111",
  9130=>"100010101",
  9131=>"010111000",
  9132=>"110101110",
  9133=>"010101110",
  9134=>"001100001",
  9135=>"100000011",
  9136=>"010010111",
  9137=>"000111100",
  9138=>"010001001",
  9139=>"101001111",
  9140=>"010101110",
  9141=>"000000011",
  9142=>"010010011",
  9143=>"110111111",
  9144=>"010011101",
  9145=>"100010100",
  9146=>"101000011",
  9147=>"000110110",
  9148=>"110101010",
  9149=>"111010111",
  9150=>"100101010",
  9151=>"010011101",
  9152=>"010101010",
  9153=>"101100000",
  9154=>"100011011",
  9155=>"101011110",
  9156=>"101110111",
  9157=>"110010011",
  9158=>"101101000",
  9159=>"000000010",
  9160=>"101101100",
  9161=>"000001111",
  9162=>"000101110",
  9163=>"111010001",
  9164=>"101100010",
  9165=>"000110011",
  9166=>"000000001",
  9167=>"100000011",
  9168=>"001100111",
  9169=>"001111111",
  9170=>"000110001",
  9171=>"101111001",
  9172=>"011011110",
  9173=>"110000001",
  9174=>"111100001",
  9175=>"101111011",
  9176=>"110000011",
  9177=>"000001010",
  9178=>"110011100",
  9179=>"100011000",
  9180=>"101101001",
  9181=>"011100100",
  9182=>"100110100",
  9183=>"101100000",
  9184=>"011010100",
  9185=>"001001101",
  9186=>"111000111",
  9187=>"101010110",
  9188=>"100110001",
  9189=>"011001111",
  9190=>"011110111",
  9191=>"001000101",
  9192=>"010001101",
  9193=>"100000010",
  9194=>"110110011",
  9195=>"001010010",
  9196=>"010000111",
  9197=>"001010011",
  9198=>"101000101",
  9199=>"111010101",
  9200=>"000000110",
  9201=>"100110000",
  9202=>"011010000",
  9203=>"111001100",
  9204=>"000000010",
  9205=>"001010000",
  9206=>"111100111",
  9207=>"010110011",
  9208=>"000101010",
  9209=>"100110010",
  9210=>"101010001",
  9211=>"111101110",
  9212=>"100110010",
  9213=>"010110010",
  9214=>"101100010",
  9215=>"011001101",
  9216=>"000100111",
  9217=>"000011100",
  9218=>"110000010",
  9219=>"001111100",
  9220=>"101100101",
  9221=>"100000100",
  9222=>"100101100",
  9223=>"111111110",
  9224=>"000001001",
  9225=>"100011001",
  9226=>"101001001",
  9227=>"110011101",
  9228=>"110101100",
  9229=>"111101100",
  9230=>"000000110",
  9231=>"000111001",
  9232=>"101100010",
  9233=>"111101110",
  9234=>"101100101",
  9235=>"011100110",
  9236=>"011111110",
  9237=>"001010011",
  9238=>"000111001",
  9239=>"101000110",
  9240=>"011011000",
  9241=>"000110110",
  9242=>"000001001",
  9243=>"001010000",
  9244=>"101000111",
  9245=>"011001101",
  9246=>"000011000",
  9247=>"100010101",
  9248=>"111100000",
  9249=>"111010001",
  9250=>"011011111",
  9251=>"010111011",
  9252=>"110001111",
  9253=>"111111100",
  9254=>"100011101",
  9255=>"011011011",
  9256=>"000000000",
  9257=>"110000101",
  9258=>"111111101",
  9259=>"100111110",
  9260=>"010010011",
  9261=>"101010010",
  9262=>"000111011",
  9263=>"111010110",
  9264=>"000010000",
  9265=>"001110100",
  9266=>"100001100",
  9267=>"000000010",
  9268=>"110101110",
  9269=>"110111111",
  9270=>"011100010",
  9271=>"110111010",
  9272=>"111001100",
  9273=>"110100010",
  9274=>"101011111",
  9275=>"111111110",
  9276=>"010011101",
  9277=>"001101101",
  9278=>"010010010",
  9279=>"010111110",
  9280=>"010011101",
  9281=>"110111101",
  9282=>"111010101",
  9283=>"010111111",
  9284=>"110110111",
  9285=>"001000111",
  9286=>"010101100",
  9287=>"100010100",
  9288=>"101110010",
  9289=>"001011010",
  9290=>"101010111",
  9291=>"111111110",
  9292=>"010100010",
  9293=>"011001011",
  9294=>"001010001",
  9295=>"001101101",
  9296=>"010001111",
  9297=>"100110111",
  9298=>"101101000",
  9299=>"001100011",
  9300=>"111000100",
  9301=>"101101101",
  9302=>"010011011",
  9303=>"101011000",
  9304=>"011010001",
  9305=>"000111100",
  9306=>"110111110",
  9307=>"111001111",
  9308=>"000000001",
  9309=>"110111110",
  9310=>"111111111",
  9311=>"111111111",
  9312=>"000011001",
  9313=>"100011101",
  9314=>"010001101",
  9315=>"001111111",
  9316=>"101000100",
  9317=>"110001110",
  9318=>"100000000",
  9319=>"000111101",
  9320=>"010001100",
  9321=>"100101010",
  9322=>"110001000",
  9323=>"111100111",
  9324=>"110101011",
  9325=>"101100011",
  9326=>"111011111",
  9327=>"000101111",
  9328=>"001101100",
  9329=>"110001001",
  9330=>"110011001",
  9331=>"011111111",
  9332=>"010100100",
  9333=>"100000100",
  9334=>"011010000",
  9335=>"100111100",
  9336=>"010111011",
  9337=>"000110000",
  9338=>"101000000",
  9339=>"101100111",
  9340=>"111000110",
  9341=>"010101001",
  9342=>"011101110",
  9343=>"000101100",
  9344=>"010011101",
  9345=>"010111110",
  9346=>"111111101",
  9347=>"110101000",
  9348=>"111111111",
  9349=>"110111101",
  9350=>"010000000",
  9351=>"100010100",
  9352=>"010101100",
  9353=>"011010011",
  9354=>"100111000",
  9355=>"101101100",
  9356=>"110111010",
  9357=>"101111000",
  9358=>"111111011",
  9359=>"111110110",
  9360=>"011000011",
  9361=>"001100011",
  9362=>"110001001",
  9363=>"010100111",
  9364=>"110010001",
  9365=>"011101111",
  9366=>"101111010",
  9367=>"000110110",
  9368=>"111110100",
  9369=>"000010110",
  9370=>"010101000",
  9371=>"010100101",
  9372=>"110000100",
  9373=>"100111000",
  9374=>"100111000",
  9375=>"000010010",
  9376=>"011101011",
  9377=>"101011010",
  9378=>"011001111",
  9379=>"100000010",
  9380=>"001100001",
  9381=>"011110011",
  9382=>"111011110",
  9383=>"110100100",
  9384=>"101100011",
  9385=>"000001100",
  9386=>"011101101",
  9387=>"101001010",
  9388=>"000111011",
  9389=>"101111100",
  9390=>"111111000",
  9391=>"001010000",
  9392=>"111101001",
  9393=>"111001101",
  9394=>"101100101",
  9395=>"110111111",
  9396=>"010010001",
  9397=>"111110101",
  9398=>"111010011",
  9399=>"100000110",
  9400=>"110010101",
  9401=>"001101000",
  9402=>"111111010",
  9403=>"111110011",
  9404=>"010110000",
  9405=>"101101100",
  9406=>"111101110",
  9407=>"010101011",
  9408=>"011111111",
  9409=>"001010001",
  9410=>"100001011",
  9411=>"101001010",
  9412=>"000000010",
  9413=>"111111010",
  9414=>"011111000",
  9415=>"110111101",
  9416=>"000100010",
  9417=>"101101101",
  9418=>"100111100",
  9419=>"001011100",
  9420=>"000000001",
  9421=>"111100101",
  9422=>"101011111",
  9423=>"101100010",
  9424=>"011010011",
  9425=>"000101100",
  9426=>"110110110",
  9427=>"001101001",
  9428=>"100011111",
  9429=>"010101100",
  9430=>"001000010",
  9431=>"101010001",
  9432=>"010111111",
  9433=>"111001100",
  9434=>"110100001",
  9435=>"011111111",
  9436=>"001001001",
  9437=>"000000001",
  9438=>"101111100",
  9439=>"001110111",
  9440=>"111110101",
  9441=>"001110001",
  9442=>"110010011",
  9443=>"110011111",
  9444=>"001110100",
  9445=>"100100100",
  9446=>"000110111",
  9447=>"111100011",
  9448=>"011011110",
  9449=>"101101010",
  9450=>"010010100",
  9451=>"100101000",
  9452=>"111101000",
  9453=>"100010111",
  9454=>"111110110",
  9455=>"001100111",
  9456=>"000000000",
  9457=>"101011010",
  9458=>"111111101",
  9459=>"011110110",
  9460=>"111110101",
  9461=>"000011000",
  9462=>"111110001",
  9463=>"100100101",
  9464=>"111110000",
  9465=>"101010001",
  9466=>"111101111",
  9467=>"001110101",
  9468=>"010100100",
  9469=>"100110001",
  9470=>"000111011",
  9471=>"001010000",
  9472=>"011101001",
  9473=>"110101010",
  9474=>"011000001",
  9475=>"110011101",
  9476=>"111010001",
  9477=>"110010001",
  9478=>"011010010",
  9479=>"000010101",
  9480=>"010111010",
  9481=>"110111110",
  9482=>"101110011",
  9483=>"110111111",
  9484=>"100111011",
  9485=>"111000101",
  9486=>"110101110",
  9487=>"111001111",
  9488=>"100001000",
  9489=>"010111000",
  9490=>"101011110",
  9491=>"010001011",
  9492=>"000011111",
  9493=>"011110011",
  9494=>"001000101",
  9495=>"111001000",
  9496=>"011010100",
  9497=>"101111010",
  9498=>"111111101",
  9499=>"001001110",
  9500=>"111110111",
  9501=>"111110110",
  9502=>"010100011",
  9503=>"111100011",
  9504=>"111110111",
  9505=>"000100111",
  9506=>"100001111",
  9507=>"111111011",
  9508=>"110110111",
  9509=>"010111001",
  9510=>"110010000",
  9511=>"010000100",
  9512=>"001100100",
  9513=>"001010000",
  9514=>"101000111",
  9515=>"011111111",
  9516=>"111011101",
  9517=>"000111111",
  9518=>"111111111",
  9519=>"111110100",
  9520=>"010001100",
  9521=>"100111100",
  9522=>"111110001",
  9523=>"011101100",
  9524=>"110011000",
  9525=>"001000111",
  9526=>"000000000",
  9527=>"101011100",
  9528=>"111110111",
  9529=>"010100001",
  9530=>"100100110",
  9531=>"110101000",
  9532=>"110100010",
  9533=>"001011001",
  9534=>"110100100",
  9535=>"111101001",
  9536=>"101101010",
  9537=>"010010101",
  9538=>"101111010",
  9539=>"010100011",
  9540=>"100111011",
  9541=>"000101110",
  9542=>"110111110",
  9543=>"001010101",
  9544=>"100011111",
  9545=>"101111111",
  9546=>"000111110",
  9547=>"111111100",
  9548=>"111110001",
  9549=>"101111101",
  9550=>"011111101",
  9551=>"101111000",
  9552=>"110110101",
  9553=>"110100111",
  9554=>"100111010",
  9555=>"110101111",
  9556=>"101000110",
  9557=>"111110100",
  9558=>"010101101",
  9559=>"101101100",
  9560=>"111011011",
  9561=>"101011011",
  9562=>"011101010",
  9563=>"000101110",
  9564=>"010110010",
  9565=>"000001001",
  9566=>"100111001",
  9567=>"111110000",
  9568=>"111101000",
  9569=>"000000100",
  9570=>"010011111",
  9571=>"111101111",
  9572=>"100101001",
  9573=>"100100100",
  9574=>"111011000",
  9575=>"001010110",
  9576=>"010000001",
  9577=>"100111100",
  9578=>"111101100",
  9579=>"110101001",
  9580=>"111011001",
  9581=>"110000010",
  9582=>"001111101",
  9583=>"000011110",
  9584=>"111001100",
  9585=>"011110011",
  9586=>"100000000",
  9587=>"100010101",
  9588=>"011101111",
  9589=>"001001110",
  9590=>"101000000",
  9591=>"110000110",
  9592=>"111111100",
  9593=>"111010010",
  9594=>"010000000",
  9595=>"101010101",
  9596=>"100100001",
  9597=>"000110011",
  9598=>"010001110",
  9599=>"101110100",
  9600=>"110101010",
  9601=>"101110001",
  9602=>"100010000",
  9603=>"011000111",
  9604=>"000011001",
  9605=>"111011011",
  9606=>"111100001",
  9607=>"110000100",
  9608=>"001010111",
  9609=>"000110100",
  9610=>"111111111",
  9611=>"011010101",
  9612=>"111111001",
  9613=>"000000111",
  9614=>"110101101",
  9615=>"101111000",
  9616=>"000101101",
  9617=>"101111111",
  9618=>"110010001",
  9619=>"110011011",
  9620=>"110100010",
  9621=>"011100111",
  9622=>"100111101",
  9623=>"001000011",
  9624=>"101100001",
  9625=>"111111111",
  9626=>"101010100",
  9627=>"010111100",
  9628=>"100010111",
  9629=>"000001100",
  9630=>"111010101",
  9631=>"111111011",
  9632=>"111101100",
  9633=>"100001110",
  9634=>"001101110",
  9635=>"111111111",
  9636=>"101100000",
  9637=>"000111101",
  9638=>"000000100",
  9639=>"101010100",
  9640=>"011100010",
  9641=>"001110100",
  9642=>"000000100",
  9643=>"111111111",
  9644=>"111111010",
  9645=>"000001000",
  9646=>"110001110",
  9647=>"110011101",
  9648=>"001110101",
  9649=>"100000101",
  9650=>"101110000",
  9651=>"101111000",
  9652=>"000011010",
  9653=>"100001111",
  9654=>"100110110",
  9655=>"001001100",
  9656=>"100101011",
  9657=>"111011111",
  9658=>"011111011",
  9659=>"100001111",
  9660=>"010111001",
  9661=>"110011101",
  9662=>"101010010",
  9663=>"011110100",
  9664=>"110011111",
  9665=>"111101010",
  9666=>"010011010",
  9667=>"101001000",
  9668=>"010111000",
  9669=>"111100000",
  9670=>"110111011",
  9671=>"101010111",
  9672=>"011000100",
  9673=>"001101101",
  9674=>"001111111",
  9675=>"101001010",
  9676=>"111011101",
  9677=>"110101010",
  9678=>"111111101",
  9679=>"000000100",
  9680=>"100000010",
  9681=>"010011100",
  9682=>"111100111",
  9683=>"011000000",
  9684=>"100001011",
  9685=>"011111111",
  9686=>"101010010",
  9687=>"111011110",
  9688=>"010111100",
  9689=>"011000011",
  9690=>"001001000",
  9691=>"011000100",
  9692=>"010000011",
  9693=>"101011100",
  9694=>"100100110",
  9695=>"111000100",
  9696=>"111000101",
  9697=>"100110011",
  9698=>"000000100",
  9699=>"010001000",
  9700=>"001001110",
  9701=>"100110001",
  9702=>"110000011",
  9703=>"010001111",
  9704=>"001101111",
  9705=>"011011011",
  9706=>"001110100",
  9707=>"011101011",
  9708=>"111111010",
  9709=>"100100011",
  9710=>"010000010",
  9711=>"000001110",
  9712=>"010110101",
  9713=>"011011001",
  9714=>"011011111",
  9715=>"010100011",
  9716=>"111100100",
  9717=>"101110011",
  9718=>"101000100",
  9719=>"010011110",
  9720=>"101001110",
  9721=>"110110011",
  9722=>"110110111",
  9723=>"101001001",
  9724=>"101100011",
  9725=>"111111000",
  9726=>"000101001",
  9727=>"010001111",
  9728=>"001110011",
  9729=>"101001100",
  9730=>"110101000",
  9731=>"000100001",
  9732=>"011101110",
  9733=>"110110011",
  9734=>"101000010",
  9735=>"000001000",
  9736=>"111111111",
  9737=>"110010011",
  9738=>"001111110",
  9739=>"101111111",
  9740=>"101011000",
  9741=>"010111001",
  9742=>"101011011",
  9743=>"010000101",
  9744=>"010111110",
  9745=>"011011111",
  9746=>"101101111",
  9747=>"111101010",
  9748=>"101111110",
  9749=>"011000010",
  9750=>"011111111",
  9751=>"010001001",
  9752=>"000011010",
  9753=>"000101001",
  9754=>"111111100",
  9755=>"011111110",
  9756=>"101011000",
  9757=>"010010101",
  9758=>"001100010",
  9759=>"111110101",
  9760=>"101100000",
  9761=>"000011010",
  9762=>"110110010",
  9763=>"100110110",
  9764=>"101011010",
  9765=>"011101111",
  9766=>"100101001",
  9767=>"010111111",
  9768=>"000001010",
  9769=>"011100000",
  9770=>"001110011",
  9771=>"110001101",
  9772=>"001110111",
  9773=>"111000110",
  9774=>"101111111",
  9775=>"110001110",
  9776=>"011101101",
  9777=>"011010101",
  9778=>"100010011",
  9779=>"110010101",
  9780=>"111101101",
  9781=>"101011111",
  9782=>"001110011",
  9783=>"110100110",
  9784=>"100011000",
  9785=>"000000100",
  9786=>"001101000",
  9787=>"011110010",
  9788=>"110100101",
  9789=>"001101001",
  9790=>"111111101",
  9791=>"100111011",
  9792=>"011111111",
  9793=>"110010011",
  9794=>"110111000",
  9795=>"101010000",
  9796=>"011011001",
  9797=>"111111110",
  9798=>"111001011",
  9799=>"111110111",
  9800=>"111011110",
  9801=>"000111001",
  9802=>"000110001",
  9803=>"101011110",
  9804=>"001001011",
  9805=>"110101111",
  9806=>"000010010",
  9807=>"000000111",
  9808=>"000010010",
  9809=>"000110001",
  9810=>"001100111",
  9811=>"101011101",
  9812=>"101001001",
  9813=>"101110111",
  9814=>"100110011",
  9815=>"011010111",
  9816=>"001000111",
  9817=>"010111001",
  9818=>"111010111",
  9819=>"111101001",
  9820=>"001110111",
  9821=>"111111001",
  9822=>"111110000",
  9823=>"110100100",
  9824=>"001110100",
  9825=>"000110000",
  9826=>"110010000",
  9827=>"110111011",
  9828=>"001010011",
  9829=>"100111010",
  9830=>"011100011",
  9831=>"100101011",
  9832=>"111011011",
  9833=>"111100111",
  9834=>"010000111",
  9835=>"001110000",
  9836=>"111101110",
  9837=>"001110001",
  9838=>"111101010",
  9839=>"001000010",
  9840=>"110011111",
  9841=>"111111011",
  9842=>"001010011",
  9843=>"110010010",
  9844=>"101010001",
  9845=>"101101111",
  9846=>"110010111",
  9847=>"110101010",
  9848=>"111111110",
  9849=>"101101010",
  9850=>"000001000",
  9851=>"011111011",
  9852=>"111011110",
  9853=>"110101110",
  9854=>"010110101",
  9855=>"011101010",
  9856=>"001000000",
  9857=>"011001000",
  9858=>"111100010",
  9859=>"111000010",
  9860=>"111011001",
  9861=>"110001111",
  9862=>"101001001",
  9863=>"000011101",
  9864=>"001010000",
  9865=>"101100110",
  9866=>"000101111",
  9867=>"111000001",
  9868=>"100100010",
  9869=>"001100000",
  9870=>"100111111",
  9871=>"101101111",
  9872=>"111100010",
  9873=>"111011001",
  9874=>"010001111",
  9875=>"101100001",
  9876=>"111111010",
  9877=>"100000100",
  9878=>"000001111",
  9879=>"101001111",
  9880=>"000000001",
  9881=>"101010110",
  9882=>"010011111",
  9883=>"001110001",
  9884=>"001011000",
  9885=>"010100100",
  9886=>"110100011",
  9887=>"000110010",
  9888=>"010000111",
  9889=>"111001011",
  9890=>"111001010",
  9891=>"100010110",
  9892=>"110101000",
  9893=>"100111011",
  9894=>"111110111",
  9895=>"101000010",
  9896=>"011010001",
  9897=>"011000011",
  9898=>"000010010",
  9899=>"100000101",
  9900=>"011110111",
  9901=>"010101111",
  9902=>"010100101",
  9903=>"101101110",
  9904=>"111110111",
  9905=>"010011111",
  9906=>"000100100",
  9907=>"010101111",
  9908=>"011110100",
  9909=>"011000011",
  9910=>"101100000",
  9911=>"000100011",
  9912=>"111111101",
  9913=>"000111110",
  9914=>"101101001",
  9915=>"011101101",
  9916=>"011110111",
  9917=>"000100011",
  9918=>"101111000",
  9919=>"111110110",
  9920=>"001000101",
  9921=>"011001010",
  9922=>"110011111",
  9923=>"001010001",
  9924=>"101010111",
  9925=>"110100100",
  9926=>"001000011",
  9927=>"001001001",
  9928=>"001001101",
  9929=>"110101010",
  9930=>"100011111",
  9931=>"101111010",
  9932=>"101110011",
  9933=>"110100000",
  9934=>"000101100",
  9935=>"111111001",
  9936=>"000000101",
  9937=>"001110010",
  9938=>"101111110",
  9939=>"010001111",
  9940=>"110100111",
  9941=>"111111001",
  9942=>"010100000",
  9943=>"101101111",
  9944=>"001111000",
  9945=>"000011100",
  9946=>"100000100",
  9947=>"000000011",
  9948=>"110100110",
  9949=>"111111010",
  9950=>"111011101",
  9951=>"101000100",
  9952=>"011011110",
  9953=>"011111100",
  9954=>"000001011",
  9955=>"011111011",
  9956=>"110110111",
  9957=>"101111011",
  9958=>"101111110",
  9959=>"111110111",
  9960=>"111101011",
  9961=>"100000111",
  9962=>"010000011",
  9963=>"001010100",
  9964=>"111011010",
  9965=>"111110100",
  9966=>"000100000",
  9967=>"101001000",
  9968=>"011001000",
  9969=>"111101100",
  9970=>"010011011",
  9971=>"100111111",
  9972=>"001100111",
  9973=>"011101111",
  9974=>"111101100",
  9975=>"110001001",
  9976=>"010010001",
  9977=>"100000110",
  9978=>"011101011",
  9979=>"111110011",
  9980=>"111100010",
  9981=>"010011110",
  9982=>"110011100",
  9983=>"010111110",
  9984=>"110111000",
  9985=>"001000010",
  9986=>"010111100",
  9987=>"111111101",
  9988=>"101001110",
  9989=>"110111111",
  9990=>"010100000",
  9991=>"011101100",
  9992=>"100111100",
  9993=>"100010001",
  9994=>"110010110",
  9995=>"111111111",
  9996=>"000110001",
  9997=>"001000000",
  9998=>"110101010",
  9999=>"011000001",
  10000=>"001111111",
  10001=>"111111110",
  10002=>"000111010",
  10003=>"000001001",
  10004=>"100011000",
  10005=>"011010001",
  10006=>"000010011",
  10007=>"010100111",
  10008=>"000101100",
  10009=>"110011110",
  10010=>"111111110",
  10011=>"010100011",
  10012=>"110011101",
  10013=>"010000001",
  10014=>"101001111",
  10015=>"001001010",
  10016=>"100001110",
  10017=>"001111111",
  10018=>"001100101",
  10019=>"100001110",
  10020=>"110010110",
  10021=>"110110000",
  10022=>"111100011",
  10023=>"101000000",
  10024=>"101110111",
  10025=>"100011001",
  10026=>"000001010",
  10027=>"001111000",
  10028=>"100001100",
  10029=>"111111101",
  10030=>"101111111",
  10031=>"101010110",
  10032=>"011111111",
  10033=>"011111111",
  10034=>"101000001",
  10035=>"010000110",
  10036=>"100000000",
  10037=>"000111111",
  10038=>"110100110",
  10039=>"010111111",
  10040=>"000110101",
  10041=>"110110101",
  10042=>"110011010",
  10043=>"101110101",
  10044=>"010110011",
  10045=>"110110110",
  10046=>"000001011",
  10047=>"010011000",
  10048=>"100101101",
  10049=>"110001000",
  10050=>"010011101",
  10051=>"000100001",
  10052=>"011111110",
  10053=>"000110010",
  10054=>"100001100",
  10055=>"110110100",
  10056=>"110010111",
  10057=>"111101101",
  10058=>"110101001",
  10059=>"110111010",
  10060=>"111101100",
  10061=>"010101000",
  10062=>"000110100",
  10063=>"110101100",
  10064=>"000100101",
  10065=>"111100001",
  10066=>"001110100",
  10067=>"001000101",
  10068=>"111000010",
  10069=>"000111000",
  10070=>"111001111",
  10071=>"110110100",
  10072=>"100000111",
  10073=>"001110011",
  10074=>"110000100",
  10075=>"110110011",
  10076=>"010101011",
  10077=>"011101001",
  10078=>"000110110",
  10079=>"111111111",
  10080=>"110111011",
  10081=>"000000110",
  10082=>"111111010",
  10083=>"111001001",
  10084=>"000001001",
  10085=>"100001011",
  10086=>"110011110",
  10087=>"110001001",
  10088=>"110110110",
  10089=>"010001001",
  10090=>"011101001",
  10091=>"011100011",
  10092=>"000111101",
  10093=>"101111001",
  10094=>"110111111",
  10095=>"111101101",
  10096=>"110011101",
  10097=>"110011011",
  10098=>"000100001",
  10099=>"111101110",
  10100=>"001111101",
  10101=>"110011111",
  10102=>"100111000",
  10103=>"111011001",
  10104=>"100011010",
  10105=>"111101110",
  10106=>"101100011",
  10107=>"010111010",
  10108=>"101110101",
  10109=>"000011111",
  10110=>"100101101",
  10111=>"000001010",
  10112=>"100000010",
  10113=>"011101110",
  10114=>"111111001",
  10115=>"110101000",
  10116=>"010011111",
  10117=>"100101111",
  10118=>"011110110",
  10119=>"110110110",
  10120=>"011100011",
  10121=>"111000001",
  10122=>"101001000",
  10123=>"100000001",
  10124=>"101000110",
  10125=>"011001010",
  10126=>"101011110",
  10127=>"110101011",
  10128=>"101110101",
  10129=>"111001011",
  10130=>"101000111",
  10131=>"101100000",
  10132=>"010000010",
  10133=>"010110101",
  10134=>"001011110",
  10135=>"010011100",
  10136=>"110101101",
  10137=>"010011111",
  10138=>"001011110",
  10139=>"111111111",
  10140=>"111000100",
  10141=>"101111100",
  10142=>"110101001",
  10143=>"100010011",
  10144=>"101010011",
  10145=>"111101100",
  10146=>"000100010",
  10147=>"001100110",
  10148=>"111111110",
  10149=>"001110101",
  10150=>"111100010",
  10151=>"111011010",
  10152=>"101010001",
  10153=>"111110010",
  10154=>"000000101",
  10155=>"001000010",
  10156=>"011100010",
  10157=>"001100000",
  10158=>"011001100",
  10159=>"111101110",
  10160=>"101000001",
  10161=>"101100011",
  10162=>"010101001",
  10163=>"011011010",
  10164=>"001101000",
  10165=>"101110111",
  10166=>"011001001",
  10167=>"011011111",
  10168=>"010111001",
  10169=>"001011101",
  10170=>"100001110",
  10171=>"001110001",
  10172=>"100000010",
  10173=>"100101000",
  10174=>"000100000",
  10175=>"100100101",
  10176=>"101000000",
  10177=>"001111100",
  10178=>"011111101",
  10179=>"111110011",
  10180=>"001000001",
  10181=>"011011101",
  10182=>"010001011",
  10183=>"000101011",
  10184=>"111111111",
  10185=>"111010011",
  10186=>"001101001",
  10187=>"100101100",
  10188=>"100011111",
  10189=>"111111110",
  10190=>"011111011",
  10191=>"100010001",
  10192=>"011100101",
  10193=>"011011100",
  10194=>"110001010",
  10195=>"101101001",
  10196=>"011100001",
  10197=>"100000111",
  10198=>"010101011",
  10199=>"100010000",
  10200=>"111111100",
  10201=>"010111001",
  10202=>"000001010",
  10203=>"100100111",
  10204=>"000101100",
  10205=>"011100000",
  10206=>"010101101",
  10207=>"111111101",
  10208=>"101101101",
  10209=>"110010100",
  10210=>"001001110",
  10211=>"000110011",
  10212=>"011111111",
  10213=>"001100111",
  10214=>"101100101",
  10215=>"101111100",
  10216=>"101111100",
  10217=>"111110100",
  10218=>"100101110",
  10219=>"001101000",
  10220=>"111010000",
  10221=>"001011111",
  10222=>"000111101",
  10223=>"101001101",
  10224=>"100010110",
  10225=>"001111000",
  10226=>"111101001",
  10227=>"010111010",
  10228=>"011110010",
  10229=>"101010000",
  10230=>"010110010",
  10231=>"010001011",
  10232=>"111011111",
  10233=>"101001011",
  10234=>"111110111",
  10235=>"001110011",
  10236=>"001001101",
  10237=>"011110001",
  10238=>"101011001",
  10239=>"111110011",
  10240=>"100101000",
  10241=>"111001000",
  10242=>"010110100",
  10243=>"101000000",
  10244=>"001110010",
  10245=>"101100010",
  10246=>"100001000",
  10247=>"010111000",
  10248=>"010010010",
  10249=>"010010100",
  10250=>"101111101",
  10251=>"001100111",
  10252=>"010000100",
  10253=>"001110101",
  10254=>"010101010",
  10255=>"111111010",
  10256=>"100001110",
  10257=>"101000100",
  10258=>"100101001",
  10259=>"010000101",
  10260=>"111111000",
  10261=>"100011000",
  10262=>"010001111",
  10263=>"111011100",
  10264=>"110100010",
  10265=>"000010110",
  10266=>"001000111",
  10267=>"111100001",
  10268=>"100111010",
  10269=>"101110010",
  10270=>"110001101",
  10271=>"011000101",
  10272=>"001010101",
  10273=>"010101111",
  10274=>"010011000",
  10275=>"110111011",
  10276=>"011111000",
  10277=>"010000110",
  10278=>"110111100",
  10279=>"100011011",
  10280=>"111001100",
  10281=>"111001000",
  10282=>"100011110",
  10283=>"001001101",
  10284=>"111110010",
  10285=>"000010101",
  10286=>"001111011",
  10287=>"111001001",
  10288=>"101101011",
  10289=>"001100010",
  10290=>"001011000",
  10291=>"011111111",
  10292=>"010010110",
  10293=>"001010110",
  10294=>"111111010",
  10295=>"100101001",
  10296=>"000001001",
  10297=>"100100000",
  10298=>"101000001",
  10299=>"111011111",
  10300=>"001101001",
  10301=>"001000000",
  10302=>"111000101",
  10303=>"100000010",
  10304=>"000111011",
  10305=>"000100110",
  10306=>"111000110",
  10307=>"000100101",
  10308=>"111000100",
  10309=>"110001111",
  10310=>"011001111",
  10311=>"010011111",
  10312=>"011111111",
  10313=>"011010100",
  10314=>"010011000",
  10315=>"110001010",
  10316=>"001110111",
  10317=>"000101101",
  10318=>"111011100",
  10319=>"011010111",
  10320=>"110110101",
  10321=>"100100100",
  10322=>"110100001",
  10323=>"010001000",
  10324=>"101110010",
  10325=>"001100010",
  10326=>"000010011",
  10327=>"001100000",
  10328=>"101110010",
  10329=>"111100011",
  10330=>"111110100",
  10331=>"111101100",
  10332=>"101001000",
  10333=>"001000101",
  10334=>"101000001",
  10335=>"100011000",
  10336=>"100000101",
  10337=>"010111111",
  10338=>"010010000",
  10339=>"000001001",
  10340=>"011010011",
  10341=>"011010010",
  10342=>"111111111",
  10343=>"001111011",
  10344=>"101101100",
  10345=>"011101011",
  10346=>"101000010",
  10347=>"101110101",
  10348=>"101001001",
  10349=>"100010001",
  10350=>"101111000",
  10351=>"101001000",
  10352=>"110000111",
  10353=>"010000000",
  10354=>"111000010",
  10355=>"111110001",
  10356=>"010000001",
  10357=>"000001010",
  10358=>"011011111",
  10359=>"011111001",
  10360=>"000011000",
  10361=>"000100011",
  10362=>"010111111",
  10363=>"100110000",
  10364=>"100101000",
  10365=>"010111010",
  10366=>"001100010",
  10367=>"010011010",
  10368=>"011110110",
  10369=>"011111111",
  10370=>"011001100",
  10371=>"000001111",
  10372=>"100010101",
  10373=>"111111100",
  10374=>"010100111",
  10375=>"001100001",
  10376=>"000011111",
  10377=>"101111100",
  10378=>"011101010",
  10379=>"111001101",
  10380=>"110001000",
  10381=>"110100000",
  10382=>"111101011",
  10383=>"110111100",
  10384=>"101100011",
  10385=>"001010001",
  10386=>"001001000",
  10387=>"000011011",
  10388=>"111111011",
  10389=>"101101001",
  10390=>"100001111",
  10391=>"000011101",
  10392=>"000000011",
  10393=>"001101000",
  10394=>"100100100",
  10395=>"011001011",
  10396=>"001100001",
  10397=>"001100111",
  10398=>"101011100",
  10399=>"011000000",
  10400=>"000011000",
  10401=>"010111111",
  10402=>"011100111",
  10403=>"011110000",
  10404=>"010000111",
  10405=>"000100110",
  10406=>"101000000",
  10407=>"110101111",
  10408=>"101110011",
  10409=>"001010000",
  10410=>"110001000",
  10411=>"010111000",
  10412=>"111110010",
  10413=>"101011101",
  10414=>"001111101",
  10415=>"010011011",
  10416=>"000010010",
  10417=>"000011000",
  10418=>"011011000",
  10419=>"010000110",
  10420=>"001110000",
  10421=>"000010000",
  10422=>"110010100",
  10423=>"101110100",
  10424=>"011010100",
  10425=>"110101010",
  10426=>"001111000",
  10427=>"101100001",
  10428=>"010001001",
  10429=>"010101011",
  10430=>"011111000",
  10431=>"000010001",
  10432=>"010011001",
  10433=>"010100111",
  10434=>"001000011",
  10435=>"000011011",
  10436=>"100111010",
  10437=>"101011010",
  10438=>"010010010",
  10439=>"000100011",
  10440=>"101011101",
  10441=>"100000011",
  10442=>"001110100",
  10443=>"110110000",
  10444=>"000000000",
  10445=>"100110100",
  10446=>"101100010",
  10447=>"110111111",
  10448=>"011100110",
  10449=>"111101001",
  10450=>"100110100",
  10451=>"000111110",
  10452=>"100101001",
  10453=>"101110001",
  10454=>"100011110",
  10455=>"000000011",
  10456=>"101100011",
  10457=>"100101101",
  10458=>"100110111",
  10459=>"000101111",
  10460=>"101010100",
  10461=>"100000110",
  10462=>"010110011",
  10463=>"110101000",
  10464=>"000011001",
  10465=>"101000010",
  10466=>"100011100",
  10467=>"000110100",
  10468=>"100000011",
  10469=>"001111001",
  10470=>"010101101",
  10471=>"101010001",
  10472=>"101111000",
  10473=>"011001010",
  10474=>"000100101",
  10475=>"100111010",
  10476=>"001100101",
  10477=>"111110101",
  10478=>"110110110",
  10479=>"001001100",
  10480=>"000111000",
  10481=>"001100110",
  10482=>"101011100",
  10483=>"010010100",
  10484=>"110011111",
  10485=>"000000011",
  10486=>"101111000",
  10487=>"100111011",
  10488=>"010001000",
  10489=>"000000000",
  10490=>"110100100",
  10491=>"010111011",
  10492=>"100101010",
  10493=>"010111100",
  10494=>"000011011",
  10495=>"010001101",
  10496=>"110100111",
  10497=>"100111111",
  10498=>"100001010",
  10499=>"001010000",
  10500=>"101110111",
  10501=>"001001000",
  10502=>"111000111",
  10503=>"101110111",
  10504=>"101111110",
  10505=>"101010001",
  10506=>"010100101",
  10507=>"101101011",
  10508=>"011001001",
  10509=>"101111110",
  10510=>"000000100",
  10511=>"101000100",
  10512=>"111110000",
  10513=>"101100000",
  10514=>"111001100",
  10515=>"111000110",
  10516=>"111111000",
  10517=>"111001101",
  10518=>"111110010",
  10519=>"011111000",
  10520=>"011011100",
  10521=>"000110111",
  10522=>"111000010",
  10523=>"010000101",
  10524=>"100010001",
  10525=>"011010100",
  10526=>"011011100",
  10527=>"011001001",
  10528=>"000011001",
  10529=>"100111111",
  10530=>"111111010",
  10531=>"010111111",
  10532=>"111001010",
  10533=>"110101000",
  10534=>"010011011",
  10535=>"101010010",
  10536=>"100001000",
  10537=>"110011001",
  10538=>"000001110",
  10539=>"110010000",
  10540=>"101101010",
  10541=>"010001100",
  10542=>"011111011",
  10543=>"111111110",
  10544=>"011101101",
  10545=>"010000001",
  10546=>"111101000",
  10547=>"011001000",
  10548=>"110100101",
  10549=>"101100010",
  10550=>"110000000",
  10551=>"011001101",
  10552=>"110111111",
  10553=>"010110000",
  10554=>"101100111",
  10555=>"101000010",
  10556=>"010001101",
  10557=>"100011101",
  10558=>"100010111",
  10559=>"110000101",
  10560=>"001000001",
  10561=>"100101000",
  10562=>"101001001",
  10563=>"010111001",
  10564=>"100100000",
  10565=>"101011001",
  10566=>"000011101",
  10567=>"011100101",
  10568=>"011011111",
  10569=>"111110111",
  10570=>"001101100",
  10571=>"001100111",
  10572=>"110001000",
  10573=>"011100110",
  10574=>"011100000",
  10575=>"010101110",
  10576=>"010111111",
  10577=>"101000010",
  10578=>"001000111",
  10579=>"010011010",
  10580=>"000000101",
  10581=>"011011100",
  10582=>"001101010",
  10583=>"100011011",
  10584=>"110111111",
  10585=>"010000001",
  10586=>"001110101",
  10587=>"011010000",
  10588=>"010000010",
  10589=>"100100010",
  10590=>"111100011",
  10591=>"110100001",
  10592=>"010100111",
  10593=>"001111101",
  10594=>"010101101",
  10595=>"101010011",
  10596=>"100011101",
  10597=>"001000010",
  10598=>"000101001",
  10599=>"010101000",
  10600=>"100011111",
  10601=>"011100000",
  10602=>"100011101",
  10603=>"000000111",
  10604=>"001011011",
  10605=>"001000111",
  10606=>"000000000",
  10607=>"110100010",
  10608=>"010010100",
  10609=>"011001000",
  10610=>"010110111",
  10611=>"001110100",
  10612=>"100000111",
  10613=>"101011101",
  10614=>"010111110",
  10615=>"101000101",
  10616=>"001101100",
  10617=>"101010111",
  10618=>"111110100",
  10619=>"110011111",
  10620=>"100111000",
  10621=>"011001001",
  10622=>"110110110",
  10623=>"010000100",
  10624=>"000110011",
  10625=>"001111010",
  10626=>"100100101",
  10627=>"001100011",
  10628=>"010111100",
  10629=>"011101110",
  10630=>"111001010",
  10631=>"010101010",
  10632=>"110101111",
  10633=>"001101111",
  10634=>"111101111",
  10635=>"000010110",
  10636=>"100011011",
  10637=>"111001011",
  10638=>"111011000",
  10639=>"111001011",
  10640=>"101100010",
  10641=>"100101000",
  10642=>"110111010",
  10643=>"001010011",
  10644=>"110110101",
  10645=>"011101110",
  10646=>"100010110",
  10647=>"101011000",
  10648=>"101110101",
  10649=>"001010011",
  10650=>"111111111",
  10651=>"000001010",
  10652=>"011101100",
  10653=>"100001100",
  10654=>"011011111",
  10655=>"001000111",
  10656=>"100101100",
  10657=>"000111001",
  10658=>"010110101",
  10659=>"001010110",
  10660=>"111001001",
  10661=>"111100000",
  10662=>"101111000",
  10663=>"000001000",
  10664=>"000110011",
  10665=>"110110110",
  10666=>"011101101",
  10667=>"110011001",
  10668=>"111001101",
  10669=>"110100010",
  10670=>"110110011",
  10671=>"010011101",
  10672=>"111100110",
  10673=>"110011000",
  10674=>"100110010",
  10675=>"110001111",
  10676=>"110010010",
  10677=>"001100000",
  10678=>"100110100",
  10679=>"011010000",
  10680=>"111010110",
  10681=>"000100010",
  10682=>"011001001",
  10683=>"111011111",
  10684=>"101010010",
  10685=>"100101010",
  10686=>"100100001",
  10687=>"000011111",
  10688=>"100010001",
  10689=>"010001101",
  10690=>"110110100",
  10691=>"100000100",
  10692=>"001110001",
  10693=>"010011001",
  10694=>"000110000",
  10695=>"000101010",
  10696=>"101101011",
  10697=>"011101101",
  10698=>"000010110",
  10699=>"010111011",
  10700=>"111110011",
  10701=>"011110110",
  10702=>"101001000",
  10703=>"101101010",
  10704=>"000101100",
  10705=>"010011100",
  10706=>"010101001",
  10707=>"100011011",
  10708=>"101011111",
  10709=>"001010101",
  10710=>"011010011",
  10711=>"001000001",
  10712=>"100101111",
  10713=>"110111011",
  10714=>"110100000",
  10715=>"001101000",
  10716=>"010111000",
  10717=>"110000110",
  10718=>"110011110",
  10719=>"110010011",
  10720=>"110001110",
  10721=>"001001011",
  10722=>"100101000",
  10723=>"000001000",
  10724=>"011000011",
  10725=>"110011111",
  10726=>"010001001",
  10727=>"110111110",
  10728=>"111011001",
  10729=>"010100100",
  10730=>"101000001",
  10731=>"111010001",
  10732=>"011111111",
  10733=>"101010100",
  10734=>"011101110",
  10735=>"100101101",
  10736=>"110011001",
  10737=>"001001100",
  10738=>"001000100",
  10739=>"101111010",
  10740=>"000001111",
  10741=>"011111100",
  10742=>"101000111",
  10743=>"101001111",
  10744=>"110000011",
  10745=>"111011111",
  10746=>"110100001",
  10747=>"001110011",
  10748=>"111000111",
  10749=>"000101010",
  10750=>"000001000",
  10751=>"110011011",
  10752=>"100011001",
  10753=>"111100011",
  10754=>"000011111",
  10755=>"110001001",
  10756=>"011010111",
  10757=>"000101010",
  10758=>"000011110",
  10759=>"001010111",
  10760=>"100001001",
  10761=>"110011000",
  10762=>"000010111",
  10763=>"010011110",
  10764=>"000001001",
  10765=>"010111101",
  10766=>"000010011",
  10767=>"000010111",
  10768=>"011011111",
  10769=>"101010101",
  10770=>"000110100",
  10771=>"010001111",
  10772=>"111000010",
  10773=>"010011001",
  10774=>"101010111",
  10775=>"010011010",
  10776=>"101011010",
  10777=>"010010100",
  10778=>"001101011",
  10779=>"100011000",
  10780=>"110101111",
  10781=>"101111101",
  10782=>"000100000",
  10783=>"000010010",
  10784=>"001100111",
  10785=>"011100100",
  10786=>"000001111",
  10787=>"000001101",
  10788=>"111010011",
  10789=>"000001000",
  10790=>"011101010",
  10791=>"100111001",
  10792=>"100000101",
  10793=>"001101100",
  10794=>"101111011",
  10795=>"100000001",
  10796=>"100110111",
  10797=>"101111011",
  10798=>"000010001",
  10799=>"011001001",
  10800=>"010110000",
  10801=>"011011001",
  10802=>"100001100",
  10803=>"011011010",
  10804=>"110111111",
  10805=>"101100110",
  10806=>"001001011",
  10807=>"001010111",
  10808=>"101001101",
  10809=>"011101110",
  10810=>"101100111",
  10811=>"111100011",
  10812=>"101111001",
  10813=>"000101010",
  10814=>"001011101",
  10815=>"100001011",
  10816=>"101101011",
  10817=>"111100100",
  10818=>"000001110",
  10819=>"111010000",
  10820=>"001100101",
  10821=>"101111001",
  10822=>"110011000",
  10823=>"001011100",
  10824=>"111110101",
  10825=>"101101101",
  10826=>"101000001",
  10827=>"000010011",
  10828=>"001011011",
  10829=>"011110110",
  10830=>"001000001",
  10831=>"001001101",
  10832=>"000011000",
  10833=>"000111011",
  10834=>"011000110",
  10835=>"011000010",
  10836=>"111001011",
  10837=>"111101001",
  10838=>"111111100",
  10839=>"111001100",
  10840=>"001001011",
  10841=>"111001101",
  10842=>"111110110",
  10843=>"000100001",
  10844=>"001100111",
  10845=>"000110010",
  10846=>"001100001",
  10847=>"011110000",
  10848=>"101100001",
  10849=>"111101100",
  10850=>"001100111",
  10851=>"100011111",
  10852=>"001010111",
  10853=>"001010010",
  10854=>"010000110",
  10855=>"101001011",
  10856=>"000101010",
  10857=>"110101110",
  10858=>"111011101",
  10859=>"110100101",
  10860=>"110100011",
  10861=>"010010111",
  10862=>"010000010",
  10863=>"001110011",
  10864=>"101000001",
  10865=>"011000101",
  10866=>"100011100",
  10867=>"110100000",
  10868=>"111010011",
  10869=>"010100000",
  10870=>"111011111",
  10871=>"111101000",
  10872=>"111010010",
  10873=>"111011100",
  10874=>"110011111",
  10875=>"110001110",
  10876=>"110000101",
  10877=>"110011000",
  10878=>"111101110",
  10879=>"000110100",
  10880=>"110100101",
  10881=>"111101100",
  10882=>"011100110",
  10883=>"000101010",
  10884=>"111000001",
  10885=>"011001001",
  10886=>"000011110",
  10887=>"110100011",
  10888=>"001001110",
  10889=>"010001010",
  10890=>"001111111",
  10891=>"011001000",
  10892=>"100011110",
  10893=>"000010000",
  10894=>"010000000",
  10895=>"101001001",
  10896=>"011011000",
  10897=>"100100000",
  10898=>"000100111",
  10899=>"111010100",
  10900=>"011110010",
  10901=>"000111010",
  10902=>"101011001",
  10903=>"111001001",
  10904=>"100011011",
  10905=>"100101011",
  10906=>"010101000",
  10907=>"000111100",
  10908=>"001001111",
  10909=>"100000010",
  10910=>"001100010",
  10911=>"110000100",
  10912=>"000011101",
  10913=>"111011101",
  10914=>"101001001",
  10915=>"100010001",
  10916=>"011110110",
  10917=>"101101100",
  10918=>"011100100",
  10919=>"100111100",
  10920=>"101110011",
  10921=>"001110010",
  10922=>"110101101",
  10923=>"011100100",
  10924=>"001000000",
  10925=>"001011000",
  10926=>"010101101",
  10927=>"110010001",
  10928=>"001100001",
  10929=>"011001111",
  10930=>"100000100",
  10931=>"000101100",
  10932=>"001001011",
  10933=>"011011011",
  10934=>"011000101",
  10935=>"011101110",
  10936=>"101111010",
  10937=>"111110001",
  10938=>"110001110",
  10939=>"010001010",
  10940=>"001010100",
  10941=>"010001010",
  10942=>"000111100",
  10943=>"010010011",
  10944=>"000110110",
  10945=>"111100111",
  10946=>"000110101",
  10947=>"100101010",
  10948=>"010001001",
  10949=>"111111100",
  10950=>"010011000",
  10951=>"110011100",
  10952=>"010110111",
  10953=>"001111010",
  10954=>"100111110",
  10955=>"100111000",
  10956=>"000110101",
  10957=>"000111111",
  10958=>"111100011",
  10959=>"110000001",
  10960=>"000001101",
  10961=>"100101011",
  10962=>"011111011",
  10963=>"001011010",
  10964=>"111010100",
  10965=>"010010111",
  10966=>"010110100",
  10967=>"001110111",
  10968=>"000010110",
  10969=>"111010100",
  10970=>"000001010",
  10971=>"100111101",
  10972=>"011001110",
  10973=>"010001010",
  10974=>"001111111",
  10975=>"001011000",
  10976=>"010011100",
  10977=>"101100110",
  10978=>"011110100",
  10979=>"010111111",
  10980=>"111100101",
  10981=>"111110001",
  10982=>"101110111",
  10983=>"111100101",
  10984=>"011111110",
  10985=>"100101011",
  10986=>"110111010",
  10987=>"010110010",
  10988=>"001000110",
  10989=>"000001011",
  10990=>"001010100",
  10991=>"010001011",
  10992=>"001011011",
  10993=>"001100101",
  10994=>"111010100",
  10995=>"101100001",
  10996=>"011010111",
  10997=>"001000001",
  10998=>"011111010",
  10999=>"001000001",
  11000=>"010001001",
  11001=>"001111000",
  11002=>"010010001",
  11003=>"001001111",
  11004=>"011100100",
  11005=>"111000011",
  11006=>"111010100",
  11007=>"001111110",
  11008=>"011011111",
  11009=>"100101101",
  11010=>"101100100",
  11011=>"111010101",
  11012=>"001111011",
  11013=>"100100101",
  11014=>"100011101",
  11015=>"011000101",
  11016=>"111101101",
  11017=>"011110111",
  11018=>"011101100",
  11019=>"101101010",
  11020=>"011011100",
  11021=>"100101100",
  11022=>"100001101",
  11023=>"000111110",
  11024=>"000001001",
  11025=>"000001100",
  11026=>"110001100",
  11027=>"111001100",
  11028=>"110001000",
  11029=>"000001000",
  11030=>"000100100",
  11031=>"001011101",
  11032=>"110111101",
  11033=>"110111001",
  11034=>"111011101",
  11035=>"011001010",
  11036=>"010100001",
  11037=>"100000000",
  11038=>"001110111",
  11039=>"010011110",
  11040=>"010001101",
  11041=>"010110011",
  11042=>"000101001",
  11043=>"000011100",
  11044=>"001010000",
  11045=>"001110111",
  11046=>"100000110",
  11047=>"101100001",
  11048=>"100111111",
  11049=>"000101001",
  11050=>"110000001",
  11051=>"011100001",
  11052=>"110101011",
  11053=>"101111111",
  11054=>"110000000",
  11055=>"001101111",
  11056=>"011011010",
  11057=>"010010100",
  11058=>"000101011",
  11059=>"101111000",
  11060=>"000001001",
  11061=>"011110000",
  11062=>"010101111",
  11063=>"000011110",
  11064=>"101010111",
  11065=>"010110101",
  11066=>"001101011",
  11067=>"000000000",
  11068=>"001000110",
  11069=>"001010101",
  11070=>"111001110",
  11071=>"110100011",
  11072=>"011011011",
  11073=>"011100010",
  11074=>"010001110",
  11075=>"111100001",
  11076=>"000111100",
  11077=>"010111010",
  11078=>"101001101",
  11079=>"010111011",
  11080=>"011000110",
  11081=>"001100100",
  11082=>"100000011",
  11083=>"000000010",
  11084=>"100110111",
  11085=>"000111011",
  11086=>"001001010",
  11087=>"101110001",
  11088=>"001100101",
  11089=>"001100100",
  11090=>"010100000",
  11091=>"000010110",
  11092=>"001101100",
  11093=>"110000100",
  11094=>"111001101",
  11095=>"101001100",
  11096=>"100000111",
  11097=>"101001001",
  11098=>"110100011",
  11099=>"000100011",
  11100=>"101001001",
  11101=>"101101100",
  11102=>"111111110",
  11103=>"011001011",
  11104=>"100111001",
  11105=>"010011100",
  11106=>"100111000",
  11107=>"111001111",
  11108=>"000001001",
  11109=>"100111110",
  11110=>"010101011",
  11111=>"111100100",
  11112=>"001000010",
  11113=>"001111001",
  11114=>"111100000",
  11115=>"011101110",
  11116=>"101110111",
  11117=>"011000111",
  11118=>"001110001",
  11119=>"001010010",
  11120=>"001110111",
  11121=>"000111101",
  11122=>"110110100",
  11123=>"000011010",
  11124=>"010111000",
  11125=>"011111110",
  11126=>"000011101",
  11127=>"100000000",
  11128=>"100010101",
  11129=>"001000001",
  11130=>"001110110",
  11131=>"011010011",
  11132=>"111110000",
  11133=>"011011100",
  11134=>"110110011",
  11135=>"001110100",
  11136=>"101010111",
  11137=>"000101111",
  11138=>"010101110",
  11139=>"111010011",
  11140=>"010001000",
  11141=>"010100000",
  11142=>"111011110",
  11143=>"110100111",
  11144=>"110110011",
  11145=>"010010011",
  11146=>"000011101",
  11147=>"100010010",
  11148=>"101001110",
  11149=>"100101011",
  11150=>"101000100",
  11151=>"110110111",
  11152=>"010000011",
  11153=>"011111100",
  11154=>"101101010",
  11155=>"010111001",
  11156=>"110110100",
  11157=>"110011111",
  11158=>"111100111",
  11159=>"001000110",
  11160=>"110000101",
  11161=>"000110000",
  11162=>"100010010",
  11163=>"101100101",
  11164=>"000100000",
  11165=>"111111100",
  11166=>"110000011",
  11167=>"000010111",
  11168=>"011000110",
  11169=>"000111111",
  11170=>"000111001",
  11171=>"000101110",
  11172=>"100111001",
  11173=>"101101001",
  11174=>"001100101",
  11175=>"000111010",
  11176=>"010111011",
  11177=>"010110001",
  11178=>"010110111",
  11179=>"111110110",
  11180=>"010001011",
  11181=>"011011000",
  11182=>"001000100",
  11183=>"111111110",
  11184=>"101001000",
  11185=>"110011101",
  11186=>"010101101",
  11187=>"000011000",
  11188=>"111001001",
  11189=>"001011001",
  11190=>"110000110",
  11191=>"111111100",
  11192=>"111110101",
  11193=>"101101111",
  11194=>"111000100",
  11195=>"110110111",
  11196=>"110100011",
  11197=>"100101000",
  11198=>"100111010",
  11199=>"100100111",
  11200=>"110011101",
  11201=>"111001111",
  11202=>"000111101",
  11203=>"100000011",
  11204=>"101000000",
  11205=>"010111010",
  11206=>"000001010",
  11207=>"100000011",
  11208=>"010101101",
  11209=>"010110011",
  11210=>"101001000",
  11211=>"101111101",
  11212=>"100101000",
  11213=>"000000100",
  11214=>"111100000",
  11215=>"010010001",
  11216=>"010000100",
  11217=>"111000001",
  11218=>"101111110",
  11219=>"101001001",
  11220=>"100001100",
  11221=>"010001010",
  11222=>"110000011",
  11223=>"000111001",
  11224=>"101000011",
  11225=>"010000110",
  11226=>"101001001",
  11227=>"001100101",
  11228=>"110111101",
  11229=>"110110101",
  11230=>"111110110",
  11231=>"100000011",
  11232=>"000110010",
  11233=>"110000010",
  11234=>"011101000",
  11235=>"011101111",
  11236=>"111000000",
  11237=>"110101100",
  11238=>"101110010",
  11239=>"100101000",
  11240=>"111011101",
  11241=>"111100010",
  11242=>"011111011",
  11243=>"101011110",
  11244=>"001010001",
  11245=>"011101101",
  11246=>"100010011",
  11247=>"111011111",
  11248=>"000011011",
  11249=>"011001011",
  11250=>"101000100",
  11251=>"100000101",
  11252=>"001000111",
  11253=>"111101011",
  11254=>"010110100",
  11255=>"010100000",
  11256=>"000010101",
  11257=>"111000001",
  11258=>"100001010",
  11259=>"000110010",
  11260=>"111010100",
  11261=>"010001001",
  11262=>"010001010",
  11263=>"110100001",
  11264=>"100011110",
  11265=>"011111111",
  11266=>"001110110",
  11267=>"011010011",
  11268=>"101001100",
  11269=>"011110011",
  11270=>"000000111",
  11271=>"010111110",
  11272=>"001000001",
  11273=>"011000000",
  11274=>"101101000",
  11275=>"010110101",
  11276=>"000001111",
  11277=>"101010010",
  11278=>"100010001",
  11279=>"110101110",
  11280=>"001001001",
  11281=>"011001110",
  11282=>"111110101",
  11283=>"110101001",
  11284=>"111010101",
  11285=>"110110101",
  11286=>"101100100",
  11287=>"001110011",
  11288=>"101001100",
  11289=>"011110010",
  11290=>"000110101",
  11291=>"101110100",
  11292=>"001101101",
  11293=>"110000110",
  11294=>"101001011",
  11295=>"001110000",
  11296=>"010110110",
  11297=>"010111001",
  11298=>"101010000",
  11299=>"001101010",
  11300=>"110111001",
  11301=>"001100101",
  11302=>"011001011",
  11303=>"101111111",
  11304=>"110011001",
  11305=>"111100100",
  11306=>"110100011",
  11307=>"100110001",
  11308=>"000111010",
  11309=>"010001100",
  11310=>"111100000",
  11311=>"010010011",
  11312=>"001000110",
  11313=>"001100001",
  11314=>"000011110",
  11315=>"000000101",
  11316=>"011010001",
  11317=>"111000011",
  11318=>"001101000",
  11319=>"101000110",
  11320=>"011101010",
  11321=>"101001000",
  11322=>"101001011",
  11323=>"111110111",
  11324=>"000010001",
  11325=>"001001000",
  11326=>"110111101",
  11327=>"110000000",
  11328=>"100100010",
  11329=>"000001011",
  11330=>"001100101",
  11331=>"010110101",
  11332=>"011101001",
  11333=>"111110000",
  11334=>"100110101",
  11335=>"101101010",
  11336=>"011110001",
  11337=>"000101010",
  11338=>"001111110",
  11339=>"011010010",
  11340=>"101110100",
  11341=>"101111111",
  11342=>"100110010",
  11343=>"011101010",
  11344=>"001110111",
  11345=>"010001110",
  11346=>"101000111",
  11347=>"111100110",
  11348=>"100010100",
  11349=>"011100010",
  11350=>"101000000",
  11351=>"110101000",
  11352=>"001110011",
  11353=>"111111011",
  11354=>"111000001",
  11355=>"000000101",
  11356=>"011101011",
  11357=>"111100001",
  11358=>"110011110",
  11359=>"100001101",
  11360=>"111110001",
  11361=>"110110100",
  11362=>"000000110",
  11363=>"110101000",
  11364=>"001000100",
  11365=>"100001101",
  11366=>"111010001",
  11367=>"001010001",
  11368=>"111101110",
  11369=>"110100011",
  11370=>"001001001",
  11371=>"011100111",
  11372=>"010100001",
  11373=>"000101101",
  11374=>"000011111",
  11375=>"001011000",
  11376=>"101000100",
  11377=>"110001000",
  11378=>"101000001",
  11379=>"101010101",
  11380=>"100111010",
  11381=>"100011100",
  11382=>"101101111",
  11383=>"101001100",
  11384=>"110101001",
  11385=>"001000010",
  11386=>"110101011",
  11387=>"100011111",
  11388=>"000101001",
  11389=>"011100010",
  11390=>"001010001",
  11391=>"101111001",
  11392=>"110111101",
  11393=>"111101111",
  11394=>"111110001",
  11395=>"111010010",
  11396=>"100101110",
  11397=>"111101010",
  11398=>"011001111",
  11399=>"010111011",
  11400=>"101010100",
  11401=>"000100010",
  11402=>"011111001",
  11403=>"000100100",
  11404=>"011111000",
  11405=>"011111000",
  11406=>"111011010",
  11407=>"111110011",
  11408=>"010101011",
  11409=>"000111010",
  11410=>"010111101",
  11411=>"110110100",
  11412=>"101110111",
  11413=>"100010101",
  11414=>"010110001",
  11415=>"001100111",
  11416=>"110101011",
  11417=>"101111010",
  11418=>"000001001",
  11419=>"101000111",
  11420=>"101000000",
  11421=>"001110010",
  11422=>"100100010",
  11423=>"010001110",
  11424=>"100100110",
  11425=>"010110100",
  11426=>"101010111",
  11427=>"011111111",
  11428=>"100001010",
  11429=>"010111111",
  11430=>"011100001",
  11431=>"111010001",
  11432=>"101010111",
  11433=>"001000100",
  11434=>"100001001",
  11435=>"000010110",
  11436=>"001000001",
  11437=>"100011001",
  11438=>"000001011",
  11439=>"000100110",
  11440=>"011101000",
  11441=>"001011011",
  11442=>"111100001",
  11443=>"010100000",
  11444=>"101100011",
  11445=>"111110000",
  11446=>"111101110",
  11447=>"110001110",
  11448=>"001011110",
  11449=>"011101110",
  11450=>"100111111",
  11451=>"011101100",
  11452=>"010111011",
  11453=>"101000100",
  11454=>"011001011",
  11455=>"100000001",
  11456=>"011011110",
  11457=>"110110100",
  11458=>"101000001",
  11459=>"010001000",
  11460=>"110111111",
  11461=>"001100110",
  11462=>"001101001",
  11463=>"010101011",
  11464=>"011100111",
  11465=>"110010011",
  11466=>"100101111",
  11467=>"101100010",
  11468=>"110010011",
  11469=>"101101110",
  11470=>"111100100",
  11471=>"000011100",
  11472=>"110100110",
  11473=>"010110101",
  11474=>"000000011",
  11475=>"010001000",
  11476=>"111111001",
  11477=>"010100111",
  11478=>"000101010",
  11479=>"000001011",
  11480=>"110100010",
  11481=>"111000101",
  11482=>"101111001",
  11483=>"001001001",
  11484=>"001010011",
  11485=>"111000100",
  11486=>"110111110",
  11487=>"100110010",
  11488=>"100111000",
  11489=>"110111100",
  11490=>"110110001",
  11491=>"101100111",
  11492=>"100110111",
  11493=>"000100000",
  11494=>"011001100",
  11495=>"110101110",
  11496=>"111100011",
  11497=>"101010111",
  11498=>"101001001",
  11499=>"101010001",
  11500=>"000010000",
  11501=>"111010010",
  11502=>"101111101",
  11503=>"000010110",
  11504=>"100110001",
  11505=>"001101001",
  11506=>"100010000",
  11507=>"000100101",
  11508=>"000110101",
  11509=>"011010010",
  11510=>"100111010",
  11511=>"111111101",
  11512=>"100111010",
  11513=>"100101100",
  11514=>"001110011",
  11515=>"100101110",
  11516=>"100010000",
  11517=>"100011100",
  11518=>"110111001",
  11519=>"001111101",
  11520=>"011100010",
  11521=>"101000001",
  11522=>"100110000",
  11523=>"000101110",
  11524=>"001000100",
  11525=>"000011011",
  11526=>"110110110",
  11527=>"110111011",
  11528=>"111100000",
  11529=>"001010000",
  11530=>"100011100",
  11531=>"010101111",
  11532=>"101111100",
  11533=>"110000001",
  11534=>"010001011",
  11535=>"111011000",
  11536=>"111110100",
  11537=>"111111111",
  11538=>"111010111",
  11539=>"110000011",
  11540=>"010101110",
  11541=>"000110101",
  11542=>"111000101",
  11543=>"101111011",
  11544=>"111100001",
  11545=>"111101001",
  11546=>"110111010",
  11547=>"111110011",
  11548=>"111000011",
  11549=>"010000100",
  11550=>"001001111",
  11551=>"100110100",
  11552=>"010110000",
  11553=>"000001011",
  11554=>"111111111",
  11555=>"001100000",
  11556=>"000000111",
  11557=>"011110001",
  11558=>"000001100",
  11559=>"000001110",
  11560=>"001010111",
  11561=>"101100111",
  11562=>"011111100",
  11563=>"100101000",
  11564=>"101001010",
  11565=>"001100111",
  11566=>"100000000",
  11567=>"110100110",
  11568=>"000100001",
  11569=>"111011010",
  11570=>"110111110",
  11571=>"101010111",
  11572=>"110111111",
  11573=>"101001111",
  11574=>"111101110",
  11575=>"100000001",
  11576=>"001101110",
  11577=>"111110001",
  11578=>"101101111",
  11579=>"001001110",
  11580=>"110000110",
  11581=>"010000100",
  11582=>"001000010",
  11583=>"011011011",
  11584=>"011011001",
  11585=>"010100101",
  11586=>"000111100",
  11587=>"100111101",
  11588=>"111110010",
  11589=>"101010101",
  11590=>"100111100",
  11591=>"100000111",
  11592=>"011111010",
  11593=>"111001010",
  11594=>"111111010",
  11595=>"111001000",
  11596=>"110001101",
  11597=>"011111110",
  11598=>"010001011",
  11599=>"110110010",
  11600=>"111011010",
  11601=>"100110100",
  11602=>"000011110",
  11603=>"010011001",
  11604=>"000110111",
  11605=>"010100110",
  11606=>"000100111",
  11607=>"010100000",
  11608=>"001000010",
  11609=>"001100101",
  11610=>"011001010",
  11611=>"111101101",
  11612=>"100010010",
  11613=>"000010110",
  11614=>"110010100",
  11615=>"011111000",
  11616=>"100111010",
  11617=>"001011010",
  11618=>"010110010",
  11619=>"001111110",
  11620=>"011111001",
  11621=>"011100001",
  11622=>"111011001",
  11623=>"001010101",
  11624=>"111001110",
  11625=>"111110110",
  11626=>"101000010",
  11627=>"010100010",
  11628=>"111001000",
  11629=>"101011000",
  11630=>"100110000",
  11631=>"010011010",
  11632=>"001101000",
  11633=>"111000011",
  11634=>"110101000",
  11635=>"101110100",
  11636=>"111100100",
  11637=>"110100111",
  11638=>"111110111",
  11639=>"000000101",
  11640=>"101001111",
  11641=>"101000111",
  11642=>"110111100",
  11643=>"011110100",
  11644=>"111010100",
  11645=>"000000110",
  11646=>"010010011",
  11647=>"000011101",
  11648=>"110010111",
  11649=>"101110101",
  11650=>"000111001",
  11651=>"011111001",
  11652=>"110000000",
  11653=>"000001100",
  11654=>"101110100",
  11655=>"000111100",
  11656=>"000010000",
  11657=>"101110001",
  11658=>"110101011",
  11659=>"011111000",
  11660=>"001011111",
  11661=>"100010010",
  11662=>"010110100",
  11663=>"011101001",
  11664=>"000000010",
  11665=>"001001111",
  11666=>"110011100",
  11667=>"110000101",
  11668=>"111010000",
  11669=>"100001100",
  11670=>"111101011",
  11671=>"100101000",
  11672=>"111000000",
  11673=>"011000001",
  11674=>"110111100",
  11675=>"011000001",
  11676=>"011101000",
  11677=>"100101010",
  11678=>"001011011",
  11679=>"011001011",
  11680=>"110011001",
  11681=>"000100010",
  11682=>"111001011",
  11683=>"110110110",
  11684=>"001111101",
  11685=>"000000011",
  11686=>"001100010",
  11687=>"000110001",
  11688=>"000111110",
  11689=>"010101101",
  11690=>"100110000",
  11691=>"000001010",
  11692=>"011111110",
  11693=>"010111110",
  11694=>"011101010",
  11695=>"110101111",
  11696=>"001001000",
  11697=>"010100110",
  11698=>"001100111",
  11699=>"010110101",
  11700=>"111011101",
  11701=>"110110110",
  11702=>"001101111",
  11703=>"011001010",
  11704=>"100000011",
  11705=>"000001010",
  11706=>"010111010",
  11707=>"011111111",
  11708=>"111011110",
  11709=>"100101111",
  11710=>"000010000",
  11711=>"001110011",
  11712=>"001001010",
  11713=>"000001111",
  11714=>"110011100",
  11715=>"111110000",
  11716=>"000001101",
  11717=>"000100011",
  11718=>"100000111",
  11719=>"001100110",
  11720=>"000010101",
  11721=>"000000101",
  11722=>"001111100",
  11723=>"011101011",
  11724=>"000111100",
  11725=>"000001101",
  11726=>"010000011",
  11727=>"010110110",
  11728=>"001011111",
  11729=>"001011010",
  11730=>"011001101",
  11731=>"010011100",
  11732=>"110011000",
  11733=>"101100001",
  11734=>"000101011",
  11735=>"101111111",
  11736=>"001110101",
  11737=>"101100101",
  11738=>"000100000",
  11739=>"011100101",
  11740=>"110010001",
  11741=>"011000001",
  11742=>"011001011",
  11743=>"001101100",
  11744=>"100100001",
  11745=>"101001011",
  11746=>"111010110",
  11747=>"101110000",
  11748=>"110110111",
  11749=>"010000100",
  11750=>"101011111",
  11751=>"110111001",
  11752=>"010001100",
  11753=>"100101101",
  11754=>"001010010",
  11755=>"010000010",
  11756=>"001001101",
  11757=>"111101101",
  11758=>"000000011",
  11759=>"110111011",
  11760=>"100001010",
  11761=>"010010101",
  11762=>"011011101",
  11763=>"111101011",
  11764=>"001001110",
  11765=>"000110001",
  11766=>"000111111",
  11767=>"000010001",
  11768=>"100100101",
  11769=>"000010001",
  11770=>"101010100",
  11771=>"110101000",
  11772=>"010000000",
  11773=>"001011001",
  11774=>"010010110",
  11775=>"011010001",
  11776=>"001000100",
  11777=>"100110010",
  11778=>"001010100",
  11779=>"110011001",
  11780=>"001110011",
  11781=>"011010110",
  11782=>"110100000",
  11783=>"100000000",
  11784=>"001010000",
  11785=>"010010110",
  11786=>"110111001",
  11787=>"111100111",
  11788=>"010000001",
  11789=>"011111100",
  11790=>"101110000",
  11791=>"010010000",
  11792=>"000010111",
  11793=>"011000000",
  11794=>"001101011",
  11795=>"011010111",
  11796=>"111010011",
  11797=>"010100111",
  11798=>"000100000",
  11799=>"001011101",
  11800=>"001001001",
  11801=>"111111011",
  11802=>"010000000",
  11803=>"110000011",
  11804=>"111111110",
  11805=>"111011111",
  11806=>"101111000",
  11807=>"000010100",
  11808=>"000111100",
  11809=>"010111110",
  11810=>"110101000",
  11811=>"101101010",
  11812=>"001111010",
  11813=>"000101100",
  11814=>"100000111",
  11815=>"101000101",
  11816=>"011110110",
  11817=>"110101011",
  11818=>"100001001",
  11819=>"101110001",
  11820=>"001111100",
  11821=>"011000101",
  11822=>"011110101",
  11823=>"011100111",
  11824=>"010101100",
  11825=>"001110011",
  11826=>"100011001",
  11827=>"010000011",
  11828=>"010110001",
  11829=>"111111110",
  11830=>"101001011",
  11831=>"011100110",
  11832=>"001011100",
  11833=>"110000111",
  11834=>"010000000",
  11835=>"101101111",
  11836=>"101001000",
  11837=>"010000000",
  11838=>"011001000",
  11839=>"011100111",
  11840=>"111111101",
  11841=>"111110011",
  11842=>"011100111",
  11843=>"010111011",
  11844=>"001001110",
  11845=>"111011111",
  11846=>"001110000",
  11847=>"111100101",
  11848=>"011011011",
  11849=>"010101011",
  11850=>"111011111",
  11851=>"011101000",
  11852=>"011010110",
  11853=>"000100000",
  11854=>"001011010",
  11855=>"110001101",
  11856=>"110101111",
  11857=>"000011110",
  11858=>"000101111",
  11859=>"100000110",
  11860=>"110110111",
  11861=>"000011110",
  11862=>"110101111",
  11863=>"011100011",
  11864=>"111010101",
  11865=>"101110000",
  11866=>"100001001",
  11867=>"011110111",
  11868=>"010000101",
  11869=>"000110000",
  11870=>"001101100",
  11871=>"110101110",
  11872=>"010010000",
  11873=>"000000001",
  11874=>"011011101",
  11875=>"000000101",
  11876=>"001000111",
  11877=>"100000011",
  11878=>"101000010",
  11879=>"011110111",
  11880=>"100110101",
  11881=>"100011000",
  11882=>"000111010",
  11883=>"100000010",
  11884=>"110001010",
  11885=>"101110011",
  11886=>"110111110",
  11887=>"010011000",
  11888=>"000010010",
  11889=>"011001000",
  11890=>"001111110",
  11891=>"101101111",
  11892=>"001000111",
  11893=>"000001010",
  11894=>"110001111",
  11895=>"000011110",
  11896=>"011010001",
  11897=>"001100101",
  11898=>"001000100",
  11899=>"000111111",
  11900=>"110011001",
  11901=>"100100001",
  11902=>"001110111",
  11903=>"100000000",
  11904=>"010111011",
  11905=>"010001000",
  11906=>"100111110",
  11907=>"000001100",
  11908=>"001001111",
  11909=>"100100011",
  11910=>"111011000",
  11911=>"001100010",
  11912=>"101101110",
  11913=>"110101011",
  11914=>"110110111",
  11915=>"110111101",
  11916=>"110010011",
  11917=>"010000010",
  11918=>"000100001",
  11919=>"100101001",
  11920=>"000010110",
  11921=>"100111010",
  11922=>"011011001",
  11923=>"001010100",
  11924=>"110100101",
  11925=>"100010111",
  11926=>"001000000",
  11927=>"110110101",
  11928=>"100111100",
  11929=>"010100010",
  11930=>"111000111",
  11931=>"000001011",
  11932=>"010110100",
  11933=>"100001111",
  11934=>"101110010",
  11935=>"110100011",
  11936=>"000000000",
  11937=>"110110011",
  11938=>"110001011",
  11939=>"001011111",
  11940=>"010110111",
  11941=>"110011000",
  11942=>"001110001",
  11943=>"010000000",
  11944=>"101001101",
  11945=>"111110110",
  11946=>"100010110",
  11947=>"001011100",
  11948=>"111111110",
  11949=>"010101111",
  11950=>"100111011",
  11951=>"110011110",
  11952=>"000111101",
  11953=>"110010101",
  11954=>"101101100",
  11955=>"111001010",
  11956=>"100100000",
  11957=>"000001010",
  11958=>"110100110",
  11959=>"001100110",
  11960=>"001101101",
  11961=>"111001100",
  11962=>"110000010",
  11963=>"010101011",
  11964=>"110101000",
  11965=>"110000010",
  11966=>"000101100",
  11967=>"000000110",
  11968=>"011110110",
  11969=>"100010000",
  11970=>"001000111",
  11971=>"100011101",
  11972=>"001101100",
  11973=>"111010100",
  11974=>"011010101",
  11975=>"000001001",
  11976=>"110101001",
  11977=>"101101111",
  11978=>"101101010",
  11979=>"110101000",
  11980=>"000100010",
  11981=>"000101011",
  11982=>"000001011",
  11983=>"000001101",
  11984=>"011001001",
  11985=>"001001111",
  11986=>"101000110",
  11987=>"110100110",
  11988=>"000011100",
  11989=>"110100101",
  11990=>"111001010",
  11991=>"111110011",
  11992=>"001001000",
  11993=>"101010011",
  11994=>"111111011",
  11995=>"001000111",
  11996=>"000100100",
  11997=>"010000110",
  11998=>"011001100",
  11999=>"001110111",
  12000=>"001010000",
  12001=>"010110010",
  12002=>"111010100",
  12003=>"000000000",
  12004=>"000101110",
  12005=>"000101000",
  12006=>"100001011",
  12007=>"100100001",
  12008=>"101001011",
  12009=>"110000001",
  12010=>"111101101",
  12011=>"000110001",
  12012=>"111111111",
  12013=>"010011101",
  12014=>"101101001",
  12015=>"010111001",
  12016=>"100101101",
  12017=>"011001110",
  12018=>"001000100",
  12019=>"000101100",
  12020=>"100010111",
  12021=>"110001000",
  12022=>"010011110",
  12023=>"100000001",
  12024=>"010010111",
  12025=>"111111010",
  12026=>"110111011",
  12027=>"101111001",
  12028=>"111000101",
  12029=>"001101100",
  12030=>"100010001",
  12031=>"011101000",
  12032=>"000010100",
  12033=>"011101111",
  12034=>"010000010",
  12035=>"100101000",
  12036=>"100011101",
  12037=>"000100110",
  12038=>"101011111",
  12039=>"101011011",
  12040=>"111001100",
  12041=>"111111111",
  12042=>"111101101",
  12043=>"101000001",
  12044=>"101100110",
  12045=>"001111101",
  12046=>"000001100",
  12047=>"010110110",
  12048=>"111100111",
  12049=>"100111111",
  12050=>"011111111",
  12051=>"101010100",
  12052=>"100110111",
  12053=>"011010010",
  12054=>"111011010",
  12055=>"111001010",
  12056=>"111101000",
  12057=>"001001010",
  12058=>"111001110",
  12059=>"100011110",
  12060=>"011000010",
  12061=>"110010111",
  12062=>"011101101",
  12063=>"111100111",
  12064=>"110010001",
  12065=>"110110101",
  12066=>"010000101",
  12067=>"111111100",
  12068=>"100101111",
  12069=>"001101111",
  12070=>"000001110",
  12071=>"010010100",
  12072=>"111010111",
  12073=>"100011010",
  12074=>"001111010",
  12075=>"010101001",
  12076=>"100111000",
  12077=>"000000000",
  12078=>"000011000",
  12079=>"110110100",
  12080=>"101110111",
  12081=>"001000011",
  12082=>"000111111",
  12083=>"000010110",
  12084=>"011100100",
  12085=>"010000001",
  12086=>"000101101",
  12087=>"000100100",
  12088=>"111001011",
  12089=>"011011101",
  12090=>"000010000",
  12091=>"100110001",
  12092=>"110011101",
  12093=>"010011110",
  12094=>"111101011",
  12095=>"001100001",
  12096=>"100111110",
  12097=>"000010111",
  12098=>"010011111",
  12099=>"010010001",
  12100=>"011000001",
  12101=>"001100000",
  12102=>"001011011",
  12103=>"111111000",
  12104=>"111110001",
  12105=>"010001001",
  12106=>"100110111",
  12107=>"000010101",
  12108=>"000010110",
  12109=>"100011011",
  12110=>"000010001",
  12111=>"100110111",
  12112=>"011001101",
  12113=>"010001010",
  12114=>"001000011",
  12115=>"001111001",
  12116=>"000100000",
  12117=>"110001000",
  12118=>"001111100",
  12119=>"001101000",
  12120=>"011110011",
  12121=>"111101001",
  12122=>"111100011",
  12123=>"100001100",
  12124=>"000010000",
  12125=>"000101111",
  12126=>"101001000",
  12127=>"000001111",
  12128=>"101000000",
  12129=>"110111010",
  12130=>"000000011",
  12131=>"001111110",
  12132=>"010100010",
  12133=>"010000101",
  12134=>"010100001",
  12135=>"011001011",
  12136=>"100000100",
  12137=>"000001110",
  12138=>"110100100",
  12139=>"011011110",
  12140=>"000100111",
  12141=>"100100110",
  12142=>"011000101",
  12143=>"111110111",
  12144=>"100010110",
  12145=>"000011110",
  12146=>"000100001",
  12147=>"010011000",
  12148=>"010111000",
  12149=>"011001011",
  12150=>"010101011",
  12151=>"011001000",
  12152=>"001001001",
  12153=>"011000111",
  12154=>"100011000",
  12155=>"111111000",
  12156=>"001111100",
  12157=>"010100111",
  12158=>"111010100",
  12159=>"100110100",
  12160=>"010010011",
  12161=>"111010001",
  12162=>"001111100",
  12163=>"010010000",
  12164=>"101010111",
  12165=>"110111001",
  12166=>"010110000",
  12167=>"000001010",
  12168=>"101111000",
  12169=>"101010100",
  12170=>"000111101",
  12171=>"000000010",
  12172=>"010111111",
  12173=>"010100110",
  12174=>"010001001",
  12175=>"011011100",
  12176=>"100011001",
  12177=>"111101000",
  12178=>"100111000",
  12179=>"011000010",
  12180=>"000001011",
  12181=>"010111100",
  12182=>"010010001",
  12183=>"011111101",
  12184=>"001011100",
  12185=>"110001011",
  12186=>"001001110",
  12187=>"001010101",
  12188=>"011000111",
  12189=>"111000100",
  12190=>"001100001",
  12191=>"001000101",
  12192=>"010000101",
  12193=>"100110111",
  12194=>"111100010",
  12195=>"111101011",
  12196=>"101110111",
  12197=>"100000111",
  12198=>"010111100",
  12199=>"011101111",
  12200=>"100101111",
  12201=>"000001000",
  12202=>"111110010",
  12203=>"101000111",
  12204=>"010110100",
  12205=>"001111111",
  12206=>"010111100",
  12207=>"110011001",
  12208=>"110011101",
  12209=>"110100011",
  12210=>"001000010",
  12211=>"000010011",
  12212=>"100001101",
  12213=>"101100111",
  12214=>"110011110",
  12215=>"001100011",
  12216=>"111100011",
  12217=>"100001001",
  12218=>"011011011",
  12219=>"011010010",
  12220=>"101011011",
  12221=>"000111011",
  12222=>"010000110",
  12223=>"111101101",
  12224=>"111110101",
  12225=>"010110011",
  12226=>"010000110",
  12227=>"101110001",
  12228=>"101010111",
  12229=>"011101000",
  12230=>"001101001",
  12231=>"110110000",
  12232=>"011011001",
  12233=>"110101011",
  12234=>"010110100",
  12235=>"000010010",
  12236=>"111101001",
  12237=>"110111100",
  12238=>"001110111",
  12239=>"011011010",
  12240=>"011000001",
  12241=>"110011100",
  12242=>"101101111",
  12243=>"000001100",
  12244=>"010111011",
  12245=>"110000100",
  12246=>"110000110",
  12247=>"001111010",
  12248=>"101110111",
  12249=>"110010010",
  12250=>"000101001",
  12251=>"100000111",
  12252=>"111000111",
  12253=>"111111101",
  12254=>"011110010",
  12255=>"001100011",
  12256=>"100000000",
  12257=>"011000000",
  12258=>"101100101",
  12259=>"000100100",
  12260=>"101000101",
  12261=>"001000000",
  12262=>"011111111",
  12263=>"000001010",
  12264=>"101011000",
  12265=>"001100000",
  12266=>"001110001",
  12267=>"001011101",
  12268=>"111011111",
  12269=>"111110111",
  12270=>"011010110",
  12271=>"010010011",
  12272=>"111001010",
  12273=>"011110100",
  12274=>"100000101",
  12275=>"101000011",
  12276=>"110110110",
  12277=>"010111101",
  12278=>"111010101",
  12279=>"010101111",
  12280=>"010001111",
  12281=>"001111100",
  12282=>"101101110",
  12283=>"111010000",
  12284=>"001010100",
  12285=>"100000011",
  12286=>"000110001",
  12287=>"001101110",
  12288=>"100101001",
  12289=>"000101011",
  12290=>"001001000",
  12291=>"111111001",
  12292=>"101001101",
  12293=>"011111110",
  12294=>"101010101",
  12295=>"111011010",
  12296=>"111100100",
  12297=>"110000001",
  12298=>"011100000",
  12299=>"011110001",
  12300=>"001111100",
  12301=>"111000010",
  12302=>"010111110",
  12303=>"011101011",
  12304=>"101000111",
  12305=>"110101011",
  12306=>"010101011",
  12307=>"001100100",
  12308=>"011101001",
  12309=>"111011001",
  12310=>"000101101",
  12311=>"100010111",
  12312=>"100111001",
  12313=>"101110111",
  12314=>"100011110",
  12315=>"010011000",
  12316=>"010111100",
  12317=>"001110001",
  12318=>"111001000",
  12319=>"101111000",
  12320=>"111111110",
  12321=>"110101001",
  12322=>"000100001",
  12323=>"010110000",
  12324=>"111001011",
  12325=>"111011000",
  12326=>"111100110",
  12327=>"110110111",
  12328=>"001011010",
  12329=>"011101001",
  12330=>"110110010",
  12331=>"101001101",
  12332=>"111101001",
  12333=>"101101110",
  12334=>"101110101",
  12335=>"001111101",
  12336=>"100110111",
  12337=>"000110110",
  12338=>"111011010",
  12339=>"100111111",
  12340=>"000111100",
  12341=>"000101011",
  12342=>"110001100",
  12343=>"011111111",
  12344=>"110110111",
  12345=>"111110011",
  12346=>"001111101",
  12347=>"100011111",
  12348=>"100110011",
  12349=>"011101100",
  12350=>"010111010",
  12351=>"110110100",
  12352=>"100101000",
  12353=>"111001100",
  12354=>"001001100",
  12355=>"001111000",
  12356=>"100000000",
  12357=>"101011101",
  12358=>"010000000",
  12359=>"000101011",
  12360=>"010100000",
  12361=>"100000100",
  12362=>"100101010",
  12363=>"111111010",
  12364=>"111110110",
  12365=>"110011110",
  12366=>"101010110",
  12367=>"010001011",
  12368=>"000000111",
  12369=>"001001000",
  12370=>"100001010",
  12371=>"011100101",
  12372=>"111100011",
  12373=>"001111011",
  12374=>"110010110",
  12375=>"011101001",
  12376=>"101011000",
  12377=>"010100010",
  12378=>"001110001",
  12379=>"110111101",
  12380=>"010111110",
  12381=>"011000011",
  12382=>"100001001",
  12383=>"000111101",
  12384=>"101100000",
  12385=>"110000010",
  12386=>"001010101",
  12387=>"000011110",
  12388=>"101100111",
  12389=>"001111110",
  12390=>"101110110",
  12391=>"001010010",
  12392=>"111101011",
  12393=>"000001000",
  12394=>"101110000",
  12395=>"001101111",
  12396=>"111001111",
  12397=>"011001010",
  12398=>"011001000",
  12399=>"111111011",
  12400=>"110101010",
  12401=>"011110100",
  12402=>"100110111",
  12403=>"111011000",
  12404=>"010011001",
  12405=>"001101001",
  12406=>"111111011",
  12407=>"001100100",
  12408=>"101000101",
  12409=>"111101011",
  12410=>"000011001",
  12411=>"100010111",
  12412=>"011110111",
  12413=>"110111000",
  12414=>"011001110",
  12415=>"100011011",
  12416=>"111011111",
  12417=>"110101010",
  12418=>"001001001",
  12419=>"010001111",
  12420=>"000110101",
  12421=>"100100010",
  12422=>"000101110",
  12423=>"101111000",
  12424=>"010101011",
  12425=>"101011100",
  12426=>"000101110",
  12427=>"011100111",
  12428=>"010011010",
  12429=>"001011011",
  12430=>"011010010",
  12431=>"010000111",
  12432=>"011010110",
  12433=>"001000110",
  12434=>"011000100",
  12435=>"011110010",
  12436=>"110100101",
  12437=>"000100111",
  12438=>"010011111",
  12439=>"001000000",
  12440=>"111101010",
  12441=>"001011100",
  12442=>"000000111",
  12443=>"101101100",
  12444=>"001010000",
  12445=>"010001100",
  12446=>"001110010",
  12447=>"010001000",
  12448=>"011111111",
  12449=>"000100111",
  12450=>"101000111",
  12451=>"110001111",
  12452=>"111100010",
  12453=>"011101001",
  12454=>"100001001",
  12455=>"011001011",
  12456=>"111001100",
  12457=>"100000100",
  12458=>"010010010",
  12459=>"100000110",
  12460=>"100101110",
  12461=>"100110000",
  12462=>"100011001",
  12463=>"000111011",
  12464=>"010001100",
  12465=>"011101111",
  12466=>"011000100",
  12467=>"000100111",
  12468=>"010100011",
  12469=>"100110101",
  12470=>"110100100",
  12471=>"001001001",
  12472=>"100001101",
  12473=>"010110010",
  12474=>"000010000",
  12475=>"000101000",
  12476=>"001100100",
  12477=>"101010100",
  12478=>"010011011",
  12479=>"010001000",
  12480=>"101100000",
  12481=>"011000100",
  12482=>"111110110",
  12483=>"110100110",
  12484=>"111101101",
  12485=>"010011101",
  12486=>"100011011",
  12487=>"101000101",
  12488=>"110000111",
  12489=>"001001101",
  12490=>"011000110",
  12491=>"010000010",
  12492=>"001110100",
  12493=>"011000010",
  12494=>"011011111",
  12495=>"111011011",
  12496=>"000111110",
  12497=>"011011101",
  12498=>"010011000",
  12499=>"101001101",
  12500=>"010011011",
  12501=>"011110010",
  12502=>"110100001",
  12503=>"000010001",
  12504=>"011111111",
  12505=>"110011001",
  12506=>"111001100",
  12507=>"111010010",
  12508=>"100001001",
  12509=>"010000110",
  12510=>"000111001",
  12511=>"111101100",
  12512=>"111110110",
  12513=>"000010001",
  12514=>"000000011",
  12515=>"111110101",
  12516=>"100001001",
  12517=>"011000100",
  12518=>"010101101",
  12519=>"001001110",
  12520=>"100010000",
  12521=>"111011011",
  12522=>"001111101",
  12523=>"101111100",
  12524=>"011100000",
  12525=>"111111001",
  12526=>"111101011",
  12527=>"010101010",
  12528=>"101110101",
  12529=>"110000110",
  12530=>"101101011",
  12531=>"000011111",
  12532=>"000101000",
  12533=>"001001000",
  12534=>"101101011",
  12535=>"110110111",
  12536=>"010000001",
  12537=>"011010111",
  12538=>"101000000",
  12539=>"010111101",
  12540=>"000000111",
  12541=>"100001010",
  12542=>"010100101",
  12543=>"110000001",
  12544=>"000001001",
  12545=>"000111010",
  12546=>"010110000",
  12547=>"101111011",
  12548=>"110100110",
  12549=>"110111100",
  12550=>"011000001",
  12551=>"101110110",
  12552=>"110101111",
  12553=>"110000111",
  12554=>"101100011",
  12555=>"110111101",
  12556=>"111011110",
  12557=>"100101100",
  12558=>"000001001",
  12559=>"110100111",
  12560=>"100101011",
  12561=>"001000110",
  12562=>"111110101",
  12563=>"100101101",
  12564=>"001110100",
  12565=>"111011100",
  12566=>"111011100",
  12567=>"010011010",
  12568=>"011110111",
  12569=>"111111000",
  12570=>"111100110",
  12571=>"111111000",
  12572=>"111111110",
  12573=>"000101100",
  12574=>"101010010",
  12575=>"001110111",
  12576=>"000010010",
  12577=>"000101010",
  12578=>"110100110",
  12579=>"111110010",
  12580=>"101110001",
  12581=>"110001001",
  12582=>"111110100",
  12583=>"000010111",
  12584=>"011100101",
  12585=>"111001000",
  12586=>"110111110",
  12587=>"011111110",
  12588=>"011100111",
  12589=>"101110010",
  12590=>"111011101",
  12591=>"110101000",
  12592=>"101011111",
  12593=>"110100101",
  12594=>"101001010",
  12595=>"100111100",
  12596=>"111010011",
  12597=>"000010000",
  12598=>"110101010",
  12599=>"001010011",
  12600=>"111100110",
  12601=>"010111011",
  12602=>"111001111",
  12603=>"000000111",
  12604=>"110110111",
  12605=>"100100110",
  12606=>"100010011",
  12607=>"110000100",
  12608=>"100110000",
  12609=>"011110011",
  12610=>"000010100",
  12611=>"011011000",
  12612=>"101110101",
  12613=>"001011101",
  12614=>"101001100",
  12615=>"010101010",
  12616=>"100010010",
  12617=>"001101101",
  12618=>"111111101",
  12619=>"000001111",
  12620=>"000001101",
  12621=>"001100100",
  12622=>"000101001",
  12623=>"011111110",
  12624=>"100010111",
  12625=>"101100101",
  12626=>"111110000",
  12627=>"001010011",
  12628=>"110100111",
  12629=>"111111000",
  12630=>"111110111",
  12631=>"001000111",
  12632=>"111011010",
  12633=>"111000101",
  12634=>"011111101",
  12635=>"011111110",
  12636=>"000110000",
  12637=>"001001000",
  12638=>"011010011",
  12639=>"100101111",
  12640=>"101001100",
  12641=>"100100110",
  12642=>"110101101",
  12643=>"111011110",
  12644=>"111001000",
  12645=>"110011000",
  12646=>"001110010",
  12647=>"111111010",
  12648=>"100000001",
  12649=>"001011110",
  12650=>"000001111",
  12651=>"100111100",
  12652=>"000100011",
  12653=>"000110111",
  12654=>"111001011",
  12655=>"010010101",
  12656=>"111100111",
  12657=>"000001101",
  12658=>"110100111",
  12659=>"010011001",
  12660=>"001110010",
  12661=>"111000101",
  12662=>"011110111",
  12663=>"110100011",
  12664=>"011110001",
  12665=>"100000111",
  12666=>"011100110",
  12667=>"000010111",
  12668=>"100110111",
  12669=>"101110001",
  12670=>"000001000",
  12671=>"010000100",
  12672=>"111010011",
  12673=>"111111110",
  12674=>"010100101",
  12675=>"100001111",
  12676=>"110100000",
  12677=>"011011111",
  12678=>"000110110",
  12679=>"110110000",
  12680=>"011111100",
  12681=>"101001111",
  12682=>"011110001",
  12683=>"011110011",
  12684=>"110110100",
  12685=>"010111111",
  12686=>"000011101",
  12687=>"000101011",
  12688=>"001000101",
  12689=>"100011101",
  12690=>"001100000",
  12691=>"101010111",
  12692=>"011100000",
  12693=>"110000011",
  12694=>"011011010",
  12695=>"010001111",
  12696=>"100100010",
  12697=>"011111011",
  12698=>"000110110",
  12699=>"100101001",
  12700=>"000001001",
  12701=>"001001100",
  12702=>"011010110",
  12703=>"110111001",
  12704=>"000100111",
  12705=>"111100000",
  12706=>"101010111",
  12707=>"111110111",
  12708=>"101000110",
  12709=>"010111011",
  12710=>"010010100",
  12711=>"111001110",
  12712=>"000101100",
  12713=>"010001010",
  12714=>"000010000",
  12715=>"111100111",
  12716=>"110111110",
  12717=>"101011101",
  12718=>"011111101",
  12719=>"101011010",
  12720=>"010110000",
  12721=>"011100101",
  12722=>"010010100",
  12723=>"010011101",
  12724=>"010010111",
  12725=>"111111010",
  12726=>"010111101",
  12727=>"100000000",
  12728=>"000101010",
  12729=>"100010111",
  12730=>"001110011",
  12731=>"101100110",
  12732=>"010100011",
  12733=>"000001010",
  12734=>"100010000",
  12735=>"110101010",
  12736=>"011010110",
  12737=>"110111000",
  12738=>"010100100",
  12739=>"101111101",
  12740=>"110001000",
  12741=>"100101000",
  12742=>"010000000",
  12743=>"100100111",
  12744=>"111011010",
  12745=>"000001110",
  12746=>"101101011",
  12747=>"110100101",
  12748=>"011001010",
  12749=>"000111011",
  12750=>"101100001",
  12751=>"101101111",
  12752=>"100011000",
  12753=>"000000110",
  12754=>"000001110",
  12755=>"011000101",
  12756=>"111011111",
  12757=>"010000111",
  12758=>"100111110",
  12759=>"100000011",
  12760=>"101011011",
  12761=>"111100011",
  12762=>"000011100",
  12763=>"011000101",
  12764=>"101111111",
  12765=>"011100010",
  12766=>"011010010",
  12767=>"000011110",
  12768=>"110011011",
  12769=>"001100111",
  12770=>"111000101",
  12771=>"101010000",
  12772=>"101110001",
  12773=>"000000100",
  12774=>"100110011",
  12775=>"111110111",
  12776=>"100010100",
  12777=>"001111111",
  12778=>"101010000",
  12779=>"011011001",
  12780=>"010001101",
  12781=>"100000000",
  12782=>"000000011",
  12783=>"010101110",
  12784=>"110010111",
  12785=>"000001010",
  12786=>"100000001",
  12787=>"000110011",
  12788=>"100000100",
  12789=>"111110011",
  12790=>"110010111",
  12791=>"000111000",
  12792=>"101101100",
  12793=>"000110000",
  12794=>"000000110",
  12795=>"101101011",
  12796=>"110000010",
  12797=>"101001000",
  12798=>"111111001",
  12799=>"111101101",
  12800=>"011101100",
  12801=>"011011001",
  12802=>"011000001",
  12803=>"001011011",
  12804=>"010000111",
  12805=>"000001010",
  12806=>"110011000",
  12807=>"101101101",
  12808=>"001111000",
  12809=>"011011011",
  12810=>"101101101",
  12811=>"010111111",
  12812=>"001101010",
  12813=>"010111111",
  12814=>"001001011",
  12815=>"101011000",
  12816=>"001100100",
  12817=>"010010110",
  12818=>"101101010",
  12819=>"011001100",
  12820=>"010011100",
  12821=>"010111001",
  12822=>"101010111",
  12823=>"001011011",
  12824=>"111000110",
  12825=>"000011100",
  12826=>"011111110",
  12827=>"010011100",
  12828=>"111101011",
  12829=>"111110011",
  12830=>"001011111",
  12831=>"011100101",
  12832=>"000001010",
  12833=>"001001010",
  12834=>"101010001",
  12835=>"111001111",
  12836=>"011001100",
  12837=>"111000110",
  12838=>"110010111",
  12839=>"010111001",
  12840=>"000111010",
  12841=>"110100001",
  12842=>"011100010",
  12843=>"100010101",
  12844=>"111010001",
  12845=>"011101101",
  12846=>"101110101",
  12847=>"000000101",
  12848=>"000110110",
  12849=>"100000010",
  12850=>"111101000",
  12851=>"000001000",
  12852=>"000111100",
  12853=>"111001111",
  12854=>"110100001",
  12855=>"100000101",
  12856=>"111111111",
  12857=>"001001111",
  12858=>"110000001",
  12859=>"110010010",
  12860=>"101100011",
  12861=>"100101011",
  12862=>"001101110",
  12863=>"111100100",
  12864=>"001000100",
  12865=>"100011101",
  12866=>"110111100",
  12867=>"001001010",
  12868=>"101001001",
  12869=>"100111111",
  12870=>"100000110",
  12871=>"000010010",
  12872=>"001000011",
  12873=>"000100100",
  12874=>"010010110",
  12875=>"000110111",
  12876=>"100011001",
  12877=>"101001111",
  12878=>"000100110",
  12879=>"000110101",
  12880=>"011101111",
  12881=>"101011010",
  12882=>"110011001",
  12883=>"111001101",
  12884=>"101111011",
  12885=>"000111100",
  12886=>"111101101",
  12887=>"110110111",
  12888=>"011101111",
  12889=>"111000010",
  12890=>"001101111",
  12891=>"011110111",
  12892=>"011011111",
  12893=>"011111010",
  12894=>"010110110",
  12895=>"101010110",
  12896=>"010000111",
  12897=>"111110110",
  12898=>"001010001",
  12899=>"001111011",
  12900=>"000000111",
  12901=>"011011001",
  12902=>"110101010",
  12903=>"000111011",
  12904=>"011111101",
  12905=>"010011101",
  12906=>"111010011",
  12907=>"011011011",
  12908=>"111011010",
  12909=>"000101011",
  12910=>"101100010",
  12911=>"000101001",
  12912=>"011001100",
  12913=>"111111100",
  12914=>"101010010",
  12915=>"101001101",
  12916=>"110100100",
  12917=>"111100101",
  12918=>"101001010",
  12919=>"111111111",
  12920=>"111101101",
  12921=>"110111010",
  12922=>"000101101",
  12923=>"111001000",
  12924=>"110010101",
  12925=>"011001001",
  12926=>"011101000",
  12927=>"000000011",
  12928=>"000000111",
  12929=>"001000000",
  12930=>"011010101",
  12931=>"111111010",
  12932=>"011100100",
  12933=>"111011111",
  12934=>"011100101",
  12935=>"111110110",
  12936=>"011110110",
  12937=>"000011101",
  12938=>"110110100",
  12939=>"011101100",
  12940=>"100111111",
  12941=>"001000000",
  12942=>"110100011",
  12943=>"111011000",
  12944=>"101100000",
  12945=>"010100000",
  12946=>"110010010",
  12947=>"011011001",
  12948=>"110010010",
  12949=>"101010101",
  12950=>"111111101",
  12951=>"011010110",
  12952=>"101001101",
  12953=>"000011011",
  12954=>"110010101",
  12955=>"011001011",
  12956=>"110110000",
  12957=>"100011101",
  12958=>"101101000",
  12959=>"101001000",
  12960=>"101101111",
  12961=>"101001110",
  12962=>"010000011",
  12963=>"101010100",
  12964=>"101010000",
  12965=>"011001010",
  12966=>"111110111",
  12967=>"111101111",
  12968=>"011011011",
  12969=>"000000011",
  12970=>"011000111",
  12971=>"100101111",
  12972=>"011111010",
  12973=>"100100011",
  12974=>"110010001",
  12975=>"000110010",
  12976=>"000110111",
  12977=>"011101100",
  12978=>"011010100",
  12979=>"100011101",
  12980=>"000001011",
  12981=>"010001101",
  12982=>"010110101",
  12983=>"010000001",
  12984=>"100100001",
  12985=>"111011100",
  12986=>"101110011",
  12987=>"011010000",
  12988=>"100100010",
  12989=>"101001110",
  12990=>"100011011",
  12991=>"011110011",
  12992=>"011011110",
  12993=>"100110000",
  12994=>"101011001",
  12995=>"100010101",
  12996=>"110100110",
  12997=>"110000011",
  12998=>"100110000",
  12999=>"010111001",
  13000=>"100000001",
  13001=>"100110000",
  13002=>"100000001",
  13003=>"110111011",
  13004=>"000101010",
  13005=>"101111010",
  13006=>"101001110",
  13007=>"010100110",
  13008=>"000010111",
  13009=>"101111101",
  13010=>"011101111",
  13011=>"111011001",
  13012=>"011000101",
  13013=>"101111101",
  13014=>"010110111",
  13015=>"101111110",
  13016=>"111111000",
  13017=>"110100000",
  13018=>"111111111",
  13019=>"011110001",
  13020=>"010010100",
  13021=>"011111110",
  13022=>"100110000",
  13023=>"010011000",
  13024=>"100101111",
  13025=>"100110010",
  13026=>"000100101",
  13027=>"001111010",
  13028=>"101011111",
  13029=>"100000100",
  13030=>"000111001",
  13031=>"001111001",
  13032=>"011111010",
  13033=>"011011100",
  13034=>"011011101",
  13035=>"000001100",
  13036=>"110111100",
  13037=>"010011111",
  13038=>"111100101",
  13039=>"001110010",
  13040=>"110101101",
  13041=>"001100110",
  13042=>"011101110",
  13043=>"010010000",
  13044=>"011000110",
  13045=>"011000110",
  13046=>"011101011",
  13047=>"111000000",
  13048=>"101000110",
  13049=>"100110110",
  13050=>"111111000",
  13051=>"101011101",
  13052=>"011111111",
  13053=>"010000011",
  13054=>"110100010",
  13055=>"100110111",
  13056=>"111010101",
  13057=>"110100101",
  13058=>"000100111",
  13059=>"010100010",
  13060=>"000001011",
  13061=>"110010001",
  13062=>"011011110",
  13063=>"000110111",
  13064=>"100100111",
  13065=>"000000100",
  13066=>"001100100",
  13067=>"001111111",
  13068=>"100101110",
  13069=>"101110111",
  13070=>"011011011",
  13071=>"000110001",
  13072=>"100011111",
  13073=>"011010010",
  13074=>"110100100",
  13075=>"001000101",
  13076=>"001011110",
  13077=>"010110110",
  13078=>"010111000",
  13079=>"111000000",
  13080=>"011011011",
  13081=>"001111001",
  13082=>"001011001",
  13083=>"111001011",
  13084=>"010001011",
  13085=>"001000010",
  13086=>"111100011",
  13087=>"100101000",
  13088=>"110100111",
  13089=>"000000011",
  13090=>"010110110",
  13091=>"101111011",
  13092=>"000011010",
  13093=>"100000100",
  13094=>"001010011",
  13095=>"110001100",
  13096=>"010100100",
  13097=>"001011001",
  13098=>"001010101",
  13099=>"010101100",
  13100=>"111001001",
  13101=>"111110010",
  13102=>"101010011",
  13103=>"001001010",
  13104=>"111010010",
  13105=>"000101001",
  13106=>"010101101",
  13107=>"010100110",
  13108=>"001000000",
  13109=>"001000010",
  13110=>"101100001",
  13111=>"111011110",
  13112=>"101011110",
  13113=>"111011011",
  13114=>"100111010",
  13115=>"010001100",
  13116=>"001001011",
  13117=>"111111100",
  13118=>"110111000",
  13119=>"101001011",
  13120=>"010110001",
  13121=>"100110000",
  13122=>"110011100",
  13123=>"001001111",
  13124=>"100110011",
  13125=>"001011101",
  13126=>"010001011",
  13127=>"001101101",
  13128=>"101101011",
  13129=>"001011100",
  13130=>"001111001",
  13131=>"001000010",
  13132=>"010110110",
  13133=>"000011010",
  13134=>"101111111",
  13135=>"101110111",
  13136=>"001101101",
  13137=>"110100011",
  13138=>"100011110",
  13139=>"011001000",
  13140=>"011111101",
  13141=>"011101011",
  13142=>"101111101",
  13143=>"111111011",
  13144=>"001000101",
  13145=>"100111011",
  13146=>"100111100",
  13147=>"111000011",
  13148=>"001110010",
  13149=>"110010010",
  13150=>"011110011",
  13151=>"111011011",
  13152=>"110011001",
  13153=>"000110101",
  13154=>"010011001",
  13155=>"001110110",
  13156=>"100011101",
  13157=>"101001111",
  13158=>"001001101",
  13159=>"001011100",
  13160=>"001110100",
  13161=>"110100011",
  13162=>"101111100",
  13163=>"110101001",
  13164=>"111000111",
  13165=>"111010001",
  13166=>"001111011",
  13167=>"111001111",
  13168=>"001100000",
  13169=>"110001110",
  13170=>"001010001",
  13171=>"110101011",
  13172=>"100110000",
  13173=>"111001110",
  13174=>"111000100",
  13175=>"101000111",
  13176=>"101111000",
  13177=>"101111011",
  13178=>"011000010",
  13179=>"000011110",
  13180=>"111011110",
  13181=>"010101111",
  13182=>"111011011",
  13183=>"110011110",
  13184=>"111111111",
  13185=>"000001111",
  13186=>"110111011",
  13187=>"100111101",
  13188=>"010101000",
  13189=>"111101110",
  13190=>"001010010",
  13191=>"001111011",
  13192=>"110111000",
  13193=>"110010110",
  13194=>"001100010",
  13195=>"110110000",
  13196=>"110111110",
  13197=>"010000111",
  13198=>"000101110",
  13199=>"101111010",
  13200=>"000110110",
  13201=>"110100110",
  13202=>"111000000",
  13203=>"110001111",
  13204=>"100000000",
  13205=>"100001100",
  13206=>"011111100",
  13207=>"111110111",
  13208=>"000110111",
  13209=>"010011000",
  13210=>"001001010",
  13211=>"110000110",
  13212=>"011101100",
  13213=>"010111111",
  13214=>"011101111",
  13215=>"111110110",
  13216=>"111100101",
  13217=>"011101100",
  13218=>"000101010",
  13219=>"001111001",
  13220=>"010010011",
  13221=>"111111111",
  13222=>"011101011",
  13223=>"110111011",
  13224=>"001110011",
  13225=>"101111100",
  13226=>"101001100",
  13227=>"000000100",
  13228=>"110011101",
  13229=>"111100011",
  13230=>"001000101",
  13231=>"101111000",
  13232=>"100011000",
  13233=>"110011001",
  13234=>"011110111",
  13235=>"000010101",
  13236=>"010001111",
  13237=>"011100110",
  13238=>"111101001",
  13239=>"011001011",
  13240=>"001100001",
  13241=>"100110110",
  13242=>"111011001",
  13243=>"101111000",
  13244=>"100000110",
  13245=>"101100000",
  13246=>"011101110",
  13247=>"001001011",
  13248=>"101111101",
  13249=>"111000111",
  13250=>"110110010",
  13251=>"101101110",
  13252=>"010110110",
  13253=>"000111000",
  13254=>"100100000",
  13255=>"010101110",
  13256=>"110111000",
  13257=>"111111111",
  13258=>"000101100",
  13259=>"101111010",
  13260=>"010011101",
  13261=>"100111011",
  13262=>"111101001",
  13263=>"101111000",
  13264=>"101011100",
  13265=>"111110101",
  13266=>"111110111",
  13267=>"010110000",
  13268=>"010011011",
  13269=>"101011001",
  13270=>"010000010",
  13271=>"100110011",
  13272=>"100010010",
  13273=>"111100000",
  13274=>"010111101",
  13275=>"011101000",
  13276=>"111010101",
  13277=>"001011100",
  13278=>"000001000",
  13279=>"100000101",
  13280=>"000100101",
  13281=>"001100110",
  13282=>"010111000",
  13283=>"010001011",
  13284=>"000001001",
  13285=>"011000110",
  13286=>"110100101",
  13287=>"000110011",
  13288=>"001101011",
  13289=>"110110000",
  13290=>"111001011",
  13291=>"011001011",
  13292=>"111110001",
  13293=>"010001101",
  13294=>"101011100",
  13295=>"110110001",
  13296=>"111010000",
  13297=>"001010000",
  13298=>"101010011",
  13299=>"011100110",
  13300=>"110011011",
  13301=>"010010110",
  13302=>"111000111",
  13303=>"000001111",
  13304=>"010010001",
  13305=>"111111011",
  13306=>"111100111",
  13307=>"000111101",
  13308=>"010000001",
  13309=>"111101111",
  13310=>"110111101",
  13311=>"001011010",
  13312=>"110011010",
  13313=>"100001100",
  13314=>"101000011",
  13315=>"101100110",
  13316=>"110011100",
  13317=>"100011110",
  13318=>"001110010",
  13319=>"110111011",
  13320=>"010000100",
  13321=>"000000000",
  13322=>"111000011",
  13323=>"011110110",
  13324=>"011011000",
  13325=>"010011011",
  13326=>"011010100",
  13327=>"100001111",
  13328=>"111101010",
  13329=>"111101001",
  13330=>"100100001",
  13331=>"100010010",
  13332=>"111011011",
  13333=>"100011011",
  13334=>"010111011",
  13335=>"001100100",
  13336=>"000001100",
  13337=>"010010011",
  13338=>"101010000",
  13339=>"110001001",
  13340=>"100111011",
  13341=>"011001001",
  13342=>"011001111",
  13343=>"100110111",
  13344=>"111100110",
  13345=>"001010001",
  13346=>"000100010",
  13347=>"001001111",
  13348=>"010101011",
  13349=>"011000110",
  13350=>"011000001",
  13351=>"101001111",
  13352=>"100110011",
  13353=>"000100110",
  13354=>"011001010",
  13355=>"100100011",
  13356=>"101011110",
  13357=>"000111000",
  13358=>"001100111",
  13359=>"010000110",
  13360=>"101010000",
  13361=>"011011011",
  13362=>"010010001",
  13363=>"100111000",
  13364=>"111010100",
  13365=>"001010010",
  13366=>"110000000",
  13367=>"011110110",
  13368=>"000010111",
  13369=>"000000101",
  13370=>"011001001",
  13371=>"111111011",
  13372=>"110111111",
  13373=>"011111001",
  13374=>"110011111",
  13375=>"010101010",
  13376=>"110111001",
  13377=>"011001001",
  13378=>"010101100",
  13379=>"001100010",
  13380=>"100000000",
  13381=>"001010011",
  13382=>"001011011",
  13383=>"111011101",
  13384=>"000111010",
  13385=>"101110010",
  13386=>"101101010",
  13387=>"101000111",
  13388=>"001101111",
  13389=>"100011100",
  13390=>"111100010",
  13391=>"000000110",
  13392=>"111101101",
  13393=>"100011100",
  13394=>"111001001",
  13395=>"101000110",
  13396=>"111110111",
  13397=>"100100000",
  13398=>"010001111",
  13399=>"000110001",
  13400=>"111010110",
  13401=>"110100000",
  13402=>"101101001",
  13403=>"001111110",
  13404=>"100110001",
  13405=>"011100100",
  13406=>"000011101",
  13407=>"010010111",
  13408=>"100000001",
  13409=>"011000011",
  13410=>"100111011",
  13411=>"110000111",
  13412=>"010110101",
  13413=>"000101100",
  13414=>"101010110",
  13415=>"111111101",
  13416=>"100000100",
  13417=>"000011000",
  13418=>"110111100",
  13419=>"010111100",
  13420=>"010010100",
  13421=>"110110110",
  13422=>"100110001",
  13423=>"000001001",
  13424=>"111001100",
  13425=>"101110001",
  13426=>"011000111",
  13427=>"001110101",
  13428=>"011101101",
  13429=>"111011011",
  13430=>"010010010",
  13431=>"110111100",
  13432=>"111010010",
  13433=>"110100110",
  13434=>"000101111",
  13435=>"100000000",
  13436=>"000010011",
  13437=>"110011111",
  13438=>"001000010",
  13439=>"110011111",
  13440=>"111011110",
  13441=>"001010111",
  13442=>"100011010",
  13443=>"100001010",
  13444=>"100010010",
  13445=>"001100011",
  13446=>"111110101",
  13447=>"000101111",
  13448=>"000011010",
  13449=>"011011100",
  13450=>"111000000",
  13451=>"001100010",
  13452=>"110000001",
  13453=>"111011010",
  13454=>"010110111",
  13455=>"010100100",
  13456=>"110000010",
  13457=>"000011000",
  13458=>"001000010",
  13459=>"101001110",
  13460=>"010100101",
  13461=>"001010100",
  13462=>"000101110",
  13463=>"001011001",
  13464=>"010110101",
  13465=>"111011101",
  13466=>"110111011",
  13467=>"101001100",
  13468=>"101100100",
  13469=>"001111000",
  13470=>"110011010",
  13471=>"110011101",
  13472=>"010111111",
  13473=>"010111000",
  13474=>"100100001",
  13475=>"101101101",
  13476=>"011100110",
  13477=>"100001101",
  13478=>"100000010",
  13479=>"000100010",
  13480=>"110110100",
  13481=>"100011111",
  13482=>"011010100",
  13483=>"110100001",
  13484=>"000010110",
  13485=>"011010111",
  13486=>"000101100",
  13487=>"000100011",
  13488=>"111110111",
  13489=>"110011001",
  13490=>"101101000",
  13491=>"001110111",
  13492=>"010001101",
  13493=>"011010000",
  13494=>"010011010",
  13495=>"001011110",
  13496=>"110000010",
  13497=>"011000001",
  13498=>"111001110",
  13499=>"000110000",
  13500=>"101101011",
  13501=>"110010011",
  13502=>"111001010",
  13503=>"011101000",
  13504=>"011101011",
  13505=>"110100000",
  13506=>"001101010",
  13507=>"010100010",
  13508=>"001100010",
  13509=>"001000011",
  13510=>"000010100",
  13511=>"110010100",
  13512=>"100110011",
  13513=>"101000111",
  13514=>"100001000",
  13515=>"001001010",
  13516=>"101011100",
  13517=>"001110111",
  13518=>"100111011",
  13519=>"101111101",
  13520=>"000100011",
  13521=>"111101000",
  13522=>"100100110",
  13523=>"000110110",
  13524=>"100010000",
  13525=>"011101001",
  13526=>"001000100",
  13527=>"101001011",
  13528=>"100001100",
  13529=>"100001111",
  13530=>"101001101",
  13531=>"111010010",
  13532=>"001011011",
  13533=>"110111110",
  13534=>"010001000",
  13535=>"011110011",
  13536=>"000100010",
  13537=>"011010100",
  13538=>"001001000",
  13539=>"110011000",
  13540=>"110111101",
  13541=>"011100111",
  13542=>"010101101",
  13543=>"110011111",
  13544=>"101010001",
  13545=>"001011101",
  13546=>"100001001",
  13547=>"000101010",
  13548=>"011110000",
  13549=>"101101101",
  13550=>"010010011",
  13551=>"000001110",
  13552=>"101010100",
  13553=>"010100101",
  13554=>"111011001",
  13555=>"001101100",
  13556=>"111010110",
  13557=>"100100011",
  13558=>"101011011",
  13559=>"111000110",
  13560=>"100011110",
  13561=>"110111000",
  13562=>"100001000",
  13563=>"110000010",
  13564=>"110111101",
  13565=>"110011001",
  13566=>"001101100",
  13567=>"001100111",
  13568=>"100101100",
  13569=>"011100000",
  13570=>"001001000",
  13571=>"011010111",
  13572=>"111011110",
  13573=>"010010000",
  13574=>"101111100",
  13575=>"110011010",
  13576=>"011011101",
  13577=>"100100011",
  13578=>"010010001",
  13579=>"101001111",
  13580=>"001010010",
  13581=>"000000001",
  13582=>"011011000",
  13583=>"111111011",
  13584=>"110011111",
  13585=>"001011100",
  13586=>"100001110",
  13587=>"110000011",
  13588=>"110000000",
  13589=>"001000000",
  13590=>"000111110",
  13591=>"001110101",
  13592=>"110110101",
  13593=>"110110111",
  13594=>"110010100",
  13595=>"010100101",
  13596=>"001100100",
  13597=>"000101000",
  13598=>"010100011",
  13599=>"010010110",
  13600=>"010010010",
  13601=>"011100110",
  13602=>"000100101",
  13603=>"001010100",
  13604=>"101011101",
  13605=>"011101110",
  13606=>"110111101",
  13607=>"011010011",
  13608=>"001001101",
  13609=>"110110010",
  13610=>"010110101",
  13611=>"111110011",
  13612=>"111101101",
  13613=>"111110111",
  13614=>"111111100",
  13615=>"001101010",
  13616=>"000111000",
  13617=>"011011010",
  13618=>"110111101",
  13619=>"111101111",
  13620=>"011101001",
  13621=>"001011110",
  13622=>"001011101",
  13623=>"110001011",
  13624=>"100000010",
  13625=>"111100111",
  13626=>"101010001",
  13627=>"101010001",
  13628=>"111000101",
  13629=>"000111101",
  13630=>"001001101",
  13631=>"000110000",
  13632=>"001001011",
  13633=>"010101101",
  13634=>"000000000",
  13635=>"110110111",
  13636=>"110010100",
  13637=>"010001101",
  13638=>"011100000",
  13639=>"010011100",
  13640=>"111100010",
  13641=>"011000000",
  13642=>"111001100",
  13643=>"110110001",
  13644=>"111101111",
  13645=>"100100000",
  13646=>"111001111",
  13647=>"101111110",
  13648=>"101000111",
  13649=>"111110101",
  13650=>"010010111",
  13651=>"001011001",
  13652=>"000101101",
  13653=>"011100101",
  13654=>"010011101",
  13655=>"111100010",
  13656=>"011111000",
  13657=>"111010100",
  13658=>"111010000",
  13659=>"110011011",
  13660=>"110001010",
  13661=>"011111000",
  13662=>"111101011",
  13663=>"010100011",
  13664=>"110000110",
  13665=>"000010011",
  13666=>"110000110",
  13667=>"010111010",
  13668=>"101110001",
  13669=>"001001011",
  13670=>"001100100",
  13671=>"101101110",
  13672=>"000111111",
  13673=>"011101100",
  13674=>"000001001",
  13675=>"010101011",
  13676=>"110110110",
  13677=>"011011011",
  13678=>"001011111",
  13679=>"011011011",
  13680=>"000001010",
  13681=>"101110111",
  13682=>"100100100",
  13683=>"101010101",
  13684=>"000001110",
  13685=>"001000010",
  13686=>"100101100",
  13687=>"110000101",
  13688=>"010000000",
  13689=>"000110010",
  13690=>"101000110",
  13691=>"100111010",
  13692=>"001101000",
  13693=>"000101000",
  13694=>"101000011",
  13695=>"010101010",
  13696=>"010000111",
  13697=>"100100100",
  13698=>"110001111",
  13699=>"011001110",
  13700=>"010111011",
  13701=>"100011000",
  13702=>"111100110",
  13703=>"100001000",
  13704=>"111001001",
  13705=>"001100101",
  13706=>"000001000",
  13707=>"000000111",
  13708=>"100001010",
  13709=>"000100011",
  13710=>"001001101",
  13711=>"001110100",
  13712=>"000000011",
  13713=>"001001000",
  13714=>"100101101",
  13715=>"100111011",
  13716=>"111101010",
  13717=>"010000101",
  13718=>"001000001",
  13719=>"001110101",
  13720=>"101110011",
  13721=>"011100010",
  13722=>"101001100",
  13723=>"010001110",
  13724=>"111111001",
  13725=>"110000111",
  13726=>"110101001",
  13727=>"111110111",
  13728=>"000000101",
  13729=>"101010111",
  13730=>"111111011",
  13731=>"000110110",
  13732=>"000100000",
  13733=>"111111101",
  13734=>"000001110",
  13735=>"010011000",
  13736=>"110110001",
  13737=>"101011011",
  13738=>"011101001",
  13739=>"100110001",
  13740=>"001100011",
  13741=>"101000000",
  13742=>"001101111",
  13743=>"001111101",
  13744=>"111100101",
  13745=>"010111000",
  13746=>"001001101",
  13747=>"011010011",
  13748=>"011110000",
  13749=>"111101000",
  13750=>"000100111",
  13751=>"011100110",
  13752=>"111011111",
  13753=>"101101100",
  13754=>"000101101",
  13755=>"110111100",
  13756=>"111101100",
  13757=>"001101010",
  13758=>"000101001",
  13759=>"000101010",
  13760=>"000000010",
  13761=>"101100000",
  13762=>"011100011",
  13763=>"100011100",
  13764=>"001011110",
  13765=>"101100101",
  13766=>"001100111",
  13767=>"001001011",
  13768=>"011101010",
  13769=>"110110010",
  13770=>"101001001",
  13771=>"111110110",
  13772=>"110111001",
  13773=>"010100100",
  13774=>"101001000",
  13775=>"001111111",
  13776=>"010101001",
  13777=>"000110001",
  13778=>"111010000",
  13779=>"110101100",
  13780=>"101111100",
  13781=>"001001001",
  13782=>"011000001",
  13783=>"010110001",
  13784=>"001110111",
  13785=>"110011100",
  13786=>"000011000",
  13787=>"001001010",
  13788=>"111010000",
  13789=>"100100110",
  13790=>"110001010",
  13791=>"111100000",
  13792=>"111011011",
  13793=>"111100111",
  13794=>"110010111",
  13795=>"001000000",
  13796=>"101110010",
  13797=>"101101000",
  13798=>"011010100",
  13799=>"010111001",
  13800=>"100111111",
  13801=>"011101111",
  13802=>"101111001",
  13803=>"110110111",
  13804=>"000010000",
  13805=>"010100100",
  13806=>"111110111",
  13807=>"000000000",
  13808=>"111111101",
  13809=>"001000110",
  13810=>"110101100",
  13811=>"010001000",
  13812=>"111000011",
  13813=>"010100100",
  13814=>"011001101",
  13815=>"101111101",
  13816=>"100111110",
  13817=>"111111111",
  13818=>"000010111",
  13819=>"010011101",
  13820=>"110001111",
  13821=>"010110110",
  13822=>"110101010",
  13823=>"011100010",
  13824=>"100001101",
  13825=>"111111000",
  13826=>"110111010",
  13827=>"011000110",
  13828=>"000010111",
  13829=>"010110101",
  13830=>"001100111",
  13831=>"111001101",
  13832=>"101111100",
  13833=>"001011111",
  13834=>"000001101",
  13835=>"110010100",
  13836=>"000101010",
  13837=>"001000100",
  13838=>"100110101",
  13839=>"011001101",
  13840=>"000010001",
  13841=>"000000101",
  13842=>"111001110",
  13843=>"100110101",
  13844=>"010001000",
  13845=>"100110100",
  13846=>"100111101",
  13847=>"101011111",
  13848=>"100110110",
  13849=>"100010010",
  13850=>"101011000",
  13851=>"111000111",
  13852=>"100100010",
  13853=>"001110001",
  13854=>"101001011",
  13855=>"011101000",
  13856=>"101000111",
  13857=>"000100001",
  13858=>"001100100",
  13859=>"010011110",
  13860=>"001001100",
  13861=>"010100001",
  13862=>"010101010",
  13863=>"001010011",
  13864=>"000010000",
  13865=>"110110100",
  13866=>"111111100",
  13867=>"001000001",
  13868=>"010110001",
  13869=>"011100100",
  13870=>"010000100",
  13871=>"100010110",
  13872=>"100110000",
  13873=>"111011111",
  13874=>"001100010",
  13875=>"001101111",
  13876=>"101011100",
  13877=>"100011100",
  13878=>"101100111",
  13879=>"000000010",
  13880=>"110000100",
  13881=>"100111111",
  13882=>"001100101",
  13883=>"101101010",
  13884=>"110101010",
  13885=>"100111001",
  13886=>"010010001",
  13887=>"111010100",
  13888=>"010011100",
  13889=>"001010001",
  13890=>"100100111",
  13891=>"100001010",
  13892=>"101010110",
  13893=>"100100101",
  13894=>"111110111",
  13895=>"100001101",
  13896=>"010011111",
  13897=>"110000001",
  13898=>"000010101",
  13899=>"001100000",
  13900=>"011110001",
  13901=>"000110100",
  13902=>"010001101",
  13903=>"100110011",
  13904=>"010111111",
  13905=>"000000000",
  13906=>"100110110",
  13907=>"011000000",
  13908=>"000001011",
  13909=>"011010000",
  13910=>"001100100",
  13911=>"010101101",
  13912=>"000010100",
  13913=>"101100010",
  13914=>"111011001",
  13915=>"101000001",
  13916=>"100010111",
  13917=>"010010011",
  13918=>"000100110",
  13919=>"001110000",
  13920=>"001101010",
  13921=>"000001010",
  13922=>"010110110",
  13923=>"010010110",
  13924=>"110000100",
  13925=>"000111110",
  13926=>"110111111",
  13927=>"011000000",
  13928=>"110000011",
  13929=>"011101111",
  13930=>"110010100",
  13931=>"011010111",
  13932=>"101110110",
  13933=>"100000110",
  13934=>"000110011",
  13935=>"111100001",
  13936=>"110011011",
  13937=>"110111110",
  13938=>"100101110",
  13939=>"101110111",
  13940=>"101100000",
  13941=>"100000010",
  13942=>"110100011",
  13943=>"011011000",
  13944=>"100101001",
  13945=>"001100101",
  13946=>"001011100",
  13947=>"101100001",
  13948=>"100110001",
  13949=>"100101000",
  13950=>"001000111",
  13951=>"011111100",
  13952=>"011011000",
  13953=>"111010010",
  13954=>"111001111",
  13955=>"111010101",
  13956=>"100001111",
  13957=>"101011110",
  13958=>"110011111",
  13959=>"010011010",
  13960=>"001000111",
  13961=>"001100010",
  13962=>"011111101",
  13963=>"100101100",
  13964=>"111101110",
  13965=>"101000000",
  13966=>"000011111",
  13967=>"111111101",
  13968=>"011111011",
  13969=>"011110110",
  13970=>"111011010",
  13971=>"100011101",
  13972=>"000010000",
  13973=>"000010011",
  13974=>"010000111",
  13975=>"110011000",
  13976=>"101110001",
  13977=>"011110101",
  13978=>"010101101",
  13979=>"000100100",
  13980=>"000110000",
  13981=>"100111010",
  13982=>"100101111",
  13983=>"011000111",
  13984=>"000001010",
  13985=>"011010110",
  13986=>"010000010",
  13987=>"001011110",
  13988=>"000110101",
  13989=>"011100010",
  13990=>"111000111",
  13991=>"001110100",
  13992=>"100100101",
  13993=>"101001100",
  13994=>"001010001",
  13995=>"111101100",
  13996=>"001000000",
  13997=>"001011010",
  13998=>"001000100",
  13999=>"101000111",
  14000=>"101100011",
  14001=>"101101110",
  14002=>"110001011",
  14003=>"111001100",
  14004=>"000100101",
  14005=>"111010111",
  14006=>"001010010",
  14007=>"010011011",
  14008=>"000001100",
  14009=>"110110111",
  14010=>"001100010",
  14011=>"111000110",
  14012=>"100001011",
  14013=>"011000111",
  14014=>"011000011",
  14015=>"010100100",
  14016=>"100111011",
  14017=>"111101011",
  14018=>"111000111",
  14019=>"101000110",
  14020=>"101101000",
  14021=>"101100111",
  14022=>"001001111",
  14023=>"010001011",
  14024=>"000010011",
  14025=>"110011111",
  14026=>"010001001",
  14027=>"011011001",
  14028=>"100001101",
  14029=>"000010110",
  14030=>"001010010",
  14031=>"101101111",
  14032=>"000001000",
  14033=>"100111100",
  14034=>"000001111",
  14035=>"100110111",
  14036=>"000110110",
  14037=>"000101111",
  14038=>"110011000",
  14039=>"100000100",
  14040=>"010000111",
  14041=>"111101000",
  14042=>"111111100",
  14043=>"000010000",
  14044=>"110100111",
  14045=>"011110000",
  14046=>"001001010",
  14047=>"101000000",
  14048=>"011101000",
  14049=>"001001111",
  14050=>"000111010",
  14051=>"000001000",
  14052=>"110100000",
  14053=>"101101001",
  14054=>"011011000",
  14055=>"011001111",
  14056=>"000000111",
  14057=>"100101000",
  14058=>"101001010",
  14059=>"101000001",
  14060=>"001011011",
  14061=>"110010111",
  14062=>"111111111",
  14063=>"001111001",
  14064=>"111100111",
  14065=>"111101001",
  14066=>"111000010",
  14067=>"010011100",
  14068=>"111110110",
  14069=>"011101011",
  14070=>"101101100",
  14071=>"010000001",
  14072=>"110000111",
  14073=>"101011100",
  14074=>"000000111",
  14075=>"001110110",
  14076=>"110010000",
  14077=>"000000001",
  14078=>"111001111",
  14079=>"101001011",
  14080=>"111111010",
  14081=>"000010110",
  14082=>"100100000",
  14083=>"010001100",
  14084=>"100110101",
  14085=>"001011010",
  14086=>"011101100",
  14087=>"001100110",
  14088=>"010010100",
  14089=>"111111101",
  14090=>"000111001",
  14091=>"011111111",
  14092=>"101001100",
  14093=>"111001110",
  14094=>"110000010",
  14095=>"111010010",
  14096=>"101110100",
  14097=>"100010000",
  14098=>"101100000",
  14099=>"111000101",
  14100=>"010010011",
  14101=>"110010101",
  14102=>"111011111",
  14103=>"101101110",
  14104=>"010010001",
  14105=>"110011011",
  14106=>"110001001",
  14107=>"011100100",
  14108=>"000110111",
  14109=>"110000111",
  14110=>"001011101",
  14111=>"011010011",
  14112=>"111000001",
  14113=>"111111000",
  14114=>"000000010",
  14115=>"011000110",
  14116=>"100011011",
  14117=>"101001011",
  14118=>"110100101",
  14119=>"001011100",
  14120=>"001000100",
  14121=>"110110010",
  14122=>"101010100",
  14123=>"111011010",
  14124=>"000100101",
  14125=>"111011001",
  14126=>"000110110",
  14127=>"001101010",
  14128=>"010011111",
  14129=>"111111111",
  14130=>"001011100",
  14131=>"110111101",
  14132=>"100110111",
  14133=>"100000101",
  14134=>"100111010",
  14135=>"011101001",
  14136=>"011001110",
  14137=>"001101000",
  14138=>"010110100",
  14139=>"110000101",
  14140=>"100001101",
  14141=>"101111010",
  14142=>"001010100",
  14143=>"101100101",
  14144=>"111000000",
  14145=>"111110100",
  14146=>"101011001",
  14147=>"011111010",
  14148=>"011000000",
  14149=>"000100100",
  14150=>"101011100",
  14151=>"111111100",
  14152=>"101111001",
  14153=>"000101010",
  14154=>"011001001",
  14155=>"101100011",
  14156=>"011111001",
  14157=>"110010100",
  14158=>"001000100",
  14159=>"110111010",
  14160=>"011011011",
  14161=>"101110010",
  14162=>"010000001",
  14163=>"010000111",
  14164=>"011001101",
  14165=>"010100011",
  14166=>"010011110",
  14167=>"110100001",
  14168=>"000111001",
  14169=>"000011011",
  14170=>"001010011",
  14171=>"100101100",
  14172=>"000011110",
  14173=>"101001101",
  14174=>"000100101",
  14175=>"010001100",
  14176=>"000110010",
  14177=>"010010111",
  14178=>"110011100",
  14179=>"011111111",
  14180=>"010001111",
  14181=>"000111000",
  14182=>"111000110",
  14183=>"101111111",
  14184=>"110101011",
  14185=>"101001101",
  14186=>"011001100",
  14187=>"000010110",
  14188=>"110110010",
  14189=>"000010111",
  14190=>"101011001",
  14191=>"100111010",
  14192=>"000111010",
  14193=>"000011101",
  14194=>"101001011",
  14195=>"000100101",
  14196=>"101111011",
  14197=>"111100000",
  14198=>"011001111",
  14199=>"000110110",
  14200=>"010011001",
  14201=>"101011001",
  14202=>"110111011",
  14203=>"000110101",
  14204=>"000001001",
  14205=>"111110111",
  14206=>"110001100",
  14207=>"101111111",
  14208=>"001100010",
  14209=>"001000101",
  14210=>"011101001",
  14211=>"000100100",
  14212=>"010011111",
  14213=>"010101101",
  14214=>"011000000",
  14215=>"101011010",
  14216=>"010001010",
  14217=>"000000011",
  14218=>"000001000",
  14219=>"110111101",
  14220=>"100001001",
  14221=>"101011101",
  14222=>"000010110",
  14223=>"100010111",
  14224=>"001110000",
  14225=>"010000110",
  14226=>"110100010",
  14227=>"001010100",
  14228=>"110100100",
  14229=>"101101001",
  14230=>"101111111",
  14231=>"100010000",
  14232=>"111011111",
  14233=>"111101010",
  14234=>"010001101",
  14235=>"100111111",
  14236=>"010101110",
  14237=>"100001001",
  14238=>"101101100",
  14239=>"000010011",
  14240=>"011101101",
  14241=>"000000111",
  14242=>"001010111",
  14243=>"000101011",
  14244=>"101000000",
  14245=>"111001101",
  14246=>"100000101",
  14247=>"010001010",
  14248=>"010000010",
  14249=>"001000111",
  14250=>"010001001",
  14251=>"010000111",
  14252=>"001010010",
  14253=>"110111111",
  14254=>"000011010",
  14255=>"011010000",
  14256=>"010101101",
  14257=>"111000011",
  14258=>"111101100",
  14259=>"111010101",
  14260=>"001001110",
  14261=>"101111101",
  14262=>"010010111",
  14263=>"000010011",
  14264=>"110100101",
  14265=>"110011101",
  14266=>"111100101",
  14267=>"101000100",
  14268=>"001010010",
  14269=>"000100000",
  14270=>"011010100",
  14271=>"111101001",
  14272=>"110110101",
  14273=>"111101101",
  14274=>"101101011",
  14275=>"010001000",
  14276=>"000000111",
  14277=>"101000010",
  14278=>"100110010",
  14279=>"000110011",
  14280=>"011100110",
  14281=>"011110111",
  14282=>"111000111",
  14283=>"100000000",
  14284=>"001001011",
  14285=>"110111010",
  14286=>"011111000",
  14287=>"001011000",
  14288=>"010101111",
  14289=>"110100101",
  14290=>"100010100",
  14291=>"111100110",
  14292=>"111001101",
  14293=>"110110110",
  14294=>"000000110",
  14295=>"011000001",
  14296=>"011011010",
  14297=>"010110111",
  14298=>"100111110",
  14299=>"110101111",
  14300=>"010101111",
  14301=>"000101000",
  14302=>"110110011",
  14303=>"101110100",
  14304=>"001001001",
  14305=>"100000001",
  14306=>"101101110",
  14307=>"100010001",
  14308=>"101100110",
  14309=>"110100000",
  14310=>"000111101",
  14311=>"001100010",
  14312=>"100101111",
  14313=>"111111101",
  14314=>"001100000",
  14315=>"010100001",
  14316=>"000101110",
  14317=>"000000101",
  14318=>"011101101",
  14319=>"001100100",
  14320=>"011010111",
  14321=>"011101111",
  14322=>"000001100",
  14323=>"000011011",
  14324=>"000100100",
  14325=>"001001110",
  14326=>"010011001",
  14327=>"100001110",
  14328=>"101111010",
  14329=>"100101101",
  14330=>"111011101",
  14331=>"111011111",
  14332=>"100010011",
  14333=>"110111111",
  14334=>"001001100",
  14335=>"100101111",
  14336=>"010100101",
  14337=>"111000000",
  14338=>"111001000",
  14339=>"000000010",
  14340=>"010000110",
  14341=>"111010011",
  14342=>"010010101",
  14343=>"110011110",
  14344=>"111011110",
  14345=>"000001000",
  14346=>"111000001",
  14347=>"111110101",
  14348=>"001001101",
  14349=>"110101010",
  14350=>"010000010",
  14351=>"100010100",
  14352=>"001010001",
  14353=>"010001100",
  14354=>"010011001",
  14355=>"111111000",
  14356=>"101001100",
  14357=>"111100001",
  14358=>"010111111",
  14359=>"000100111",
  14360=>"100010100",
  14361=>"011010000",
  14362=>"010101001",
  14363=>"010100010",
  14364=>"011101101",
  14365=>"110010000",
  14366=>"110100101",
  14367=>"101100100",
  14368=>"101000110",
  14369=>"010110001",
  14370=>"110101010",
  14371=>"110111111",
  14372=>"100110000",
  14373=>"011100000",
  14374=>"100011010",
  14375=>"000111011",
  14376=>"101100101",
  14377=>"101000001",
  14378=>"011111110",
  14379=>"100010110",
  14380=>"000011011",
  14381=>"001001101",
  14382=>"101011101",
  14383=>"111001101",
  14384=>"001001111",
  14385=>"110110110",
  14386=>"000010010",
  14387=>"001110001",
  14388=>"111100111",
  14389=>"101110000",
  14390=>"011110110",
  14391=>"010110001",
  14392=>"011010010",
  14393=>"110100110",
  14394=>"001000110",
  14395=>"000010101",
  14396=>"101001110",
  14397=>"000000101",
  14398=>"111110011",
  14399=>"011001101",
  14400=>"001101100",
  14401=>"001010100",
  14402=>"111110101",
  14403=>"011101010",
  14404=>"111001101",
  14405=>"110011000",
  14406=>"010000111",
  14407=>"100100000",
  14408=>"101000111",
  14409=>"000110010",
  14410=>"001000100",
  14411=>"100000011",
  14412=>"111111100",
  14413=>"100110111",
  14414=>"110001000",
  14415=>"110111100",
  14416=>"111110110",
  14417=>"010011000",
  14418=>"010010011",
  14419=>"001110110",
  14420=>"101110101",
  14421=>"110111001",
  14422=>"010000110",
  14423=>"001001001",
  14424=>"001111100",
  14425=>"001000001",
  14426=>"000011101",
  14427=>"101101011",
  14428=>"001100011",
  14429=>"100101101",
  14430=>"001111000",
  14431=>"001000110",
  14432=>"001100010",
  14433=>"111001111",
  14434=>"000100000",
  14435=>"000101101",
  14436=>"100110000",
  14437=>"010110000",
  14438=>"001000011",
  14439=>"101111011",
  14440=>"101101100",
  14441=>"001111111",
  14442=>"101101001",
  14443=>"100010011",
  14444=>"111010100",
  14445=>"101110000",
  14446=>"000101011",
  14447=>"010110100",
  14448=>"011001001",
  14449=>"000100101",
  14450=>"110010010",
  14451=>"010110101",
  14452=>"111010001",
  14453=>"101101001",
  14454=>"011100010",
  14455=>"011000011",
  14456=>"000101101",
  14457=>"110000110",
  14458=>"001101111",
  14459=>"111101001",
  14460=>"100110000",
  14461=>"010010001",
  14462=>"101100111",
  14463=>"001011101",
  14464=>"101111011",
  14465=>"000010010",
  14466=>"100111000",
  14467=>"011010101",
  14468=>"111011101",
  14469=>"111001100",
  14470=>"011100001",
  14471=>"000010101",
  14472=>"100011100",
  14473=>"110011101",
  14474=>"000010010",
  14475=>"111101111",
  14476=>"001000000",
  14477=>"001000011",
  14478=>"111100010",
  14479=>"101000001",
  14480=>"111110110",
  14481=>"111011101",
  14482=>"000100111",
  14483=>"111000011",
  14484=>"001111000",
  14485=>"110001100",
  14486=>"001111000",
  14487=>"010010001",
  14488=>"110100010",
  14489=>"101101111",
  14490=>"110011111",
  14491=>"101010101",
  14492=>"000000001",
  14493=>"100110101",
  14494=>"001111000",
  14495=>"011100111",
  14496=>"001100011",
  14497=>"010010100",
  14498=>"110100100",
  14499=>"100000000",
  14500=>"000001011",
  14501=>"110100000",
  14502=>"011001011",
  14503=>"011000001",
  14504=>"001100111",
  14505=>"011000001",
  14506=>"111111111",
  14507=>"110111011",
  14508=>"001111001",
  14509=>"100100011",
  14510=>"100001011",
  14511=>"100101000",
  14512=>"011111111",
  14513=>"110011000",
  14514=>"110110101",
  14515=>"011110011",
  14516=>"010100101",
  14517=>"010101011",
  14518=>"110001001",
  14519=>"010101000",
  14520=>"000010001",
  14521=>"101100001",
  14522=>"101010111",
  14523=>"111100010",
  14524=>"101001001",
  14525=>"100001011",
  14526=>"100101010",
  14527=>"001110010",
  14528=>"100100010",
  14529=>"100101111",
  14530=>"111100111",
  14531=>"110011010",
  14532=>"011011000",
  14533=>"001011111",
  14534=>"101111010",
  14535=>"100110111",
  14536=>"100100110",
  14537=>"001001110",
  14538=>"111010110",
  14539=>"111010101",
  14540=>"111100100",
  14541=>"000110101",
  14542=>"011000011",
  14543=>"100010010",
  14544=>"000111010",
  14545=>"011011101",
  14546=>"010100010",
  14547=>"011010110",
  14548=>"011010100",
  14549=>"010000010",
  14550=>"111100100",
  14551=>"001000100",
  14552=>"001010111",
  14553=>"000010000",
  14554=>"001101110",
  14555=>"011110000",
  14556=>"101100001",
  14557=>"111000100",
  14558=>"100101111",
  14559=>"011011001",
  14560=>"010010110",
  14561=>"101011010",
  14562=>"010110011",
  14563=>"000101000",
  14564=>"001110100",
  14565=>"110101100",
  14566=>"000100101",
  14567=>"010110110",
  14568=>"101111100",
  14569=>"110001100",
  14570=>"011100000",
  14571=>"001000100",
  14572=>"101000101",
  14573=>"010111010",
  14574=>"110000011",
  14575=>"010001100",
  14576=>"001001000",
  14577=>"010111011",
  14578=>"001100001",
  14579=>"100110111",
  14580=>"001111100",
  14581=>"000000000",
  14582=>"101010110",
  14583=>"000110111",
  14584=>"001111100",
  14585=>"101011010",
  14586=>"000111110",
  14587=>"000011000",
  14588=>"100011010",
  14589=>"010101100",
  14590=>"100000000",
  14591=>"011111011",
  14592=>"100000001",
  14593=>"100010010",
  14594=>"000101000",
  14595=>"111011000",
  14596=>"110100110",
  14597=>"000010010",
  14598=>"111010111",
  14599=>"100010110",
  14600=>"000001000",
  14601=>"000100111",
  14602=>"001001111",
  14603=>"000101001",
  14604=>"001110011",
  14605=>"000001100",
  14606=>"011101011",
  14607=>"111011011",
  14608=>"011000000",
  14609=>"011000100",
  14610=>"110100010",
  14611=>"110101110",
  14612=>"101100011",
  14613=>"011100111",
  14614=>"010011000",
  14615=>"111101111",
  14616=>"001100110",
  14617=>"000100110",
  14618=>"100110000",
  14619=>"110100010",
  14620=>"010110011",
  14621=>"000001101",
  14622=>"111111111",
  14623=>"010000000",
  14624=>"001100011",
  14625=>"000001100",
  14626=>"001001011",
  14627=>"000000001",
  14628=>"100111010",
  14629=>"010111111",
  14630=>"011000011",
  14631=>"101010111",
  14632=>"111001110",
  14633=>"000110110",
  14634=>"111001011",
  14635=>"011011011",
  14636=>"100011000",
  14637=>"011011010",
  14638=>"010101111",
  14639=>"010101011",
  14640=>"011001001",
  14641=>"110001000",
  14642=>"011110111",
  14643=>"010011101",
  14644=>"101000000",
  14645=>"010001101",
  14646=>"110100100",
  14647=>"100111001",
  14648=>"000100010",
  14649=>"000101011",
  14650=>"110110100",
  14651=>"110111111",
  14652=>"000001101",
  14653=>"101110101",
  14654=>"001010000",
  14655=>"101100010",
  14656=>"100000010",
  14657=>"101010010",
  14658=>"011001000",
  14659=>"000111101",
  14660=>"110101111",
  14661=>"101111000",
  14662=>"000110100",
  14663=>"001111111",
  14664=>"100101111",
  14665=>"000100001",
  14666=>"110100110",
  14667=>"111000110",
  14668=>"000111011",
  14669=>"010001001",
  14670=>"101111111",
  14671=>"000110110",
  14672=>"001111001",
  14673=>"000010111",
  14674=>"001001011",
  14675=>"101100100",
  14676=>"001001001",
  14677=>"100001010",
  14678=>"011000111",
  14679=>"001110001",
  14680=>"010001110",
  14681=>"011110001",
  14682=>"010101110",
  14683=>"001110111",
  14684=>"100001111",
  14685=>"000110000",
  14686=>"101001101",
  14687=>"011111100",
  14688=>"100100101",
  14689=>"101100100",
  14690=>"100100110",
  14691=>"001000000",
  14692=>"101001011",
  14693=>"000100011",
  14694=>"011110100",
  14695=>"100011101",
  14696=>"000011001",
  14697=>"101010001",
  14698=>"000101100",
  14699=>"010110111",
  14700=>"100011001",
  14701=>"111111101",
  14702=>"011110011",
  14703=>"001011111",
  14704=>"111000111",
  14705=>"001111101",
  14706=>"101110010",
  14707=>"001011111",
  14708=>"010111100",
  14709=>"000001001",
  14710=>"010111010",
  14711=>"110101101",
  14712=>"010100011",
  14713=>"011110000",
  14714=>"110011010",
  14715=>"010000000",
  14716=>"011110010",
  14717=>"011000010",
  14718=>"101010111",
  14719=>"110001011",
  14720=>"000101010",
  14721=>"100001100",
  14722=>"010100110",
  14723=>"110010011",
  14724=>"110011100",
  14725=>"010100100",
  14726=>"010001110",
  14727=>"111011111",
  14728=>"000010111",
  14729=>"111011001",
  14730=>"011000010",
  14731=>"101100001",
  14732=>"111010010",
  14733=>"010111100",
  14734=>"001000110",
  14735=>"111111001",
  14736=>"101110001",
  14737=>"011010000",
  14738=>"010011000",
  14739=>"111111001",
  14740=>"001111111",
  14741=>"001001000",
  14742=>"001101010",
  14743=>"011110111",
  14744=>"111011100",
  14745=>"000101101",
  14746=>"110110111",
  14747=>"111000101",
  14748=>"100111011",
  14749=>"110101010",
  14750=>"011000101",
  14751=>"001100100",
  14752=>"001001111",
  14753=>"001010000",
  14754=>"101001000",
  14755=>"000000001",
  14756=>"101101010",
  14757=>"010001010",
  14758=>"110100110",
  14759=>"111110000",
  14760=>"000110001",
  14761=>"001010011",
  14762=>"110000011",
  14763=>"001110011",
  14764=>"010010100",
  14765=>"010111101",
  14766=>"101111010",
  14767=>"100101111",
  14768=>"001001001",
  14769=>"011110001",
  14770=>"101011000",
  14771=>"111111100",
  14772=>"010110010",
  14773=>"101011010",
  14774=>"001011110",
  14775=>"100110100",
  14776=>"111100110",
  14777=>"010100000",
  14778=>"000111111",
  14779=>"101001100",
  14780=>"011001011",
  14781=>"100110000",
  14782=>"011110111",
  14783=>"010010000",
  14784=>"010000011",
  14785=>"100010001",
  14786=>"101011001",
  14787=>"001110100",
  14788=>"100000000",
  14789=>"101011000",
  14790=>"101010001",
  14791=>"111000000",
  14792=>"000111100",
  14793=>"111000001",
  14794=>"011000000",
  14795=>"111011110",
  14796=>"000101001",
  14797=>"111000011",
  14798=>"110110001",
  14799=>"010111011",
  14800=>"100111111",
  14801=>"001011110",
  14802=>"111011001",
  14803=>"101111110",
  14804=>"101011111",
  14805=>"000001110",
  14806=>"101111011",
  14807=>"110111110",
  14808=>"011000110",
  14809=>"111011101",
  14810=>"101010001",
  14811=>"010000111",
  14812=>"010110000",
  14813=>"100011111",
  14814=>"111011100",
  14815=>"101000000",
  14816=>"100100111",
  14817=>"100010100",
  14818=>"111110110",
  14819=>"011000010",
  14820=>"011101001",
  14821=>"100110011",
  14822=>"000100100",
  14823=>"101010010",
  14824=>"001111101",
  14825=>"110101001",
  14826=>"010001010",
  14827=>"101101010",
  14828=>"111000101",
  14829=>"011001110",
  14830=>"100010100",
  14831=>"100001110",
  14832=>"100111001",
  14833=>"111001101",
  14834=>"000000111",
  14835=>"101001011",
  14836=>"111111001",
  14837=>"111111100",
  14838=>"011001000",
  14839=>"110111000",
  14840=>"111011001",
  14841=>"100001100",
  14842=>"000101001",
  14843=>"000110101",
  14844=>"000000001",
  14845=>"000100111",
  14846=>"000000110",
  14847=>"001010111",
  14848=>"110111101",
  14849=>"010001011",
  14850=>"000101010",
  14851=>"011111010",
  14852=>"100010111",
  14853=>"101000101",
  14854=>"111110110",
  14855=>"001110001",
  14856=>"101001011",
  14857=>"001000101",
  14858=>"010100000",
  14859=>"101111000",
  14860=>"001000010",
  14861=>"110110000",
  14862=>"110000100",
  14863=>"001110011",
  14864=>"011010010",
  14865=>"011111000",
  14866=>"111111011",
  14867=>"101001000",
  14868=>"011101110",
  14869=>"111110001",
  14870=>"001011011",
  14871=>"011110000",
  14872=>"000110011",
  14873=>"111100110",
  14874=>"010010101",
  14875=>"100000001",
  14876=>"011011001",
  14877=>"010000001",
  14878=>"101000011",
  14879=>"001010010",
  14880=>"110000111",
  14881=>"101111000",
  14882=>"001110101",
  14883=>"000011101",
  14884=>"000001101",
  14885=>"001111111",
  14886=>"101010111",
  14887=>"000011010",
  14888=>"000111000",
  14889=>"100010111",
  14890=>"010010001",
  14891=>"001110011",
  14892=>"111001000",
  14893=>"001000100",
  14894=>"100100001",
  14895=>"000100000",
  14896=>"111100111",
  14897=>"000000001",
  14898=>"111001101",
  14899=>"100101101",
  14900=>"110010001",
  14901=>"011101100",
  14902=>"000010000",
  14903=>"001011101",
  14904=>"101110011",
  14905=>"101010011",
  14906=>"100111110",
  14907=>"000101011",
  14908=>"000001101",
  14909=>"000001100",
  14910=>"010101010",
  14911=>"111111001",
  14912=>"010111001",
  14913=>"110011100",
  14914=>"111011110",
  14915=>"000101111",
  14916=>"011010100",
  14917=>"011000001",
  14918=>"111001011",
  14919=>"111000111",
  14920=>"000011000",
  14921=>"000000100",
  14922=>"111001110",
  14923=>"011000011",
  14924=>"111000111",
  14925=>"000101001",
  14926=>"100100100",
  14927=>"111101000",
  14928=>"100100101",
  14929=>"101101101",
  14930=>"110010001",
  14931=>"100000111",
  14932=>"011010100",
  14933=>"000010101",
  14934=>"000100000",
  14935=>"100000000",
  14936=>"011111111",
  14937=>"000111101",
  14938=>"010100011",
  14939=>"111111010",
  14940=>"010000111",
  14941=>"010011000",
  14942=>"011011100",
  14943=>"111001001",
  14944=>"110111010",
  14945=>"000000001",
  14946=>"001100001",
  14947=>"011110010",
  14948=>"010001111",
  14949=>"010111001",
  14950=>"110010011",
  14951=>"100100111",
  14952=>"001000000",
  14953=>"000000000",
  14954=>"010011111",
  14955=>"110011100",
  14956=>"000011110",
  14957=>"011110111",
  14958=>"001100000",
  14959=>"000101111",
  14960=>"101001011",
  14961=>"000111001",
  14962=>"110100011",
  14963=>"010110000",
  14964=>"001110001",
  14965=>"010100100",
  14966=>"000111100",
  14967=>"011001000",
  14968=>"100100111",
  14969=>"000111100",
  14970=>"101010100",
  14971=>"111001000",
  14972=>"101110001",
  14973=>"101000101",
  14974=>"001110010",
  14975=>"001100000",
  14976=>"101000100",
  14977=>"101111111",
  14978=>"110101111",
  14979=>"101010110",
  14980=>"010010100",
  14981=>"101001111",
  14982=>"101000101",
  14983=>"101111000",
  14984=>"011010000",
  14985=>"110111110",
  14986=>"111101101",
  14987=>"110010100",
  14988=>"101000111",
  14989=>"011000110",
  14990=>"001100011",
  14991=>"100100011",
  14992=>"100101110",
  14993=>"110111011",
  14994=>"111011100",
  14995=>"111000111",
  14996=>"010101101",
  14997=>"000010101",
  14998=>"110001001",
  14999=>"001001100",
  15000=>"110001100",
  15001=>"101110101",
  15002=>"000001010",
  15003=>"011010010",
  15004=>"111001101",
  15005=>"011111100",
  15006=>"000001111",
  15007=>"011010010",
  15008=>"111011010",
  15009=>"100111110",
  15010=>"111111010",
  15011=>"011110101",
  15012=>"001001000",
  15013=>"001101111",
  15014=>"010111000",
  15015=>"000101100",
  15016=>"010100000",
  15017=>"001100000",
  15018=>"100000001",
  15019=>"011001010",
  15020=>"100101101",
  15021=>"100100011",
  15022=>"010100000",
  15023=>"010001111",
  15024=>"000000001",
  15025=>"111011000",
  15026=>"011100100",
  15027=>"010000001",
  15028=>"101101010",
  15029=>"100000000",
  15030=>"001001011",
  15031=>"100101110",
  15032=>"000010100",
  15033=>"010101000",
  15034=>"001000010",
  15035=>"000000110",
  15036=>"001000111",
  15037=>"000101011",
  15038=>"101000011",
  15039=>"111000111",
  15040=>"011111100",
  15041=>"110010001",
  15042=>"001001000",
  15043=>"000101011",
  15044=>"111001000",
  15045=>"000011000",
  15046=>"001011001",
  15047=>"011111111",
  15048=>"000111111",
  15049=>"101001110",
  15050=>"101111110",
  15051=>"001100010",
  15052=>"011011010",
  15053=>"110001110",
  15054=>"001100111",
  15055=>"100100110",
  15056=>"011101111",
  15057=>"000001001",
  15058=>"010101001",
  15059=>"000111110",
  15060=>"000110010",
  15061=>"100101001",
  15062=>"100111110",
  15063=>"110100010",
  15064=>"100100011",
  15065=>"101100111",
  15066=>"010100100",
  15067=>"000010011",
  15068=>"011001100",
  15069=>"011001011",
  15070=>"110000110",
  15071=>"011001111",
  15072=>"110110110",
  15073=>"000011000",
  15074=>"111101100",
  15075=>"101111011",
  15076=>"000011000",
  15077=>"011100100",
  15078=>"011011001",
  15079=>"111111111",
  15080=>"101111101",
  15081=>"111111001",
  15082=>"101001010",
  15083=>"110100111",
  15084=>"010101011",
  15085=>"011110001",
  15086=>"000100110",
  15087=>"000011001",
  15088=>"011101010",
  15089=>"100001101",
  15090=>"011001100",
  15091=>"000010100",
  15092=>"011000111",
  15093=>"101001011",
  15094=>"101100010",
  15095=>"011111000",
  15096=>"001010100",
  15097=>"100000010",
  15098=>"101011011",
  15099=>"101011101",
  15100=>"001111010",
  15101=>"000010001",
  15102=>"100001001",
  15103=>"101101110",
  15104=>"000100100",
  15105=>"011101011",
  15106=>"111100000",
  15107=>"111001110",
  15108=>"011010100",
  15109=>"010010000",
  15110=>"000100010",
  15111=>"101100011",
  15112=>"000010101",
  15113=>"001110001",
  15114=>"010001110",
  15115=>"111100000",
  15116=>"010101101",
  15117=>"001111001",
  15118=>"101100001",
  15119=>"110110011",
  15120=>"100011001",
  15121=>"111000000",
  15122=>"111110101",
  15123=>"011110001",
  15124=>"010111100",
  15125=>"101011001",
  15126=>"000000111",
  15127=>"110100100",
  15128=>"111111111",
  15129=>"000000110",
  15130=>"111111000",
  15131=>"000111110",
  15132=>"010000011",
  15133=>"101111110",
  15134=>"011111110",
  15135=>"001101101",
  15136=>"010101111",
  15137=>"101100110",
  15138=>"111111100",
  15139=>"100100000",
  15140=>"001111111",
  15141=>"100111110",
  15142=>"010100001",
  15143=>"110110011",
  15144=>"010111011",
  15145=>"101010001",
  15146=>"000011000",
  15147=>"111001100",
  15148=>"101111010",
  15149=>"111000001",
  15150=>"010001001",
  15151=>"111001110",
  15152=>"100010000",
  15153=>"110001001",
  15154=>"000100001",
  15155=>"101010001",
  15156=>"110010000",
  15157=>"111110100",
  15158=>"000000000",
  15159=>"011010101",
  15160=>"110001111",
  15161=>"111000000",
  15162=>"101011100",
  15163=>"110101000",
  15164=>"100111001",
  15165=>"100000000",
  15166=>"000101010",
  15167=>"001010000",
  15168=>"010111110",
  15169=>"011111011",
  15170=>"011001101",
  15171=>"010110011",
  15172=>"001011100",
  15173=>"101101011",
  15174=>"000110001",
  15175=>"000011010",
  15176=>"100001010",
  15177=>"110101110",
  15178=>"100111010",
  15179=>"110011101",
  15180=>"111101011",
  15181=>"110011111",
  15182=>"011110101",
  15183=>"010001110",
  15184=>"000001101",
  15185=>"100100101",
  15186=>"001011111",
  15187=>"011101101",
  15188=>"110110111",
  15189=>"000011110",
  15190=>"100011010",
  15191=>"000000001",
  15192=>"100001100",
  15193=>"000011000",
  15194=>"000011010",
  15195=>"010110110",
  15196=>"110010100",
  15197=>"010011100",
  15198=>"010000011",
  15199=>"011000010",
  15200=>"001111000",
  15201=>"011100111",
  15202=>"010100101",
  15203=>"001111001",
  15204=>"111011111",
  15205=>"000100001",
  15206=>"001001101",
  15207=>"100001000",
  15208=>"101100011",
  15209=>"000000111",
  15210=>"101100101",
  15211=>"001100110",
  15212=>"111001000",
  15213=>"101100000",
  15214=>"011100110",
  15215=>"110101100",
  15216=>"110001010",
  15217=>"110100010",
  15218=>"100101001",
  15219=>"100010101",
  15220=>"000100001",
  15221=>"011100111",
  15222=>"110000110",
  15223=>"111010010",
  15224=>"100100111",
  15225=>"010001110",
  15226=>"011100011",
  15227=>"101111010",
  15228=>"001001011",
  15229=>"000011110",
  15230=>"011101100",
  15231=>"110010011",
  15232=>"101100111",
  15233=>"100101100",
  15234=>"100001111",
  15235=>"100011110",
  15236=>"001100001",
  15237=>"010010111",
  15238=>"010100010",
  15239=>"011010010",
  15240=>"011010000",
  15241=>"011101000",
  15242=>"001111000",
  15243=>"011111111",
  15244=>"111101001",
  15245=>"001010001",
  15246=>"111110110",
  15247=>"010001110",
  15248=>"101101010",
  15249=>"111101111",
  15250=>"000000000",
  15251=>"000110111",
  15252=>"110101111",
  15253=>"001111011",
  15254=>"000101010",
  15255=>"101011111",
  15256=>"001000010",
  15257=>"101111000",
  15258=>"111010001",
  15259=>"111100000",
  15260=>"110111110",
  15261=>"110111011",
  15262=>"011000000",
  15263=>"111111100",
  15264=>"100111110",
  15265=>"000111100",
  15266=>"010110101",
  15267=>"001111111",
  15268=>"000101100",
  15269=>"111100011",
  15270=>"001110001",
  15271=>"111011111",
  15272=>"000110010",
  15273=>"011010001",
  15274=>"011000110",
  15275=>"001010000",
  15276=>"001110101",
  15277=>"100000011",
  15278=>"111101111",
  15279=>"110101011",
  15280=>"001001110",
  15281=>"000101001",
  15282=>"000101001",
  15283=>"100101010",
  15284=>"010110101",
  15285=>"001010010",
  15286=>"111110000",
  15287=>"001001100",
  15288=>"111001100",
  15289=>"011001000",
  15290=>"000011000",
  15291=>"000000110",
  15292=>"101100111",
  15293=>"000001100",
  15294=>"010011100",
  15295=>"111000001",
  15296=>"001001101",
  15297=>"010100001",
  15298=>"011010001",
  15299=>"000110001",
  15300=>"011101010",
  15301=>"001001111",
  15302=>"001011111",
  15303=>"101101101",
  15304=>"100011100",
  15305=>"111100111",
  15306=>"100000001",
  15307=>"110110011",
  15308=>"011001100",
  15309=>"111000100",
  15310=>"010101011",
  15311=>"011010011",
  15312=>"010000111",
  15313=>"100100110",
  15314=>"110101001",
  15315=>"101100110",
  15316=>"011101011",
  15317=>"010110100",
  15318=>"001000011",
  15319=>"010110111",
  15320=>"111100110",
  15321=>"000111001",
  15322=>"101110100",
  15323=>"011001111",
  15324=>"111111011",
  15325=>"101111010",
  15326=>"110000101",
  15327=>"110001111",
  15328=>"110011111",
  15329=>"100011111",
  15330=>"011101110",
  15331=>"101011101",
  15332=>"110010010",
  15333=>"100101110",
  15334=>"111101111",
  15335=>"111001000",
  15336=>"010000101",
  15337=>"010000101",
  15338=>"111100111",
  15339=>"111000011",
  15340=>"001001110",
  15341=>"110100001",
  15342=>"101111111",
  15343=>"010100101",
  15344=>"110111010",
  15345=>"101000110",
  15346=>"101001000",
  15347=>"111001111",
  15348=>"000110110",
  15349=>"011000000",
  15350=>"011110011",
  15351=>"001111100",
  15352=>"000011000",
  15353=>"110000100",
  15354=>"101100111",
  15355=>"110011000",
  15356=>"011011111",
  15357=>"101100011",
  15358=>"001011000",
  15359=>"100100101",
  15360=>"010010000",
  15361=>"000000000",
  15362=>"110010101",
  15363=>"000000001",
  15364=>"100011000",
  15365=>"001110011",
  15366=>"010010010",
  15367=>"001010011",
  15368=>"101110011",
  15369=>"101010000",
  15370=>"100010111",
  15371=>"011111101",
  15372=>"110101001",
  15373=>"111101111",
  15374=>"110110001",
  15375=>"101000010",
  15376=>"111100011",
  15377=>"000100101",
  15378=>"110110000",
  15379=>"101001111",
  15380=>"011010111",
  15381=>"101000010",
  15382=>"111111111",
  15383=>"111110010",
  15384=>"101001000",
  15385=>"111001100",
  15386=>"011000110",
  15387=>"100011101",
  15388=>"101101101",
  15389=>"010011000",
  15390=>"110110111",
  15391=>"010101111",
  15392=>"011010010",
  15393=>"010001011",
  15394=>"110111101",
  15395=>"101100100",
  15396=>"000000110",
  15397=>"000000011",
  15398=>"010110110",
  15399=>"111010101",
  15400=>"011101111",
  15401=>"111110110",
  15402=>"110001111",
  15403=>"011111100",
  15404=>"101110011",
  15405=>"101101010",
  15406=>"000101111",
  15407=>"111111011",
  15408=>"010001101",
  15409=>"100101000",
  15410=>"110000001",
  15411=>"100100000",
  15412=>"101100000",
  15413=>"001111100",
  15414=>"110100001",
  15415=>"000101101",
  15416=>"101011101",
  15417=>"110111110",
  15418=>"010100001",
  15419=>"000110100",
  15420=>"100111101",
  15421=>"100100101",
  15422=>"011111111",
  15423=>"000000010",
  15424=>"011101010",
  15425=>"011110110",
  15426=>"110110110",
  15427=>"010011110",
  15428=>"110001101",
  15429=>"101100111",
  15430=>"000100100",
  15431=>"100001000",
  15432=>"001111101",
  15433=>"000110000",
  15434=>"100101101",
  15435=>"100000100",
  15436=>"101110001",
  15437=>"111011110",
  15438=>"011000011",
  15439=>"111101100",
  15440=>"111100011",
  15441=>"010001101",
  15442=>"010101000",
  15443=>"001000101",
  15444=>"001001011",
  15445=>"101100001",
  15446=>"011110001",
  15447=>"001011010",
  15448=>"101111111",
  15449=>"011111101",
  15450=>"110100000",
  15451=>"001000100",
  15452=>"111000110",
  15453=>"101001001",
  15454=>"100101110",
  15455=>"100010110",
  15456=>"010111110",
  15457=>"000011110",
  15458=>"011110110",
  15459=>"000010011",
  15460=>"000010000",
  15461=>"000011001",
  15462=>"100101011",
  15463=>"000101001",
  15464=>"010110100",
  15465=>"110101000",
  15466=>"101111001",
  15467=>"110110010",
  15468=>"111010101",
  15469=>"100101111",
  15470=>"001000110",
  15471=>"110101010",
  15472=>"111101100",
  15473=>"111000010",
  15474=>"111001000",
  15475=>"110001110",
  15476=>"011000011",
  15477=>"010111010",
  15478=>"011000100",
  15479=>"100011110",
  15480=>"100111101",
  15481=>"110011100",
  15482=>"101011110",
  15483=>"000101110",
  15484=>"110011011",
  15485=>"011111111",
  15486=>"100111101",
  15487=>"001111110",
  15488=>"000111100",
  15489=>"110101100",
  15490=>"101111000",
  15491=>"110000000",
  15492=>"101011000",
  15493=>"100110001",
  15494=>"111010001",
  15495=>"111111111",
  15496=>"011010101",
  15497=>"110111010",
  15498=>"100111010",
  15499=>"100010011",
  15500=>"000000011",
  15501=>"001110101",
  15502=>"101000010",
  15503=>"001011001",
  15504=>"111111011",
  15505=>"000001110",
  15506=>"000001010",
  15507=>"000011101",
  15508=>"110001010",
  15509=>"011011000",
  15510=>"101000001",
  15511=>"110010000",
  15512=>"011011000",
  15513=>"001001010",
  15514=>"101000000",
  15515=>"110110101",
  15516=>"000100011",
  15517=>"010110101",
  15518=>"110001001",
  15519=>"111100111",
  15520=>"001100000",
  15521=>"110010010",
  15522=>"101111001",
  15523=>"011010110",
  15524=>"100010011",
  15525=>"010110101",
  15526=>"001001011",
  15527=>"000100101",
  15528=>"111100100",
  15529=>"110001000",
  15530=>"011110001",
  15531=>"001000111",
  15532=>"011110000",
  15533=>"111010011",
  15534=>"010111110",
  15535=>"011101000",
  15536=>"100001111",
  15537=>"110110011",
  15538=>"110110111",
  15539=>"001010110",
  15540=>"001000000",
  15541=>"100001111",
  15542=>"011101110",
  15543=>"100011010",
  15544=>"100001101",
  15545=>"101101011",
  15546=>"101000110",
  15547=>"000100011",
  15548=>"111000001",
  15549=>"100101001",
  15550=>"001001001",
  15551=>"100011000",
  15552=>"001111000",
  15553=>"101011000",
  15554=>"110000000",
  15555=>"010011111",
  15556=>"111010100",
  15557=>"000111100",
  15558=>"011010000",
  15559=>"011111111",
  15560=>"000010101",
  15561=>"001100000",
  15562=>"110100111",
  15563=>"011010011",
  15564=>"000010011",
  15565=>"101111111",
  15566=>"001100000",
  15567=>"111010110",
  15568=>"001111101",
  15569=>"100101101",
  15570=>"010001111",
  15571=>"011111010",
  15572=>"111001110",
  15573=>"010110010",
  15574=>"100111001",
  15575=>"100111110",
  15576=>"100101000",
  15577=>"011110000",
  15578=>"101111110",
  15579=>"100001000",
  15580=>"001000000",
  15581=>"100000110",
  15582=>"111010011",
  15583=>"001000100",
  15584=>"010000000",
  15585=>"100100111",
  15586=>"011111011",
  15587=>"010000011",
  15588=>"000111010",
  15589=>"110110001",
  15590=>"101101110",
  15591=>"001101001",
  15592=>"111100010",
  15593=>"010011000",
  15594=>"101000100",
  15595=>"101110110",
  15596=>"011001010",
  15597=>"110110111",
  15598=>"111011011",
  15599=>"000100100",
  15600=>"010011111",
  15601=>"000110101",
  15602=>"000111000",
  15603=>"000110101",
  15604=>"110011010",
  15605=>"100101101",
  15606=>"101100001",
  15607=>"001011011",
  15608=>"100000111",
  15609=>"010101110",
  15610=>"000101110",
  15611=>"010111011",
  15612=>"000011001",
  15613=>"001001100",
  15614=>"001011010",
  15615=>"010111111",
  15616=>"101000001",
  15617=>"010100000",
  15618=>"011111110",
  15619=>"111010000",
  15620=>"111011101",
  15621=>"001001011",
  15622=>"011010110",
  15623=>"010001011",
  15624=>"000001010",
  15625=>"010110001",
  15626=>"101100111",
  15627=>"101101000",
  15628=>"001001101",
  15629=>"111101011",
  15630=>"010001111",
  15631=>"000100111",
  15632=>"101001011",
  15633=>"011000101",
  15634=>"101011010",
  15635=>"101000011",
  15636=>"000110010",
  15637=>"101011100",
  15638=>"101100110",
  15639=>"110010111",
  15640=>"111001101",
  15641=>"001111111",
  15642=>"100000100",
  15643=>"000101001",
  15644=>"000110101",
  15645=>"000100010",
  15646=>"001000100",
  15647=>"011111110",
  15648=>"001111101",
  15649=>"011101000",
  15650=>"010111011",
  15651=>"100011001",
  15652=>"100101011",
  15653=>"000010010",
  15654=>"010110000",
  15655=>"001001110",
  15656=>"101100011",
  15657=>"010100000",
  15658=>"100111001",
  15659=>"001011110",
  15660=>"111101000",
  15661=>"000111010",
  15662=>"110000100",
  15663=>"011110011",
  15664=>"000010000",
  15665=>"011011101",
  15666=>"111101111",
  15667=>"000101110",
  15668=>"001000000",
  15669=>"010100100",
  15670=>"110111010",
  15671=>"101000110",
  15672=>"011010111",
  15673=>"110001001",
  15674=>"010000011",
  15675=>"010010100",
  15676=>"001000000",
  15677=>"000101100",
  15678=>"001101011",
  15679=>"010000001",
  15680=>"110110110",
  15681=>"100111111",
  15682=>"110000010",
  15683=>"011110100",
  15684=>"001000101",
  15685=>"110011011",
  15686=>"100100001",
  15687=>"100111011",
  15688=>"111011010",
  15689=>"000110001",
  15690=>"010011000",
  15691=>"100010001",
  15692=>"001001001",
  15693=>"100110101",
  15694=>"101100010",
  15695=>"000100011",
  15696=>"101011110",
  15697=>"100111110",
  15698=>"111110000",
  15699=>"111001001",
  15700=>"110010100",
  15701=>"011110111",
  15702=>"110100110",
  15703=>"000000110",
  15704=>"001000110",
  15705=>"001010001",
  15706=>"011110111",
  15707=>"001101110",
  15708=>"010011011",
  15709=>"000000011",
  15710=>"010100111",
  15711=>"000111001",
  15712=>"101011100",
  15713=>"100010010",
  15714=>"101001101",
  15715=>"011011100",
  15716=>"000111101",
  15717=>"110101101",
  15718=>"010000101",
  15719=>"100010000",
  15720=>"001010010",
  15721=>"101010001",
  15722=>"110110011",
  15723=>"100110110",
  15724=>"110011101",
  15725=>"011001100",
  15726=>"001001010",
  15727=>"111101101",
  15728=>"001011001",
  15729=>"111000101",
  15730=>"101010010",
  15731=>"111000001",
  15732=>"110101010",
  15733=>"110011110",
  15734=>"111011101",
  15735=>"110101110",
  15736=>"101100111",
  15737=>"000100100",
  15738=>"001000011",
  15739=>"100001111",
  15740=>"110100011",
  15741=>"011100000",
  15742=>"100101001",
  15743=>"101101111",
  15744=>"011100101",
  15745=>"000011110",
  15746=>"000001011",
  15747=>"110100011",
  15748=>"110010101",
  15749=>"011010101",
  15750=>"000010000",
  15751=>"100011101",
  15752=>"001000000",
  15753=>"111011100",
  15754=>"010001001",
  15755=>"001010011",
  15756=>"100001011",
  15757=>"111011001",
  15758=>"010101011",
  15759=>"010111011",
  15760=>"111110000",
  15761=>"111011101",
  15762=>"101001000",
  15763=>"001001101",
  15764=>"011010101",
  15765=>"000010111",
  15766=>"001000100",
  15767=>"101101000",
  15768=>"001011010",
  15769=>"100011001",
  15770=>"000010111",
  15771=>"111110011",
  15772=>"110001111",
  15773=>"001000011",
  15774=>"110000011",
  15775=>"000010001",
  15776=>"110100101",
  15777=>"111100110",
  15778=>"000010010",
  15779=>"110010100",
  15780=>"100011000",
  15781=>"000010001",
  15782=>"111101110",
  15783=>"011001111",
  15784=>"010110100",
  15785=>"010001110",
  15786=>"111111101",
  15787=>"010000010",
  15788=>"111110101",
  15789=>"011100010",
  15790=>"000100000",
  15791=>"100111010",
  15792=>"000010101",
  15793=>"010010100",
  15794=>"110011000",
  15795=>"100010110",
  15796=>"001110011",
  15797=>"010010011",
  15798=>"011110111",
  15799=>"011110001",
  15800=>"001000111",
  15801=>"101001000",
  15802=>"010001010",
  15803=>"001001010",
  15804=>"011010100",
  15805=>"000110101",
  15806=>"001001000",
  15807=>"101111010",
  15808=>"110101011",
  15809=>"111010000",
  15810=>"101111000",
  15811=>"110100000",
  15812=>"110000010",
  15813=>"010000000",
  15814=>"111000000",
  15815=>"101100001",
  15816=>"101101000",
  15817=>"100100000",
  15818=>"000110010",
  15819=>"111100001",
  15820=>"101100010",
  15821=>"001101101",
  15822=>"000100110",
  15823=>"001111110",
  15824=>"110110111",
  15825=>"001110011",
  15826=>"001111001",
  15827=>"000010010",
  15828=>"101110000",
  15829=>"110101000",
  15830=>"101111001",
  15831=>"010010001",
  15832=>"010100100",
  15833=>"111010110",
  15834=>"100010011",
  15835=>"100101001",
  15836=>"000010011",
  15837=>"010011101",
  15838=>"111111110",
  15839=>"010011101",
  15840=>"101110110",
  15841=>"000101011",
  15842=>"010001011",
  15843=>"001010101",
  15844=>"010000100",
  15845=>"010010011",
  15846=>"010110110",
  15847=>"111001011",
  15848=>"100010011",
  15849=>"001010001",
  15850=>"011111011",
  15851=>"000101000",
  15852=>"110111010",
  15853=>"110000000",
  15854=>"011110010",
  15855=>"011001010",
  15856=>"011000101",
  15857=>"010011010",
  15858=>"010100110",
  15859=>"100101101",
  15860=>"001000001",
  15861=>"100010010",
  15862=>"011101101",
  15863=>"110000101",
  15864=>"001110101",
  15865=>"111010100",
  15866=>"000010110",
  15867=>"010111101",
  15868=>"101000101",
  15869=>"110001110",
  15870=>"010111111",
  15871=>"000110100",
  15872=>"101101100",
  15873=>"101000010",
  15874=>"001111011",
  15875=>"000100100",
  15876=>"111100001",
  15877=>"100011011",
  15878=>"111100101",
  15879=>"111000110",
  15880=>"001100100",
  15881=>"111011101",
  15882=>"101011100",
  15883=>"010010011",
  15884=>"010001010",
  15885=>"110111111",
  15886=>"011010100",
  15887=>"001110101",
  15888=>"000101010",
  15889=>"110000111",
  15890=>"111010101",
  15891=>"001110001",
  15892=>"000010100",
  15893=>"110011010",
  15894=>"111001010",
  15895=>"001101011",
  15896=>"111101010",
  15897=>"100011100",
  15898=>"101110010",
  15899=>"010110101",
  15900=>"000101100",
  15901=>"111101101",
  15902=>"110010011",
  15903=>"001010101",
  15904=>"010110011",
  15905=>"001101100",
  15906=>"101010011",
  15907=>"111011000",
  15908=>"100000001",
  15909=>"111110101",
  15910=>"111000011",
  15911=>"110010100",
  15912=>"010100000",
  15913=>"111010111",
  15914=>"010010001",
  15915=>"110011100",
  15916=>"111000101",
  15917=>"100010111",
  15918=>"101101000",
  15919=>"111000111",
  15920=>"100001111",
  15921=>"100100111",
  15922=>"111111100",
  15923=>"111010101",
  15924=>"010110010",
  15925=>"100010010",
  15926=>"100110101",
  15927=>"011101111",
  15928=>"000011101",
  15929=>"100001001",
  15930=>"101000010",
  15931=>"010110001",
  15932=>"011110100",
  15933=>"101000100",
  15934=>"110101011",
  15935=>"001101001",
  15936=>"011100111",
  15937=>"101011011",
  15938=>"011000010",
  15939=>"000000111",
  15940=>"000100100",
  15941=>"110000000",
  15942=>"000101000",
  15943=>"101100000",
  15944=>"100000010",
  15945=>"010100001",
  15946=>"110100100",
  15947=>"101100001",
  15948=>"110100101",
  15949=>"001101000",
  15950=>"110111111",
  15951=>"100001100",
  15952=>"010101001",
  15953=>"001011100",
  15954=>"010010101",
  15955=>"101101101",
  15956=>"011110101",
  15957=>"110100101",
  15958=>"000100111",
  15959=>"011010010",
  15960=>"010001010",
  15961=>"011010000",
  15962=>"100001111",
  15963=>"010000000",
  15964=>"000111011",
  15965=>"100010110",
  15966=>"110010110",
  15967=>"000011000",
  15968=>"010000111",
  15969=>"101010101",
  15970=>"101101101",
  15971=>"111110101",
  15972=>"111011101",
  15973=>"111111001",
  15974=>"000110011",
  15975=>"100100010",
  15976=>"100100011",
  15977=>"000000110",
  15978=>"110101111",
  15979=>"000000011",
  15980=>"101001100",
  15981=>"000111101",
  15982=>"101101101",
  15983=>"010001111",
  15984=>"100010100",
  15985=>"111101000",
  15986=>"010111000",
  15987=>"111110100",
  15988=>"000000101",
  15989=>"000101101",
  15990=>"111001111",
  15991=>"111110011",
  15992=>"011001110",
  15993=>"011010011",
  15994=>"010111101",
  15995=>"000100010",
  15996=>"110111101",
  15997=>"111010111",
  15998=>"101010101",
  15999=>"111000010",
  16000=>"000101000",
  16001=>"000011000",
  16002=>"010111100",
  16003=>"101100000",
  16004=>"111001011",
  16005=>"111101001",
  16006=>"011010001",
  16007=>"001100111",
  16008=>"110011010",
  16009=>"010011100",
  16010=>"000001100",
  16011=>"111101111",
  16012=>"110101101",
  16013=>"000110010",
  16014=>"001001001",
  16015=>"110100101",
  16016=>"111110101",
  16017=>"101000011",
  16018=>"111100111",
  16019=>"001110101",
  16020=>"111100011",
  16021=>"000111010",
  16022=>"110111000",
  16023=>"001010001",
  16024=>"001110010",
  16025=>"001110101",
  16026=>"000110010",
  16027=>"111101100",
  16028=>"100100011",
  16029=>"011011100",
  16030=>"010000000",
  16031=>"000011011",
  16032=>"111000111",
  16033=>"100001011",
  16034=>"001101011",
  16035=>"100010111",
  16036=>"010100101",
  16037=>"100011011",
  16038=>"001001000",
  16039=>"101000101",
  16040=>"000100010",
  16041=>"111100000",
  16042=>"001000011",
  16043=>"100000000",
  16044=>"000001000",
  16045=>"110110101",
  16046=>"001001010",
  16047=>"101001010",
  16048=>"010110111",
  16049=>"101100011",
  16050=>"100011100",
  16051=>"111101010",
  16052=>"101001010",
  16053=>"110010111",
  16054=>"010001011",
  16055=>"100111101",
  16056=>"010100111",
  16057=>"001001000",
  16058=>"110100000",
  16059=>"111000001",
  16060=>"110000101",
  16061=>"100101110",
  16062=>"101100111",
  16063=>"101011101",
  16064=>"011110111",
  16065=>"111101010",
  16066=>"101001011",
  16067=>"111010000",
  16068=>"110100000",
  16069=>"000001010",
  16070=>"010111000",
  16071=>"101000111",
  16072=>"101100001",
  16073=>"111001010",
  16074=>"100001010",
  16075=>"101001100",
  16076=>"001001101",
  16077=>"101010000",
  16078=>"000010011",
  16079=>"111011101",
  16080=>"100010110",
  16081=>"100010110",
  16082=>"111011001",
  16083=>"111101111",
  16084=>"000001010",
  16085=>"000000110",
  16086=>"010110111",
  16087=>"010111000",
  16088=>"000101001",
  16089=>"001110110",
  16090=>"001101101",
  16091=>"110100100",
  16092=>"101101111",
  16093=>"011011000",
  16094=>"101011110",
  16095=>"100010111",
  16096=>"010100111",
  16097=>"100000010",
  16098=>"101110100",
  16099=>"010101000",
  16100=>"010001111",
  16101=>"010011011",
  16102=>"101110101",
  16103=>"101000001",
  16104=>"001100010",
  16105=>"111111000",
  16106=>"101111010",
  16107=>"101111001",
  16108=>"101101000",
  16109=>"000101010",
  16110=>"100011111",
  16111=>"000001000",
  16112=>"111110011",
  16113=>"110110010",
  16114=>"111011001",
  16115=>"000011110",
  16116=>"111001101",
  16117=>"000011101",
  16118=>"010011001",
  16119=>"110011110",
  16120=>"100000001",
  16121=>"110110110",
  16122=>"110011010",
  16123=>"010001000",
  16124=>"101110001",
  16125=>"011001110",
  16126=>"010011001",
  16127=>"000010000",
  16128=>"000000101",
  16129=>"010100000",
  16130=>"110101001",
  16131=>"000010010",
  16132=>"110000001",
  16133=>"110101111",
  16134=>"010101010",
  16135=>"000000110",
  16136=>"001110111",
  16137=>"101111011",
  16138=>"111010110",
  16139=>"111010010",
  16140=>"111001101",
  16141=>"001001110",
  16142=>"100111101",
  16143=>"011000111",
  16144=>"010100101",
  16145=>"011101100",
  16146=>"001000011",
  16147=>"101110110",
  16148=>"110000010",
  16149=>"110001000",
  16150=>"010010100",
  16151=>"111010111",
  16152=>"011010111",
  16153=>"101000000",
  16154=>"101000101",
  16155=>"011101100",
  16156=>"010100001",
  16157=>"110001011",
  16158=>"001001101",
  16159=>"000101110",
  16160=>"001000001",
  16161=>"111101001",
  16162=>"011010010",
  16163=>"010111011",
  16164=>"100101011",
  16165=>"000100100",
  16166=>"111011010",
  16167=>"000110110",
  16168=>"110000011",
  16169=>"101010000",
  16170=>"001110100",
  16171=>"001111101",
  16172=>"110111101",
  16173=>"101110101",
  16174=>"100000100",
  16175=>"000000000",
  16176=>"000100110",
  16177=>"111010011",
  16178=>"101010110",
  16179=>"101001001",
  16180=>"111111010",
  16181=>"000101101",
  16182=>"111110111",
  16183=>"000111000",
  16184=>"010011111",
  16185=>"110001001",
  16186=>"000011110",
  16187=>"101001110",
  16188=>"000001000",
  16189=>"000010000",
  16190=>"101010000",
  16191=>"010101001",
  16192=>"111111001",
  16193=>"000010000",
  16194=>"000111010",
  16195=>"010011101",
  16196=>"011101101",
  16197=>"010000101",
  16198=>"001000111",
  16199=>"100011010",
  16200=>"010110001",
  16201=>"000000111",
  16202=>"010100010",
  16203=>"011010010",
  16204=>"110001101",
  16205=>"100101100",
  16206=>"001001001",
  16207=>"010010001",
  16208=>"100100100",
  16209=>"000001010",
  16210=>"010100000",
  16211=>"110010100",
  16212=>"011000011",
  16213=>"101110100",
  16214=>"011001010",
  16215=>"101111100",
  16216=>"011100111",
  16217=>"101001001",
  16218=>"011100000",
  16219=>"100101100",
  16220=>"011011000",
  16221=>"001000100",
  16222=>"001001101",
  16223=>"000000011",
  16224=>"101000101",
  16225=>"101000110",
  16226=>"001001010",
  16227=>"001010011",
  16228=>"101000001",
  16229=>"000100011",
  16230=>"100111000",
  16231=>"100011000",
  16232=>"011111110",
  16233=>"101010101",
  16234=>"011100111",
  16235=>"110101011",
  16236=>"110101111",
  16237=>"110101011",
  16238=>"110011100",
  16239=>"011111110",
  16240=>"100111110",
  16241=>"111101110",
  16242=>"101101010",
  16243=>"001000000",
  16244=>"000010001",
  16245=>"110100101",
  16246=>"111010100",
  16247=>"010000110",
  16248=>"011111010",
  16249=>"100100001",
  16250=>"100011110",
  16251=>"011111101",
  16252=>"000100011",
  16253=>"101010111",
  16254=>"000001000",
  16255=>"011110100",
  16256=>"011111101",
  16257=>"010111011",
  16258=>"101011110",
  16259=>"101000000",
  16260=>"010100011",
  16261=>"001100001",
  16262=>"000101001",
  16263=>"000100000",
  16264=>"110010100",
  16265=>"011011011",
  16266=>"111110101",
  16267=>"101010001",
  16268=>"111101001",
  16269=>"001001011",
  16270=>"011110110",
  16271=>"100110011",
  16272=>"000101100",
  16273=>"010111010",
  16274=>"100001110",
  16275=>"100000011",
  16276=>"000011101",
  16277=>"010010001",
  16278=>"000101101",
  16279=>"011100111",
  16280=>"110000001",
  16281=>"110001011",
  16282=>"110111000",
  16283=>"101000001",
  16284=>"110101100",
  16285=>"001010000",
  16286=>"011010010",
  16287=>"101000111",
  16288=>"111101001",
  16289=>"110011110",
  16290=>"000111000",
  16291=>"100101001",
  16292=>"010111110",
  16293=>"111001100",
  16294=>"111101100",
  16295=>"100110101",
  16296=>"001101001",
  16297=>"101111011",
  16298=>"110000010",
  16299=>"110011011",
  16300=>"010000111",
  16301=>"000010011",
  16302=>"100101011",
  16303=>"101100100",
  16304=>"100110110",
  16305=>"000011111",
  16306=>"101111001",
  16307=>"000110101",
  16308=>"011111111",
  16309=>"111101011",
  16310=>"101111101",
  16311=>"001001101",
  16312=>"100010001",
  16313=>"111011000",
  16314=>"001111010",
  16315=>"000100111",
  16316=>"110001110",
  16317=>"110001110",
  16318=>"001010000",
  16319=>"000001110",
  16320=>"010000000",
  16321=>"101011110",
  16322=>"001101110",
  16323=>"000110001",
  16324=>"100100101",
  16325=>"101111100",
  16326=>"011100111",
  16327=>"010110101",
  16328=>"001010111",
  16329=>"101111101",
  16330=>"100101100",
  16331=>"011101101",
  16332=>"101011110",
  16333=>"101100011",
  16334=>"100010001",
  16335=>"011001101",
  16336=>"000110010",
  16337=>"011100011",
  16338=>"110011010",
  16339=>"110001011",
  16340=>"100100101",
  16341=>"000000010",
  16342=>"011011101",
  16343=>"111001100",
  16344=>"110010010",
  16345=>"100101100",
  16346=>"001010010",
  16347=>"110000101",
  16348=>"111001000",
  16349=>"011001111",
  16350=>"110010010",
  16351=>"001000101",
  16352=>"100101010",
  16353=>"001000101",
  16354=>"111011101",
  16355=>"010111000",
  16356=>"111110001",
  16357=>"101001001",
  16358=>"101101000",
  16359=>"100100111",
  16360=>"000000010",
  16361=>"011011001",
  16362=>"010000100",
  16363=>"100101111",
  16364=>"011001000",
  16365=>"110101100",
  16366=>"111011000",
  16367=>"001000111",
  16368=>"001101111",
  16369=>"101001111",
  16370=>"101100010",
  16371=>"111011001",
  16372=>"100010011",
  16373=>"010100010",
  16374=>"100001110",
  16375=>"011001111",
  16376=>"011111011",
  16377=>"101110101",
  16378=>"110001100",
  16379=>"111101100",
  16380=>"001000110",
  16381=>"000111100",
  16382=>"111111111",
  16383=>"000111011",
  16384=>"110101111",
  16385=>"111011101",
  16386=>"010001110",
  16387=>"000000010",
  16388=>"010100101",
  16389=>"111011100",
  16390=>"011110110",
  16391=>"101000101",
  16392=>"100010000",
  16393=>"100001111",
  16394=>"000001010",
  16395=>"101111001",
  16396=>"101100001",
  16397=>"001000111",
  16398=>"010100100",
  16399=>"001001001",
  16400=>"010010110",
  16401=>"101010011",
  16402=>"101010101",
  16403=>"001010110",
  16404=>"111100100",
  16405=>"101100010",
  16406=>"100100000",
  16407=>"101011010",
  16408=>"000100110",
  16409=>"100101111",
  16410=>"000100000",
  16411=>"000010100",
  16412=>"100001111",
  16413=>"010001101",
  16414=>"111110111",
  16415=>"001100001",
  16416=>"010000110",
  16417=>"011000001",
  16418=>"000011111",
  16419=>"000100000",
  16420=>"001101001",
  16421=>"000111010",
  16422=>"110110111",
  16423=>"110000111",
  16424=>"010001110",
  16425=>"000111111",
  16426=>"000010000",
  16427=>"111101100",
  16428=>"001110110",
  16429=>"111110010",
  16430=>"001011101",
  16431=>"010001011",
  16432=>"010011111",
  16433=>"111101100",
  16434=>"011011001",
  16435=>"001110010",
  16436=>"111101011",
  16437=>"000010001",
  16438=>"110010101",
  16439=>"111111111",
  16440=>"001101111",
  16441=>"101111110",
  16442=>"001000000",
  16443=>"110000111",
  16444=>"110001001",
  16445=>"110000100",
  16446=>"000110101",
  16447=>"111100011",
  16448=>"011100000",
  16449=>"001110001",
  16450=>"110111000",
  16451=>"010101110",
  16452=>"000111010",
  16453=>"101010000",
  16454=>"010110110",
  16455=>"000100110",
  16456=>"100110100",
  16457=>"001110010",
  16458=>"000110110",
  16459=>"110100111",
  16460=>"001110110",
  16461=>"010101111",
  16462=>"100010000",
  16463=>"000000010",
  16464=>"111011101",
  16465=>"000111111",
  16466=>"110111001",
  16467=>"011110110",
  16468=>"101001101",
  16469=>"010110011",
  16470=>"011000100",
  16471=>"001011011",
  16472=>"111111110",
  16473=>"010011010",
  16474=>"110111101",
  16475=>"000100011",
  16476=>"010010000",
  16477=>"111101001",
  16478=>"111000100",
  16479=>"100111010",
  16480=>"011111101",
  16481=>"000001010",
  16482=>"000101101",
  16483=>"111011101",
  16484=>"011100101",
  16485=>"110011001",
  16486=>"000000100",
  16487=>"101000001",
  16488=>"000101100",
  16489=>"110100101",
  16490=>"101010111",
  16491=>"111100110",
  16492=>"110000001",
  16493=>"111011010",
  16494=>"100101110",
  16495=>"111101110",
  16496=>"110010111",
  16497=>"100010011",
  16498=>"000000000",
  16499=>"110001100",
  16500=>"100011110",
  16501=>"111000000",
  16502=>"101100001",
  16503=>"111001010",
  16504=>"110110100",
  16505=>"110001001",
  16506=>"001111110",
  16507=>"000111010",
  16508=>"100100110",
  16509=>"010100000",
  16510=>"010101110",
  16511=>"001100000",
  16512=>"010000000",
  16513=>"111110101",
  16514=>"011100001",
  16515=>"101010101",
  16516=>"111011110",
  16517=>"010110101",
  16518=>"011100010",
  16519=>"001110100",
  16520=>"011001111",
  16521=>"111011001",
  16522=>"111111011",
  16523=>"111111101",
  16524=>"011111100",
  16525=>"011001110",
  16526=>"000011011",
  16527=>"001010010",
  16528=>"101000011",
  16529=>"000110011",
  16530=>"011100101",
  16531=>"000110010",
  16532=>"110100000",
  16533=>"010010100",
  16534=>"111111000",
  16535=>"110110001",
  16536=>"000111010",
  16537=>"111101000",
  16538=>"101111000",
  16539=>"010101000",
  16540=>"111011110",
  16541=>"000111100",
  16542=>"011000110",
  16543=>"100011001",
  16544=>"011011111",
  16545=>"100001110",
  16546=>"110100001",
  16547=>"111111000",
  16548=>"111011110",
  16549=>"111100110",
  16550=>"011010001",
  16551=>"011111011",
  16552=>"001011001",
  16553=>"110010111",
  16554=>"100101110",
  16555=>"000001001",
  16556=>"111001100",
  16557=>"111110011",
  16558=>"000011101",
  16559=>"000111000",
  16560=>"010010001",
  16561=>"111110101",
  16562=>"010000100",
  16563=>"110110010",
  16564=>"000001101",
  16565=>"011100000",
  16566=>"001110000",
  16567=>"111111000",
  16568=>"001111001",
  16569=>"101011111",
  16570=>"011010000",
  16571=>"000011101",
  16572=>"010111011",
  16573=>"011111110",
  16574=>"111010100",
  16575=>"111000111",
  16576=>"001100111",
  16577=>"001100100",
  16578=>"101111101",
  16579=>"111101010",
  16580=>"101010000",
  16581=>"111011011",
  16582=>"111111011",
  16583=>"011011011",
  16584=>"001101110",
  16585=>"001011111",
  16586=>"010000100",
  16587=>"011111111",
  16588=>"100010011",
  16589=>"110100100",
  16590=>"111001111",
  16591=>"010001111",
  16592=>"111010101",
  16593=>"111110100",
  16594=>"010000011",
  16595=>"010100111",
  16596=>"010100101",
  16597=>"101011110",
  16598=>"001100001",
  16599=>"001010011",
  16600=>"001000111",
  16601=>"111111100",
  16602=>"111011101",
  16603=>"000111110",
  16604=>"111100011",
  16605=>"000011111",
  16606=>"111110011",
  16607=>"001010011",
  16608=>"010110101",
  16609=>"101110010",
  16610=>"111111001",
  16611=>"101010101",
  16612=>"101000010",
  16613=>"001010000",
  16614=>"000000101",
  16615=>"010011011",
  16616=>"000001110",
  16617=>"011101101",
  16618=>"110001110",
  16619=>"000110001",
  16620=>"000100100",
  16621=>"111100111",
  16622=>"101111101",
  16623=>"011111000",
  16624=>"110100100",
  16625=>"010001000",
  16626=>"001100101",
  16627=>"000001100",
  16628=>"110010100",
  16629=>"101001010",
  16630=>"000010101",
  16631=>"000110101",
  16632=>"110010101",
  16633=>"100101110",
  16634=>"001111101",
  16635=>"101101011",
  16636=>"010100011",
  16637=>"110011110",
  16638=>"101110001",
  16639=>"010010001",
  16640=>"111000000",
  16641=>"011110111",
  16642=>"110010011",
  16643=>"001111100",
  16644=>"001000011",
  16645=>"111000001",
  16646=>"111010111",
  16647=>"100010111",
  16648=>"111110111",
  16649=>"110000011",
  16650=>"001000000",
  16651=>"101001100",
  16652=>"011100111",
  16653=>"110101000",
  16654=>"001100001",
  16655=>"000001001",
  16656=>"000000111",
  16657=>"001110100",
  16658=>"111110101",
  16659=>"100010100",
  16660=>"010001001",
  16661=>"010110001",
  16662=>"001010011",
  16663=>"010111010",
  16664=>"100000101",
  16665=>"111100101",
  16666=>"111101100",
  16667=>"101101011",
  16668=>"010010111",
  16669=>"011000101",
  16670=>"100010101",
  16671=>"111110011",
  16672=>"001001100",
  16673=>"100010110",
  16674=>"111011100",
  16675=>"100111000",
  16676=>"110010010",
  16677=>"111100101",
  16678=>"010110000",
  16679=>"111111010",
  16680=>"110010110",
  16681=>"101110000",
  16682=>"001100101",
  16683=>"010000111",
  16684=>"101101001",
  16685=>"111101011",
  16686=>"100001110",
  16687=>"001010110",
  16688=>"100010010",
  16689=>"110101110",
  16690=>"001000110",
  16691=>"001011111",
  16692=>"000110100",
  16693=>"111111011",
  16694=>"110111000",
  16695=>"000000000",
  16696=>"111101010",
  16697=>"001011010",
  16698=>"001101111",
  16699=>"010000010",
  16700=>"111000010",
  16701=>"101001110",
  16702=>"000011110",
  16703=>"101011101",
  16704=>"000011101",
  16705=>"111000111",
  16706=>"000100000",
  16707=>"001001011",
  16708=>"001100011",
  16709=>"000111011",
  16710=>"100000101",
  16711=>"110011010",
  16712=>"111100100",
  16713=>"001001011",
  16714=>"110000111",
  16715=>"011110101",
  16716=>"011100001",
  16717=>"111110111",
  16718=>"100110011",
  16719=>"110110001",
  16720=>"011000011",
  16721=>"111001101",
  16722=>"100101111",
  16723=>"010101001",
  16724=>"011110011",
  16725=>"100110111",
  16726=>"100001010",
  16727=>"100111010",
  16728=>"011101111",
  16729=>"111010011",
  16730=>"000001010",
  16731=>"101100101",
  16732=>"111001010",
  16733=>"011100111",
  16734=>"111011101",
  16735=>"011001010",
  16736=>"111101111",
  16737=>"010111010",
  16738=>"010010001",
  16739=>"111100101",
  16740=>"000011101",
  16741=>"000111011",
  16742=>"011010101",
  16743=>"000100101",
  16744=>"111000011",
  16745=>"111000001",
  16746=>"110010011",
  16747=>"100011000",
  16748=>"100000110",
  16749=>"000010010",
  16750=>"100011101",
  16751=>"011000111",
  16752=>"110000110",
  16753=>"100100010",
  16754=>"001110110",
  16755=>"111001110",
  16756=>"001010000",
  16757=>"011110011",
  16758=>"101100101",
  16759=>"101001100",
  16760=>"111010111",
  16761=>"010110110",
  16762=>"010010111",
  16763=>"010011010",
  16764=>"010010111",
  16765=>"001110110",
  16766=>"011110000",
  16767=>"101011101",
  16768=>"111110011",
  16769=>"111110100",
  16770=>"111000100",
  16771=>"100011101",
  16772=>"111110101",
  16773=>"111111010",
  16774=>"110111110",
  16775=>"100100001",
  16776=>"010100011",
  16777=>"001111100",
  16778=>"001000010",
  16779=>"111101101",
  16780=>"100111100",
  16781=>"111110000",
  16782=>"011111000",
  16783=>"100000100",
  16784=>"111100000",
  16785=>"110111111",
  16786=>"101011011",
  16787=>"100111011",
  16788=>"100111111",
  16789=>"010110100",
  16790=>"011110011",
  16791=>"110100010",
  16792=>"101011100",
  16793=>"001011011",
  16794=>"000100001",
  16795=>"000101111",
  16796=>"000000111",
  16797=>"010111111",
  16798=>"111000100",
  16799=>"111010101",
  16800=>"111111010",
  16801=>"001110000",
  16802=>"001000000",
  16803=>"011011111",
  16804=>"001101101",
  16805=>"101110000",
  16806=>"101011100",
  16807=>"110000111",
  16808=>"001000011",
  16809=>"011000010",
  16810=>"001001011",
  16811=>"100011011",
  16812=>"111110101",
  16813=>"000001101",
  16814=>"000010001",
  16815=>"100010111",
  16816=>"011101011",
  16817=>"011000000",
  16818=>"100101011",
  16819=>"011011011",
  16820=>"000000010",
  16821=>"000011101",
  16822=>"110111110",
  16823=>"001110011",
  16824=>"001101101",
  16825=>"000011011",
  16826=>"111111000",
  16827=>"111100010",
  16828=>"110101001",
  16829=>"000101001",
  16830=>"010010111",
  16831=>"101011111",
  16832=>"001000000",
  16833=>"011110000",
  16834=>"001001110",
  16835=>"000010001",
  16836=>"110111111",
  16837=>"011011000",
  16838=>"111000000",
  16839=>"100011100",
  16840=>"011001111",
  16841=>"111101111",
  16842=>"100111000",
  16843=>"101110101",
  16844=>"100111110",
  16845=>"001001101",
  16846=>"001110110",
  16847=>"000100100",
  16848=>"101110101",
  16849=>"010011111",
  16850=>"000000101",
  16851=>"110111111",
  16852=>"001110100",
  16853=>"100010010",
  16854=>"000010011",
  16855=>"010011010",
  16856=>"101111110",
  16857=>"000001111",
  16858=>"001100010",
  16859=>"111000111",
  16860=>"011000111",
  16861=>"111101001",
  16862=>"110000100",
  16863=>"000100111",
  16864=>"110101100",
  16865=>"011110011",
  16866=>"000110111",
  16867=>"110011110",
  16868=>"000100111",
  16869=>"100000111",
  16870=>"100100111",
  16871=>"100111001",
  16872=>"011011001",
  16873=>"011010101",
  16874=>"110100110",
  16875=>"000011110",
  16876=>"001110000",
  16877=>"011110110",
  16878=>"001000111",
  16879=>"110101111",
  16880=>"011011100",
  16881=>"001000011",
  16882=>"011100010",
  16883=>"011100000",
  16884=>"100001000",
  16885=>"000010111",
  16886=>"001000110",
  16887=>"011011010",
  16888=>"000111111",
  16889=>"010110000",
  16890=>"110110111",
  16891=>"101111001",
  16892=>"101100010",
  16893=>"100010111",
  16894=>"101110010",
  16895=>"000100001",
  16896=>"110100010",
  16897=>"001001011",
  16898=>"001001100",
  16899=>"011100001",
  16900=>"110101111",
  16901=>"000001010",
  16902=>"010010111",
  16903=>"100010110",
  16904=>"001010111",
  16905=>"110111011",
  16906=>"010000100",
  16907=>"111110110",
  16908=>"011100100",
  16909=>"100011010",
  16910=>"000010111",
  16911=>"110110000",
  16912=>"110101110",
  16913=>"100101000",
  16914=>"000011110",
  16915=>"100000101",
  16916=>"100000010",
  16917=>"100011110",
  16918=>"110100001",
  16919=>"011001100",
  16920=>"001000000",
  16921=>"000111011",
  16922=>"111110010",
  16923=>"000001001",
  16924=>"100110111",
  16925=>"000010100",
  16926=>"011111000",
  16927=>"110001011",
  16928=>"000011011",
  16929=>"101011111",
  16930=>"111011111",
  16931=>"000011010",
  16932=>"001100100",
  16933=>"001100101",
  16934=>"010000101",
  16935=>"001100111",
  16936=>"111100100",
  16937=>"001110010",
  16938=>"100100000",
  16939=>"111001001",
  16940=>"011111010",
  16941=>"011101000",
  16942=>"111100001",
  16943=>"001111101",
  16944=>"100010111",
  16945=>"111000100",
  16946=>"111011101",
  16947=>"101010110",
  16948=>"011011111",
  16949=>"001101010",
  16950=>"011101001",
  16951=>"100100101",
  16952=>"111111100",
  16953=>"101101011",
  16954=>"000101001",
  16955=>"010101000",
  16956=>"001011101",
  16957=>"111110010",
  16958=>"000100001",
  16959=>"100010101",
  16960=>"101110111",
  16961=>"010011100",
  16962=>"001100001",
  16963=>"010000111",
  16964=>"000000111",
  16965=>"111101001",
  16966=>"001001011",
  16967=>"000011110",
  16968=>"000011100",
  16969=>"000010110",
  16970=>"100100000",
  16971=>"111111011",
  16972=>"100100111",
  16973=>"001101101",
  16974=>"000000011",
  16975=>"010111010",
  16976=>"011010111",
  16977=>"001001111",
  16978=>"011111011",
  16979=>"000010010",
  16980=>"011110000",
  16981=>"110011011",
  16982=>"100110011",
  16983=>"110001111",
  16984=>"001011010",
  16985=>"110011100",
  16986=>"101000001",
  16987=>"001100111",
  16988=>"011111100",
  16989=>"001001000",
  16990=>"001001100",
  16991=>"110011001",
  16992=>"101111111",
  16993=>"000000101",
  16994=>"110111001",
  16995=>"110111111",
  16996=>"011011001",
  16997=>"110100101",
  16998=>"110101101",
  16999=>"110000101",
  17000=>"111001010",
  17001=>"001010101",
  17002=>"001001111",
  17003=>"100111000",
  17004=>"001010101",
  17005=>"110001000",
  17006=>"111110001",
  17007=>"100001110",
  17008=>"111111011",
  17009=>"101101010",
  17010=>"000001000",
  17011=>"010111010",
  17012=>"110000000",
  17013=>"100110011",
  17014=>"011001110",
  17015=>"001101100",
  17016=>"100001010",
  17017=>"101101011",
  17018=>"001110000",
  17019=>"111110110",
  17020=>"001100110",
  17021=>"010010011",
  17022=>"100111000",
  17023=>"010001000",
  17024=>"000100111",
  17025=>"010000011",
  17026=>"000100110",
  17027=>"101110100",
  17028=>"101100110",
  17029=>"110110110",
  17030=>"001111101",
  17031=>"011010101",
  17032=>"111101111",
  17033=>"111011000",
  17034=>"001100000",
  17035=>"100101111",
  17036=>"011010100",
  17037=>"111011100",
  17038=>"011101101",
  17039=>"010000010",
  17040=>"101000100",
  17041=>"110100110",
  17042=>"000010101",
  17043=>"110101011",
  17044=>"101101000",
  17045=>"001110001",
  17046=>"110011110",
  17047=>"011110110",
  17048=>"100110011",
  17049=>"001010110",
  17050=>"101101101",
  17051=>"010000110",
  17052=>"001111110",
  17053=>"110100100",
  17054=>"000000111",
  17055=>"111111111",
  17056=>"111010000",
  17057=>"000101001",
  17058=>"111010101",
  17059=>"111100000",
  17060=>"011101010",
  17061=>"101011000",
  17062=>"001001111",
  17063=>"000011011",
  17064=>"111010000",
  17065=>"100010101",
  17066=>"000001011",
  17067=>"010010011",
  17068=>"010001000",
  17069=>"101101100",
  17070=>"011000101",
  17071=>"101100011",
  17072=>"101001110",
  17073=>"101110101",
  17074=>"111111000",
  17075=>"111110011",
  17076=>"110101100",
  17077=>"011100000",
  17078=>"111000010",
  17079=>"010101110",
  17080=>"000101010",
  17081=>"110111110",
  17082=>"111011100",
  17083=>"001111111",
  17084=>"010000111",
  17085=>"001000011",
  17086=>"011011011",
  17087=>"111101010",
  17088=>"011100000",
  17089=>"110111101",
  17090=>"101100010",
  17091=>"010100110",
  17092=>"101010100",
  17093=>"010111101",
  17094=>"110000101",
  17095=>"100011011",
  17096=>"110011101",
  17097=>"010110100",
  17098=>"111011001",
  17099=>"111000101",
  17100=>"111001101",
  17101=>"111011101",
  17102=>"000001110",
  17103=>"110000000",
  17104=>"000110111",
  17105=>"101101100",
  17106=>"011010110",
  17107=>"101011110",
  17108=>"100001111",
  17109=>"111111100",
  17110=>"110011100",
  17111=>"111011010",
  17112=>"111111110",
  17113=>"000100110",
  17114=>"110100001",
  17115=>"001011011",
  17116=>"001111111",
  17117=>"111000000",
  17118=>"111010100",
  17119=>"101111100",
  17120=>"011011101",
  17121=>"111011101",
  17122=>"001010011",
  17123=>"001101111",
  17124=>"101010010",
  17125=>"110010000",
  17126=>"001110111",
  17127=>"000000101",
  17128=>"001001111",
  17129=>"110001101",
  17130=>"111110110",
  17131=>"000001011",
  17132=>"111111101",
  17133=>"001101100",
  17134=>"110101010",
  17135=>"011001101",
  17136=>"010001111",
  17137=>"110100001",
  17138=>"011110011",
  17139=>"100001010",
  17140=>"111111101",
  17141=>"010011101",
  17142=>"011110011",
  17143=>"001010010",
  17144=>"110011111",
  17145=>"010011110",
  17146=>"111110010",
  17147=>"011010010",
  17148=>"010001001",
  17149=>"110111100",
  17150=>"110110111",
  17151=>"101100010",
  17152=>"110000001",
  17153=>"011000100",
  17154=>"110010111",
  17155=>"110101000",
  17156=>"000110101",
  17157=>"111110111",
  17158=>"001001011",
  17159=>"011110011",
  17160=>"001011100",
  17161=>"001000000",
  17162=>"011101011",
  17163=>"010001101",
  17164=>"110100101",
  17165=>"111111111",
  17166=>"101010011",
  17167=>"110101110",
  17168=>"110001001",
  17169=>"100111000",
  17170=>"001101011",
  17171=>"101100010",
  17172=>"011111001",
  17173=>"101010110",
  17174=>"011000100",
  17175=>"100000101",
  17176=>"011000001",
  17177=>"100011000",
  17178=>"010111110",
  17179=>"111100111",
  17180=>"100101011",
  17181=>"111010101",
  17182=>"101100101",
  17183=>"010010001",
  17184=>"110111111",
  17185=>"000101000",
  17186=>"011101000",
  17187=>"101001011",
  17188=>"101010101",
  17189=>"111000011",
  17190=>"100011000",
  17191=>"110100010",
  17192=>"111000110",
  17193=>"010001101",
  17194=>"101001001",
  17195=>"111000011",
  17196=>"100001110",
  17197=>"111010010",
  17198=>"101101011",
  17199=>"010101000",
  17200=>"101110010",
  17201=>"110110001",
  17202=>"110000001",
  17203=>"001100001",
  17204=>"000000000",
  17205=>"100110011",
  17206=>"001000000",
  17207=>"000011000",
  17208=>"111011001",
  17209=>"101011011",
  17210=>"001110011",
  17211=>"001001100",
  17212=>"111111000",
  17213=>"000111110",
  17214=>"000011011",
  17215=>"110110001",
  17216=>"000111101",
  17217=>"011101000",
  17218=>"010101000",
  17219=>"001010001",
  17220=>"110001010",
  17221=>"111010011",
  17222=>"011101100",
  17223=>"010010011",
  17224=>"000100011",
  17225=>"011010011",
  17226=>"010111110",
  17227=>"001101011",
  17228=>"000011110",
  17229=>"010000010",
  17230=>"110110011",
  17231=>"111101110",
  17232=>"110100101",
  17233=>"000000011",
  17234=>"110100011",
  17235=>"101010011",
  17236=>"001101011",
  17237=>"000011100",
  17238=>"101010010",
  17239=>"101000111",
  17240=>"100100101",
  17241=>"011000001",
  17242=>"111001110",
  17243=>"001101101",
  17244=>"011011010",
  17245=>"011001001",
  17246=>"000001111",
  17247=>"100010001",
  17248=>"101001110",
  17249=>"000101111",
  17250=>"101011101",
  17251=>"001101000",
  17252=>"000010111",
  17253=>"110110000",
  17254=>"000101111",
  17255=>"101101010",
  17256=>"100001000",
  17257=>"011001110",
  17258=>"001111010",
  17259=>"001110110",
  17260=>"101001111",
  17261=>"011110100",
  17262=>"100100100",
  17263=>"100100101",
  17264=>"111000101",
  17265=>"011011001",
  17266=>"110000001",
  17267=>"110101101",
  17268=>"101101100",
  17269=>"111000011",
  17270=>"110110111",
  17271=>"011010111",
  17272=>"111101010",
  17273=>"111111111",
  17274=>"101001001",
  17275=>"000011011",
  17276=>"100110100",
  17277=>"001111000",
  17278=>"000101110",
  17279=>"100110011",
  17280=>"100100110",
  17281=>"100101010",
  17282=>"110011110",
  17283=>"111101100",
  17284=>"110000010",
  17285=>"110011011",
  17286=>"101111101",
  17287=>"000000001",
  17288=>"111111010",
  17289=>"101000001",
  17290=>"111111110",
  17291=>"101111010",
  17292=>"110010111",
  17293=>"101100000",
  17294=>"111101100",
  17295=>"000101101",
  17296=>"101101100",
  17297=>"100101000",
  17298=>"000011001",
  17299=>"011110101",
  17300=>"011011111",
  17301=>"011001000",
  17302=>"110000000",
  17303=>"111101100",
  17304=>"001101110",
  17305=>"010110101",
  17306=>"011001011",
  17307=>"100000011",
  17308=>"111101101",
  17309=>"011010000",
  17310=>"100101011",
  17311=>"111010001",
  17312=>"111011001",
  17313=>"101000011",
  17314=>"110101110",
  17315=>"011100111",
  17316=>"000000000",
  17317=>"011111101",
  17318=>"101111000",
  17319=>"010000001",
  17320=>"011011111",
  17321=>"000010111",
  17322=>"110100100",
  17323=>"000100111",
  17324=>"000100110",
  17325=>"000010010",
  17326=>"010100111",
  17327=>"001101100",
  17328=>"100100000",
  17329=>"010001011",
  17330=>"110010001",
  17331=>"010110111",
  17332=>"110011001",
  17333=>"111100011",
  17334=>"010011001",
  17335=>"010010110",
  17336=>"010101010",
  17337=>"101011110",
  17338=>"101010101",
  17339=>"010111110",
  17340=>"100110001",
  17341=>"010000000",
  17342=>"010001110",
  17343=>"101101110",
  17344=>"000111100",
  17345=>"100110010",
  17346=>"111010110",
  17347=>"100000000",
  17348=>"000100101",
  17349=>"101010110",
  17350=>"011111100",
  17351=>"001100110",
  17352=>"110100000",
  17353=>"000000000",
  17354=>"100111101",
  17355=>"111110000",
  17356=>"101000011",
  17357=>"111111111",
  17358=>"001001100",
  17359=>"101000001",
  17360=>"010000110",
  17361=>"100011001",
  17362=>"110110101",
  17363=>"100011001",
  17364=>"111001111",
  17365=>"111001001",
  17366=>"111111111",
  17367=>"000101110",
  17368=>"101111011",
  17369=>"110111000",
  17370=>"010100100",
  17371=>"111101110",
  17372=>"011011001",
  17373=>"001111111",
  17374=>"100000111",
  17375=>"100010111",
  17376=>"110011001",
  17377=>"111111111",
  17378=>"011111110",
  17379=>"111000000",
  17380=>"000101110",
  17381=>"000001101",
  17382=>"110111001",
  17383=>"011111011",
  17384=>"101010011",
  17385=>"001111111",
  17386=>"101101111",
  17387=>"111100111",
  17388=>"110010001",
  17389=>"000111111",
  17390=>"101011011",
  17391=>"010101111",
  17392=>"000100110",
  17393=>"100001011",
  17394=>"110110011",
  17395=>"011101101",
  17396=>"010001111",
  17397=>"010001001",
  17398=>"100011100",
  17399=>"101100101",
  17400=>"100110110",
  17401=>"101100011",
  17402=>"001100010",
  17403=>"111101010",
  17404=>"011111111",
  17405=>"111110110",
  17406=>"111110111",
  17407=>"010111110",
  17408=>"001000100",
  17409=>"110100001",
  17410=>"110111101",
  17411=>"110000010",
  17412=>"000000010",
  17413=>"111110110",
  17414=>"000000001",
  17415=>"110100100",
  17416=>"110001110",
  17417=>"110111011",
  17418=>"100001111",
  17419=>"110011010",
  17420=>"011010110",
  17421=>"000000111",
  17422=>"111000011",
  17423=>"011111001",
  17424=>"110010010",
  17425=>"100100001",
  17426=>"110101111",
  17427=>"001111011",
  17428=>"101001110",
  17429=>"101111111",
  17430=>"110000010",
  17431=>"110100011",
  17432=>"001001011",
  17433=>"000111111",
  17434=>"011011001",
  17435=>"111011101",
  17436=>"110010010",
  17437=>"001011111",
  17438=>"001000100",
  17439=>"101111111",
  17440=>"000001001",
  17441=>"100000110",
  17442=>"111111001",
  17443=>"010110111",
  17444=>"010010111",
  17445=>"110011110",
  17446=>"101000100",
  17447=>"010100001",
  17448=>"000011001",
  17449=>"000011000",
  17450=>"110111111",
  17451=>"110100100",
  17452=>"100010000",
  17453=>"010001011",
  17454=>"011010000",
  17455=>"101100111",
  17456=>"011010100",
  17457=>"000010000",
  17458=>"111001111",
  17459=>"111100111",
  17460=>"101010110",
  17461=>"000001000",
  17462=>"001001110",
  17463=>"001110101",
  17464=>"100001010",
  17465=>"011011001",
  17466=>"010001001",
  17467=>"010100100",
  17468=>"110011001",
  17469=>"100101010",
  17470=>"010111110",
  17471=>"101010110",
  17472=>"010111110",
  17473=>"011011001",
  17474=>"100001100",
  17475=>"110000111",
  17476=>"101100100",
  17477=>"111010011",
  17478=>"000010011",
  17479=>"110010011",
  17480=>"110101111",
  17481=>"101001100",
  17482=>"111000100",
  17483=>"110001000",
  17484=>"001111001",
  17485=>"100011001",
  17486=>"010111110",
  17487=>"101111101",
  17488=>"000110010",
  17489=>"010001000",
  17490=>"001111110",
  17491=>"101000100",
  17492=>"000010011",
  17493=>"101001000",
  17494=>"010100001",
  17495=>"110001110",
  17496=>"010100110",
  17497=>"000110101",
  17498=>"111001011",
  17499=>"000011000",
  17500=>"001100011",
  17501=>"011000111",
  17502=>"110011000",
  17503=>"011001001",
  17504=>"000110100",
  17505=>"111001111",
  17506=>"001110001",
  17507=>"111111011",
  17508=>"101001010",
  17509=>"100010010",
  17510=>"100111011",
  17511=>"000011111",
  17512=>"101110000",
  17513=>"111111001",
  17514=>"100001100",
  17515=>"010000010",
  17516=>"001100000",
  17517=>"000001010",
  17518=>"101001001",
  17519=>"000101011",
  17520=>"101010000",
  17521=>"101000100",
  17522=>"000111001",
  17523=>"011101101",
  17524=>"101010110",
  17525=>"010101100",
  17526=>"011010011",
  17527=>"011001101",
  17528=>"000000101",
  17529=>"011100000",
  17530=>"111000001",
  17531=>"100000111",
  17532=>"100011000",
  17533=>"011000011",
  17534=>"010000011",
  17535=>"110101010",
  17536=>"101001100",
  17537=>"000011001",
  17538=>"111010100",
  17539=>"100010010",
  17540=>"000010010",
  17541=>"101110100",
  17542=>"111011101",
  17543=>"010011101",
  17544=>"101011110",
  17545=>"000110111",
  17546=>"010101001",
  17547=>"111110001",
  17548=>"110001010",
  17549=>"000011101",
  17550=>"000000101",
  17551=>"001001100",
  17552=>"011010100",
  17553=>"000001010",
  17554=>"110111111",
  17555=>"100100100",
  17556=>"111101000",
  17557=>"000010000",
  17558=>"001000000",
  17559=>"001001100",
  17560=>"111011001",
  17561=>"110000001",
  17562=>"001110111",
  17563=>"010100011",
  17564=>"000010100",
  17565=>"100110001",
  17566=>"111100111",
  17567=>"000110010",
  17568=>"001001100",
  17569=>"110110000",
  17570=>"101001101",
  17571=>"000111010",
  17572=>"000011100",
  17573=>"111001111",
  17574=>"110010111",
  17575=>"010001111",
  17576=>"001100001",
  17577=>"001000010",
  17578=>"111101001",
  17579=>"110001100",
  17580=>"011111100",
  17581=>"110101100",
  17582=>"100000100",
  17583=>"101100001",
  17584=>"010011110",
  17585=>"000100111",
  17586=>"111100010",
  17587=>"001100010",
  17588=>"101010000",
  17589=>"100111111",
  17590=>"000101001",
  17591=>"111100111",
  17592=>"011111100",
  17593=>"010000111",
  17594=>"000011001",
  17595=>"010100001",
  17596=>"101010001",
  17597=>"101111111",
  17598=>"011101010",
  17599=>"011011001",
  17600=>"110100011",
  17601=>"100000010",
  17602=>"010111011",
  17603=>"001100110",
  17604=>"010011000",
  17605=>"001101010",
  17606=>"111111011",
  17607=>"011111001",
  17608=>"111000001",
  17609=>"100000110",
  17610=>"110111011",
  17611=>"011111001",
  17612=>"100001101",
  17613=>"100010010",
  17614=>"111111110",
  17615=>"110111101",
  17616=>"011111011",
  17617=>"011110111",
  17618=>"000010101",
  17619=>"111001010",
  17620=>"000010101",
  17621=>"011111001",
  17622=>"010110100",
  17623=>"100000010",
  17624=>"100110110",
  17625=>"100110111",
  17626=>"000011110",
  17627=>"001000011",
  17628=>"101000010",
  17629=>"011100111",
  17630=>"001101000",
  17631=>"010011011",
  17632=>"101110111",
  17633=>"110100110",
  17634=>"101011000",
  17635=>"101011010",
  17636=>"101101010",
  17637=>"001100000",
  17638=>"011001111",
  17639=>"111101100",
  17640=>"001011001",
  17641=>"111110000",
  17642=>"010110111",
  17643=>"001010010",
  17644=>"100011011",
  17645=>"101101000",
  17646=>"000110001",
  17647=>"101000000",
  17648=>"010000001",
  17649=>"101111111",
  17650=>"000101101",
  17651=>"100011000",
  17652=>"000001010",
  17653=>"111011001",
  17654=>"011011110",
  17655=>"101111111",
  17656=>"000010011",
  17657=>"000010111",
  17658=>"000111110",
  17659=>"000000011",
  17660=>"000000000",
  17661=>"011100111",
  17662=>"011101000",
  17663=>"000010110",
  17664=>"011001101",
  17665=>"110110000",
  17666=>"010101110",
  17667=>"001101101",
  17668=>"101000100",
  17669=>"111010000",
  17670=>"100110000",
  17671=>"011110110",
  17672=>"001100111",
  17673=>"101000001",
  17674=>"110111110",
  17675=>"101010111",
  17676=>"010001011",
  17677=>"100011000",
  17678=>"100111111",
  17679=>"000111100",
  17680=>"110111110",
  17681=>"001100110",
  17682=>"111111110",
  17683=>"111101111",
  17684=>"001100100",
  17685=>"100110111",
  17686=>"111100000",
  17687=>"100010001",
  17688=>"001111011",
  17689=>"001011100",
  17690=>"010110111",
  17691=>"000100000",
  17692=>"001110000",
  17693=>"000001010",
  17694=>"111111100",
  17695=>"000010000",
  17696=>"110000000",
  17697=>"000111010",
  17698=>"101100111",
  17699=>"110110110",
  17700=>"111011000",
  17701=>"011100001",
  17702=>"110000110",
  17703=>"111110110",
  17704=>"101110001",
  17705=>"001010001",
  17706=>"011110111",
  17707=>"011110001",
  17708=>"001101001",
  17709=>"100001101",
  17710=>"010010100",
  17711=>"100010000",
  17712=>"000100111",
  17713=>"100011111",
  17714=>"110011100",
  17715=>"000001110",
  17716=>"111110110",
  17717=>"111111010",
  17718=>"100010100",
  17719=>"000000001",
  17720=>"000010111",
  17721=>"010011110",
  17722=>"000111000",
  17723=>"000100010",
  17724=>"100101010",
  17725=>"110111000",
  17726=>"110011011",
  17727=>"111001001",
  17728=>"000101001",
  17729=>"110111100",
  17730=>"111111010",
  17731=>"001101000",
  17732=>"011100011",
  17733=>"110001001",
  17734=>"011001100",
  17735=>"101011111",
  17736=>"011000001",
  17737=>"010101001",
  17738=>"101010001",
  17739=>"000001100",
  17740=>"011110111",
  17741=>"111010010",
  17742=>"000000111",
  17743=>"100111111",
  17744=>"000001011",
  17745=>"110100111",
  17746=>"001110011",
  17747=>"100001110",
  17748=>"101011011",
  17749=>"111111011",
  17750=>"010011101",
  17751=>"011111011",
  17752=>"000000010",
  17753=>"111001101",
  17754=>"011001010",
  17755=>"000100000",
  17756=>"100110000",
  17757=>"000100111",
  17758=>"101011010",
  17759=>"101011101",
  17760=>"111100101",
  17761=>"101101100",
  17762=>"010110000",
  17763=>"101011011",
  17764=>"100001111",
  17765=>"101111001",
  17766=>"100101000",
  17767=>"111001101",
  17768=>"101011010",
  17769=>"011110010",
  17770=>"000100001",
  17771=>"001010100",
  17772=>"100000101",
  17773=>"100000111",
  17774=>"100110011",
  17775=>"100100001",
  17776=>"111111011",
  17777=>"000111100",
  17778=>"111100100",
  17779=>"011111100",
  17780=>"010111101",
  17781=>"000101010",
  17782=>"011101111",
  17783=>"110111011",
  17784=>"000001101",
  17785=>"001011001",
  17786=>"101010110",
  17787=>"000001011",
  17788=>"010001011",
  17789=>"111101011",
  17790=>"101011011",
  17791=>"111110111",
  17792=>"010100111",
  17793=>"101111011",
  17794=>"010010001",
  17795=>"111000100",
  17796=>"110010110",
  17797=>"000000001",
  17798=>"110100010",
  17799=>"001100110",
  17800=>"111111111",
  17801=>"000000000",
  17802=>"001100010",
  17803=>"111100010",
  17804=>"110110101",
  17805=>"101011010",
  17806=>"010110111",
  17807=>"100100110",
  17808=>"000101010",
  17809=>"011101111",
  17810=>"000001111",
  17811=>"010111110",
  17812=>"101111101",
  17813=>"000101011",
  17814=>"010100010",
  17815=>"111000101",
  17816=>"010011111",
  17817=>"001001100",
  17818=>"101111110",
  17819=>"010000100",
  17820=>"000000111",
  17821=>"101101111",
  17822=>"000100111",
  17823=>"000000001",
  17824=>"100010100",
  17825=>"111001101",
  17826=>"100010010",
  17827=>"000000000",
  17828=>"100000111",
  17829=>"011010001",
  17830=>"011110110",
  17831=>"001000110",
  17832=>"011101100",
  17833=>"111101100",
  17834=>"110010000",
  17835=>"101001101",
  17836=>"111110000",
  17837=>"001001000",
  17838=>"010001000",
  17839=>"100101001",
  17840=>"010111001",
  17841=>"110011111",
  17842=>"100110111",
  17843=>"010010100",
  17844=>"000100001",
  17845=>"111101111",
  17846=>"010100111",
  17847=>"100011011",
  17848=>"111111100",
  17849=>"000001100",
  17850=>"001000010",
  17851=>"001100110",
  17852=>"101111110",
  17853=>"111110101",
  17854=>"001110110",
  17855=>"010000100",
  17856=>"100011111",
  17857=>"001001111",
  17858=>"010010001",
  17859=>"101001011",
  17860=>"100010010",
  17861=>"111110111",
  17862=>"100001001",
  17863=>"010111010",
  17864=>"101110000",
  17865=>"000000011",
  17866=>"010111110",
  17867=>"010100000",
  17868=>"000011010",
  17869=>"100101001",
  17870=>"111010001",
  17871=>"011010101",
  17872=>"101100101",
  17873=>"101100000",
  17874=>"000000110",
  17875=>"111100001",
  17876=>"101010010",
  17877=>"011010101",
  17878=>"111100101",
  17879=>"111000001",
  17880=>"000011101",
  17881=>"101100000",
  17882=>"111000010",
  17883=>"011011000",
  17884=>"101001010",
  17885=>"001011000",
  17886=>"001111001",
  17887=>"110100011",
  17888=>"000000011",
  17889=>"110100110",
  17890=>"111010101",
  17891=>"100101110",
  17892=>"110110000",
  17893=>"100111010",
  17894=>"111000110",
  17895=>"000000101",
  17896=>"101011011",
  17897=>"000001010",
  17898=>"000110001",
  17899=>"101101100",
  17900=>"110000100",
  17901=>"101110101",
  17902=>"100011101",
  17903=>"001000111",
  17904=>"010101100",
  17905=>"100101010",
  17906=>"110010001",
  17907=>"011000110",
  17908=>"110000001",
  17909=>"000111011",
  17910=>"000001110",
  17911=>"100101001",
  17912=>"111011111",
  17913=>"101001100",
  17914=>"001110100",
  17915=>"001010100",
  17916=>"111000000",
  17917=>"110100101",
  17918=>"110001001",
  17919=>"101111100",
  17920=>"111100101",
  17921=>"001001111",
  17922=>"110000010",
  17923=>"001100001",
  17924=>"000100110",
  17925=>"000110011",
  17926=>"011111000",
  17927=>"111111111",
  17928=>"111011010",
  17929=>"110110110",
  17930=>"101010101",
  17931=>"001100001",
  17932=>"111000010",
  17933=>"111111011",
  17934=>"001111101",
  17935=>"001100011",
  17936=>"000011001",
  17937=>"000100101",
  17938=>"000101101",
  17939=>"001111000",
  17940=>"100001101",
  17941=>"010000111",
  17942=>"010011101",
  17943=>"010011110",
  17944=>"010010010",
  17945=>"010101000",
  17946=>"100011010",
  17947=>"110111010",
  17948=>"000110010",
  17949=>"101000111",
  17950=>"011100101",
  17951=>"101010011",
  17952=>"011111000",
  17953=>"111000111",
  17954=>"111000010",
  17955=>"101011100",
  17956=>"110100010",
  17957=>"100011001",
  17958=>"011010001",
  17959=>"011111100",
  17960=>"101011000",
  17961=>"000101111",
  17962=>"011001110",
  17963=>"110110000",
  17964=>"101111000",
  17965=>"011001000",
  17966=>"100101111",
  17967=>"011010111",
  17968=>"000001010",
  17969=>"010001001",
  17970=>"011001100",
  17971=>"011110000",
  17972=>"110101011",
  17973=>"000001110",
  17974=>"011110111",
  17975=>"110011001",
  17976=>"010011010",
  17977=>"111001110",
  17978=>"100101011",
  17979=>"010111011",
  17980=>"111010011",
  17981=>"000001001",
  17982=>"000100110",
  17983=>"100110001",
  17984=>"101001101",
  17985=>"010011111",
  17986=>"111101011",
  17987=>"011010110",
  17988=>"010011011",
  17989=>"100000001",
  17990=>"010010011",
  17991=>"001110010",
  17992=>"000001110",
  17993=>"010001000",
  17994=>"101110111",
  17995=>"111010010",
  17996=>"101111011",
  17997=>"010001000",
  17998=>"011011010",
  17999=>"001001100",
  18000=>"110011100",
  18001=>"111101110",
  18002=>"010010000",
  18003=>"001010100",
  18004=>"010100100",
  18005=>"011000111",
  18006=>"110000000",
  18007=>"101100101",
  18008=>"000000010",
  18009=>"000000110",
  18010=>"111101110",
  18011=>"011011000",
  18012=>"000110110",
  18013=>"111000000",
  18014=>"111011111",
  18015=>"110000010",
  18016=>"010101100",
  18017=>"010001010",
  18018=>"000000000",
  18019=>"100101010",
  18020=>"000011000",
  18021=>"101010010",
  18022=>"110110000",
  18023=>"000011010",
  18024=>"100000100",
  18025=>"000010001",
  18026=>"011101011",
  18027=>"110111001",
  18028=>"000100001",
  18029=>"101000101",
  18030=>"100000110",
  18031=>"010010000",
  18032=>"111101000",
  18033=>"000001100",
  18034=>"011110110",
  18035=>"001100010",
  18036=>"011111000",
  18037=>"000000001",
  18038=>"111101111",
  18039=>"101101111",
  18040=>"011111000",
  18041=>"110000010",
  18042=>"000010111",
  18043=>"100011101",
  18044=>"001100010",
  18045=>"110011001",
  18046=>"010100011",
  18047=>"000111111",
  18048=>"000100001",
  18049=>"110001100",
  18050=>"001010011",
  18051=>"001001101",
  18052=>"100111101",
  18053=>"101000000",
  18054=>"011000101",
  18055=>"111100110",
  18056=>"010010011",
  18057=>"110101000",
  18058=>"001111101",
  18059=>"111100000",
  18060=>"111101111",
  18061=>"010100000",
  18062=>"000110110",
  18063=>"001000000",
  18064=>"100110101",
  18065=>"011011111",
  18066=>"101110110",
  18067=>"011101100",
  18068=>"011101010",
  18069=>"001100111",
  18070=>"101100011",
  18071=>"011111111",
  18072=>"100101101",
  18073=>"011011110",
  18074=>"100101111",
  18075=>"010001001",
  18076=>"010000101",
  18077=>"100101111",
  18078=>"100111011",
  18079=>"111100101",
  18080=>"010010110",
  18081=>"010100011",
  18082=>"100010100",
  18083=>"010000110",
  18084=>"001000001",
  18085=>"101101000",
  18086=>"000010100",
  18087=>"000000000",
  18088=>"111011001",
  18089=>"110010101",
  18090=>"101011000",
  18091=>"100000000",
  18092=>"100010100",
  18093=>"001011000",
  18094=>"100000010",
  18095=>"000110000",
  18096=>"000101000",
  18097=>"101000101",
  18098=>"111011111",
  18099=>"110111001",
  18100=>"100001111",
  18101=>"101100011",
  18102=>"000110011",
  18103=>"111000000",
  18104=>"100000011",
  18105=>"110011111",
  18106=>"110101100",
  18107=>"100001011",
  18108=>"111111011",
  18109=>"110001000",
  18110=>"010001000",
  18111=>"101101111",
  18112=>"011100110",
  18113=>"111111000",
  18114=>"000001000",
  18115=>"110001011",
  18116=>"000100011",
  18117=>"100100011",
  18118=>"001001001",
  18119=>"000100010",
  18120=>"000010011",
  18121=>"100001010",
  18122=>"110100001",
  18123=>"000001101",
  18124=>"110011011",
  18125=>"000000111",
  18126=>"001111000",
  18127=>"111011000",
  18128=>"011110000",
  18129=>"110010111",
  18130=>"111101110",
  18131=>"000001011",
  18132=>"011000110",
  18133=>"010101100",
  18134=>"011110111",
  18135=>"110011100",
  18136=>"000101101",
  18137=>"100101100",
  18138=>"000111101",
  18139=>"010100110",
  18140=>"110100101",
  18141=>"010110110",
  18142=>"000111110",
  18143=>"011001111",
  18144=>"001000010",
  18145=>"100101101",
  18146=>"100100111",
  18147=>"000111111",
  18148=>"001111110",
  18149=>"000001001",
  18150=>"100001000",
  18151=>"000000100",
  18152=>"010000000",
  18153=>"101011110",
  18154=>"001111111",
  18155=>"001011101",
  18156=>"100000100",
  18157=>"100000000",
  18158=>"001101101",
  18159=>"010011111",
  18160=>"010010001",
  18161=>"000100010",
  18162=>"000000001",
  18163=>"011010000",
  18164=>"100001011",
  18165=>"001100010",
  18166=>"001011111",
  18167=>"011000110",
  18168=>"001100100",
  18169=>"010111111",
  18170=>"011010101",
  18171=>"011011010",
  18172=>"011010010",
  18173=>"000001111",
  18174=>"111011001",
  18175=>"000110110",
  18176=>"001001101",
  18177=>"100011101",
  18178=>"111110010",
  18179=>"001000001",
  18180=>"000110100",
  18181=>"101000010",
  18182=>"010000011",
  18183=>"100110000",
  18184=>"001110101",
  18185=>"000111100",
  18186=>"001100111",
  18187=>"011001101",
  18188=>"100011100",
  18189=>"100101111",
  18190=>"111010011",
  18191=>"010010001",
  18192=>"110101001",
  18193=>"111000101",
  18194=>"001110011",
  18195=>"110001100",
  18196=>"000101001",
  18197=>"000001110",
  18198=>"000110110",
  18199=>"111000100",
  18200=>"001011101",
  18201=>"111101010",
  18202=>"010110010",
  18203=>"000111011",
  18204=>"001111111",
  18205=>"101101010",
  18206=>"001010011",
  18207=>"100000000",
  18208=>"111101000",
  18209=>"101000111",
  18210=>"111111000",
  18211=>"000000011",
  18212=>"011010010",
  18213=>"011000000",
  18214=>"001001111",
  18215=>"111110100",
  18216=>"101010011",
  18217=>"100010101",
  18218=>"110010100",
  18219=>"010011110",
  18220=>"011010000",
  18221=>"000010001",
  18222=>"100111010",
  18223=>"111011010",
  18224=>"011100101",
  18225=>"010000101",
  18226=>"111100110",
  18227=>"111001000",
  18228=>"000000101",
  18229=>"011110011",
  18230=>"000100101",
  18231=>"011011100",
  18232=>"010110111",
  18233=>"001010100",
  18234=>"011011101",
  18235=>"101101001",
  18236=>"000000000",
  18237=>"000001011",
  18238=>"100001010",
  18239=>"010100001",
  18240=>"110111001",
  18241=>"000001011",
  18242=>"001011110",
  18243=>"110111110",
  18244=>"110011011",
  18245=>"111110111",
  18246=>"100100111",
  18247=>"110011111",
  18248=>"001100011",
  18249=>"111000001",
  18250=>"100110010",
  18251=>"011101011",
  18252=>"111001110",
  18253=>"000110100",
  18254=>"001011001",
  18255=>"011011111",
  18256=>"110110100",
  18257=>"101110110",
  18258=>"000000101",
  18259=>"100011101",
  18260=>"011011010",
  18261=>"110100010",
  18262=>"011101011",
  18263=>"001101001",
  18264=>"001100110",
  18265=>"110000000",
  18266=>"101100011",
  18267=>"000001110",
  18268=>"111111110",
  18269=>"110010101",
  18270=>"011111010",
  18271=>"010001000",
  18272=>"011011011",
  18273=>"111110010",
  18274=>"010101100",
  18275=>"110110111",
  18276=>"001101111",
  18277=>"000001111",
  18278=>"010100011",
  18279=>"011001000",
  18280=>"101010001",
  18281=>"011010111",
  18282=>"111100011",
  18283=>"011010000",
  18284=>"000010100",
  18285=>"111110000",
  18286=>"001001100",
  18287=>"010101001",
  18288=>"110111111",
  18289=>"111001111",
  18290=>"000100100",
  18291=>"100100101",
  18292=>"110010011",
  18293=>"101000011",
  18294=>"011010110",
  18295=>"100001000",
  18296=>"011111100",
  18297=>"100000001",
  18298=>"001011001",
  18299=>"000110001",
  18300=>"101011000",
  18301=>"010010110",
  18302=>"001010101",
  18303=>"110111010",
  18304=>"010001100",
  18305=>"100100111",
  18306=>"110111101",
  18307=>"011011100",
  18308=>"111101000",
  18309=>"011000100",
  18310=>"100101000",
  18311=>"001011011",
  18312=>"011011010",
  18313=>"000100100",
  18314=>"101000111",
  18315=>"001111100",
  18316=>"000011011",
  18317=>"001101101",
  18318=>"101111001",
  18319=>"011000100",
  18320=>"011000100",
  18321=>"011011100",
  18322=>"111011001",
  18323=>"010001000",
  18324=>"000100111",
  18325=>"000101011",
  18326=>"111000010",
  18327=>"001011110",
  18328=>"001110000",
  18329=>"011101110",
  18330=>"100001010",
  18331=>"101000001",
  18332=>"000110100",
  18333=>"010110110",
  18334=>"100100001",
  18335=>"101111011",
  18336=>"010110111",
  18337=>"101011011",
  18338=>"110110001",
  18339=>"101100011",
  18340=>"011111001",
  18341=>"000000011",
  18342=>"100011110",
  18343=>"010011111",
  18344=>"101110111",
  18345=>"110010110",
  18346=>"111111010",
  18347=>"101011000",
  18348=>"011101110",
  18349=>"001000001",
  18350=>"101101111",
  18351=>"111001111",
  18352=>"100001101",
  18353=>"000000110",
  18354=>"111101001",
  18355=>"100100000",
  18356=>"111100110",
  18357=>"100001011",
  18358=>"100000110",
  18359=>"011000001",
  18360=>"110110011",
  18361=>"111111111",
  18362=>"010110001",
  18363=>"111001000",
  18364=>"100010101",
  18365=>"001100100",
  18366=>"101110010",
  18367=>"101011001",
  18368=>"110101010",
  18369=>"010011000",
  18370=>"100000000",
  18371=>"001011101",
  18372=>"000100010",
  18373=>"010101101",
  18374=>"101111111",
  18375=>"011100001",
  18376=>"100111000",
  18377=>"000010110",
  18378=>"001101101",
  18379=>"111110100",
  18380=>"101011111",
  18381=>"111011011",
  18382=>"111000011",
  18383=>"010011010",
  18384=>"100101101",
  18385=>"010101110",
  18386=>"100100110",
  18387=>"011000101",
  18388=>"000001101",
  18389=>"110110000",
  18390=>"010011000",
  18391=>"111101110",
  18392=>"010100001",
  18393=>"001011000",
  18394=>"111011100",
  18395=>"110111010",
  18396=>"111001011",
  18397=>"010111000",
  18398=>"110001101",
  18399=>"000010101",
  18400=>"110110100",
  18401=>"010101110",
  18402=>"100111001",
  18403=>"101100000",
  18404=>"110001110",
  18405=>"101100111",
  18406=>"100010110",
  18407=>"001001100",
  18408=>"001100000",
  18409=>"110101001",
  18410=>"100110100",
  18411=>"110101101",
  18412=>"010110010",
  18413=>"110100100",
  18414=>"100110110",
  18415=>"011010000",
  18416=>"111000101",
  18417=>"110000010",
  18418=>"000111010",
  18419=>"001000011",
  18420=>"101111101",
  18421=>"000011101",
  18422=>"111010101",
  18423=>"100000000",
  18424=>"000111101",
  18425=>"100111111",
  18426=>"110101111",
  18427=>"010010111",
  18428=>"000010001",
  18429=>"010010100",
  18430=>"001101011",
  18431=>"000011000",
  18432=>"010000101",
  18433=>"010100100",
  18434=>"110010000",
  18435=>"011010001",
  18436=>"000000000",
  18437=>"010101100",
  18438=>"011110000",
  18439=>"100010011",
  18440=>"111101100",
  18441=>"101011100",
  18442=>"001011011",
  18443=>"100011111",
  18444=>"111100001",
  18445=>"101001101",
  18446=>"111001011",
  18447=>"000001111",
  18448=>"110010111",
  18449=>"110000000",
  18450=>"110101101",
  18451=>"101101101",
  18452=>"100100011",
  18453=>"010110000",
  18454=>"001000110",
  18455=>"001100010",
  18456=>"100001101",
  18457=>"111010010",
  18458=>"001111111",
  18459=>"101001100",
  18460=>"011010011",
  18461=>"001110100",
  18462=>"001010100",
  18463=>"111000100",
  18464=>"110110111",
  18465=>"110100100",
  18466=>"000000000",
  18467=>"111110110",
  18468=>"101011101",
  18469=>"100001001",
  18470=>"011101110",
  18471=>"010100000",
  18472=>"111111010",
  18473=>"101100100",
  18474=>"000110100",
  18475=>"010011010",
  18476=>"010010000",
  18477=>"111000101",
  18478=>"100000101",
  18479=>"000110101",
  18480=>"000000111",
  18481=>"101100010",
  18482=>"011011111",
  18483=>"111110010",
  18484=>"111010001",
  18485=>"011100100",
  18486=>"001111111",
  18487=>"000111100",
  18488=>"000111011",
  18489=>"000010100",
  18490=>"100011111",
  18491=>"101000000",
  18492=>"000010011",
  18493=>"000100010",
  18494=>"001000001",
  18495=>"010111010",
  18496=>"000011000",
  18497=>"110101011",
  18498=>"110001101",
  18499=>"001101101",
  18500=>"110011000",
  18501=>"111100101",
  18502=>"110000101",
  18503=>"100010010",
  18504=>"001000011",
  18505=>"110100110",
  18506=>"100101000",
  18507=>"010011001",
  18508=>"110101100",
  18509=>"111010110",
  18510=>"011111000",
  18511=>"011110000",
  18512=>"100100111",
  18513=>"111010110",
  18514=>"001111100",
  18515=>"001000101",
  18516=>"110011000",
  18517=>"000011100",
  18518=>"101101110",
  18519=>"110010001",
  18520=>"100011111",
  18521=>"011100000",
  18522=>"011011110",
  18523=>"110011110",
  18524=>"010110111",
  18525=>"100001110",
  18526=>"110100011",
  18527=>"111110010",
  18528=>"101000110",
  18529=>"001000000",
  18530=>"111100000",
  18531=>"001100011",
  18532=>"100111110",
  18533=>"100010000",
  18534=>"111100110",
  18535=>"101010101",
  18536=>"101100011",
  18537=>"110001101",
  18538=>"110100110",
  18539=>"111110100",
  18540=>"011001101",
  18541=>"000011011",
  18542=>"001001000",
  18543=>"010100110",
  18544=>"101111110",
  18545=>"000001000",
  18546=>"100111110",
  18547=>"111101000",
  18548=>"010010100",
  18549=>"100110010",
  18550=>"001011110",
  18551=>"100001001",
  18552=>"011101001",
  18553=>"000001011",
  18554=>"100001011",
  18555=>"001101100",
  18556=>"001001000",
  18557=>"101101101",
  18558=>"001011010",
  18559=>"100010111",
  18560=>"101000110",
  18561=>"000101001",
  18562=>"000001100",
  18563=>"000111111",
  18564=>"110000001",
  18565=>"010110101",
  18566=>"001100001",
  18567=>"100000000",
  18568=>"101011001",
  18569=>"111101111",
  18570=>"111000100",
  18571=>"110001100",
  18572=>"011111111",
  18573=>"110000010",
  18574=>"001100100",
  18575=>"101111100",
  18576=>"001101000",
  18577=>"001110100",
  18578=>"100010010",
  18579=>"011111011",
  18580=>"010101011",
  18581=>"000000010",
  18582=>"101110001",
  18583=>"010000010",
  18584=>"100010101",
  18585=>"011000101",
  18586=>"011111010",
  18587=>"011010000",
  18588=>"101100101",
  18589=>"001110100",
  18590=>"101101011",
  18591=>"100000110",
  18592=>"001111100",
  18593=>"001000011",
  18594=>"101101101",
  18595=>"111001100",
  18596=>"111000110",
  18597=>"110111001",
  18598=>"001001101",
  18599=>"100010110",
  18600=>"011110100",
  18601=>"010101101",
  18602=>"101110110",
  18603=>"110101010",
  18604=>"101011011",
  18605=>"100010000",
  18606=>"000010010",
  18607=>"100000000",
  18608=>"101000010",
  18609=>"111101100",
  18610=>"011111101",
  18611=>"000010100",
  18612=>"011001001",
  18613=>"010001011",
  18614=>"001001010",
  18615=>"111110111",
  18616=>"001101011",
  18617=>"010111000",
  18618=>"101010100",
  18619=>"111000101",
  18620=>"000000100",
  18621=>"000101010",
  18622=>"101001101",
  18623=>"000101000",
  18624=>"010000101",
  18625=>"000011011",
  18626=>"000011101",
  18627=>"100111100",
  18628=>"100011111",
  18629=>"011000001",
  18630=>"000010011",
  18631=>"110000001",
  18632=>"001110111",
  18633=>"100101101",
  18634=>"111100110",
  18635=>"000100011",
  18636=>"111100101",
  18637=>"110111100",
  18638=>"011111010",
  18639=>"010011001",
  18640=>"001111100",
  18641=>"101111110",
  18642=>"000010000",
  18643=>"100111101",
  18644=>"001010011",
  18645=>"010110011",
  18646=>"100101010",
  18647=>"111001001",
  18648=>"111011110",
  18649=>"111111101",
  18650=>"111101010",
  18651=>"011000010",
  18652=>"001100111",
  18653=>"010001001",
  18654=>"111000100",
  18655=>"100110011",
  18656=>"100010001",
  18657=>"110101000",
  18658=>"000001011",
  18659=>"000111001",
  18660=>"001001011",
  18661=>"000011111",
  18662=>"011001111",
  18663=>"001010010",
  18664=>"110101001",
  18665=>"110101000",
  18666=>"000110001",
  18667=>"101011111",
  18668=>"111111100",
  18669=>"000101100",
  18670=>"011011111",
  18671=>"000101100",
  18672=>"111110001",
  18673=>"100010111",
  18674=>"000100000",
  18675=>"100000111",
  18676=>"001101010",
  18677=>"000011100",
  18678=>"001100100",
  18679=>"000101001",
  18680=>"000010111",
  18681=>"111110010",
  18682=>"011110101",
  18683=>"011011000",
  18684=>"100011001",
  18685=>"011100010",
  18686=>"110000110",
  18687=>"010001110",
  18688=>"101111101",
  18689=>"000010111",
  18690=>"110000101",
  18691=>"101111001",
  18692=>"101110010",
  18693=>"100110111",
  18694=>"001001011",
  18695=>"001100111",
  18696=>"110001000",
  18697=>"001001010",
  18698=>"101000000",
  18699=>"110010111",
  18700=>"101101101",
  18701=>"001001010",
  18702=>"101001010",
  18703=>"010000011",
  18704=>"101100110",
  18705=>"110100001",
  18706=>"000010011",
  18707=>"100011011",
  18708=>"000100110",
  18709=>"111110010",
  18710=>"000000110",
  18711=>"010000001",
  18712=>"111110100",
  18713=>"100101101",
  18714=>"000010011",
  18715=>"100010000",
  18716=>"011110110",
  18717=>"111011111",
  18718=>"100001110",
  18719=>"000111001",
  18720=>"000001110",
  18721=>"100101001",
  18722=>"110011100",
  18723=>"100000010",
  18724=>"011010100",
  18725=>"000100100",
  18726=>"110101010",
  18727=>"010011101",
  18728=>"111000001",
  18729=>"000011001",
  18730=>"000010001",
  18731=>"011111100",
  18732=>"010010011",
  18733=>"000101001",
  18734=>"010010011",
  18735=>"111110010",
  18736=>"001001100",
  18737=>"011110110",
  18738=>"110111111",
  18739=>"010001101",
  18740=>"111000110",
  18741=>"010011101",
  18742=>"000000100",
  18743=>"011001001",
  18744=>"110111101",
  18745=>"110100101",
  18746=>"100000001",
  18747=>"101001011",
  18748=>"110011000",
  18749=>"111011011",
  18750=>"000000010",
  18751=>"100111110",
  18752=>"010101000",
  18753=>"000111001",
  18754=>"000101110",
  18755=>"101011100",
  18756=>"010111111",
  18757=>"100110000",
  18758=>"100010010",
  18759=>"101110000",
  18760=>"000010010",
  18761=>"111111110",
  18762=>"011010110",
  18763=>"111111101",
  18764=>"000010010",
  18765=>"010111100",
  18766=>"000011101",
  18767=>"001010101",
  18768=>"100110100",
  18769=>"101001000",
  18770=>"011000111",
  18771=>"100111010",
  18772=>"011110000",
  18773=>"111001001",
  18774=>"100101110",
  18775=>"000011000",
  18776=>"000100000",
  18777=>"110100011",
  18778=>"001101110",
  18779=>"000111101",
  18780=>"100000010",
  18781=>"111100001",
  18782=>"010001110",
  18783=>"011000110",
  18784=>"100100111",
  18785=>"001111111",
  18786=>"010001010",
  18787=>"000010110",
  18788=>"000110011",
  18789=>"110001001",
  18790=>"000111100",
  18791=>"110000111",
  18792=>"101000100",
  18793=>"011000110",
  18794=>"110001111",
  18795=>"100010100",
  18796=>"001111011",
  18797=>"111100000",
  18798=>"001110100",
  18799=>"011111100",
  18800=>"101000001",
  18801=>"000011011",
  18802=>"001010110",
  18803=>"000011000",
  18804=>"100101111",
  18805=>"001100001",
  18806=>"110111010",
  18807=>"010010011",
  18808=>"000110000",
  18809=>"110101100",
  18810=>"001011111",
  18811=>"100001110",
  18812=>"000010001",
  18813=>"001110111",
  18814=>"001010100",
  18815=>"010101001",
  18816=>"010011000",
  18817=>"011000001",
  18818=>"000110100",
  18819=>"000111111",
  18820=>"011011011",
  18821=>"001011000",
  18822=>"011011111",
  18823=>"101111001",
  18824=>"001000000",
  18825=>"110001001",
  18826=>"111010101",
  18827=>"011010001",
  18828=>"010101001",
  18829=>"100101010",
  18830=>"000011011",
  18831=>"000101100",
  18832=>"101001010",
  18833=>"011010111",
  18834=>"111001111",
  18835=>"010100010",
  18836=>"101101111",
  18837=>"100100011",
  18838=>"100100011",
  18839=>"000011101",
  18840=>"011111011",
  18841=>"010010111",
  18842=>"110001101",
  18843=>"010000101",
  18844=>"000111111",
  18845=>"000100000",
  18846=>"101101111",
  18847=>"111111111",
  18848=>"101010100",
  18849=>"111100010",
  18850=>"100001000",
  18851=>"001110111",
  18852=>"011001010",
  18853=>"000101111",
  18854=>"111111011",
  18855=>"111110000",
  18856=>"101010001",
  18857=>"000100110",
  18858=>"011111110",
  18859=>"010111111",
  18860=>"101100100",
  18861=>"110011110",
  18862=>"001111000",
  18863=>"111011000",
  18864=>"000101001",
  18865=>"011000000",
  18866=>"111100100",
  18867=>"111101011",
  18868=>"001001011",
  18869=>"000000101",
  18870=>"000011111",
  18871=>"000101000",
  18872=>"100010111",
  18873=>"010100110",
  18874=>"000100001",
  18875=>"000011010",
  18876=>"100100110",
  18877=>"011000101",
  18878=>"110011001",
  18879=>"010000000",
  18880=>"000000110",
  18881=>"000100011",
  18882=>"000101110",
  18883=>"110001100",
  18884=>"100101000",
  18885=>"001001000",
  18886=>"111111001",
  18887=>"011000011",
  18888=>"101011110",
  18889=>"110010110",
  18890=>"100001001",
  18891=>"111010111",
  18892=>"010100100",
  18893=>"001010100",
  18894=>"101111110",
  18895=>"110011000",
  18896=>"111010001",
  18897=>"100101110",
  18898=>"010101101",
  18899=>"000111110",
  18900=>"011000000",
  18901=>"110001111",
  18902=>"001100010",
  18903=>"101011100",
  18904=>"111000011",
  18905=>"100001000",
  18906=>"111100000",
  18907=>"100001000",
  18908=>"101101100",
  18909=>"101010000",
  18910=>"011111110",
  18911=>"100101111",
  18912=>"100000000",
  18913=>"000111101",
  18914=>"100110010",
  18915=>"111100111",
  18916=>"010001101",
  18917=>"110010010",
  18918=>"110010001",
  18919=>"000001110",
  18920=>"100000100",
  18921=>"011001100",
  18922=>"111011101",
  18923=>"100101011",
  18924=>"001011001",
  18925=>"100111001",
  18926=>"101110100",
  18927=>"011110101",
  18928=>"000110000",
  18929=>"111011000",
  18930=>"111100100",
  18931=>"010001001",
  18932=>"111101010",
  18933=>"101011111",
  18934=>"000100100",
  18935=>"000111101",
  18936=>"011101000",
  18937=>"101110010",
  18938=>"111110010",
  18939=>"101110001",
  18940=>"010000011",
  18941=>"101110110",
  18942=>"011000100",
  18943=>"011010101",
  18944=>"100111110",
  18945=>"111010111",
  18946=>"011000000",
  18947=>"001111001",
  18948=>"101101000",
  18949=>"100011011",
  18950=>"100100001",
  18951=>"001011010",
  18952=>"100111000",
  18953=>"110110000",
  18954=>"111101101",
  18955=>"001111011",
  18956=>"110110111",
  18957=>"110011110",
  18958=>"101111001",
  18959=>"111001110",
  18960=>"100101111",
  18961=>"011110011",
  18962=>"010101111",
  18963=>"010011000",
  18964=>"100111100",
  18965=>"111111100",
  18966=>"000100011",
  18967=>"000100110",
  18968=>"110011000",
  18969=>"101000000",
  18970=>"010011001",
  18971=>"111101011",
  18972=>"011110111",
  18973=>"110101111",
  18974=>"010010011",
  18975=>"001110101",
  18976=>"110010000",
  18977=>"011111100",
  18978=>"010001110",
  18979=>"010100010",
  18980=>"000010101",
  18981=>"010101000",
  18982=>"101101001",
  18983=>"001000111",
  18984=>"111101101",
  18985=>"100110111",
  18986=>"001011000",
  18987=>"011110101",
  18988=>"111111101",
  18989=>"001101011",
  18990=>"011011010",
  18991=>"111001000",
  18992=>"011101101",
  18993=>"101010010",
  18994=>"100011100",
  18995=>"000100000",
  18996=>"111111011",
  18997=>"101010110",
  18998=>"111101010",
  18999=>"100010110",
  19000=>"101011101",
  19001=>"101111011",
  19002=>"001011111",
  19003=>"011000000",
  19004=>"000100110",
  19005=>"001011101",
  19006=>"110001100",
  19007=>"101110100",
  19008=>"000001100",
  19009=>"100011001",
  19010=>"111110001",
  19011=>"000100111",
  19012=>"010100110",
  19013=>"001110100",
  19014=>"101100111",
  19015=>"011000001",
  19016=>"110011000",
  19017=>"101010110",
  19018=>"011101000",
  19019=>"100100110",
  19020=>"011111011",
  19021=>"000000000",
  19022=>"010001111",
  19023=>"110000111",
  19024=>"100101111",
  19025=>"000001001",
  19026=>"011000110",
  19027=>"000110001",
  19028=>"100100111",
  19029=>"011010101",
  19030=>"110011011",
  19031=>"110101110",
  19032=>"111111010",
  19033=>"110000001",
  19034=>"111110100",
  19035=>"000001010",
  19036=>"000111011",
  19037=>"001001110",
  19038=>"111001011",
  19039=>"011001101",
  19040=>"100011010",
  19041=>"101000101",
  19042=>"110010101",
  19043=>"100000111",
  19044=>"011011000",
  19045=>"100010110",
  19046=>"110011100",
  19047=>"111100010",
  19048=>"000010100",
  19049=>"011001101",
  19050=>"010110010",
  19051=>"100111001",
  19052=>"001001001",
  19053=>"010001010",
  19054=>"000100111",
  19055=>"000010111",
  19056=>"001011000",
  19057=>"110001110",
  19058=>"110101101",
  19059=>"001101100",
  19060=>"111010001",
  19061=>"111011101",
  19062=>"000001001",
  19063=>"010010011",
  19064=>"000101110",
  19065=>"000111000",
  19066=>"100100011",
  19067=>"011100100",
  19068=>"011110011",
  19069=>"110010001",
  19070=>"100110010",
  19071=>"001010000",
  19072=>"001001010",
  19073=>"100011100",
  19074=>"000010100",
  19075=>"001010001",
  19076=>"000011100",
  19077=>"000001101",
  19078=>"101001100",
  19079=>"111100111",
  19080=>"000010100",
  19081=>"011110111",
  19082=>"111000110",
  19083=>"110111001",
  19084=>"001001000",
  19085=>"000011110",
  19086=>"111000000",
  19087=>"101001010",
  19088=>"000111010",
  19089=>"010011010",
  19090=>"100000111",
  19091=>"101101011",
  19092=>"011110111",
  19093=>"101110111",
  19094=>"010100100",
  19095=>"110011101",
  19096=>"001011010",
  19097=>"001101001",
  19098=>"000111111",
  19099=>"011100001",
  19100=>"010011010",
  19101=>"111101000",
  19102=>"101100100",
  19103=>"101100000",
  19104=>"111011011",
  19105=>"010110000",
  19106=>"111101101",
  19107=>"000010000",
  19108=>"101001000",
  19109=>"101110011",
  19110=>"001011111",
  19111=>"011000010",
  19112=>"111111001",
  19113=>"100011000",
  19114=>"100100010",
  19115=>"111100001",
  19116=>"010101100",
  19117=>"111011000",
  19118=>"011110111",
  19119=>"001000100",
  19120=>"011110111",
  19121=>"111100000",
  19122=>"010101010",
  19123=>"100010001",
  19124=>"100110110",
  19125=>"000100100",
  19126=>"110111000",
  19127=>"001001001",
  19128=>"001101110",
  19129=>"000000101",
  19130=>"111110011",
  19131=>"100110000",
  19132=>"000001110",
  19133=>"010101111",
  19134=>"010011100",
  19135=>"111011000",
  19136=>"100001001",
  19137=>"000110011",
  19138=>"110001100",
  19139=>"101001000",
  19140=>"110111010",
  19141=>"010011011",
  19142=>"010111111",
  19143=>"000010110",
  19144=>"001010010",
  19145=>"100101101",
  19146=>"001001010",
  19147=>"111111011",
  19148=>"110110101",
  19149=>"111011100",
  19150=>"001110101",
  19151=>"010100110",
  19152=>"011000011",
  19153=>"001110110",
  19154=>"111100000",
  19155=>"010101001",
  19156=>"111111111",
  19157=>"101001111",
  19158=>"000100100",
  19159=>"101010100",
  19160=>"010011111",
  19161=>"111000010",
  19162=>"010101010",
  19163=>"111001000",
  19164=>"100010000",
  19165=>"111100000",
  19166=>"100011001",
  19167=>"110101011",
  19168=>"001101011",
  19169=>"001110000",
  19170=>"101010111",
  19171=>"011101101",
  19172=>"011011011",
  19173=>"111110101",
  19174=>"000100000",
  19175=>"011000000",
  19176=>"000110111",
  19177=>"110010111",
  19178=>"000010010",
  19179=>"011100110",
  19180=>"111111100",
  19181=>"100100111",
  19182=>"001011101",
  19183=>"001000010",
  19184=>"110000001",
  19185=>"000000001",
  19186=>"100101001",
  19187=>"100001100",
  19188=>"000110101",
  19189=>"101100111",
  19190=>"011100000",
  19191=>"000001111",
  19192=>"001101111",
  19193=>"010110111",
  19194=>"101001111",
  19195=>"110001100",
  19196=>"000001011",
  19197=>"001111111",
  19198=>"010100001",
  19199=>"011001100",
  19200=>"111010010",
  19201=>"100001100",
  19202=>"010110101",
  19203=>"101100110",
  19204=>"110110101",
  19205=>"001000100",
  19206=>"000010000",
  19207=>"101001010",
  19208=>"001011101",
  19209=>"000010101",
  19210=>"011110101",
  19211=>"000101001",
  19212=>"100101000",
  19213=>"001011100",
  19214=>"011110010",
  19215=>"110111011",
  19216=>"011010001",
  19217=>"000000111",
  19218=>"111010111",
  19219=>"001100100",
  19220=>"100100101",
  19221=>"110110010",
  19222=>"100100010",
  19223=>"111100000",
  19224=>"001100011",
  19225=>"100001010",
  19226=>"100011111",
  19227=>"010110110",
  19228=>"000100001",
  19229=>"011011011",
  19230=>"011111001",
  19231=>"001000010",
  19232=>"100010011",
  19233=>"111100001",
  19234=>"110110110",
  19235=>"101111000",
  19236=>"110001100",
  19237=>"101110011",
  19238=>"011111000",
  19239=>"011100001",
  19240=>"101001111",
  19241=>"011100100",
  19242=>"001111101",
  19243=>"100000011",
  19244=>"100000110",
  19245=>"000101101",
  19246=>"000101001",
  19247=>"101001011",
  19248=>"000010001",
  19249=>"011010011",
  19250=>"111100000",
  19251=>"000111110",
  19252=>"001111010",
  19253=>"111111101",
  19254=>"101011100",
  19255=>"001000011",
  19256=>"100010011",
  19257=>"100000101",
  19258=>"010010000",
  19259=>"010100010",
  19260=>"010000100",
  19261=>"011100111",
  19262=>"010001000",
  19263=>"100011000",
  19264=>"010000011",
  19265=>"010010100",
  19266=>"010111111",
  19267=>"100100000",
  19268=>"000000000",
  19269=>"100110011",
  19270=>"000000001",
  19271=>"000110101",
  19272=>"010000101",
  19273=>"100011111",
  19274=>"001110010",
  19275=>"000101111",
  19276=>"001010001",
  19277=>"001111100",
  19278=>"011010001",
  19279=>"001101111",
  19280=>"101100000",
  19281=>"001100100",
  19282=>"001000101",
  19283=>"110000000",
  19284=>"101011100",
  19285=>"001101000",
  19286=>"110111010",
  19287=>"100001001",
  19288=>"000110000",
  19289=>"100100011",
  19290=>"011000110",
  19291=>"111001000",
  19292=>"011101001",
  19293=>"000010010",
  19294=>"011011101",
  19295=>"110011000",
  19296=>"011100011",
  19297=>"011111000",
  19298=>"000011110",
  19299=>"000101100",
  19300=>"111001010",
  19301=>"100111100",
  19302=>"110100001",
  19303=>"010000010",
  19304=>"110111000",
  19305=>"100011010",
  19306=>"110110010",
  19307=>"000010111",
  19308=>"101011110",
  19309=>"001101110",
  19310=>"100000110",
  19311=>"101101101",
  19312=>"011101111",
  19313=>"011011010",
  19314=>"101011011",
  19315=>"010110110",
  19316=>"001011010",
  19317=>"000000000",
  19318=>"000011101",
  19319=>"011101110",
  19320=>"011111110",
  19321=>"111011000",
  19322=>"011101011",
  19323=>"001010110",
  19324=>"101100000",
  19325=>"110011011",
  19326=>"111110001",
  19327=>"011010000",
  19328=>"000101111",
  19329=>"010100001",
  19330=>"001011010",
  19331=>"000100101",
  19332=>"110000101",
  19333=>"101111100",
  19334=>"000000001",
  19335=>"011110001",
  19336=>"011100111",
  19337=>"001000101",
  19338=>"101011101",
  19339=>"001011001",
  19340=>"011000011",
  19341=>"010000111",
  19342=>"001100101",
  19343=>"010010101",
  19344=>"000011000",
  19345=>"011001011",
  19346=>"110011000",
  19347=>"101010110",
  19348=>"101010010",
  19349=>"011000000",
  19350=>"001110000",
  19351=>"101100000",
  19352=>"000010100",
  19353=>"111011000",
  19354=>"111010000",
  19355=>"011011111",
  19356=>"110011000",
  19357=>"111010011",
  19358=>"111011111",
  19359=>"111000110",
  19360=>"011100010",
  19361=>"001011011",
  19362=>"000101001",
  19363=>"101100001",
  19364=>"100110100",
  19365=>"000111011",
  19366=>"100111001",
  19367=>"010111111",
  19368=>"001101101",
  19369=>"000110000",
  19370=>"101111100",
  19371=>"001110001",
  19372=>"000011111",
  19373=>"110000100",
  19374=>"010001101",
  19375=>"110000100",
  19376=>"011111010",
  19377=>"110110000",
  19378=>"000010011",
  19379=>"110111111",
  19380=>"110110011",
  19381=>"001101000",
  19382=>"110000011",
  19383=>"001101000",
  19384=>"001010001",
  19385=>"111001111",
  19386=>"111100110",
  19387=>"000111110",
  19388=>"111011001",
  19389=>"100100010",
  19390=>"100110010",
  19391=>"000001011",
  19392=>"110111011",
  19393=>"010111100",
  19394=>"010111101",
  19395=>"000000110",
  19396=>"111001010",
  19397=>"011100101",
  19398=>"011000010",
  19399=>"110110011",
  19400=>"001011101",
  19401=>"001101110",
  19402=>"111111010",
  19403=>"000101000",
  19404=>"101001000",
  19405=>"010100000",
  19406=>"101011111",
  19407=>"001111000",
  19408=>"011010100",
  19409=>"001001100",
  19410=>"111101001",
  19411=>"100001110",
  19412=>"001011111",
  19413=>"111000110",
  19414=>"110111100",
  19415=>"000101111",
  19416=>"000000000",
  19417=>"100000110",
  19418=>"110010110",
  19419=>"100001101",
  19420=>"110110110",
  19421=>"000011111",
  19422=>"111101100",
  19423=>"011011000",
  19424=>"101010010",
  19425=>"000100011",
  19426=>"111100100",
  19427=>"011111010",
  19428=>"100101111",
  19429=>"001111011",
  19430=>"101011100",
  19431=>"010100100",
  19432=>"010010010",
  19433=>"101000000",
  19434=>"110001010",
  19435=>"010101011",
  19436=>"111111101",
  19437=>"001001011",
  19438=>"011001001",
  19439=>"000011100",
  19440=>"110110110",
  19441=>"000101100",
  19442=>"010000111",
  19443=>"010000000",
  19444=>"010110110",
  19445=>"000110110",
  19446=>"110111000",
  19447=>"000010001",
  19448=>"111111111",
  19449=>"111010000",
  19450=>"011110111",
  19451=>"101101000",
  19452=>"001101110",
  19453=>"001000011",
  19454=>"011111100",
  19455=>"111011010",
  19456=>"011000110",
  19457=>"000100101",
  19458=>"100111101",
  19459=>"110111101",
  19460=>"110010011",
  19461=>"011000001",
  19462=>"010101111",
  19463=>"011101111",
  19464=>"111000011",
  19465=>"011010011",
  19466=>"001100111",
  19467=>"110000001",
  19468=>"100010010",
  19469=>"010010110",
  19470=>"011001111",
  19471=>"010110011",
  19472=>"100111111",
  19473=>"110001000",
  19474=>"111111110",
  19475=>"010100000",
  19476=>"100001100",
  19477=>"100101111",
  19478=>"110110011",
  19479=>"110110100",
  19480=>"101111010",
  19481=>"000101001",
  19482=>"000000011",
  19483=>"111111011",
  19484=>"111001011",
  19485=>"011000000",
  19486=>"110000001",
  19487=>"011101011",
  19488=>"001011011",
  19489=>"000110011",
  19490=>"001001100",
  19491=>"101100111",
  19492=>"111101010",
  19493=>"011101101",
  19494=>"101110111",
  19495=>"110011111",
  19496=>"111010111",
  19497=>"000001001",
  19498=>"010100010",
  19499=>"101110000",
  19500=>"110001011",
  19501=>"110101011",
  19502=>"101100010",
  19503=>"100100100",
  19504=>"101100100",
  19505=>"000110100",
  19506=>"111101001",
  19507=>"000011001",
  19508=>"111110001",
  19509=>"101011001",
  19510=>"011111100",
  19511=>"001010010",
  19512=>"011101100",
  19513=>"101001101",
  19514=>"101000111",
  19515=>"010011110",
  19516=>"001000001",
  19517=>"011011101",
  19518=>"101101010",
  19519=>"110000100",
  19520=>"010000101",
  19521=>"101000001",
  19522=>"100000000",
  19523=>"011010010",
  19524=>"011010000",
  19525=>"110011111",
  19526=>"100010110",
  19527=>"100010000",
  19528=>"010001100",
  19529=>"110101100",
  19530=>"110011001",
  19531=>"101100001",
  19532=>"001011111",
  19533=>"000000000",
  19534=>"110110100",
  19535=>"010110101",
  19536=>"010010111",
  19537=>"001111110",
  19538=>"001011101",
  19539=>"101100010",
  19540=>"100010010",
  19541=>"111000100",
  19542=>"100100111",
  19543=>"100100100",
  19544=>"011011011",
  19545=>"111001001",
  19546=>"011110110",
  19547=>"011010000",
  19548=>"001011111",
  19549=>"000011000",
  19550=>"000101011",
  19551=>"101101101",
  19552=>"010000011",
  19553=>"011100110",
  19554=>"100010000",
  19555=>"000100101",
  19556=>"000100101",
  19557=>"111011101",
  19558=>"000110000",
  19559=>"101000100",
  19560=>"001001101",
  19561=>"111001110",
  19562=>"110000101",
  19563=>"100111011",
  19564=>"101000111",
  19565=>"000101000",
  19566=>"101001100",
  19567=>"011100000",
  19568=>"110001101",
  19569=>"100110000",
  19570=>"011100011",
  19571=>"100000110",
  19572=>"000110100",
  19573=>"001100011",
  19574=>"100101101",
  19575=>"110011110",
  19576=>"011011100",
  19577=>"010111010",
  19578=>"101000100",
  19579=>"011110100",
  19580=>"001100100",
  19581=>"111100111",
  19582=>"001000111",
  19583=>"001010100",
  19584=>"011110010",
  19585=>"101000111",
  19586=>"111110011",
  19587=>"000111100",
  19588=>"110101100",
  19589=>"110101010",
  19590=>"000101000",
  19591=>"111100101",
  19592=>"101010001",
  19593=>"001011100",
  19594=>"010000001",
  19595=>"000000000",
  19596=>"010000100",
  19597=>"101100110",
  19598=>"010101011",
  19599=>"001111001",
  19600=>"001111101",
  19601=>"001000100",
  19602=>"001110101",
  19603=>"100010101",
  19604=>"011111000",
  19605=>"110101010",
  19606=>"110100111",
  19607=>"000101111",
  19608=>"110101000",
  19609=>"101011101",
  19610=>"100101100",
  19611=>"101111110",
  19612=>"001001000",
  19613=>"111110111",
  19614=>"011100010",
  19615=>"000110000",
  19616=>"001100110",
  19617=>"011100111",
  19618=>"100110100",
  19619=>"110001001",
  19620=>"111000111",
  19621=>"000111010",
  19622=>"111111011",
  19623=>"101101101",
  19624=>"110001101",
  19625=>"100011110",
  19626=>"001010110",
  19627=>"100000111",
  19628=>"011011011",
  19629=>"010010010",
  19630=>"010110101",
  19631=>"111010111",
  19632=>"000011010",
  19633=>"010001011",
  19634=>"101000100",
  19635=>"100011010",
  19636=>"101001110",
  19637=>"001000011",
  19638=>"101011100",
  19639=>"010001011",
  19640=>"101110100",
  19641=>"110010010",
  19642=>"100001110",
  19643=>"011000000",
  19644=>"001101000",
  19645=>"100001111",
  19646=>"111100101",
  19647=>"100110100",
  19648=>"110011001",
  19649=>"111000001",
  19650=>"011100001",
  19651=>"111111111",
  19652=>"101111000",
  19653=>"000101000",
  19654=>"100110001",
  19655=>"000110110",
  19656=>"010001001",
  19657=>"010010100",
  19658=>"100000100",
  19659=>"100110010",
  19660=>"101100010",
  19661=>"100110000",
  19662=>"001011110",
  19663=>"011110011",
  19664=>"110010111",
  19665=>"101010100",
  19666=>"001101011",
  19667=>"010000011",
  19668=>"110001100",
  19669=>"001000111",
  19670=>"101010111",
  19671=>"111100111",
  19672=>"010110010",
  19673=>"110010100",
  19674=>"111011010",
  19675=>"001100000",
  19676=>"011111000",
  19677=>"110100001",
  19678=>"010111010",
  19679=>"111110010",
  19680=>"010000010",
  19681=>"001010110",
  19682=>"111111101",
  19683=>"010010010",
  19684=>"100100111",
  19685=>"001001010",
  19686=>"111010011",
  19687=>"101011011",
  19688=>"111110000",
  19689=>"010001110",
  19690=>"111001110",
  19691=>"010000100",
  19692=>"011110111",
  19693=>"111100001",
  19694=>"001101100",
  19695=>"000001000",
  19696=>"010100010",
  19697=>"101001010",
  19698=>"100101100",
  19699=>"000100100",
  19700=>"010100101",
  19701=>"000001000",
  19702=>"101010101",
  19703=>"101001000",
  19704=>"111001111",
  19705=>"111010000",
  19706=>"011111000",
  19707=>"000000111",
  19708=>"111000010",
  19709=>"111111000",
  19710=>"010001100",
  19711=>"100111011",
  19712=>"100011111",
  19713=>"101000000",
  19714=>"011011111",
  19715=>"011101001",
  19716=>"011011011",
  19717=>"100010111",
  19718=>"100000000",
  19719=>"011111101",
  19720=>"001111111",
  19721=>"110101000",
  19722=>"101100101",
  19723=>"101000100",
  19724=>"101001100",
  19725=>"111101010",
  19726=>"011000101",
  19727=>"100000001",
  19728=>"100011100",
  19729=>"111000100",
  19730=>"101001001",
  19731=>"100100101",
  19732=>"000100001",
  19733=>"000111101",
  19734=>"010001001",
  19735=>"100111001",
  19736=>"111101111",
  19737=>"011011000",
  19738=>"011101000",
  19739=>"101111101",
  19740=>"111010010",
  19741=>"100101100",
  19742=>"111111111",
  19743=>"000011101",
  19744=>"111000001",
  19745=>"110001101",
  19746=>"100100110",
  19747=>"001000101",
  19748=>"000101110",
  19749=>"101011100",
  19750=>"111001101",
  19751=>"010011010",
  19752=>"001000110",
  19753=>"000100111",
  19754=>"010001101",
  19755=>"000001011",
  19756=>"101110001",
  19757=>"110110000",
  19758=>"010001100",
  19759=>"001010011",
  19760=>"000111010",
  19761=>"111111010",
  19762=>"110001100",
  19763=>"010010010",
  19764=>"001011001",
  19765=>"100001001",
  19766=>"111111111",
  19767=>"111011100",
  19768=>"000101000",
  19769=>"011010001",
  19770=>"010010110",
  19771=>"100111010",
  19772=>"001000000",
  19773=>"010000111",
  19774=>"000001011",
  19775=>"000001000",
  19776=>"100010000",
  19777=>"011000100",
  19778=>"010010100",
  19779=>"111100010",
  19780=>"000100000",
  19781=>"000101111",
  19782=>"101000011",
  19783=>"001101011",
  19784=>"001101011",
  19785=>"010111100",
  19786=>"000010111",
  19787=>"010001100",
  19788=>"000001101",
  19789=>"111101111",
  19790=>"000010101",
  19791=>"101110010",
  19792=>"010110001",
  19793=>"000001110",
  19794=>"011001100",
  19795=>"000011000",
  19796=>"111000000",
  19797=>"110010010",
  19798=>"111001000",
  19799=>"011010010",
  19800=>"001100110",
  19801=>"110010010",
  19802=>"110110100",
  19803=>"010110101",
  19804=>"100000011",
  19805=>"110110001",
  19806=>"110101110",
  19807=>"000001001",
  19808=>"111111000",
  19809=>"110010100",
  19810=>"111011000",
  19811=>"111001010",
  19812=>"101101010",
  19813=>"111001001",
  19814=>"010110110",
  19815=>"111111110",
  19816=>"000011111",
  19817=>"000011100",
  19818=>"001011100",
  19819=>"100000010",
  19820=>"110100110",
  19821=>"110011110",
  19822=>"011111010",
  19823=>"011111111",
  19824=>"001000000",
  19825=>"100011100",
  19826=>"101111100",
  19827=>"110001000",
  19828=>"100101101",
  19829=>"101010111",
  19830=>"100011000",
  19831=>"000001010",
  19832=>"111111111",
  19833=>"110101001",
  19834=>"011010010",
  19835=>"000100111",
  19836=>"000010100",
  19837=>"111011010",
  19838=>"000110000",
  19839=>"011001111",
  19840=>"100010111",
  19841=>"011001000",
  19842=>"101111111",
  19843=>"000001000",
  19844=>"101101011",
  19845=>"111100001",
  19846=>"111100000",
  19847=>"011011000",
  19848=>"101101111",
  19849=>"101010111",
  19850=>"001000011",
  19851=>"010111010",
  19852=>"000010100",
  19853=>"000000110",
  19854=>"111001100",
  19855=>"011111101",
  19856=>"011101101",
  19857=>"110000110",
  19858=>"111110000",
  19859=>"000101100",
  19860=>"010111000",
  19861=>"000011101",
  19862=>"011010010",
  19863=>"101011101",
  19864=>"111001100",
  19865=>"001000010",
  19866=>"000010111",
  19867=>"000000100",
  19868=>"101011001",
  19869=>"010001001",
  19870=>"111100000",
  19871=>"000100000",
  19872=>"001110000",
  19873=>"000010010",
  19874=>"111001100",
  19875=>"101000101",
  19876=>"010000100",
  19877=>"111001100",
  19878=>"110111111",
  19879=>"010011101",
  19880=>"110110110",
  19881=>"111101001",
  19882=>"100100100",
  19883=>"011001101",
  19884=>"000000001",
  19885=>"010111001",
  19886=>"111101000",
  19887=>"001111100",
  19888=>"001001000",
  19889=>"000110011",
  19890=>"001010000",
  19891=>"110001010",
  19892=>"000001011",
  19893=>"101010001",
  19894=>"001011111",
  19895=>"100100011",
  19896=>"101001001",
  19897=>"010101110",
  19898=>"000001100",
  19899=>"000000011",
  19900=>"010010110",
  19901=>"101111111",
  19902=>"101111111",
  19903=>"010000000",
  19904=>"001000001",
  19905=>"100011111",
  19906=>"111000100",
  19907=>"011010010",
  19908=>"010110010",
  19909=>"111101011",
  19910=>"110001001",
  19911=>"010001000",
  19912=>"100100111",
  19913=>"001011011",
  19914=>"011100110",
  19915=>"010001111",
  19916=>"111100011",
  19917=>"111111010",
  19918=>"101100010",
  19919=>"000001110",
  19920=>"101111111",
  19921=>"100110011",
  19922=>"100101111",
  19923=>"100100010",
  19924=>"101001101",
  19925=>"101000110",
  19926=>"111000111",
  19927=>"101010100",
  19928=>"110001011",
  19929=>"011110010",
  19930=>"101001001",
  19931=>"000111100",
  19932=>"110010111",
  19933=>"101101100",
  19934=>"010011001",
  19935=>"000111110",
  19936=>"101110010",
  19937=>"000010100",
  19938=>"111011000",
  19939=>"011111111",
  19940=>"111111001",
  19941=>"101111000",
  19942=>"000011100",
  19943=>"111101000",
  19944=>"001001010",
  19945=>"101100100",
  19946=>"100000010",
  19947=>"100001101",
  19948=>"011100010",
  19949=>"011101010",
  19950=>"100000110",
  19951=>"011000010",
  19952=>"000001001",
  19953=>"011011111",
  19954=>"100010010",
  19955=>"000100100",
  19956=>"011011110",
  19957=>"111011101",
  19958=>"001011001",
  19959=>"010110101",
  19960=>"001010000",
  19961=>"010100001",
  19962=>"000110010",
  19963=>"000010100",
  19964=>"100100100",
  19965=>"001100001",
  19966=>"011010011",
  19967=>"111001000",
  19968=>"100011101",
  19969=>"000101111",
  19970=>"111000001",
  19971=>"110011000",
  19972=>"000000101",
  19973=>"011101010",
  19974=>"110110010",
  19975=>"110000010",
  19976=>"101100001",
  19977=>"000110111",
  19978=>"010010111",
  19979=>"000001010",
  19980=>"000000111",
  19981=>"010010100",
  19982=>"111011101",
  19983=>"111001110",
  19984=>"110111001",
  19985=>"010000010",
  19986=>"011001111",
  19987=>"101010000",
  19988=>"110001100",
  19989=>"110101101",
  19990=>"111110010",
  19991=>"111000010",
  19992=>"001101001",
  19993=>"110011000",
  19994=>"001000101",
  19995=>"011001010",
  19996=>"110011100",
  19997=>"110111000",
  19998=>"100101000",
  19999=>"011001111",
  20000=>"111101001",
  20001=>"011001001",
  20002=>"000111100",
  20003=>"010001010",
  20004=>"101001001",
  20005=>"110000110",
  20006=>"100100101",
  20007=>"111011011",
  20008=>"010110000",
  20009=>"000000101",
  20010=>"100111010",
  20011=>"100100101",
  20012=>"100001011",
  20013=>"101001011",
  20014=>"010111100",
  20015=>"100101011",
  20016=>"111001010",
  20017=>"111101111",
  20018=>"101100000",
  20019=>"100100001",
  20020=>"011000011",
  20021=>"110011011",
  20022=>"010101001",
  20023=>"100101011",
  20024=>"111011100",
  20025=>"001001011",
  20026=>"100011010",
  20027=>"010011101",
  20028=>"010101101",
  20029=>"010001010",
  20030=>"101101000",
  20031=>"100110110",
  20032=>"001000111",
  20033=>"010000001",
  20034=>"101000101",
  20035=>"110001100",
  20036=>"111000111",
  20037=>"000101101",
  20038=>"011100011",
  20039=>"001101000",
  20040=>"100100100",
  20041=>"000000001",
  20042=>"111001010",
  20043=>"001101100",
  20044=>"011001101",
  20045=>"001001111",
  20046=>"111110011",
  20047=>"001101011",
  20048=>"110111111",
  20049=>"010001010",
  20050=>"101011100",
  20051=>"001000100",
  20052=>"010001111",
  20053=>"001110001",
  20054=>"111000100",
  20055=>"011001001",
  20056=>"000010100",
  20057=>"001101010",
  20058=>"110011100",
  20059=>"011101101",
  20060=>"100101101",
  20061=>"100101001",
  20062=>"000010110",
  20063=>"111000011",
  20064=>"101100001",
  20065=>"100001110",
  20066=>"101011101",
  20067=>"100001110",
  20068=>"011110111",
  20069=>"100101101",
  20070=>"010111010",
  20071=>"011011001",
  20072=>"000001001",
  20073=>"111001101",
  20074=>"000001011",
  20075=>"000000101",
  20076=>"010011110",
  20077=>"100010000",
  20078=>"110110111",
  20079=>"000110011",
  20080=>"011010010",
  20081=>"110011001",
  20082=>"011100110",
  20083=>"000111111",
  20084=>"000001101",
  20085=>"101001001",
  20086=>"001000001",
  20087=>"001101010",
  20088=>"100011000",
  20089=>"000111110",
  20090=>"111111011",
  20091=>"010011100",
  20092=>"011011010",
  20093=>"100101011",
  20094=>"100111011",
  20095=>"111001011",
  20096=>"111011011",
  20097=>"011110111",
  20098=>"011011001",
  20099=>"100001100",
  20100=>"101111100",
  20101=>"111001100",
  20102=>"010111111",
  20103=>"001101110",
  20104=>"000101100",
  20105=>"001110111",
  20106=>"000111110",
  20107=>"000011011",
  20108=>"100100011",
  20109=>"111101001",
  20110=>"011010001",
  20111=>"100000001",
  20112=>"101111001",
  20113=>"011111011",
  20114=>"101000111",
  20115=>"100100011",
  20116=>"000101100",
  20117=>"110101011",
  20118=>"111001010",
  20119=>"100100100",
  20120=>"100111000",
  20121=>"110111110",
  20122=>"001001010",
  20123=>"100111010",
  20124=>"101001010",
  20125=>"000011011",
  20126=>"000011010",
  20127=>"110010010",
  20128=>"100101010",
  20129=>"110110100",
  20130=>"010111101",
  20131=>"001011010",
  20132=>"110010001",
  20133=>"000010111",
  20134=>"111011111",
  20135=>"101100000",
  20136=>"000001101",
  20137=>"101000000",
  20138=>"100000111",
  20139=>"011010101",
  20140=>"110010101",
  20141=>"000000001",
  20142=>"010011101",
  20143=>"010110011",
  20144=>"011010000",
  20145=>"000110001",
  20146=>"100101100",
  20147=>"011110100",
  20148=>"100001111",
  20149=>"001011010",
  20150=>"111010110",
  20151=>"110100000",
  20152=>"100000000",
  20153=>"100001110",
  20154=>"100001000",
  20155=>"101001010",
  20156=>"111010011",
  20157=>"011110111",
  20158=>"001010010",
  20159=>"100001111",
  20160=>"001100010",
  20161=>"110000010",
  20162=>"110011010",
  20163=>"111110010",
  20164=>"100101111",
  20165=>"001010111",
  20166=>"110111111",
  20167=>"011000100",
  20168=>"110110000",
  20169=>"011101011",
  20170=>"100101010",
  20171=>"010110101",
  20172=>"000010011",
  20173=>"111111101",
  20174=>"111110010",
  20175=>"010011001",
  20176=>"101000111",
  20177=>"010101100",
  20178=>"000001000",
  20179=>"010101011",
  20180=>"100101101",
  20181=>"011100100",
  20182=>"111000111",
  20183=>"000000111",
  20184=>"011011011",
  20185=>"111111111",
  20186=>"111001010",
  20187=>"110001111",
  20188=>"011100101",
  20189=>"000001100",
  20190=>"101000000",
  20191=>"101011110",
  20192=>"000100101",
  20193=>"101101101",
  20194=>"000101110",
  20195=>"000011101",
  20196=>"111000110",
  20197=>"100111001",
  20198=>"110001010",
  20199=>"100000001",
  20200=>"010110011",
  20201=>"110011010",
  20202=>"001101000",
  20203=>"010100010",
  20204=>"101011010",
  20205=>"000111001",
  20206=>"101011111",
  20207=>"001111101",
  20208=>"110101010",
  20209=>"101000111",
  20210=>"110001001",
  20211=>"111000101",
  20212=>"100000001",
  20213=>"101010111",
  20214=>"001000001",
  20215=>"100001111",
  20216=>"011001110",
  20217=>"001011111",
  20218=>"010001011",
  20219=>"110000001",
  20220=>"000111010",
  20221=>"110101100",
  20222=>"010000010",
  20223=>"101100001",
  20224=>"111011001",
  20225=>"111110011",
  20226=>"000101110",
  20227=>"110101110",
  20228=>"000110001",
  20229=>"100011001",
  20230=>"000111010",
  20231=>"100010011",
  20232=>"100101010",
  20233=>"001001101",
  20234=>"101000010",
  20235=>"101011101",
  20236=>"101100101",
  20237=>"100111011",
  20238=>"111111000",
  20239=>"011010110",
  20240=>"001111100",
  20241=>"001011011",
  20242=>"000110011",
  20243=>"110110011",
  20244=>"001010010",
  20245=>"001011100",
  20246=>"000111111",
  20247=>"100000001",
  20248=>"111100101",
  20249=>"001100000",
  20250=>"000101111",
  20251=>"000010010",
  20252=>"000111000",
  20253=>"110110011",
  20254=>"000010000",
  20255=>"111011001",
  20256=>"110111001",
  20257=>"110010010",
  20258=>"101111100",
  20259=>"101010001",
  20260=>"010001101",
  20261=>"010111000",
  20262=>"010101011",
  20263=>"110110010",
  20264=>"101101100",
  20265=>"111110001",
  20266=>"010110010",
  20267=>"010111100",
  20268=>"010001000",
  20269=>"000010101",
  20270=>"100110001",
  20271=>"101001000",
  20272=>"000101011",
  20273=>"000011001",
  20274=>"010010010",
  20275=>"001010111",
  20276=>"101011000",
  20277=>"001010000",
  20278=>"000010100",
  20279=>"011101011",
  20280=>"001110001",
  20281=>"100011010",
  20282=>"011010001",
  20283=>"011110100",
  20284=>"110000110",
  20285=>"000101000",
  20286=>"010000010",
  20287=>"011111100",
  20288=>"011000101",
  20289=>"111001011",
  20290=>"111010001",
  20291=>"101001110",
  20292=>"001110100",
  20293=>"101010000",
  20294=>"101000000",
  20295=>"000101011",
  20296=>"001001001",
  20297=>"110000001",
  20298=>"001111100",
  20299=>"001010100",
  20300=>"111100110",
  20301=>"101010100",
  20302=>"101000110",
  20303=>"010010100",
  20304=>"000010010",
  20305=>"011001011",
  20306=>"111110100",
  20307=>"101000100",
  20308=>"011111100",
  20309=>"101011100",
  20310=>"000000010",
  20311=>"000011000",
  20312=>"111010110",
  20313=>"111110100",
  20314=>"001110011",
  20315=>"100000001",
  20316=>"101101101",
  20317=>"111100111",
  20318=>"101100100",
  20319=>"100010111",
  20320=>"101111100",
  20321=>"101101111",
  20322=>"000111000",
  20323=>"100100010",
  20324=>"001011001",
  20325=>"101111010",
  20326=>"110000010",
  20327=>"100010100",
  20328=>"101111111",
  20329=>"111011011",
  20330=>"101100001",
  20331=>"011011000",
  20332=>"011010000",
  20333=>"010100101",
  20334=>"101011100",
  20335=>"100000111",
  20336=>"000101100",
  20337=>"011100011",
  20338=>"011001110",
  20339=>"111001011",
  20340=>"000110000",
  20341=>"011001111",
  20342=>"100100111",
  20343=>"110101001",
  20344=>"000010000",
  20345=>"001011011",
  20346=>"000110001",
  20347=>"111000000",
  20348=>"010101010",
  20349=>"000001101",
  20350=>"000100110",
  20351=>"111100011",
  20352=>"101011001",
  20353=>"011110011",
  20354=>"000111110",
  20355=>"110110110",
  20356=>"100010011",
  20357=>"010100010",
  20358=>"001101010",
  20359=>"010010111",
  20360=>"110101101",
  20361=>"001011101",
  20362=>"001110100",
  20363=>"011111000",
  20364=>"000001100",
  20365=>"101010001",
  20366=>"100100101",
  20367=>"101111110",
  20368=>"010100010",
  20369=>"101010010",
  20370=>"010001000",
  20371=>"011000101",
  20372=>"111101111",
  20373=>"100010111",
  20374=>"001001101",
  20375=>"100111010",
  20376=>"001101000",
  20377=>"000100000",
  20378=>"001000111",
  20379=>"000000001",
  20380=>"100000101",
  20381=>"000111101",
  20382=>"101011100",
  20383=>"000001010",
  20384=>"100101000",
  20385=>"111111101",
  20386=>"010011100",
  20387=>"001000111",
  20388=>"011101100",
  20389=>"110111101",
  20390=>"001101111",
  20391=>"100110101",
  20392=>"000011100",
  20393=>"101101100",
  20394=>"001100111",
  20395=>"100110001",
  20396=>"110010100",
  20397=>"101101101",
  20398=>"110110101",
  20399=>"001001000",
  20400=>"111111000",
  20401=>"110011100",
  20402=>"001100111",
  20403=>"111011010",
  20404=>"110110100",
  20405=>"111011110",
  20406=>"010100011",
  20407=>"110100001",
  20408=>"000101101",
  20409=>"000001110",
  20410=>"001110011",
  20411=>"011000010",
  20412=>"010110111",
  20413=>"111111000",
  20414=>"100010010",
  20415=>"101100110",
  20416=>"101010110",
  20417=>"010111111",
  20418=>"110101111",
  20419=>"010101001",
  20420=>"100000011",
  20421=>"010110111",
  20422=>"110010101",
  20423=>"111111100",
  20424=>"001111001",
  20425=>"000010111",
  20426=>"110100000",
  20427=>"000101100",
  20428=>"000110000",
  20429=>"000001110",
  20430=>"100010101",
  20431=>"011101011",
  20432=>"100110110",
  20433=>"111111110",
  20434=>"011100010",
  20435=>"010001000",
  20436=>"100011100",
  20437=>"000110000",
  20438=>"011111100",
  20439=>"101111100",
  20440=>"101000011",
  20441=>"110101111",
  20442=>"110100111",
  20443=>"000000001",
  20444=>"011101111",
  20445=>"111010000",
  20446=>"110001101",
  20447=>"001110010",
  20448=>"010000110",
  20449=>"001111001",
  20450=>"110001101",
  20451=>"011110111",
  20452=>"011001000",
  20453=>"000100000",
  20454=>"100111001",
  20455=>"111001011",
  20456=>"000000000",
  20457=>"101100111",
  20458=>"101000111",
  20459=>"000000000",
  20460=>"110101111",
  20461=>"110010101",
  20462=>"010101001",
  20463=>"000000100",
  20464=>"000101111",
  20465=>"011011111",
  20466=>"010001011",
  20467=>"000101100",
  20468=>"011000100",
  20469=>"000011011",
  20470=>"001011001",
  20471=>"001011010",
  20472=>"011100111",
  20473=>"101011111",
  20474=>"000000000",
  20475=>"010011010",
  20476=>"001001010",
  20477=>"010000101",
  20478=>"000011101",
  20479=>"010000011",
  20480=>"011110111",
  20481=>"001010111",
  20482=>"000111000",
  20483=>"011010110",
  20484=>"011000001",
  20485=>"011001101",
  20486=>"000111001",
  20487=>"100000100",
  20488=>"011110001",
  20489=>"000000000",
  20490=>"101101100",
  20491=>"001001100",
  20492=>"000011010",
  20493=>"000110000",
  20494=>"101101111",
  20495=>"101000100",
  20496=>"000110010",
  20497=>"000111000",
  20498=>"111111010",
  20499=>"111111011",
  20500=>"000010110",
  20501=>"010010101",
  20502=>"111000000",
  20503=>"010010101",
  20504=>"000001100",
  20505=>"101100101",
  20506=>"110000011",
  20507=>"001001111",
  20508=>"100110000",
  20509=>"111110011",
  20510=>"000000011",
  20511=>"100110110",
  20512=>"111001010",
  20513=>"100011111",
  20514=>"111000111",
  20515=>"001000110",
  20516=>"011100001",
  20517=>"011010001",
  20518=>"001000000",
  20519=>"110111001",
  20520=>"101111011",
  20521=>"011101000",
  20522=>"010100011",
  20523=>"111001011",
  20524=>"000100100",
  20525=>"110111111",
  20526=>"010110001",
  20527=>"011011011",
  20528=>"100011011",
  20529=>"010110011",
  20530=>"111000000",
  20531=>"110101101",
  20532=>"111110001",
  20533=>"010110100",
  20534=>"010000100",
  20535=>"111000000",
  20536=>"000000100",
  20537=>"100011100",
  20538=>"110000001",
  20539=>"101110011",
  20540=>"100001000",
  20541=>"000110101",
  20542=>"011110100",
  20543=>"100100100",
  20544=>"011001011",
  20545=>"110001001",
  20546=>"010111001",
  20547=>"010001100",
  20548=>"100011000",
  20549=>"100111111",
  20550=>"001011010",
  20551=>"000111101",
  20552=>"001000000",
  20553=>"110001010",
  20554=>"001010100",
  20555=>"110001001",
  20556=>"111011110",
  20557=>"001010011",
  20558=>"111001110",
  20559=>"000000000",
  20560=>"100000011",
  20561=>"000101111",
  20562=>"110110011",
  20563=>"101111000",
  20564=>"001000000",
  20565=>"000001101",
  20566=>"011011011",
  20567=>"001001000",
  20568=>"010010101",
  20569=>"001001010",
  20570=>"101100010",
  20571=>"111000010",
  20572=>"000101000",
  20573=>"010000001",
  20574=>"000110111",
  20575=>"010000010",
  20576=>"111011000",
  20577=>"001010101",
  20578=>"010100010",
  20579=>"000011000",
  20580=>"101011101",
  20581=>"010111000",
  20582=>"110010000",
  20583=>"000000000",
  20584=>"010110111",
  20585=>"100111001",
  20586=>"000000110",
  20587=>"100000111",
  20588=>"111001101",
  20589=>"001110101",
  20590=>"110101001",
  20591=>"011000101",
  20592=>"110100110",
  20593=>"101000010",
  20594=>"010011010",
  20595=>"110000001",
  20596=>"111010100",
  20597=>"000010100",
  20598=>"100111100",
  20599=>"000101100",
  20600=>"101001010",
  20601=>"100101100",
  20602=>"110011111",
  20603=>"001100000",
  20604=>"101000010",
  20605=>"111000000",
  20606=>"011100111",
  20607=>"100111101",
  20608=>"101101101",
  20609=>"110011101",
  20610=>"001001111",
  20611=>"001000100",
  20612=>"001101100",
  20613=>"101111011",
  20614=>"001110100",
  20615=>"000100101",
  20616=>"000011100",
  20617=>"100101000",
  20618=>"001001000",
  20619=>"111011111",
  20620=>"110011011",
  20621=>"101000011",
  20622=>"001110101",
  20623=>"011011011",
  20624=>"110010001",
  20625=>"011111110",
  20626=>"100100111",
  20627=>"010010000",
  20628=>"100111011",
  20629=>"100110010",
  20630=>"001010010",
  20631=>"100101010",
  20632=>"010000000",
  20633=>"011001000",
  20634=>"001001101",
  20635=>"100011010",
  20636=>"001000000",
  20637=>"101001011",
  20638=>"111110111",
  20639=>"100001111",
  20640=>"101001110",
  20641=>"110010001",
  20642=>"001001100",
  20643=>"000000100",
  20644=>"001011000",
  20645=>"010001111",
  20646=>"001101101",
  20647=>"110100100",
  20648=>"011000101",
  20649=>"010000011",
  20650=>"001111011",
  20651=>"000111110",
  20652=>"100111100",
  20653=>"011101111",
  20654=>"010001100",
  20655=>"011011001",
  20656=>"011010001",
  20657=>"010101011",
  20658=>"110001010",
  20659=>"100010000",
  20660=>"101011101",
  20661=>"000000011",
  20662=>"110100001",
  20663=>"110101010",
  20664=>"000001000",
  20665=>"101000000",
  20666=>"101010111",
  20667=>"000101101",
  20668=>"110101111",
  20669=>"101011101",
  20670=>"001001111",
  20671=>"010000000",
  20672=>"001110000",
  20673=>"001001111",
  20674=>"000010010",
  20675=>"101001011",
  20676=>"001111010",
  20677=>"001111000",
  20678=>"011110110",
  20679=>"001000001",
  20680=>"000011011",
  20681=>"001111111",
  20682=>"101101110",
  20683=>"100001101",
  20684=>"110010000",
  20685=>"011101101",
  20686=>"000001110",
  20687=>"001111011",
  20688=>"011111011",
  20689=>"001111011",
  20690=>"000101000",
  20691=>"001111111",
  20692=>"011011100",
  20693=>"000000111",
  20694=>"101101110",
  20695=>"001001101",
  20696=>"110000011",
  20697=>"001101001",
  20698=>"000000000",
  20699=>"000000101",
  20700=>"000011100",
  20701=>"000001011",
  20702=>"011001001",
  20703=>"011111000",
  20704=>"110111110",
  20705=>"111101101",
  20706=>"110011011",
  20707=>"011011110",
  20708=>"100100010",
  20709=>"110101111",
  20710=>"100000010",
  20711=>"011000010",
  20712=>"011110000",
  20713=>"110100000",
  20714=>"011000100",
  20715=>"011001011",
  20716=>"110111011",
  20717=>"100000110",
  20718=>"000000000",
  20719=>"010100101",
  20720=>"111111011",
  20721=>"001001010",
  20722=>"000110110",
  20723=>"110101011",
  20724=>"101100010",
  20725=>"010000110",
  20726=>"010011101",
  20727=>"000001000",
  20728=>"001111101",
  20729=>"000100011",
  20730=>"100111101",
  20731=>"000010000",
  20732=>"100001101",
  20733=>"100101101",
  20734=>"000011001",
  20735=>"010110001",
  20736=>"110111010",
  20737=>"101111111",
  20738=>"111001010",
  20739=>"110101001",
  20740=>"100001110",
  20741=>"001010011",
  20742=>"111110111",
  20743=>"110100010",
  20744=>"110000100",
  20745=>"110000110",
  20746=>"011000001",
  20747=>"010111111",
  20748=>"010001111",
  20749=>"100000111",
  20750=>"000111000",
  20751=>"010000111",
  20752=>"010110011",
  20753=>"001110000",
  20754=>"101011111",
  20755=>"101001111",
  20756=>"111001011",
  20757=>"010010111",
  20758=>"000000000",
  20759=>"011100110",
  20760=>"111001011",
  20761=>"100001010",
  20762=>"011010101",
  20763=>"001000010",
  20764=>"001111011",
  20765=>"101110010",
  20766=>"111111101",
  20767=>"111001010",
  20768=>"100100000",
  20769=>"111111011",
  20770=>"001000110",
  20771=>"010100101",
  20772=>"110001101",
  20773=>"111010010",
  20774=>"110111100",
  20775=>"011011110",
  20776=>"111100010",
  20777=>"010101111",
  20778=>"101011100",
  20779=>"110111000",
  20780=>"101111111",
  20781=>"111011100",
  20782=>"000000101",
  20783=>"111100100",
  20784=>"101010111",
  20785=>"011001110",
  20786=>"111001000",
  20787=>"000110001",
  20788=>"111010100",
  20789=>"111011001",
  20790=>"110100100",
  20791=>"011110011",
  20792=>"010000010",
  20793=>"110101100",
  20794=>"000100101",
  20795=>"001110001",
  20796=>"010010101",
  20797=>"101111000",
  20798=>"100010110",
  20799=>"111000100",
  20800=>"111011111",
  20801=>"111100100",
  20802=>"011111111",
  20803=>"101111000",
  20804=>"011111101",
  20805=>"000011011",
  20806=>"000001011",
  20807=>"001111000",
  20808=>"011010001",
  20809=>"000101011",
  20810=>"101100010",
  20811=>"101010110",
  20812=>"111100110",
  20813=>"010010001",
  20814=>"111110011",
  20815=>"010000100",
  20816=>"110010001",
  20817=>"101010001",
  20818=>"011010101",
  20819=>"101010110",
  20820=>"100100000",
  20821=>"011010110",
  20822=>"000100110",
  20823=>"100000011",
  20824=>"111000000",
  20825=>"010000111",
  20826=>"000001101",
  20827=>"111010001",
  20828=>"101011011",
  20829=>"111001010",
  20830=>"101100011",
  20831=>"001101101",
  20832=>"000101010",
  20833=>"010010101",
  20834=>"110111011",
  20835=>"001000100",
  20836=>"100100111",
  20837=>"000100000",
  20838=>"110000110",
  20839=>"110000101",
  20840=>"001110000",
  20841=>"000000100",
  20842=>"000111100",
  20843=>"000001000",
  20844=>"001110101",
  20845=>"110010010",
  20846=>"010000001",
  20847=>"101010011",
  20848=>"000000010",
  20849=>"011001110",
  20850=>"011110101",
  20851=>"100101100",
  20852=>"011011000",
  20853=>"111011111",
  20854=>"111011101",
  20855=>"000100101",
  20856=>"110001100",
  20857=>"100010000",
  20858=>"111111010",
  20859=>"001000011",
  20860=>"100011010",
  20861=>"101101110",
  20862=>"001000001",
  20863=>"001001100",
  20864=>"000011011",
  20865=>"101001011",
  20866=>"000111011",
  20867=>"010100010",
  20868=>"010010101",
  20869=>"101011111",
  20870=>"011101011",
  20871=>"111100100",
  20872=>"001010101",
  20873=>"110110110",
  20874=>"001011101",
  20875=>"000110010",
  20876=>"111011100",
  20877=>"110000000",
  20878=>"011000110",
  20879=>"010110101",
  20880=>"011001110",
  20881=>"101010111",
  20882=>"001000101",
  20883=>"011101101",
  20884=>"111111010",
  20885=>"111010101",
  20886=>"101111111",
  20887=>"000000110",
  20888=>"000111101",
  20889=>"100001000",
  20890=>"010101001",
  20891=>"001111111",
  20892=>"100000001",
  20893=>"011011110",
  20894=>"011001110",
  20895=>"111100110",
  20896=>"011000000",
  20897=>"001010101",
  20898=>"011111011",
  20899=>"111101100",
  20900=>"111011110",
  20901=>"000000010",
  20902=>"110101001",
  20903=>"010011110",
  20904=>"001010101",
  20905=>"111000010",
  20906=>"000110010",
  20907=>"111110100",
  20908=>"010110001",
  20909=>"010111010",
  20910=>"110100001",
  20911=>"101101001",
  20912=>"001111000",
  20913=>"101010001",
  20914=>"010100100",
  20915=>"001011111",
  20916=>"101100100",
  20917=>"110100111",
  20918=>"101010110",
  20919=>"010000100",
  20920=>"101000000",
  20921=>"110001010",
  20922=>"010101100",
  20923=>"100101100",
  20924=>"010111010",
  20925=>"100011010",
  20926=>"011011110",
  20927=>"100100101",
  20928=>"101001000",
  20929=>"000100000",
  20930=>"011010011",
  20931=>"010111011",
  20932=>"011100101",
  20933=>"000110110",
  20934=>"001011110",
  20935=>"001101101",
  20936=>"101000000",
  20937=>"001000011",
  20938=>"100100001",
  20939=>"011000000",
  20940=>"011100110",
  20941=>"100001100",
  20942=>"010111111",
  20943=>"110000111",
  20944=>"101011000",
  20945=>"100001000",
  20946=>"110110101",
  20947=>"010111110",
  20948=>"001101101",
  20949=>"111111001",
  20950=>"011101101",
  20951=>"010111000",
  20952=>"011000101",
  20953=>"110110000",
  20954=>"100010101",
  20955=>"011010011",
  20956=>"011110000",
  20957=>"011001110",
  20958=>"111100110",
  20959=>"010110110",
  20960=>"010010101",
  20961=>"010001001",
  20962=>"001100000",
  20963=>"001000100",
  20964=>"101100111",
  20965=>"100110011",
  20966=>"110100110",
  20967=>"001001000",
  20968=>"010000001",
  20969=>"110111111",
  20970=>"100100110",
  20971=>"011001110",
  20972=>"100100000",
  20973=>"001111011",
  20974=>"000010011",
  20975=>"010000101",
  20976=>"000001000",
  20977=>"110000001",
  20978=>"111010101",
  20979=>"010000111",
  20980=>"110001010",
  20981=>"000110100",
  20982=>"100111101",
  20983=>"100111110",
  20984=>"010110011",
  20985=>"101101111",
  20986=>"101111111",
  20987=>"100111100",
  20988=>"100111111",
  20989=>"100000010",
  20990=>"011101101",
  20991=>"101110010",
  20992=>"100110100",
  20993=>"000001010",
  20994=>"010100100",
  20995=>"101010000",
  20996=>"110011001",
  20997=>"001001101",
  20998=>"111010011",
  20999=>"000010010",
  21000=>"100100011",
  21001=>"101000000",
  21002=>"000110101",
  21003=>"101001100",
  21004=>"011110100",
  21005=>"011110111",
  21006=>"101100111",
  21007=>"110110001",
  21008=>"000101011",
  21009=>"001000001",
  21010=>"110101111",
  21011=>"000010001",
  21012=>"011100011",
  21013=>"100000111",
  21014=>"110011110",
  21015=>"100100000",
  21016=>"110100010",
  21017=>"000111111",
  21018=>"001011000",
  21019=>"110000000",
  21020=>"110111110",
  21021=>"111111001",
  21022=>"111100000",
  21023=>"010101001",
  21024=>"001010000",
  21025=>"010000100",
  21026=>"000011110",
  21027=>"000000100",
  21028=>"011000100",
  21029=>"100011101",
  21030=>"100110101",
  21031=>"110101010",
  21032=>"010100000",
  21033=>"011100001",
  21034=>"101001011",
  21035=>"001100101",
  21036=>"001000001",
  21037=>"011101100",
  21038=>"010000110",
  21039=>"111111000",
  21040=>"101000000",
  21041=>"011101101",
  21042=>"101000010",
  21043=>"100011101",
  21044=>"101010111",
  21045=>"111010000",
  21046=>"100100000",
  21047=>"100100101",
  21048=>"101110011",
  21049=>"111011110",
  21050=>"110111001",
  21051=>"010011101",
  21052=>"100100111",
  21053=>"001010111",
  21054=>"010000101",
  21055=>"000001010",
  21056=>"001001111",
  21057=>"101101010",
  21058=>"011000000",
  21059=>"000110101",
  21060=>"110101101",
  21061=>"111110100",
  21062=>"111100101",
  21063=>"000101010",
  21064=>"111100010",
  21065=>"001011011",
  21066=>"010011011",
  21067=>"111110110",
  21068=>"010101010",
  21069=>"100101001",
  21070=>"100000010",
  21071=>"010101100",
  21072=>"010010000",
  21073=>"010011100",
  21074=>"000100111",
  21075=>"111100000",
  21076=>"111111110",
  21077=>"111110110",
  21078=>"100000000",
  21079=>"101111010",
  21080=>"000000000",
  21081=>"111000110",
  21082=>"110101110",
  21083=>"011111011",
  21084=>"000011001",
  21085=>"100110110",
  21086=>"000011011",
  21087=>"111000111",
  21088=>"101110000",
  21089=>"001000000",
  21090=>"001001110",
  21091=>"101100101",
  21092=>"000010010",
  21093=>"001110111",
  21094=>"000001000",
  21095=>"010000110",
  21096=>"011001010",
  21097=>"101011011",
  21098=>"000010111",
  21099=>"101000110",
  21100=>"101110011",
  21101=>"101101010",
  21102=>"000010111",
  21103=>"100011011",
  21104=>"010111010",
  21105=>"000110000",
  21106=>"111011111",
  21107=>"000100000",
  21108=>"100000001",
  21109=>"110100001",
  21110=>"101111010",
  21111=>"010111111",
  21112=>"110111001",
  21113=>"000000001",
  21114=>"000010111",
  21115=>"001001100",
  21116=>"111111010",
  21117=>"010011100",
  21118=>"111101110",
  21119=>"001010101",
  21120=>"101011000",
  21121=>"111000001",
  21122=>"101111000",
  21123=>"100111011",
  21124=>"100000100",
  21125=>"101100011",
  21126=>"001111101",
  21127=>"010011001",
  21128=>"011010110",
  21129=>"110111000",
  21130=>"011101111",
  21131=>"111111001",
  21132=>"000101111",
  21133=>"001111110",
  21134=>"011111101",
  21135=>"010000010",
  21136=>"011111000",
  21137=>"001101011",
  21138=>"010101111",
  21139=>"011110000",
  21140=>"100011001",
  21141=>"111111111",
  21142=>"011010110",
  21143=>"001011100",
  21144=>"101000011",
  21145=>"111100000",
  21146=>"000110010",
  21147=>"010111001",
  21148=>"001010110",
  21149=>"011010111",
  21150=>"111111111",
  21151=>"001111111",
  21152=>"100001111",
  21153=>"100111001",
  21154=>"101100001",
  21155=>"010011010",
  21156=>"001001001",
  21157=>"000100111",
  21158=>"001011010",
  21159=>"100011110",
  21160=>"000001001",
  21161=>"001101100",
  21162=>"101011011",
  21163=>"000011110",
  21164=>"000001110",
  21165=>"111001100",
  21166=>"000010000",
  21167=>"010010101",
  21168=>"001011101",
  21169=>"110111011",
  21170=>"010000100",
  21171=>"010010100",
  21172=>"101111110",
  21173=>"000000110",
  21174=>"111010000",
  21175=>"100010100",
  21176=>"001010100",
  21177=>"010001011",
  21178=>"101110011",
  21179=>"000100010",
  21180=>"000101100",
  21181=>"000010001",
  21182=>"000000000",
  21183=>"100101000",
  21184=>"000110110",
  21185=>"100100000",
  21186=>"001101001",
  21187=>"101110001",
  21188=>"011001110",
  21189=>"101101100",
  21190=>"100001001",
  21191=>"101100011",
  21192=>"011011000",
  21193=>"001101010",
  21194=>"010110111",
  21195=>"110100101",
  21196=>"011100010",
  21197=>"011010011",
  21198=>"101011111",
  21199=>"101001101",
  21200=>"111110100",
  21201=>"010010110",
  21202=>"011011100",
  21203=>"100001001",
  21204=>"011101110",
  21205=>"000011100",
  21206=>"101100010",
  21207=>"010100101",
  21208=>"001001000",
  21209=>"000101101",
  21210=>"100011001",
  21211=>"001100010",
  21212=>"001011000",
  21213=>"100101100",
  21214=>"001010000",
  21215=>"010000000",
  21216=>"011001011",
  21217=>"001110100",
  21218=>"111011100",
  21219=>"001000000",
  21220=>"101111011",
  21221=>"101110101",
  21222=>"000101101",
  21223=>"010001110",
  21224=>"011101001",
  21225=>"010000000",
  21226=>"101110000",
  21227=>"000111100",
  21228=>"010000100",
  21229=>"100000111",
  21230=>"101010101",
  21231=>"001101111",
  21232=>"111000100",
  21233=>"110010011",
  21234=>"100110101",
  21235=>"001100000",
  21236=>"100100011",
  21237=>"001000111",
  21238=>"100000000",
  21239=>"011100100",
  21240=>"000110011",
  21241=>"011000011",
  21242=>"101111010",
  21243=>"010101110",
  21244=>"100011001",
  21245=>"001101100",
  21246=>"000010110",
  21247=>"001101010",
  21248=>"100101001",
  21249=>"001010101",
  21250=>"010101101",
  21251=>"101011010",
  21252=>"001100001",
  21253=>"111001110",
  21254=>"010000110",
  21255=>"111111110",
  21256=>"100110000",
  21257=>"000000010",
  21258=>"011111011",
  21259=>"000010010",
  21260=>"010101110",
  21261=>"010001111",
  21262=>"010110110",
  21263=>"011011100",
  21264=>"001000110",
  21265=>"001101011",
  21266=>"110111101",
  21267=>"010000101",
  21268=>"011000010",
  21269=>"110000100",
  21270=>"100110000",
  21271=>"000000000",
  21272=>"011010011",
  21273=>"001001010",
  21274=>"111111011",
  21275=>"010101010",
  21276=>"011010110",
  21277=>"000000111",
  21278=>"010000010",
  21279=>"010001101",
  21280=>"000100101",
  21281=>"001110000",
  21282=>"000010010",
  21283=>"011101011",
  21284=>"000011110",
  21285=>"010011110",
  21286=>"100000110",
  21287=>"011010110",
  21288=>"101001110",
  21289=>"010100110",
  21290=>"110100101",
  21291=>"010011010",
  21292=>"111011010",
  21293=>"011111110",
  21294=>"101100110",
  21295=>"010111111",
  21296=>"011011100",
  21297=>"011110000",
  21298=>"000111100",
  21299=>"101000101",
  21300=>"100010010",
  21301=>"010101100",
  21302=>"101110000",
  21303=>"001010110",
  21304=>"110101010",
  21305=>"100010000",
  21306=>"000010000",
  21307=>"110110000",
  21308=>"001010000",
  21309=>"100000111",
  21310=>"000101000",
  21311=>"000101110",
  21312=>"111111010",
  21313=>"000011001",
  21314=>"000100011",
  21315=>"100100001",
  21316=>"111101111",
  21317=>"100111101",
  21318=>"110111101",
  21319=>"100011011",
  21320=>"110100111",
  21321=>"000001110",
  21322=>"000000001",
  21323=>"000100100",
  21324=>"010100100",
  21325=>"000100110",
  21326=>"011110011",
  21327=>"011111101",
  21328=>"000110111",
  21329=>"001000000",
  21330=>"001000001",
  21331=>"000011101",
  21332=>"110110101",
  21333=>"011000011",
  21334=>"000000101",
  21335=>"111111011",
  21336=>"001010001",
  21337=>"100000011",
  21338=>"100010111",
  21339=>"111001011",
  21340=>"101111100",
  21341=>"000000000",
  21342=>"101110011",
  21343=>"000000111",
  21344=>"011100100",
  21345=>"001111001",
  21346=>"101101000",
  21347=>"010001000",
  21348=>"011101011",
  21349=>"010100001",
  21350=>"100011011",
  21351=>"010000110",
  21352=>"110000010",
  21353=>"101100101",
  21354=>"011010000",
  21355=>"010110110",
  21356=>"001110110",
  21357=>"101100010",
  21358=>"110000011",
  21359=>"011011011",
  21360=>"000100010",
  21361=>"100000000",
  21362=>"100010100",
  21363=>"101010010",
  21364=>"000000001",
  21365=>"011000111",
  21366=>"101000110",
  21367=>"001010010",
  21368=>"111000000",
  21369=>"101100001",
  21370=>"100100100",
  21371=>"100000110",
  21372=>"000001000",
  21373=>"011001001",
  21374=>"100000011",
  21375=>"000001010",
  21376=>"011001110",
  21377=>"000010101",
  21378=>"000110111",
  21379=>"100100100",
  21380=>"000010100",
  21381=>"000101010",
  21382=>"110000100",
  21383=>"101100111",
  21384=>"000000000",
  21385=>"010000001",
  21386=>"100100011",
  21387=>"110011110",
  21388=>"000000110",
  21389=>"111101111",
  21390=>"111111101",
  21391=>"000011000",
  21392=>"001000011",
  21393=>"000101110",
  21394=>"010100010",
  21395=>"111001110",
  21396=>"001100010",
  21397=>"001101001",
  21398=>"001101001",
  21399=>"001011111",
  21400=>"100001011",
  21401=>"110100010",
  21402=>"101100011",
  21403=>"101001111",
  21404=>"011011010",
  21405=>"111011000",
  21406=>"111001010",
  21407=>"111101000",
  21408=>"011011010",
  21409=>"001010110",
  21410=>"110011000",
  21411=>"110010110",
  21412=>"011011000",
  21413=>"010110111",
  21414=>"110111010",
  21415=>"110100100",
  21416=>"100010001",
  21417=>"001001000",
  21418=>"011110001",
  21419=>"100111010",
  21420=>"101010000",
  21421=>"111010110",
  21422=>"001111111",
  21423=>"100001110",
  21424=>"001110000",
  21425=>"000101111",
  21426=>"110000111",
  21427=>"110010100",
  21428=>"001010110",
  21429=>"000001010",
  21430=>"011000010",
  21431=>"111010000",
  21432=>"011010001",
  21433=>"010101100",
  21434=>"111010110",
  21435=>"101001101",
  21436=>"011001001",
  21437=>"010001111",
  21438=>"111111111",
  21439=>"110000000",
  21440=>"101101111",
  21441=>"100010101",
  21442=>"110001111",
  21443=>"101100111",
  21444=>"001000011",
  21445=>"010101001",
  21446=>"001011010",
  21447=>"001110101",
  21448=>"101100101",
  21449=>"100110010",
  21450=>"010101110",
  21451=>"111111000",
  21452=>"000011000",
  21453=>"110011101",
  21454=>"111101100",
  21455=>"100111010",
  21456=>"001010100",
  21457=>"001000010",
  21458=>"111100001",
  21459=>"111011111",
  21460=>"001011100",
  21461=>"101001011",
  21462=>"011010111",
  21463=>"111010001",
  21464=>"010010000",
  21465=>"100110101",
  21466=>"101000001",
  21467=>"011011011",
  21468=>"001111110",
  21469=>"101100010",
  21470=>"011000111",
  21471=>"001001111",
  21472=>"110100110",
  21473=>"100100111",
  21474=>"100101101",
  21475=>"000011010",
  21476=>"100100111",
  21477=>"001100111",
  21478=>"001000101",
  21479=>"111111001",
  21480=>"111010000",
  21481=>"000011111",
  21482=>"110101010",
  21483=>"000010011",
  21484=>"011100000",
  21485=>"001101011",
  21486=>"101110010",
  21487=>"111001110",
  21488=>"011011011",
  21489=>"101001111",
  21490=>"011100000",
  21491=>"100001111",
  21492=>"011011110",
  21493=>"011001110",
  21494=>"100010010",
  21495=>"010000101",
  21496=>"101110010",
  21497=>"010110110",
  21498=>"111001101",
  21499=>"101001100",
  21500=>"100100011",
  21501=>"001000011",
  21502=>"001110100",
  21503=>"101100000",
  21504=>"111011000",
  21505=>"101110001",
  21506=>"101110011",
  21507=>"010001101",
  21508=>"111010101",
  21509=>"110100100",
  21510=>"111010011",
  21511=>"111111011",
  21512=>"011011101",
  21513=>"000010100",
  21514=>"010110101",
  21515=>"001110111",
  21516=>"001001011",
  21517=>"101011010",
  21518=>"110011110",
  21519=>"000000110",
  21520=>"011110110",
  21521=>"001000111",
  21522=>"000010011",
  21523=>"110010011",
  21524=>"001101010",
  21525=>"111000110",
  21526=>"001100010",
  21527=>"011101000",
  21528=>"010001110",
  21529=>"001000001",
  21530=>"110111011",
  21531=>"100100111",
  21532=>"110010111",
  21533=>"010001111",
  21534=>"111110111",
  21535=>"000101010",
  21536=>"110010100",
  21537=>"110100111",
  21538=>"000001101",
  21539=>"001010000",
  21540=>"100110011",
  21541=>"100111100",
  21542=>"111011001",
  21543=>"110100000",
  21544=>"001111001",
  21545=>"101000110",
  21546=>"110111101",
  21547=>"000011011",
  21548=>"010011101",
  21549=>"011010001",
  21550=>"000101010",
  21551=>"010000101",
  21552=>"100101011",
  21553=>"001001110",
  21554=>"001011111",
  21555=>"100100101",
  21556=>"101011000",
  21557=>"010011100",
  21558=>"110110111",
  21559=>"101100011",
  21560=>"010001100",
  21561=>"100110000",
  21562=>"011011010",
  21563=>"001001011",
  21564=>"000010110",
  21565=>"110100010",
  21566=>"001111000",
  21567=>"111010010",
  21568=>"100111011",
  21569=>"000000001",
  21570=>"011000001",
  21571=>"101101111",
  21572=>"100011000",
  21573=>"111010000",
  21574=>"111110000",
  21575=>"100110011",
  21576=>"001100000",
  21577=>"111000111",
  21578=>"110010110",
  21579=>"110110100",
  21580=>"011001101",
  21581=>"011011101",
  21582=>"110111101",
  21583=>"000101101",
  21584=>"001101000",
  21585=>"010110111",
  21586=>"110110110",
  21587=>"001001010",
  21588=>"111010110",
  21589=>"000111000",
  21590=>"000110010",
  21591=>"100011101",
  21592=>"000101101",
  21593=>"001100111",
  21594=>"101101000",
  21595=>"111010000",
  21596=>"000100101",
  21597=>"111101001",
  21598=>"011101101",
  21599=>"110100000",
  21600=>"100110011",
  21601=>"110110110",
  21602=>"001011011",
  21603=>"101011001",
  21604=>"110100010",
  21605=>"011110001",
  21606=>"101001101",
  21607=>"100011110",
  21608=>"001100111",
  21609=>"101110011",
  21610=>"010010000",
  21611=>"110100110",
  21612=>"000000110",
  21613=>"000011011",
  21614=>"011111111",
  21615=>"111011010",
  21616=>"111110011",
  21617=>"101010010",
  21618=>"101100001",
  21619=>"111000000",
  21620=>"010010100",
  21621=>"000001011",
  21622=>"000011100",
  21623=>"000000010",
  21624=>"111111010",
  21625=>"010000000",
  21626=>"000100000",
  21627=>"011100001",
  21628=>"001011011",
  21629=>"100110001",
  21630=>"001010001",
  21631=>"110111111",
  21632=>"001111110",
  21633=>"111011001",
  21634=>"111111110",
  21635=>"011010111",
  21636=>"111111010",
  21637=>"000101100",
  21638=>"001000010",
  21639=>"010011100",
  21640=>"100110101",
  21641=>"001000111",
  21642=>"000101101",
  21643=>"111110111",
  21644=>"000101110",
  21645=>"100000001",
  21646=>"110001111",
  21647=>"000100000",
  21648=>"110011000",
  21649=>"010000000",
  21650=>"101000001",
  21651=>"011101100",
  21652=>"111100001",
  21653=>"000110001",
  21654=>"100001110",
  21655=>"011100000",
  21656=>"100000000",
  21657=>"111101111",
  21658=>"000111011",
  21659=>"010100010",
  21660=>"100000011",
  21661=>"100001110",
  21662=>"011000101",
  21663=>"011001111",
  21664=>"001010100",
  21665=>"101111100",
  21666=>"011010101",
  21667=>"101101011",
  21668=>"110101110",
  21669=>"110010011",
  21670=>"010011001",
  21671=>"000100000",
  21672=>"100111000",
  21673=>"000011000",
  21674=>"101100000",
  21675=>"000010110",
  21676=>"011011001",
  21677=>"011111001",
  21678=>"001000111",
  21679=>"001000000",
  21680=>"110011000",
  21681=>"100101111",
  21682=>"111111000",
  21683=>"101000010",
  21684=>"011111000",
  21685=>"100101010",
  21686=>"000000100",
  21687=>"000010100",
  21688=>"111000000",
  21689=>"100100100",
  21690=>"001101101",
  21691=>"100101100",
  21692=>"100001010",
  21693=>"110001111",
  21694=>"110011111",
  21695=>"001110100",
  21696=>"000110000",
  21697=>"011100011",
  21698=>"100111110",
  21699=>"110000110",
  21700=>"001100000",
  21701=>"011100001",
  21702=>"100000111",
  21703=>"000111110",
  21704=>"110001000",
  21705=>"010111000",
  21706=>"110001011",
  21707=>"001000100",
  21708=>"100101000",
  21709=>"011101101",
  21710=>"110111000",
  21711=>"010101000",
  21712=>"110111010",
  21713=>"000001000",
  21714=>"000010111",
  21715=>"110101011",
  21716=>"111001000",
  21717=>"100001101",
  21718=>"011101000",
  21719=>"101101000",
  21720=>"001101010",
  21721=>"100000001",
  21722=>"101101100",
  21723=>"110001011",
  21724=>"110011000",
  21725=>"101000000",
  21726=>"001010000",
  21727=>"100011001",
  21728=>"001000010",
  21729=>"110110100",
  21730=>"100000010",
  21731=>"000101111",
  21732=>"100110000",
  21733=>"000000100",
  21734=>"110010011",
  21735=>"000111100",
  21736=>"010000010",
  21737=>"000101001",
  21738=>"110101110",
  21739=>"111100000",
  21740=>"011100101",
  21741=>"111000100",
  21742=>"100101010",
  21743=>"100000010",
  21744=>"111000011",
  21745=>"111010110",
  21746=>"110100011",
  21747=>"000111110",
  21748=>"001111111",
  21749=>"100001000",
  21750=>"110010100",
  21751=>"100100001",
  21752=>"111011101",
  21753=>"110111101",
  21754=>"011000010",
  21755=>"100000111",
  21756=>"101000000",
  21757=>"000000000",
  21758=>"010011111",
  21759=>"110110001",
  21760=>"111001000",
  21761=>"001111010",
  21762=>"110000111",
  21763=>"000101000",
  21764=>"011001010",
  21765=>"100011001",
  21766=>"010001111",
  21767=>"100001111",
  21768=>"111011000",
  21769=>"111101010",
  21770=>"010110111",
  21771=>"111000100",
  21772=>"111110010",
  21773=>"000101110",
  21774=>"011100010",
  21775=>"111110000",
  21776=>"011101011",
  21777=>"111011010",
  21778=>"111101010",
  21779=>"001010111",
  21780=>"111110110",
  21781=>"011101111",
  21782=>"011010001",
  21783=>"000010111",
  21784=>"001100111",
  21785=>"100000000",
  21786=>"100011100",
  21787=>"001100100",
  21788=>"011111011",
  21789=>"101111011",
  21790=>"111011110",
  21791=>"010000001",
  21792=>"111001001",
  21793=>"101100000",
  21794=>"000100110",
  21795=>"011110001",
  21796=>"101100000",
  21797=>"111011000",
  21798=>"001001000",
  21799=>"011001101",
  21800=>"011010010",
  21801=>"111111101",
  21802=>"101010111",
  21803=>"100111011",
  21804=>"000100001",
  21805=>"111100101",
  21806=>"000001000",
  21807=>"010000100",
  21808=>"110100111",
  21809=>"101010010",
  21810=>"010010010",
  21811=>"100001100",
  21812=>"111101110",
  21813=>"000010001",
  21814=>"111100001",
  21815=>"011001000",
  21816=>"001101011",
  21817=>"001010111",
  21818=>"100001001",
  21819=>"110110101",
  21820=>"111111000",
  21821=>"000110010",
  21822=>"101110110",
  21823=>"000111000",
  21824=>"111110011",
  21825=>"011111111",
  21826=>"000011111",
  21827=>"011010100",
  21828=>"100100101",
  21829=>"010111001",
  21830=>"110010001",
  21831=>"000111101",
  21832=>"011101011",
  21833=>"001110010",
  21834=>"111001100",
  21835=>"101001111",
  21836=>"101000011",
  21837=>"001111100",
  21838=>"010110110",
  21839=>"010000001",
  21840=>"000011110",
  21841=>"000010101",
  21842=>"110001010",
  21843=>"100001111",
  21844=>"011100011",
  21845=>"010010111",
  21846=>"101111100",
  21847=>"010100100",
  21848=>"100100011",
  21849=>"001111111",
  21850=>"010100111",
  21851=>"111010101",
  21852=>"111010110",
  21853=>"001101011",
  21854=>"111000011",
  21855=>"010011111",
  21856=>"100110111",
  21857=>"010011111",
  21858=>"001001100",
  21859=>"001000010",
  21860=>"011011110",
  21861=>"010100001",
  21862=>"000100001",
  21863=>"110111111",
  21864=>"101000001",
  21865=>"110100100",
  21866=>"011111011",
  21867=>"010110010",
  21868=>"101000111",
  21869=>"111001000",
  21870=>"100000111",
  21871=>"000001011",
  21872=>"000000010",
  21873=>"100000011",
  21874=>"001101010",
  21875=>"010101000",
  21876=>"111111010",
  21877=>"101000100",
  21878=>"011111111",
  21879=>"110111011",
  21880=>"010000011",
  21881=>"001101111",
  21882=>"110010001",
  21883=>"000111110",
  21884=>"011100110",
  21885=>"010111011",
  21886=>"001100111",
  21887=>"111110001",
  21888=>"000100100",
  21889=>"101010000",
  21890=>"010011101",
  21891=>"010110011",
  21892=>"100011011",
  21893=>"110101001",
  21894=>"100111101",
  21895=>"010100001",
  21896=>"010111111",
  21897=>"110000101",
  21898=>"010001001",
  21899=>"100110001",
  21900=>"110111010",
  21901=>"000010110",
  21902=>"000101010",
  21903=>"000101010",
  21904=>"111100011",
  21905=>"101100001",
  21906=>"100100001",
  21907=>"110000101",
  21908=>"000111111",
  21909=>"101000100",
  21910=>"001100001",
  21911=>"101000100",
  21912=>"000011000",
  21913=>"011100111",
  21914=>"110001110",
  21915=>"000111100",
  21916=>"101011001",
  21917=>"111000001",
  21918=>"010011111",
  21919=>"011100001",
  21920=>"110100111",
  21921=>"101000100",
  21922=>"101000010",
  21923=>"111010101",
  21924=>"111100110",
  21925=>"010110010",
  21926=>"101100000",
  21927=>"101110111",
  21928=>"111011010",
  21929=>"011100011",
  21930=>"110110100",
  21931=>"010101101",
  21932=>"110010100",
  21933=>"111001001",
  21934=>"011111110",
  21935=>"111111111",
  21936=>"101010111",
  21937=>"101100100",
  21938=>"011000110",
  21939=>"001110111",
  21940=>"011111000",
  21941=>"111010111",
  21942=>"000110110",
  21943=>"100010001",
  21944=>"111001000",
  21945=>"110011010",
  21946=>"101110011",
  21947=>"000111110",
  21948=>"011100000",
  21949=>"111101100",
  21950=>"000000000",
  21951=>"100010110",
  21952=>"011000001",
  21953=>"100011111",
  21954=>"110011011",
  21955=>"000111100",
  21956=>"000101110",
  21957=>"001001100",
  21958=>"010111011",
  21959=>"001000100",
  21960=>"000110101",
  21961=>"111100000",
  21962=>"000101100",
  21963=>"001110000",
  21964=>"010001100",
  21965=>"000110001",
  21966=>"100010111",
  21967=>"001011010",
  21968=>"010101110",
  21969=>"110100111",
  21970=>"000101110",
  21971=>"110101111",
  21972=>"111011011",
  21973=>"111011000",
  21974=>"101011001",
  21975=>"001010110",
  21976=>"011000111",
  21977=>"111110111",
  21978=>"000000111",
  21979=>"101111110",
  21980=>"101001101",
  21981=>"111001000",
  21982=>"111000001",
  21983=>"001000010",
  21984=>"100111001",
  21985=>"010000011",
  21986=>"110010101",
  21987=>"100000010",
  21988=>"000001001",
  21989=>"010001001",
  21990=>"000100101",
  21991=>"001001001",
  21992=>"110101100",
  21993=>"100011111",
  21994=>"000100011",
  21995=>"010101000",
  21996=>"000001111",
  21997=>"100000000",
  21998=>"111101100",
  21999=>"101100011",
  22000=>"000111100",
  22001=>"011011101",
  22002=>"101110100",
  22003=>"010011100",
  22004=>"101001110",
  22005=>"001001101",
  22006=>"110011011",
  22007=>"100100001",
  22008=>"000001000",
  22009=>"101110100",
  22010=>"101011111",
  22011=>"101101010",
  22012=>"100011101",
  22013=>"111000000",
  22014=>"111011010",
  22015=>"011100100",
  22016=>"000001000",
  22017=>"010000010",
  22018=>"001011100",
  22019=>"011000000",
  22020=>"011101010",
  22021=>"110010110",
  22022=>"011010001",
  22023=>"111101111",
  22024=>"100010011",
  22025=>"111100010",
  22026=>"000110101",
  22027=>"010001011",
  22028=>"010000111",
  22029=>"010001100",
  22030=>"110000100",
  22031=>"000111011",
  22032=>"111000001",
  22033=>"001001100",
  22034=>"101011100",
  22035=>"010001101",
  22036=>"010001101",
  22037=>"101110101",
  22038=>"010000111",
  22039=>"001001111",
  22040=>"100000110",
  22041=>"001011001",
  22042=>"110001000",
  22043=>"110110000",
  22044=>"110001010",
  22045=>"111100000",
  22046=>"000000001",
  22047=>"000000101",
  22048=>"000101011",
  22049=>"110100010",
  22050=>"010000111",
  22051=>"100000101",
  22052=>"100111110",
  22053=>"111001111",
  22054=>"111011000",
  22055=>"100010000",
  22056=>"010011001",
  22057=>"111101000",
  22058=>"010000010",
  22059=>"100000000",
  22060=>"100101000",
  22061=>"011010100",
  22062=>"011011111",
  22063=>"000001110",
  22064=>"000100011",
  22065=>"010111000",
  22066=>"010011010",
  22067=>"100101010",
  22068=>"011000010",
  22069=>"000101100",
  22070=>"101001100",
  22071=>"010110000",
  22072=>"100011101",
  22073=>"010011100",
  22074=>"111000000",
  22075=>"010101000",
  22076=>"000101011",
  22077=>"110000111",
  22078=>"011001001",
  22079=>"100110001",
  22080=>"011100011",
  22081=>"110111110",
  22082=>"000100000",
  22083=>"100100011",
  22084=>"001000010",
  22085=>"011010000",
  22086=>"111000001",
  22087=>"001010110",
  22088=>"010011000",
  22089=>"001111000",
  22090=>"100111011",
  22091=>"000100100",
  22092=>"000010000",
  22093=>"100001010",
  22094=>"010100011",
  22095=>"111111101",
  22096=>"011000111",
  22097=>"101001110",
  22098=>"000001001",
  22099=>"000111101",
  22100=>"010110100",
  22101=>"010110011",
  22102=>"001111011",
  22103=>"001110100",
  22104=>"010100101",
  22105=>"101100111",
  22106=>"010111010",
  22107=>"110011100",
  22108=>"111111100",
  22109=>"111101101",
  22110=>"010001111",
  22111=>"001101010",
  22112=>"011101010",
  22113=>"001110100",
  22114=>"111000000",
  22115=>"110010000",
  22116=>"110010110",
  22117=>"000011011",
  22118=>"001100101",
  22119=>"000100101",
  22120=>"111001000",
  22121=>"011100010",
  22122=>"000011101",
  22123=>"111101011",
  22124=>"100001001",
  22125=>"011000001",
  22126=>"001110111",
  22127=>"011111010",
  22128=>"111110000",
  22129=>"011111011",
  22130=>"100111010",
  22131=>"011001101",
  22132=>"101111101",
  22133=>"010101100",
  22134=>"000111110",
  22135=>"110110111",
  22136=>"000001010",
  22137=>"010101110",
  22138=>"100111010",
  22139=>"101101110",
  22140=>"110101001",
  22141=>"001010111",
  22142=>"111010101",
  22143=>"101110110",
  22144=>"111101111",
  22145=>"000100100",
  22146=>"101100111",
  22147=>"110010101",
  22148=>"100001100",
  22149=>"011011000",
  22150=>"001101100",
  22151=>"000111001",
  22152=>"001011110",
  22153=>"110001110",
  22154=>"111111111",
  22155=>"010101010",
  22156=>"110010010",
  22157=>"110001110",
  22158=>"110110000",
  22159=>"001100110",
  22160=>"110001010",
  22161=>"101000100",
  22162=>"110110100",
  22163=>"011111110",
  22164=>"000101000",
  22165=>"101011010",
  22166=>"001101010",
  22167=>"010000000",
  22168=>"111111011",
  22169=>"110000111",
  22170=>"011110111",
  22171=>"001110101",
  22172=>"010010010",
  22173=>"000000101",
  22174=>"110000011",
  22175=>"100011110",
  22176=>"111000111",
  22177=>"101100111",
  22178=>"010101011",
  22179=>"100000001",
  22180=>"000100001",
  22181=>"000000100",
  22182=>"001100000",
  22183=>"100101111",
  22184=>"000111100",
  22185=>"010111111",
  22186=>"110110000",
  22187=>"011001111",
  22188=>"011011111",
  22189=>"011111001",
  22190=>"001001001",
  22191=>"011101101",
  22192=>"010110000",
  22193=>"111010111",
  22194=>"111010010",
  22195=>"101010101",
  22196=>"100010011",
  22197=>"001001001",
  22198=>"110010000",
  22199=>"000001100",
  22200=>"111110101",
  22201=>"011011110",
  22202=>"000101011",
  22203=>"100000000",
  22204=>"011100101",
  22205=>"011111000",
  22206=>"110101100",
  22207=>"000000100",
  22208=>"111110101",
  22209=>"000001000",
  22210=>"011000101",
  22211=>"101001110",
  22212=>"100101110",
  22213=>"000101101",
  22214=>"001100100",
  22215=>"011111000",
  22216=>"111101110",
  22217=>"101001001",
  22218=>"010001000",
  22219=>"101000110",
  22220=>"110010100",
  22221=>"101000010",
  22222=>"000111001",
  22223=>"001111000",
  22224=>"011101011",
  22225=>"000100000",
  22226=>"000110011",
  22227=>"000000000",
  22228=>"100010110",
  22229=>"001001111",
  22230=>"101111010",
  22231=>"010111100",
  22232=>"110010100",
  22233=>"100011010",
  22234=>"111101100",
  22235=>"011111001",
  22236=>"111100101",
  22237=>"110010000",
  22238=>"000010100",
  22239=>"010110111",
  22240=>"111010100",
  22241=>"100001100",
  22242=>"100101000",
  22243=>"011101110",
  22244=>"111011100",
  22245=>"010101100",
  22246=>"110111111",
  22247=>"010110010",
  22248=>"000001100",
  22249=>"101100100",
  22250=>"100111011",
  22251=>"000000011",
  22252=>"110100011",
  22253=>"010111010",
  22254=>"000010001",
  22255=>"100010100",
  22256=>"100110110",
  22257=>"101100011",
  22258=>"101101010",
  22259=>"001111011",
  22260=>"111100000",
  22261=>"001101110",
  22262=>"011110010",
  22263=>"011000110",
  22264=>"011110110",
  22265=>"111110110",
  22266=>"111111111",
  22267=>"111110100",
  22268=>"001001101",
  22269=>"011011010",
  22270=>"100100111",
  22271=>"010011011",
  22272=>"101001011",
  22273=>"010100011",
  22274=>"010110000",
  22275=>"011000011",
  22276=>"110000000",
  22277=>"000101101",
  22278=>"000010011",
  22279=>"000101010",
  22280=>"000100010",
  22281=>"010111101",
  22282=>"000010111",
  22283=>"100100100",
  22284=>"000001111",
  22285=>"110001111",
  22286=>"011101111",
  22287=>"011010110",
  22288=>"010001110",
  22289=>"100000100",
  22290=>"010011000",
  22291=>"011001011",
  22292=>"001011100",
  22293=>"110100001",
  22294=>"000010000",
  22295=>"010011101",
  22296=>"001000111",
  22297=>"000001111",
  22298=>"001000000",
  22299=>"100110001",
  22300=>"110111100",
  22301=>"111001110",
  22302=>"011111101",
  22303=>"001000101",
  22304=>"011011011",
  22305=>"011010101",
  22306=>"101010100",
  22307=>"101111000",
  22308=>"000001111",
  22309=>"110000001",
  22310=>"100001110",
  22311=>"000101100",
  22312=>"011010001",
  22313=>"101101000",
  22314=>"101111011",
  22315=>"011001000",
  22316=>"010110100",
  22317=>"111100000",
  22318=>"110111100",
  22319=>"001111100",
  22320=>"001000111",
  22321=>"111010010",
  22322=>"100000111",
  22323=>"111011101",
  22324=>"111101110",
  22325=>"001010110",
  22326=>"111111000",
  22327=>"010011110",
  22328=>"010110101",
  22329=>"111001000",
  22330=>"111100000",
  22331=>"000010110",
  22332=>"100111010",
  22333=>"110011010",
  22334=>"001010100",
  22335=>"111101111",
  22336=>"100100001",
  22337=>"110011000",
  22338=>"110101000",
  22339=>"010111011",
  22340=>"111110010",
  22341=>"101000100",
  22342=>"010100100",
  22343=>"011101100",
  22344=>"000110001",
  22345=>"010101010",
  22346=>"010101011",
  22347=>"111000011",
  22348=>"010001101",
  22349=>"101111101",
  22350=>"000000001",
  22351=>"000010000",
  22352=>"010000100",
  22353=>"000101111",
  22354=>"100000010",
  22355=>"000000111",
  22356=>"011011110",
  22357=>"100100101",
  22358=>"000001000",
  22359=>"111010000",
  22360=>"010100101",
  22361=>"011110010",
  22362=>"010100011",
  22363=>"111111000",
  22364=>"011010110",
  22365=>"000111111",
  22366=>"001111100",
  22367=>"110000000",
  22368=>"111001110",
  22369=>"000000101",
  22370=>"001100110",
  22371=>"001001111",
  22372=>"100000001",
  22373=>"100110001",
  22374=>"111100000",
  22375=>"111100110",
  22376=>"011001000",
  22377=>"110001010",
  22378=>"001100010",
  22379=>"011111110",
  22380=>"011101111",
  22381=>"011010101",
  22382=>"110000011",
  22383=>"101101110",
  22384=>"000010110",
  22385=>"011100000",
  22386=>"110101001",
  22387=>"011011110",
  22388=>"010111010",
  22389=>"111110101",
  22390=>"010000010",
  22391=>"001111101",
  22392=>"000000111",
  22393=>"110011100",
  22394=>"100111101",
  22395=>"111001100",
  22396=>"100101101",
  22397=>"001000001",
  22398=>"111001111",
  22399=>"110101111",
  22400=>"111010010",
  22401=>"000100101",
  22402=>"001000000",
  22403=>"110011010",
  22404=>"011000111",
  22405=>"110110011",
  22406=>"010010110",
  22407=>"011011001",
  22408=>"011011000",
  22409=>"100010101",
  22410=>"110110100",
  22411=>"100010110",
  22412=>"100011000",
  22413=>"101001101",
  22414=>"111111011",
  22415=>"110111010",
  22416=>"111001011",
  22417=>"101011000",
  22418=>"001101010",
  22419=>"000011001",
  22420=>"111100110",
  22421=>"001100110",
  22422=>"000000010",
  22423=>"010010111",
  22424=>"011011101",
  22425=>"011010101",
  22426=>"111111101",
  22427=>"100000010",
  22428=>"111110100",
  22429=>"100100001",
  22430=>"110000010",
  22431=>"101000110",
  22432=>"010011100",
  22433=>"100100110",
  22434=>"100011101",
  22435=>"011000111",
  22436=>"000100100",
  22437=>"110011110",
  22438=>"000110001",
  22439=>"010001110",
  22440=>"000001011",
  22441=>"110011101",
  22442=>"000110000",
  22443=>"101100001",
  22444=>"011110111",
  22445=>"001110000",
  22446=>"110111001",
  22447=>"100001100",
  22448=>"111011000",
  22449=>"111100011",
  22450=>"001110011",
  22451=>"100001110",
  22452=>"001010010",
  22453=>"010110110",
  22454=>"011010011",
  22455=>"011001011",
  22456=>"110000110",
  22457=>"110110111",
  22458=>"001001101",
  22459=>"111000000",
  22460=>"110110011",
  22461=>"001011111",
  22462=>"010000110",
  22463=>"001110110",
  22464=>"110111111",
  22465=>"011010111",
  22466=>"100100000",
  22467=>"111111010",
  22468=>"000111001",
  22469=>"111010001",
  22470=>"101111111",
  22471=>"101001000",
  22472=>"111000100",
  22473=>"001111101",
  22474=>"110000111",
  22475=>"000111110",
  22476=>"001011001",
  22477=>"111000101",
  22478=>"001001000",
  22479=>"010111000",
  22480=>"000110111",
  22481=>"000010111",
  22482=>"010001011",
  22483=>"101110010",
  22484=>"100001110",
  22485=>"010001000",
  22486=>"101101100",
  22487=>"110100000",
  22488=>"010101100",
  22489=>"100001010",
  22490=>"011000001",
  22491=>"011111001",
  22492=>"001010110",
  22493=>"011110000",
  22494=>"100011011",
  22495=>"010111110",
  22496=>"111101101",
  22497=>"110001111",
  22498=>"100101101",
  22499=>"011100100",
  22500=>"010011000",
  22501=>"010110101",
  22502=>"111010011",
  22503=>"000101111",
  22504=>"101101100",
  22505=>"000111001",
  22506=>"100100111",
  22507=>"011001001",
  22508=>"111011010",
  22509=>"000111010",
  22510=>"100111000",
  22511=>"010100000",
  22512=>"101011111",
  22513=>"010100100",
  22514=>"101000001",
  22515=>"101100100",
  22516=>"001111011",
  22517=>"011100101",
  22518=>"111010010",
  22519=>"000101000",
  22520=>"101110111",
  22521=>"101000000",
  22522=>"011001110",
  22523=>"110010100",
  22524=>"000101101",
  22525=>"100001111",
  22526=>"111100011",
  22527=>"111111010",
  22528=>"001100001",
  22529=>"101101010",
  22530=>"101110100",
  22531=>"000000100",
  22532=>"011000010",
  22533=>"101101111",
  22534=>"000111100",
  22535=>"111100010",
  22536=>"110101001",
  22537=>"010011100",
  22538=>"110000100",
  22539=>"011100101",
  22540=>"101000110",
  22541=>"110101000",
  22542=>"000100110",
  22543=>"111101010",
  22544=>"110111000",
  22545=>"000110000",
  22546=>"101101010",
  22547=>"011111111",
  22548=>"111110010",
  22549=>"011101111",
  22550=>"011011010",
  22551=>"001100100",
  22552=>"001001001",
  22553=>"101110101",
  22554=>"000001000",
  22555=>"100011010",
  22556=>"111110011",
  22557=>"000000111",
  22558=>"011100000",
  22559=>"100001111",
  22560=>"110100100",
  22561=>"011001100",
  22562=>"000101001",
  22563=>"001001001",
  22564=>"111111001",
  22565=>"101010100",
  22566=>"010100001",
  22567=>"111111011",
  22568=>"001010001",
  22569=>"011110111",
  22570=>"111111110",
  22571=>"110100000",
  22572=>"111011011",
  22573=>"111100110",
  22574=>"101111011",
  22575=>"110101111",
  22576=>"011000100",
  22577=>"010000000",
  22578=>"101011010",
  22579=>"110101000",
  22580=>"000101010",
  22581=>"100000000",
  22582=>"111010000",
  22583=>"001011010",
  22584=>"010000110",
  22585=>"010010111",
  22586=>"000101111",
  22587=>"111111101",
  22588=>"100001000",
  22589=>"100101111",
  22590=>"100011001",
  22591=>"100100100",
  22592=>"110001111",
  22593=>"000101100",
  22594=>"000000010",
  22595=>"011110010",
  22596=>"100001101",
  22597=>"110000110",
  22598=>"100011100",
  22599=>"100111100",
  22600=>"111100111",
  22601=>"001001011",
  22602=>"000001111",
  22603=>"000010100",
  22604=>"001100011",
  22605=>"010100010",
  22606=>"011001011",
  22607=>"000000001",
  22608=>"110000011",
  22609=>"001101001",
  22610=>"000011000",
  22611=>"101001100",
  22612=>"001111000",
  22613=>"010011011",
  22614=>"001010100",
  22615=>"110101110",
  22616=>"111110110",
  22617=>"000001100",
  22618=>"000000100",
  22619=>"110011111",
  22620=>"001110010",
  22621=>"111111000",
  22622=>"110000101",
  22623=>"100011100",
  22624=>"100001101",
  22625=>"111101010",
  22626=>"001011110",
  22627=>"101101000",
  22628=>"000111111",
  22629=>"010000101",
  22630=>"010101001",
  22631=>"000000000",
  22632=>"110100110",
  22633=>"010000110",
  22634=>"000001000",
  22635=>"010110101",
  22636=>"100000000",
  22637=>"110000111",
  22638=>"010000101",
  22639=>"111011110",
  22640=>"100010000",
  22641=>"010011000",
  22642=>"010111101",
  22643=>"101101001",
  22644=>"001110100",
  22645=>"100110110",
  22646=>"100001101",
  22647=>"100001001",
  22648=>"101110011",
  22649=>"111110000",
  22650=>"100110001",
  22651=>"100101101",
  22652=>"100010111",
  22653=>"001010010",
  22654=>"110100000",
  22655=>"100001000",
  22656=>"100000010",
  22657=>"100100011",
  22658=>"100111001",
  22659=>"110011110",
  22660=>"000000110",
  22661=>"100110010",
  22662=>"110100011",
  22663=>"101000010",
  22664=>"110110110",
  22665=>"011000101",
  22666=>"100100101",
  22667=>"101010001",
  22668=>"110100100",
  22669=>"111010110",
  22670=>"000001110",
  22671=>"000000010",
  22672=>"001011101",
  22673=>"110001000",
  22674=>"001010110",
  22675=>"010111100",
  22676=>"110010001",
  22677=>"011110111",
  22678=>"010101001",
  22679=>"111001111",
  22680=>"101000010",
  22681=>"011101000",
  22682=>"000000011",
  22683=>"011011100",
  22684=>"000001000",
  22685=>"001011100",
  22686=>"100000100",
  22687=>"110010001",
  22688=>"111111000",
  22689=>"011001100",
  22690=>"001000100",
  22691=>"011100111",
  22692=>"000101011",
  22693=>"001000010",
  22694=>"101100011",
  22695=>"000011000",
  22696=>"011011100",
  22697=>"011010100",
  22698=>"101000001",
  22699=>"111000100",
  22700=>"101101101",
  22701=>"110011101",
  22702=>"010010110",
  22703=>"101001011",
  22704=>"100101101",
  22705=>"110101100",
  22706=>"011110000",
  22707=>"000001011",
  22708=>"011011000",
  22709=>"000010100",
  22710=>"100011111",
  22711=>"001000101",
  22712=>"110110001",
  22713=>"001000000",
  22714=>"110110000",
  22715=>"011111100",
  22716=>"010111100",
  22717=>"000101101",
  22718=>"001101101",
  22719=>"000101001",
  22720=>"101110001",
  22721=>"001001010",
  22722=>"000100000",
  22723=>"001101100",
  22724=>"000101001",
  22725=>"110110001",
  22726=>"111010110",
  22727=>"100111000",
  22728=>"001011110",
  22729=>"011110100",
  22730=>"111000100",
  22731=>"111101101",
  22732=>"000000110",
  22733=>"010010111",
  22734=>"010000100",
  22735=>"100100100",
  22736=>"010101001",
  22737=>"000000111",
  22738=>"100100010",
  22739=>"110100010",
  22740=>"111000111",
  22741=>"100101110",
  22742=>"101111011",
  22743=>"110100011",
  22744=>"101100000",
  22745=>"110010100",
  22746=>"111000000",
  22747=>"111011000",
  22748=>"000000100",
  22749=>"111001111",
  22750=>"010001010",
  22751=>"101000111",
  22752=>"000001100",
  22753=>"001000011",
  22754=>"111011111",
  22755=>"001000010",
  22756=>"001010010",
  22757=>"100011100",
  22758=>"000001000",
  22759=>"010101111",
  22760=>"110000000",
  22761=>"100111111",
  22762=>"100100110",
  22763=>"101000101",
  22764=>"101001110",
  22765=>"000010111",
  22766=>"110000110",
  22767=>"010011100",
  22768=>"101010110",
  22769=>"001001100",
  22770=>"100100000",
  22771=>"001001010",
  22772=>"010000001",
  22773=>"111101101",
  22774=>"010011000",
  22775=>"001000101",
  22776=>"001000001",
  22777=>"001101000",
  22778=>"111111100",
  22779=>"010010101",
  22780=>"010110110",
  22781=>"011110010",
  22782=>"110001100",
  22783=>"101101111",
  22784=>"100000000",
  22785=>"100101100",
  22786=>"111010000",
  22787=>"100001101",
  22788=>"101000010",
  22789=>"111111010",
  22790=>"101010000",
  22791=>"111110110",
  22792=>"111011010",
  22793=>"110011111",
  22794=>"001110011",
  22795=>"001000000",
  22796=>"101101010",
  22797=>"111001111",
  22798=>"111101001",
  22799=>"100001100",
  22800=>"001001000",
  22801=>"001011110",
  22802=>"010010111",
  22803=>"111111101",
  22804=>"000110111",
  22805=>"100110010",
  22806=>"011001101",
  22807=>"011111010",
  22808=>"001000011",
  22809=>"101110110",
  22810=>"010110011",
  22811=>"111100100",
  22812=>"110100010",
  22813=>"101010000",
  22814=>"111001101",
  22815=>"001000111",
  22816=>"000011110",
  22817=>"001000001",
  22818=>"000100110",
  22819=>"001000100",
  22820=>"100011001",
  22821=>"010010001",
  22822=>"100100111",
  22823=>"111000011",
  22824=>"111000001",
  22825=>"110000011",
  22826=>"110011010",
  22827=>"010001010",
  22828=>"001010001",
  22829=>"001100001",
  22830=>"000000101",
  22831=>"010010110",
  22832=>"100101101",
  22833=>"100101111",
  22834=>"101001110",
  22835=>"010000101",
  22836=>"011010110",
  22837=>"100010001",
  22838=>"101001111",
  22839=>"011001010",
  22840=>"010110111",
  22841=>"000000010",
  22842=>"100010000",
  22843=>"000101110",
  22844=>"010001111",
  22845=>"111000110",
  22846=>"100000011",
  22847=>"001111101",
  22848=>"000010101",
  22849=>"010001001",
  22850=>"111010001",
  22851=>"110100110",
  22852=>"000001110",
  22853=>"010010001",
  22854=>"001011001",
  22855=>"100101110",
  22856=>"110100010",
  22857=>"000010100",
  22858=>"011001100",
  22859=>"000110010",
  22860=>"101111011",
  22861=>"111100011",
  22862=>"001111010",
  22863=>"010011010",
  22864=>"110001100",
  22865=>"101110000",
  22866=>"101010111",
  22867=>"011111111",
  22868=>"001000011",
  22869=>"010111111",
  22870=>"000010101",
  22871=>"010101110",
  22872=>"100111001",
  22873=>"001000111",
  22874=>"000110010",
  22875=>"000000010",
  22876=>"000100111",
  22877=>"100111111",
  22878=>"110001001",
  22879=>"111001001",
  22880=>"111000111",
  22881=>"000100010",
  22882=>"101001001",
  22883=>"101110100",
  22884=>"010001100",
  22885=>"101011101",
  22886=>"110001110",
  22887=>"101010001",
  22888=>"111110110",
  22889=>"010101101",
  22890=>"011010010",
  22891=>"100010111",
  22892=>"001000111",
  22893=>"111111011",
  22894=>"101111011",
  22895=>"010011100",
  22896=>"000111111",
  22897=>"101111000",
  22898=>"101010110",
  22899=>"011010110",
  22900=>"001101100",
  22901=>"001000001",
  22902=>"100011111",
  22903=>"010011110",
  22904=>"010111001",
  22905=>"000010000",
  22906=>"000101100",
  22907=>"010101010",
  22908=>"101101001",
  22909=>"111101111",
  22910=>"001111110",
  22911=>"110010101",
  22912=>"000000110",
  22913=>"001010000",
  22914=>"111010010",
  22915=>"000010011",
  22916=>"110111100",
  22917=>"101110110",
  22918=>"000011110",
  22919=>"110101101",
  22920=>"011101101",
  22921=>"101001000",
  22922=>"101011000",
  22923=>"000011010",
  22924=>"001000100",
  22925=>"111001001",
  22926=>"110001000",
  22927=>"011110111",
  22928=>"110011001",
  22929=>"100101100",
  22930=>"100101101",
  22931=>"010100101",
  22932=>"001000110",
  22933=>"010100000",
  22934=>"101110110",
  22935=>"000110111",
  22936=>"111001110",
  22937=>"111010101",
  22938=>"101001100",
  22939=>"010011011",
  22940=>"110000011",
  22941=>"110110111",
  22942=>"001101100",
  22943=>"011010011",
  22944=>"101011001",
  22945=>"000001001",
  22946=>"000001000",
  22947=>"000100011",
  22948=>"100110001",
  22949=>"010000001",
  22950=>"010111110",
  22951=>"010000000",
  22952=>"100110110",
  22953=>"101100000",
  22954=>"101100100",
  22955=>"011000101",
  22956=>"010000001",
  22957=>"010000000",
  22958=>"101001110",
  22959=>"110101111",
  22960=>"010001010",
  22961=>"001011000",
  22962=>"010000010",
  22963=>"010011010",
  22964=>"011100000",
  22965=>"000101111",
  22966=>"000110111",
  22967=>"111111011",
  22968=>"100100111",
  22969=>"110000111",
  22970=>"101010000",
  22971=>"111100100",
  22972=>"010110100",
  22973=>"011010100",
  22974=>"010110111",
  22975=>"001111000",
  22976=>"101111100",
  22977=>"011011010",
  22978=>"100011110",
  22979=>"111000101",
  22980=>"001111111",
  22981=>"001110001",
  22982=>"000110010",
  22983=>"111001010",
  22984=>"001011011",
  22985=>"011000101",
  22986=>"001110000",
  22987=>"010001001",
  22988=>"110101101",
  22989=>"111000000",
  22990=>"011110100",
  22991=>"101000100",
  22992=>"011000011",
  22993=>"001100110",
  22994=>"111000111",
  22995=>"001110010",
  22996=>"111101111",
  22997=>"001100001",
  22998=>"100011110",
  22999=>"101011011",
  23000=>"100101001",
  23001=>"010000100",
  23002=>"011111101",
  23003=>"010111000",
  23004=>"111100111",
  23005=>"000110010",
  23006=>"001100001",
  23007=>"010111101",
  23008=>"000110000",
  23009=>"111011110",
  23010=>"001000001",
  23011=>"010010001",
  23012=>"000001001",
  23013=>"000100010",
  23014=>"100100010",
  23015=>"101000010",
  23016=>"001100010",
  23017=>"000101001",
  23018=>"000010001",
  23019=>"010001001",
  23020=>"001000011",
  23021=>"011100010",
  23022=>"110010010",
  23023=>"100011001",
  23024=>"111011010",
  23025=>"011000100",
  23026=>"100010100",
  23027=>"000000100",
  23028=>"101110100",
  23029=>"000100100",
  23030=>"010101001",
  23031=>"001111001",
  23032=>"011010000",
  23033=>"100110100",
  23034=>"110010011",
  23035=>"110010111",
  23036=>"000001010",
  23037=>"111100001",
  23038=>"000011011",
  23039=>"011011111",
  23040=>"001110010",
  23041=>"110100100",
  23042=>"011000001",
  23043=>"000011111",
  23044=>"110100010",
  23045=>"101010011",
  23046=>"110111110",
  23047=>"110011100",
  23048=>"011000111",
  23049=>"011101111",
  23050=>"000100111",
  23051=>"001010001",
  23052=>"100000111",
  23053=>"110110000",
  23054=>"001110110",
  23055=>"010000110",
  23056=>"010110000",
  23057=>"001111101",
  23058=>"000000111",
  23059=>"100100011",
  23060=>"000111010",
  23061=>"001001010",
  23062=>"000000011",
  23063=>"101110100",
  23064=>"000101010",
  23065=>"111100000",
  23066=>"110100001",
  23067=>"010000001",
  23068=>"000010010",
  23069=>"000000111",
  23070=>"101111100",
  23071=>"100100110",
  23072=>"100010100",
  23073=>"010010000",
  23074=>"110010000",
  23075=>"101000000",
  23076=>"100010010",
  23077=>"100110100",
  23078=>"001101000",
  23079=>"101000101",
  23080=>"111101001",
  23081=>"001100000",
  23082=>"010011011",
  23083=>"100011010",
  23084=>"101111000",
  23085=>"011110001",
  23086=>"110110100",
  23087=>"000010000",
  23088=>"110001101",
  23089=>"101000010",
  23090=>"100110000",
  23091=>"111111011",
  23092=>"000101101",
  23093=>"011010000",
  23094=>"111100011",
  23095=>"100001111",
  23096=>"111011010",
  23097=>"001000111",
  23098=>"000010100",
  23099=>"000111100",
  23100=>"000001011",
  23101=>"000101001",
  23102=>"111001010",
  23103=>"001111110",
  23104=>"011100101",
  23105=>"010101001",
  23106=>"011100011",
  23107=>"010010011",
  23108=>"100001011",
  23109=>"000000100",
  23110=>"000101011",
  23111=>"000000001",
  23112=>"100110000",
  23113=>"001101010",
  23114=>"010101010",
  23115=>"100001001",
  23116=>"001111010",
  23117=>"011101010",
  23118=>"000010111",
  23119=>"001001100",
  23120=>"110100100",
  23121=>"011110001",
  23122=>"111100001",
  23123=>"000111110",
  23124=>"010011000",
  23125=>"001010001",
  23126=>"010000000",
  23127=>"000001101",
  23128=>"000000100",
  23129=>"101010111",
  23130=>"111001001",
  23131=>"001110110",
  23132=>"111100011",
  23133=>"101001011",
  23134=>"000111100",
  23135=>"110011010",
  23136=>"100011011",
  23137=>"111001000",
  23138=>"101101100",
  23139=>"101010000",
  23140=>"101110001",
  23141=>"101111011",
  23142=>"110011010",
  23143=>"000000110",
  23144=>"000001001",
  23145=>"110110101",
  23146=>"001111011",
  23147=>"111101001",
  23148=>"100000101",
  23149=>"110100100",
  23150=>"100011010",
  23151=>"001100011",
  23152=>"001001001",
  23153=>"111001010",
  23154=>"011000000",
  23155=>"101000110",
  23156=>"110011010",
  23157=>"011111100",
  23158=>"110000011",
  23159=>"010100101",
  23160=>"100001101",
  23161=>"110010000",
  23162=>"100001111",
  23163=>"110011110",
  23164=>"111111010",
  23165=>"010010101",
  23166=>"001001110",
  23167=>"111001100",
  23168=>"101101011",
  23169=>"111000010",
  23170=>"110101110",
  23171=>"100110111",
  23172=>"111000011",
  23173=>"010101100",
  23174=>"101111111",
  23175=>"011010110",
  23176=>"001010101",
  23177=>"001010101",
  23178=>"101100011",
  23179=>"011011110",
  23180=>"001111110",
  23181=>"111111110",
  23182=>"111111110",
  23183=>"010101110",
  23184=>"000010001",
  23185=>"110001001",
  23186=>"100010010",
  23187=>"000101011",
  23188=>"010010011",
  23189=>"110100000",
  23190=>"110001011",
  23191=>"010100101",
  23192=>"100110110",
  23193=>"011011111",
  23194=>"011011111",
  23195=>"100100001",
  23196=>"010100101",
  23197=>"000011111",
  23198=>"010011000",
  23199=>"000000100",
  23200=>"011001100",
  23201=>"000111110",
  23202=>"000010111",
  23203=>"111111011",
  23204=>"000001010",
  23205=>"000010100",
  23206=>"101011111",
  23207=>"000001010",
  23208=>"100111001",
  23209=>"110101110",
  23210=>"000110001",
  23211=>"001010111",
  23212=>"011001001",
  23213=>"110111010",
  23214=>"101101001",
  23215=>"000000101",
  23216=>"110111101",
  23217=>"000110110",
  23218=>"011101000",
  23219=>"101110100",
  23220=>"000111001",
  23221=>"010101000",
  23222=>"001000111",
  23223=>"011001100",
  23224=>"101001001",
  23225=>"011100110",
  23226=>"100100110",
  23227=>"100101101",
  23228=>"000111001",
  23229=>"110111000",
  23230=>"101110011",
  23231=>"101000111",
  23232=>"000010111",
  23233=>"001011011",
  23234=>"100000110",
  23235=>"001010000",
  23236=>"000011000",
  23237=>"111110110",
  23238=>"110100100",
  23239=>"100101011",
  23240=>"100001110",
  23241=>"000100100",
  23242=>"100011010",
  23243=>"010110010",
  23244=>"010110101",
  23245=>"011011110",
  23246=>"110001001",
  23247=>"100001011",
  23248=>"010100101",
  23249=>"000110010",
  23250=>"001110110",
  23251=>"110000110",
  23252=>"101001101",
  23253=>"001101101",
  23254=>"101011000",
  23255=>"111111100",
  23256=>"000011100",
  23257=>"100110011",
  23258=>"110110011",
  23259=>"000010001",
  23260=>"001011011",
  23261=>"111010000",
  23262=>"111110010",
  23263=>"000110110",
  23264=>"101010011",
  23265=>"000001011",
  23266=>"111110011",
  23267=>"001111000",
  23268=>"110011101",
  23269=>"100110111",
  23270=>"010001011",
  23271=>"001010100",
  23272=>"100110111",
  23273=>"110110100",
  23274=>"100000011",
  23275=>"000010100",
  23276=>"011111100",
  23277=>"100001001",
  23278=>"001011001",
  23279=>"111101111",
  23280=>"011001101",
  23281=>"010011110",
  23282=>"100110010",
  23283=>"110011111",
  23284=>"010010011",
  23285=>"101000010",
  23286=>"100011011",
  23287=>"101110010",
  23288=>"010111111",
  23289=>"011000011",
  23290=>"111111000",
  23291=>"110010010",
  23292=>"001000011",
  23293=>"001011100",
  23294=>"111010000",
  23295=>"111000111",
  23296=>"000011110",
  23297=>"011100011",
  23298=>"100110010",
  23299=>"100010010",
  23300=>"101011101",
  23301=>"110100000",
  23302=>"010111100",
  23303=>"000011000",
  23304=>"110100001",
  23305=>"100101110",
  23306=>"000101111",
  23307=>"011100001",
  23308=>"111001110",
  23309=>"001110011",
  23310=>"110100000",
  23311=>"101100011",
  23312=>"010101111",
  23313=>"100010100",
  23314=>"111011000",
  23315=>"000110001",
  23316=>"011111001",
  23317=>"000100001",
  23318=>"011000100",
  23319=>"001100000",
  23320=>"110110110",
  23321=>"001001011",
  23322=>"010101000",
  23323=>"100101011",
  23324=>"100000011",
  23325=>"101011011",
  23326=>"101010111",
  23327=>"001110001",
  23328=>"000000110",
  23329=>"111010011",
  23330=>"001001101",
  23331=>"001100010",
  23332=>"011100100",
  23333=>"111100101",
  23334=>"001010101",
  23335=>"100010010",
  23336=>"100001001",
  23337=>"011100101",
  23338=>"001001101",
  23339=>"110010010",
  23340=>"011101111",
  23341=>"100010000",
  23342=>"100101011",
  23343=>"000101101",
  23344=>"001001111",
  23345=>"001100100",
  23346=>"101010110",
  23347=>"011011111",
  23348=>"111001000",
  23349=>"101110100",
  23350=>"101000010",
  23351=>"100110000",
  23352=>"011001001",
  23353=>"000000101",
  23354=>"100000000",
  23355=>"000100010",
  23356=>"000010101",
  23357=>"101111111",
  23358=>"000000111",
  23359=>"101010101",
  23360=>"111001010",
  23361=>"111010101",
  23362=>"011010111",
  23363=>"001110101",
  23364=>"100110101",
  23365=>"110011011",
  23366=>"010111101",
  23367=>"111000101",
  23368=>"111111100",
  23369=>"101001100",
  23370=>"111110100",
  23371=>"101010001",
  23372=>"101000010",
  23373=>"110000101",
  23374=>"000110100",
  23375=>"111110110",
  23376=>"110011110",
  23377=>"111111110",
  23378=>"001110010",
  23379=>"010100011",
  23380=>"001100010",
  23381=>"101011111",
  23382=>"011100101",
  23383=>"001100101",
  23384=>"000001101",
  23385=>"100011100",
  23386=>"101100100",
  23387=>"000101101",
  23388=>"000010011",
  23389=>"000001000",
  23390=>"100100110",
  23391=>"010001100",
  23392=>"010011000",
  23393=>"011011110",
  23394=>"100001110",
  23395=>"101001000",
  23396=>"011000101",
  23397=>"111100110",
  23398=>"101000001",
  23399=>"110010100",
  23400=>"100101000",
  23401=>"001110010",
  23402=>"010011011",
  23403=>"111101000",
  23404=>"010010000",
  23405=>"011001001",
  23406=>"110100001",
  23407=>"011110100",
  23408=>"000011001",
  23409=>"111111000",
  23410=>"010100111",
  23411=>"011011010",
  23412=>"110011000",
  23413=>"011000010",
  23414=>"110110111",
  23415=>"101001011",
  23416=>"000111011",
  23417=>"111000100",
  23418=>"110110111",
  23419=>"001100111",
  23420=>"000000011",
  23421=>"100000000",
  23422=>"110110010",
  23423=>"010011101",
  23424=>"110111111",
  23425=>"111010110",
  23426=>"110001000",
  23427=>"010111100",
  23428=>"001110100",
  23429=>"011001011",
  23430=>"000111111",
  23431=>"001111010",
  23432=>"011110001",
  23433=>"011010001",
  23434=>"010110000",
  23435=>"011000110",
  23436=>"001000010",
  23437=>"010110001",
  23438=>"010010010",
  23439=>"110000100",
  23440=>"100111001",
  23441=>"001011110",
  23442=>"000101111",
  23443=>"000101110",
  23444=>"101011010",
  23445=>"100011011",
  23446=>"000110000",
  23447=>"100100001",
  23448=>"111011011",
  23449=>"000101100",
  23450=>"001100100",
  23451=>"101100101",
  23452=>"000000100",
  23453=>"111001010",
  23454=>"000100001",
  23455=>"110000011",
  23456=>"111000100",
  23457=>"110100111",
  23458=>"000110001",
  23459=>"111000111",
  23460=>"000001011",
  23461=>"111110011",
  23462=>"110011110",
  23463=>"011110101",
  23464=>"100101111",
  23465=>"010100110",
  23466=>"111101111",
  23467=>"111000100",
  23468=>"011001110",
  23469=>"100110110",
  23470=>"011110011",
  23471=>"011001011",
  23472=>"011100111",
  23473=>"101000110",
  23474=>"000001011",
  23475=>"101100000",
  23476=>"011010111",
  23477=>"010000010",
  23478=>"010110011",
  23479=>"101111100",
  23480=>"010100111",
  23481=>"010110110",
  23482=>"001010111",
  23483=>"110011100",
  23484=>"011101010",
  23485=>"010100100",
  23486=>"111111110",
  23487=>"110100000",
  23488=>"110011011",
  23489=>"011111100",
  23490=>"010001000",
  23491=>"001000000",
  23492=>"001011100",
  23493=>"111010001",
  23494=>"111000000",
  23495=>"110011110",
  23496=>"000000100",
  23497=>"010111110",
  23498=>"111010111",
  23499=>"011110011",
  23500=>"100001000",
  23501=>"010000111",
  23502=>"001100001",
  23503=>"010011010",
  23504=>"000100011",
  23505=>"000010111",
  23506=>"011001000",
  23507=>"011010010",
  23508=>"111000101",
  23509=>"100111111",
  23510=>"000111111",
  23511=>"101100110",
  23512=>"001100011",
  23513=>"101110111",
  23514=>"110100001",
  23515=>"111011011",
  23516=>"111001100",
  23517=>"000111011",
  23518=>"111011000",
  23519=>"000111000",
  23520=>"010000010",
  23521=>"101011001",
  23522=>"101000000",
  23523=>"010000100",
  23524=>"000110000",
  23525=>"000001000",
  23526=>"001111101",
  23527=>"011000100",
  23528=>"110001000",
  23529=>"010111011",
  23530=>"100110011",
  23531=>"100101010",
  23532=>"111100011",
  23533=>"011110001",
  23534=>"111000001",
  23535=>"000100010",
  23536=>"001001110",
  23537=>"111100011",
  23538=>"001010000",
  23539=>"000100101",
  23540=>"100100010",
  23541=>"011000001",
  23542=>"100110011",
  23543=>"110001011",
  23544=>"010101111",
  23545=>"111100101",
  23546=>"001010110",
  23547=>"001111000",
  23548=>"100111110",
  23549=>"111101101",
  23550=>"010110111",
  23551=>"010110100",
  23552=>"101010111",
  23553=>"001000001",
  23554=>"110010101",
  23555=>"101011100",
  23556=>"100110101",
  23557=>"111101010",
  23558=>"011011101",
  23559=>"000110111",
  23560=>"111011011",
  23561=>"011100111",
  23562=>"000111100",
  23563=>"011111110",
  23564=>"001100100",
  23565=>"001101100",
  23566=>"001100110",
  23567=>"011110011",
  23568=>"001011111",
  23569=>"101110101",
  23570=>"110110100",
  23571=>"011111110",
  23572=>"000111110",
  23573=>"001101101",
  23574=>"001000000",
  23575=>"111001100",
  23576=>"110010011",
  23577=>"101010001",
  23578=>"001100111",
  23579=>"111001010",
  23580=>"111011000",
  23581=>"001100111",
  23582=>"010101000",
  23583=>"001111101",
  23584=>"001110000",
  23585=>"010111001",
  23586=>"110001000",
  23587=>"101010010",
  23588=>"101101101",
  23589=>"110111110",
  23590=>"111010010",
  23591=>"001011000",
  23592=>"001010100",
  23593=>"100011011",
  23594=>"111111001",
  23595=>"011110111",
  23596=>"100000001",
  23597=>"001110100",
  23598=>"111010000",
  23599=>"000001011",
  23600=>"100100000",
  23601=>"101011111",
  23602=>"000100111",
  23603=>"110011111",
  23604=>"110000011",
  23605=>"001111000",
  23606=>"001011000",
  23607=>"111111111",
  23608=>"100001001",
  23609=>"001010111",
  23610=>"010111110",
  23611=>"100100111",
  23612=>"110010010",
  23613=>"111110100",
  23614=>"001100111",
  23615=>"100000111",
  23616=>"011001111",
  23617=>"000110100",
  23618=>"011110110",
  23619=>"101111101",
  23620=>"000111110",
  23621=>"100010001",
  23622=>"101100111",
  23623=>"111110001",
  23624=>"110010100",
  23625=>"101101000",
  23626=>"111101111",
  23627=>"010011010",
  23628=>"111111101",
  23629=>"111101110",
  23630=>"001010010",
  23631=>"010101000",
  23632=>"101111111",
  23633=>"101111100",
  23634=>"000110111",
  23635=>"100010110",
  23636=>"011001001",
  23637=>"111000111",
  23638=>"000101101",
  23639=>"010000100",
  23640=>"101000011",
  23641=>"011100001",
  23642=>"101101111",
  23643=>"100000011",
  23644=>"100111111",
  23645=>"111011100",
  23646=>"110111000",
  23647=>"110111100",
  23648=>"111011100",
  23649=>"110000110",
  23650=>"101110001",
  23651=>"100111111",
  23652=>"011101000",
  23653=>"101110111",
  23654=>"110000000",
  23655=>"010011100",
  23656=>"101101001",
  23657=>"110100111",
  23658=>"100010001",
  23659=>"000111011",
  23660=>"001001111",
  23661=>"001101000",
  23662=>"000111001",
  23663=>"000110101",
  23664=>"010011100",
  23665=>"110110111",
  23666=>"001100000",
  23667=>"111100100",
  23668=>"011010010",
  23669=>"011011110",
  23670=>"010110111",
  23671=>"110101100",
  23672=>"000011010",
  23673=>"010011000",
  23674=>"111000111",
  23675=>"000100110",
  23676=>"111010010",
  23677=>"100111111",
  23678=>"100110111",
  23679=>"100110110",
  23680=>"001001101",
  23681=>"101010101",
  23682=>"001100001",
  23683=>"111100110",
  23684=>"000000110",
  23685=>"100001001",
  23686=>"100101000",
  23687=>"100111001",
  23688=>"111111000",
  23689=>"111110100",
  23690=>"101011111",
  23691=>"110000010",
  23692=>"111011000",
  23693=>"000101101",
  23694=>"110000111",
  23695=>"011110001",
  23696=>"000011111",
  23697=>"000011100",
  23698=>"110100011",
  23699=>"001000001",
  23700=>"110110010",
  23701=>"011001101",
  23702=>"000011011",
  23703=>"000111110",
  23704=>"010111000",
  23705=>"100111010",
  23706=>"101100001",
  23707=>"101000000",
  23708=>"110101000",
  23709=>"100101111",
  23710=>"110111110",
  23711=>"010010111",
  23712=>"011000110",
  23713=>"011011001",
  23714=>"110110000",
  23715=>"011000011",
  23716=>"001010011",
  23717=>"000101010",
  23718=>"101111011",
  23719=>"110111000",
  23720=>"000010110",
  23721=>"010100111",
  23722=>"110010001",
  23723=>"101010001",
  23724=>"110100000",
  23725=>"011011011",
  23726=>"011111011",
  23727=>"101001101",
  23728=>"101110101",
  23729=>"101111111",
  23730=>"001011000",
  23731=>"101100101",
  23732=>"011000101",
  23733=>"010011110",
  23734=>"111010110",
  23735=>"110100011",
  23736=>"110110111",
  23737=>"000101001",
  23738=>"110110001",
  23739=>"110001000",
  23740=>"001100010",
  23741=>"001100000",
  23742=>"100001000",
  23743=>"111001001",
  23744=>"000100110",
  23745=>"000010110",
  23746=>"111101011",
  23747=>"111000000",
  23748=>"110110010",
  23749=>"001110011",
  23750=>"110011000",
  23751=>"101110011",
  23752=>"111100101",
  23753=>"010000001",
  23754=>"011011011",
  23755=>"110101100",
  23756=>"110100100",
  23757=>"000100010",
  23758=>"101000001",
  23759=>"001000100",
  23760=>"101000111",
  23761=>"101110110",
  23762=>"001111111",
  23763=>"010011011",
  23764=>"000001101",
  23765=>"110101100",
  23766=>"111111100",
  23767=>"001111010",
  23768=>"010011110",
  23769=>"000011011",
  23770=>"101100001",
  23771=>"001010111",
  23772=>"110010100",
  23773=>"000001101",
  23774=>"001100100",
  23775=>"000011001",
  23776=>"001000101",
  23777=>"111110000",
  23778=>"100101010",
  23779=>"101101110",
  23780=>"101000010",
  23781=>"011111000",
  23782=>"111110000",
  23783=>"011101000",
  23784=>"010110001",
  23785=>"000001010",
  23786=>"000101110",
  23787=>"100010001",
  23788=>"000000011",
  23789=>"101010000",
  23790=>"000011111",
  23791=>"100100111",
  23792=>"111011010",
  23793=>"001101000",
  23794=>"000101101",
  23795=>"110100011",
  23796=>"011001010",
  23797=>"101000110",
  23798=>"000000111",
  23799=>"101101111",
  23800=>"000010001",
  23801=>"010101101",
  23802=>"010000101",
  23803=>"001110010",
  23804=>"110010100",
  23805=>"000110001",
  23806=>"110000111",
  23807=>"000010001",
  23808=>"011100011",
  23809=>"111111011",
  23810=>"011011110",
  23811=>"001111001",
  23812=>"011100110",
  23813=>"011011010",
  23814=>"100011100",
  23815=>"111110010",
  23816=>"110111010",
  23817=>"001110010",
  23818=>"111100010",
  23819=>"011111101",
  23820=>"010101101",
  23821=>"000000111",
  23822=>"100010101",
  23823=>"100001110",
  23824=>"000010010",
  23825=>"110001111",
  23826=>"111111111",
  23827=>"100111010",
  23828=>"100011101",
  23829=>"111000001",
  23830=>"000101101",
  23831=>"101011001",
  23832=>"111100111",
  23833=>"000100010",
  23834=>"010100000",
  23835=>"110010011",
  23836=>"101010100",
  23837=>"110111110",
  23838=>"011000101",
  23839=>"000110101",
  23840=>"011110100",
  23841=>"000010100",
  23842=>"000001111",
  23843=>"110001011",
  23844=>"101110000",
  23845=>"000100001",
  23846=>"000010000",
  23847=>"010101100",
  23848=>"010010111",
  23849=>"001111111",
  23850=>"110001111",
  23851=>"011010110",
  23852=>"000100000",
  23853=>"110001010",
  23854=>"101101101",
  23855=>"111111100",
  23856=>"110100101",
  23857=>"101101110",
  23858=>"000110110",
  23859=>"111110010",
  23860=>"110101011",
  23861=>"011110011",
  23862=>"110110010",
  23863=>"011000100",
  23864=>"000011001",
  23865=>"001100010",
  23866=>"110101110",
  23867=>"110000010",
  23868=>"010011110",
  23869=>"101011011",
  23870=>"100010011",
  23871=>"101001001",
  23872=>"001011011",
  23873=>"010010010",
  23874=>"101101101",
  23875=>"110100000",
  23876=>"010110000",
  23877=>"110110001",
  23878=>"010011001",
  23879=>"110110110",
  23880=>"110111010",
  23881=>"111110101",
  23882=>"110001110",
  23883=>"100000001",
  23884=>"001011100",
  23885=>"111100000",
  23886=>"100001000",
  23887=>"010111110",
  23888=>"010010100",
  23889=>"111000101",
  23890=>"111100010",
  23891=>"110001100",
  23892=>"000001010",
  23893=>"011111111",
  23894=>"011000110",
  23895=>"111010001",
  23896=>"000011000",
  23897=>"001100111",
  23898=>"101001000",
  23899=>"000100111",
  23900=>"100000101",
  23901=>"000000110",
  23902=>"000011111",
  23903=>"100111111",
  23904=>"001111010",
  23905=>"001110101",
  23906=>"011011110",
  23907=>"001111110",
  23908=>"111100111",
  23909=>"110111111",
  23910=>"110010001",
  23911=>"000001011",
  23912=>"100001010",
  23913=>"110111101",
  23914=>"010000110",
  23915=>"100101111",
  23916=>"101010000",
  23917=>"000011010",
  23918=>"100100011",
  23919=>"110101000",
  23920=>"110101011",
  23921=>"100011011",
  23922=>"110000100",
  23923=>"101011000",
  23924=>"101001101",
  23925=>"010110101",
  23926=>"101010011",
  23927=>"100001110",
  23928=>"101001100",
  23929=>"010010000",
  23930=>"000000001",
  23931=>"000000000",
  23932=>"010000001",
  23933=>"001010010",
  23934=>"101100110",
  23935=>"100101101",
  23936=>"110111110",
  23937=>"111111010",
  23938=>"001000000",
  23939=>"001000011",
  23940=>"110111000",
  23941=>"000111010",
  23942=>"000101101",
  23943=>"110010101",
  23944=>"011100100",
  23945=>"110100001",
  23946=>"010010101",
  23947=>"010001000",
  23948=>"111100001",
  23949=>"000011101",
  23950=>"001110011",
  23951=>"000011110",
  23952=>"010000011",
  23953=>"010100101",
  23954=>"100001000",
  23955=>"001000011",
  23956=>"011011001",
  23957=>"111100010",
  23958=>"101001110",
  23959=>"010000011",
  23960=>"100100111",
  23961=>"100001110",
  23962=>"111111001",
  23963=>"000111101",
  23964=>"101000100",
  23965=>"100111110",
  23966=>"011100001",
  23967=>"011000010",
  23968=>"110100100",
  23969=>"011111011",
  23970=>"101000000",
  23971=>"110111010",
  23972=>"100011110",
  23973=>"100110001",
  23974=>"010000110",
  23975=>"011111110",
  23976=>"111100010",
  23977=>"000100101",
  23978=>"010100111",
  23979=>"000111110",
  23980=>"110100001",
  23981=>"111101100",
  23982=>"111110000",
  23983=>"010000001",
  23984=>"000010111",
  23985=>"111111110",
  23986=>"111010001",
  23987=>"101110111",
  23988=>"111101111",
  23989=>"100000100",
  23990=>"100111110",
  23991=>"100101010",
  23992=>"001010110",
  23993=>"111000011",
  23994=>"101100010",
  23995=>"101001001",
  23996=>"101101000",
  23997=>"001010010",
  23998=>"010010010",
  23999=>"011100010",
  24000=>"100100110",
  24001=>"010100100",
  24002=>"000101100",
  24003=>"100000011",
  24004=>"111111111",
  24005=>"111100101",
  24006=>"101100000",
  24007=>"110111111",
  24008=>"010100101",
  24009=>"010111110",
  24010=>"111111110",
  24011=>"101100011",
  24012=>"000010111",
  24013=>"100100100",
  24014=>"101011110",
  24015=>"010011001",
  24016=>"010000010",
  24017=>"101011111",
  24018=>"110001001",
  24019=>"011110100",
  24020=>"000100001",
  24021=>"111111111",
  24022=>"011000110",
  24023=>"111011011",
  24024=>"110111000",
  24025=>"111101001",
  24026=>"111110001",
  24027=>"100100111",
  24028=>"000000010",
  24029=>"110000100",
  24030=>"001001000",
  24031=>"101110111",
  24032=>"010011110",
  24033=>"110111111",
  24034=>"101110111",
  24035=>"111110111",
  24036=>"110101101",
  24037=>"010000001",
  24038=>"110111100",
  24039=>"010101010",
  24040=>"011101010",
  24041=>"110000000",
  24042=>"110110111",
  24043=>"010000000",
  24044=>"100101110",
  24045=>"001010100",
  24046=>"101011111",
  24047=>"111110100",
  24048=>"000000000",
  24049=>"101111100",
  24050=>"010001010",
  24051=>"001110111",
  24052=>"010110010",
  24053=>"011111110",
  24054=>"010101000",
  24055=>"111011001",
  24056=>"110111100",
  24057=>"111101011",
  24058=>"111111101",
  24059=>"000111000",
  24060=>"100010011",
  24061=>"110111011",
  24062=>"101000001",
  24063=>"110000110",
  24064=>"010110001",
  24065=>"010001111",
  24066=>"100001110",
  24067=>"100011011",
  24068=>"000111100",
  24069=>"101010101",
  24070=>"011010010",
  24071=>"011110111",
  24072=>"001100110",
  24073=>"101111111",
  24074=>"010001011",
  24075=>"010111101",
  24076=>"011001010",
  24077=>"101011011",
  24078=>"010101000",
  24079=>"010001011",
  24080=>"010010011",
  24081=>"111001101",
  24082=>"000101110",
  24083=>"011010100",
  24084=>"101011001",
  24085=>"100111111",
  24086=>"100100110",
  24087=>"000111111",
  24088=>"011011000",
  24089=>"001000001",
  24090=>"000101011",
  24091=>"100001100",
  24092=>"100011110",
  24093=>"000110011",
  24094=>"010100110",
  24095=>"111101101",
  24096=>"000101001",
  24097=>"000010011",
  24098=>"111111101",
  24099=>"011000110",
  24100=>"101110110",
  24101=>"011001101",
  24102=>"011101111",
  24103=>"011111101",
  24104=>"100001110",
  24105=>"101000001",
  24106=>"111111110",
  24107=>"100000001",
  24108=>"000011110",
  24109=>"000000100",
  24110=>"111111111",
  24111=>"001001010",
  24112=>"000010010",
  24113=>"010000011",
  24114=>"111100000",
  24115=>"000101011",
  24116=>"000100010",
  24117=>"100011010",
  24118=>"000111011",
  24119=>"110000001",
  24120=>"011101111",
  24121=>"100111010",
  24122=>"010000000",
  24123=>"000101000",
  24124=>"010110010",
  24125=>"111011100",
  24126=>"101101100",
  24127=>"110110101",
  24128=>"010110111",
  24129=>"100100010",
  24130=>"001010101",
  24131=>"000000110",
  24132=>"101111111",
  24133=>"011111010",
  24134=>"111010111",
  24135=>"101001111",
  24136=>"111110101",
  24137=>"101110001",
  24138=>"111110010",
  24139=>"010000110",
  24140=>"110101010",
  24141=>"101101110",
  24142=>"110010010",
  24143=>"001110100",
  24144=>"110110101",
  24145=>"010111110",
  24146=>"100011010",
  24147=>"110111011",
  24148=>"001111000",
  24149=>"111011001",
  24150=>"100111101",
  24151=>"100011111",
  24152=>"001001001",
  24153=>"011101100",
  24154=>"101100010",
  24155=>"010101001",
  24156=>"000100011",
  24157=>"010110111",
  24158=>"111011011",
  24159=>"101000111",
  24160=>"001001010",
  24161=>"000101001",
  24162=>"100001111",
  24163=>"001000101",
  24164=>"000001001",
  24165=>"000000001",
  24166=>"100100101",
  24167=>"101010111",
  24168=>"111110110",
  24169=>"001111111",
  24170=>"001000001",
  24171=>"100011111",
  24172=>"010010000",
  24173=>"001010000",
  24174=>"101101011",
  24175=>"101111100",
  24176=>"111111110",
  24177=>"010111001",
  24178=>"010011011",
  24179=>"101000000",
  24180=>"001100000",
  24181=>"110011111",
  24182=>"100011000",
  24183=>"100110011",
  24184=>"110100011",
  24185=>"001100000",
  24186=>"010000110",
  24187=>"001010010",
  24188=>"100110111",
  24189=>"000111101",
  24190=>"011011011",
  24191=>"010101010",
  24192=>"000010011",
  24193=>"101001101",
  24194=>"110100001",
  24195=>"101111000",
  24196=>"010010001",
  24197=>"100011111",
  24198=>"011001101",
  24199=>"110110100",
  24200=>"000111100",
  24201=>"101100010",
  24202=>"000100010",
  24203=>"000000100",
  24204=>"001111100",
  24205=>"010011111",
  24206=>"010101111",
  24207=>"001011011",
  24208=>"001100110",
  24209=>"011110001",
  24210=>"001101011",
  24211=>"011011100",
  24212=>"000111001",
  24213=>"110010100",
  24214=>"111101101",
  24215=>"000100110",
  24216=>"110111101",
  24217=>"100001011",
  24218=>"000110011",
  24219=>"100100011",
  24220=>"011111101",
  24221=>"101110100",
  24222=>"111000010",
  24223=>"100000101",
  24224=>"111100101",
  24225=>"011011111",
  24226=>"011110010",
  24227=>"011011100",
  24228=>"000100101",
  24229=>"001100011",
  24230=>"011101001",
  24231=>"101001001",
  24232=>"000000001",
  24233=>"101011011",
  24234=>"111110110",
  24235=>"001011101",
  24236=>"100010011",
  24237=>"110110110",
  24238=>"111110100",
  24239=>"010000001",
  24240=>"011001111",
  24241=>"111101101",
  24242=>"111110010",
  24243=>"110101011",
  24244=>"101110111",
  24245=>"101000000",
  24246=>"101111100",
  24247=>"001000011",
  24248=>"000101110",
  24249=>"011011001",
  24250=>"000011010",
  24251=>"111100100",
  24252=>"111001100",
  24253=>"100110100",
  24254=>"000101110",
  24255=>"110100111",
  24256=>"001100101",
  24257=>"000111101",
  24258=>"100111110",
  24259=>"000110100",
  24260=>"101100110",
  24261=>"111010110",
  24262=>"101010010",
  24263=>"111010010",
  24264=>"100111101",
  24265=>"100101110",
  24266=>"101011011",
  24267=>"101000000",
  24268=>"011110000",
  24269=>"110100111",
  24270=>"001111110",
  24271=>"001100001",
  24272=>"000111110",
  24273=>"110110011",
  24274=>"010111011",
  24275=>"010100100",
  24276=>"101111101",
  24277=>"110111010",
  24278=>"110101011",
  24279=>"111101111",
  24280=>"011010100",
  24281=>"000010001",
  24282=>"111110000",
  24283=>"111001010",
  24284=>"001011001",
  24285=>"110101010",
  24286=>"010010010",
  24287=>"110010100",
  24288=>"110111101",
  24289=>"000101110",
  24290=>"001111101",
  24291=>"001010000",
  24292=>"110111000",
  24293=>"001001011",
  24294=>"111110111",
  24295=>"110010110",
  24296=>"010011111",
  24297=>"111000001",
  24298=>"000001001",
  24299=>"001111110",
  24300=>"011101110",
  24301=>"101111111",
  24302=>"000111100",
  24303=>"010000000",
  24304=>"110011100",
  24305=>"011011010",
  24306=>"100110111",
  24307=>"111010111",
  24308=>"110011001",
  24309=>"000001010",
  24310=>"100001100",
  24311=>"000011001",
  24312=>"111010100",
  24313=>"000110001",
  24314=>"110001001",
  24315=>"111110100",
  24316=>"100111111",
  24317=>"001001111",
  24318=>"010110110",
  24319=>"010000101",
  24320=>"110000101",
  24321=>"110101001",
  24322=>"010001110",
  24323=>"010100000",
  24324=>"101111111",
  24325=>"111001111",
  24326=>"000101101",
  24327=>"100100110",
  24328=>"010101111",
  24329=>"100011101",
  24330=>"011000101",
  24331=>"001100100",
  24332=>"111001111",
  24333=>"000010011",
  24334=>"100010100",
  24335=>"101010000",
  24336=>"101100111",
  24337=>"001100101",
  24338=>"101001101",
  24339=>"101100010",
  24340=>"010011011",
  24341=>"000000010",
  24342=>"001110000",
  24343=>"111001001",
  24344=>"100100101",
  24345=>"100001100",
  24346=>"001111011",
  24347=>"110111110",
  24348=>"000001001",
  24349=>"001111100",
  24350=>"011101111",
  24351=>"011100001",
  24352=>"110110111",
  24353=>"000000111",
  24354=>"000010000",
  24355=>"000110010",
  24356=>"001001011",
  24357=>"110011100",
  24358=>"100100000",
  24359=>"101110101",
  24360=>"010100000",
  24361=>"100010011",
  24362=>"110110110",
  24363=>"001100001",
  24364=>"010010111",
  24365=>"100110111",
  24366=>"011111110",
  24367=>"111100001",
  24368=>"100011100",
  24369=>"110101010",
  24370=>"110001111",
  24371=>"101111000",
  24372=>"101010010",
  24373=>"101000010",
  24374=>"000000110",
  24375=>"001111001",
  24376=>"101101010",
  24377=>"101001010",
  24378=>"111111001",
  24379=>"010110001",
  24380=>"011001101",
  24381=>"111101100",
  24382=>"111110111",
  24383=>"010011001",
  24384=>"000001110",
  24385=>"110001111",
  24386=>"001000011",
  24387=>"000010000",
  24388=>"000011111",
  24389=>"010001001",
  24390=>"010011100",
  24391=>"100100010",
  24392=>"110011110",
  24393=>"001101111",
  24394=>"000011110",
  24395=>"010011000",
  24396=>"010110011",
  24397=>"100100010",
  24398=>"010111011",
  24399=>"101111010",
  24400=>"100100111",
  24401=>"111001011",
  24402=>"010111101",
  24403=>"111001111",
  24404=>"001010100",
  24405=>"000101000",
  24406=>"111100010",
  24407=>"000010110",
  24408=>"000010111",
  24409=>"111100111",
  24410=>"010101100",
  24411=>"111110101",
  24412=>"010111110",
  24413=>"101001111",
  24414=>"100101011",
  24415=>"110110111",
  24416=>"110111000",
  24417=>"011100101",
  24418=>"100100101",
  24419=>"011001000",
  24420=>"000000001",
  24421=>"100011111",
  24422=>"011111100",
  24423=>"010011000",
  24424=>"000111101",
  24425=>"110000010",
  24426=>"100001111",
  24427=>"011011011",
  24428=>"010101011",
  24429=>"111110000",
  24430=>"111111001",
  24431=>"000100001",
  24432=>"110110100",
  24433=>"010100100",
  24434=>"000001000",
  24435=>"100000101",
  24436=>"110101110",
  24437=>"111101001",
  24438=>"110111011",
  24439=>"011001101",
  24440=>"101111001",
  24441=>"010011000",
  24442=>"111001000",
  24443=>"010000110",
  24444=>"110100101",
  24445=>"000011000",
  24446=>"100110011",
  24447=>"110100010",
  24448=>"001001011",
  24449=>"000011111",
  24450=>"010111000",
  24451=>"111011100",
  24452=>"101111111",
  24453=>"101000101",
  24454=>"110011111",
  24455=>"001000101",
  24456=>"000001000",
  24457=>"011000001",
  24458=>"110110011",
  24459=>"000111000",
  24460=>"111111010",
  24461=>"010110001",
  24462=>"001010100",
  24463=>"100101000",
  24464=>"100110110",
  24465=>"000001110",
  24466=>"101010000",
  24467=>"110000010",
  24468=>"011101100",
  24469=>"100000100",
  24470=>"000010111",
  24471=>"000010000",
  24472=>"000101101",
  24473=>"000011111",
  24474=>"100001111",
  24475=>"001000010",
  24476=>"100011111",
  24477=>"111000011",
  24478=>"010111101",
  24479=>"000110100",
  24480=>"001010110",
  24481=>"000101011",
  24482=>"111011101",
  24483=>"001111011",
  24484=>"000100000",
  24485=>"100001111",
  24486=>"101111000",
  24487=>"001110001",
  24488=>"011101111",
  24489=>"110101110",
  24490=>"100010111",
  24491=>"111111000",
  24492=>"111010111",
  24493=>"000000100",
  24494=>"101100010",
  24495=>"000110001",
  24496=>"010011101",
  24497=>"110110110",
  24498=>"000010111",
  24499=>"110100011",
  24500=>"110000000",
  24501=>"111010000",
  24502=>"010000000",
  24503=>"110101110",
  24504=>"010001011",
  24505=>"011001010",
  24506=>"101010000",
  24507=>"110111011",
  24508=>"010100100",
  24509=>"110100010",
  24510=>"011110101",
  24511=>"110000000",
  24512=>"101111011",
  24513=>"011100011",
  24514=>"110001100",
  24515=>"011010011",
  24516=>"011000111",
  24517=>"000010000",
  24518=>"111011001",
  24519=>"111011111",
  24520=>"111010111",
  24521=>"001110010",
  24522=>"111101100",
  24523=>"000010011",
  24524=>"000111111",
  24525=>"111111111",
  24526=>"000110110",
  24527=>"011110011",
  24528=>"001110111",
  24529=>"010010011",
  24530=>"100110101",
  24531=>"000011111",
  24532=>"111111111",
  24533=>"000011010",
  24534=>"011010010",
  24535=>"010001010",
  24536=>"110111100",
  24537=>"100011100",
  24538=>"010001101",
  24539=>"101000010",
  24540=>"110101111",
  24541=>"101010001",
  24542=>"101110010",
  24543=>"110101100",
  24544=>"000111110",
  24545=>"100000010",
  24546=>"001011000",
  24547=>"010001110",
  24548=>"000111111",
  24549=>"001111010",
  24550=>"100100000",
  24551=>"110000110",
  24552=>"101010100",
  24553=>"110100100",
  24554=>"000000110",
  24555=>"011100000",
  24556=>"100010000",
  24557=>"111010110",
  24558=>"010111101",
  24559=>"110001100",
  24560=>"111010111",
  24561=>"011100111",
  24562=>"101001111",
  24563=>"001101110",
  24564=>"111011101",
  24565=>"011101110",
  24566=>"011111110",
  24567=>"101101111",
  24568=>"011010101",
  24569=>"110111111",
  24570=>"110101111",
  24571=>"101101000",
  24572=>"100010110",
  24573=>"100001111",
  24574=>"100000100",
  24575=>"011111001",
  24576=>"000111101",
  24577=>"010101010",
  24578=>"001110100",
  24579=>"110000111",
  24580=>"011111010",
  24581=>"001010100",
  24582=>"000010110",
  24583=>"100111101",
  24584=>"111111100",
  24585=>"110100000",
  24586=>"011100000",
  24587=>"111100000",
  24588=>"110110000",
  24589=>"100100101",
  24590=>"001001111",
  24591=>"001111010",
  24592=>"000100011",
  24593=>"010000100",
  24594=>"000000100",
  24595=>"000100101",
  24596=>"001110110",
  24597=>"000110010",
  24598=>"110100011",
  24599=>"111010101",
  24600=>"011110111",
  24601=>"011001001",
  24602=>"101000000",
  24603=>"001001000",
  24604=>"011001011",
  24605=>"110111011",
  24606=>"001110100",
  24607=>"010110000",
  24608=>"101111110",
  24609=>"010000110",
  24610=>"101010001",
  24611=>"111110100",
  24612=>"001011011",
  24613=>"011110011",
  24614=>"000000001",
  24615=>"010110010",
  24616=>"101101000",
  24617=>"000011111",
  24618=>"110101111",
  24619=>"101111010",
  24620=>"110001010",
  24621=>"010010101",
  24622=>"011101000",
  24623=>"110111011",
  24624=>"110010101",
  24625=>"011111110",
  24626=>"011110100",
  24627=>"000001000",
  24628=>"101010010",
  24629=>"011010111",
  24630=>"101011010",
  24631=>"100011000",
  24632=>"001011011",
  24633=>"000000100",
  24634=>"100100010",
  24635=>"000010000",
  24636=>"110011001",
  24637=>"110010011",
  24638=>"111000110",
  24639=>"110011001",
  24640=>"101101100",
  24641=>"010100100",
  24642=>"110000010",
  24643=>"001001111",
  24644=>"000100100",
  24645=>"111011010",
  24646=>"101010010",
  24647=>"000010111",
  24648=>"110011111",
  24649=>"010011010",
  24650=>"110111010",
  24651=>"000011000",
  24652=>"011101000",
  24653=>"010001000",
  24654=>"100010010",
  24655=>"100000110",
  24656=>"101001111",
  24657=>"001101001",
  24658=>"111101101",
  24659=>"101000110",
  24660=>"001011111",
  24661=>"100011110",
  24662=>"001010000",
  24663=>"011000000",
  24664=>"000010000",
  24665=>"001010100",
  24666=>"100011010",
  24667=>"000000100",
  24668=>"011010001",
  24669=>"000011100",
  24670=>"101101000",
  24671=>"111000000",
  24672=>"000110100",
  24673=>"010000001",
  24674=>"000010110",
  24675=>"001000011",
  24676=>"010100111",
  24677=>"000001011",
  24678=>"011011010",
  24679=>"000011000",
  24680=>"000110111",
  24681=>"001001100",
  24682=>"100100000",
  24683=>"011000001",
  24684=>"111101000",
  24685=>"100000011",
  24686=>"111011101",
  24687=>"111110111",
  24688=>"001000110",
  24689=>"110110100",
  24690=>"010111100",
  24691=>"000111111",
  24692=>"100100010",
  24693=>"000000100",
  24694=>"111101011",
  24695=>"100110110",
  24696=>"011000100",
  24697=>"111001101",
  24698=>"000011000",
  24699=>"101101111",
  24700=>"100000000",
  24701=>"110000100",
  24702=>"000010111",
  24703=>"000001010",
  24704=>"001101010",
  24705=>"111111000",
  24706=>"001010011",
  24707=>"000111010",
  24708=>"111110100",
  24709=>"001111110",
  24710=>"100101110",
  24711=>"011010011",
  24712=>"100000111",
  24713=>"011111101",
  24714=>"001010000",
  24715=>"111111111",
  24716=>"001010100",
  24717=>"000011100",
  24718=>"000000110",
  24719=>"110011010",
  24720=>"000111110",
  24721=>"110101101",
  24722=>"111010001",
  24723=>"100001111",
  24724=>"010001101",
  24725=>"000011101",
  24726=>"001000000",
  24727=>"000100110",
  24728=>"100100010",
  24729=>"100111110",
  24730=>"101111100",
  24731=>"101100111",
  24732=>"001000111",
  24733=>"100001111",
  24734=>"111100001",
  24735=>"110011001",
  24736=>"100101011",
  24737=>"100001100",
  24738=>"101000000",
  24739=>"101011000",
  24740=>"101000110",
  24741=>"110101110",
  24742=>"011111010",
  24743=>"000001001",
  24744=>"001110110",
  24745=>"101100011",
  24746=>"110000001",
  24747=>"011010111",
  24748=>"111101100",
  24749=>"110010110",
  24750=>"101000000",
  24751=>"001000011",
  24752=>"001101110",
  24753=>"101101000",
  24754=>"010101100",
  24755=>"101100110",
  24756=>"101001101",
  24757=>"010100010",
  24758=>"111101010",
  24759=>"000100000",
  24760=>"111111111",
  24761=>"111001010",
  24762=>"101000010",
  24763=>"100000011",
  24764=>"110111100",
  24765=>"111111110",
  24766=>"100011001",
  24767=>"001011000",
  24768=>"001000001",
  24769=>"010110110",
  24770=>"101011011",
  24771=>"110010101",
  24772=>"011111011",
  24773=>"100000001",
  24774=>"111000010",
  24775=>"101010010",
  24776=>"111111111",
  24777=>"010011111",
  24778=>"100011001",
  24779=>"011111101",
  24780=>"011100100",
  24781=>"110010010",
  24782=>"001000001",
  24783=>"000110000",
  24784=>"100101100",
  24785=>"010010101",
  24786=>"001010010",
  24787=>"000011011",
  24788=>"000100010",
  24789=>"001010010",
  24790=>"101101011",
  24791=>"100101001",
  24792=>"000101010",
  24793=>"010001011",
  24794=>"000010011",
  24795=>"111111000",
  24796=>"000111000",
  24797=>"110110100",
  24798=>"001001000",
  24799=>"010111111",
  24800=>"101111101",
  24801=>"100010111",
  24802=>"111110000",
  24803=>"000110110",
  24804=>"000101000",
  24805=>"001111110",
  24806=>"101001011",
  24807=>"000011111",
  24808=>"000011000",
  24809=>"100000001",
  24810=>"011110101",
  24811=>"000001110",
  24812=>"011000110",
  24813=>"010010100",
  24814=>"111111000",
  24815=>"101001010",
  24816=>"011101000",
  24817=>"011000100",
  24818=>"000011000",
  24819=>"000110000",
  24820=>"000101010",
  24821=>"000111000",
  24822=>"010011100",
  24823=>"110111111",
  24824=>"110000010",
  24825=>"101000110",
  24826=>"101101010",
  24827=>"111010111",
  24828=>"000101011",
  24829=>"001011111",
  24830=>"011101110",
  24831=>"000111111",
  24832=>"010011001",
  24833=>"101100001",
  24834=>"111010010",
  24835=>"001100000",
  24836=>"100010110",
  24837=>"000100000",
  24838=>"111110011",
  24839=>"110110001",
  24840=>"001101001",
  24841=>"100101101",
  24842=>"010110101",
  24843=>"100100001",
  24844=>"010001000",
  24845=>"010101010",
  24846=>"000001000",
  24847=>"101110110",
  24848=>"100100110",
  24849=>"110101010",
  24850=>"000001110",
  24851=>"010000100",
  24852=>"010110000",
  24853=>"101100110",
  24854=>"111011100",
  24855=>"101111001",
  24856=>"010100101",
  24857=>"101110110",
  24858=>"100110011",
  24859=>"110101011",
  24860=>"110100011",
  24861=>"101000110",
  24862=>"100100110",
  24863=>"111100101",
  24864=>"100011001",
  24865=>"111011001",
  24866=>"101111100",
  24867=>"000110000",
  24868=>"001001011",
  24869=>"001110110",
  24870=>"010111010",
  24871=>"101101111",
  24872=>"110011011",
  24873=>"000001110",
  24874=>"010110001",
  24875=>"010011100",
  24876=>"100001111",
  24877=>"010100011",
  24878=>"000000000",
  24879=>"010010001",
  24880=>"110111111",
  24881=>"011001100",
  24882=>"000010000",
  24883=>"010011001",
  24884=>"101011010",
  24885=>"010010110",
  24886=>"000011011",
  24887=>"001111001",
  24888=>"001000110",
  24889=>"110010011",
  24890=>"010101111",
  24891=>"101001100",
  24892=>"011010010",
  24893=>"101111011",
  24894=>"011101010",
  24895=>"011111001",
  24896=>"110001101",
  24897=>"100011000",
  24898=>"101010111",
  24899=>"001000101",
  24900=>"101010101",
  24901=>"100101100",
  24902=>"000111101",
  24903=>"010010011",
  24904=>"111110110",
  24905=>"000101101",
  24906=>"001011000",
  24907=>"000010001",
  24908=>"010011000",
  24909=>"100101110",
  24910=>"010101000",
  24911=>"011010100",
  24912=>"011011100",
  24913=>"011101000",
  24914=>"000010011",
  24915=>"000001110",
  24916=>"100101100",
  24917=>"100100010",
  24918=>"011000001",
  24919=>"000100100",
  24920=>"101110001",
  24921=>"111110101",
  24922=>"110101110",
  24923=>"010100000",
  24924=>"000101011",
  24925=>"110011100",
  24926=>"001000111",
  24927=>"010001001",
  24928=>"111001011",
  24929=>"000000000",
  24930=>"111101000",
  24931=>"100101111",
  24932=>"010110001",
  24933=>"010101101",
  24934=>"100101111",
  24935=>"000000011",
  24936=>"110111100",
  24937=>"100111101",
  24938=>"110101100",
  24939=>"111110000",
  24940=>"100111010",
  24941=>"110100011",
  24942=>"110010111",
  24943=>"111110110",
  24944=>"001000001",
  24945=>"101101110",
  24946=>"100001100",
  24947=>"011010001",
  24948=>"111110101",
  24949=>"100111001",
  24950=>"111100110",
  24951=>"010110011",
  24952=>"111100101",
  24953=>"000111111",
  24954=>"010010100",
  24955=>"100111011",
  24956=>"000000000",
  24957=>"010011000",
  24958=>"111010000",
  24959=>"111111011",
  24960=>"010010011",
  24961=>"001111010",
  24962=>"100110011",
  24963=>"011100011",
  24964=>"000111100",
  24965=>"010100010",
  24966=>"100001110",
  24967=>"101100001",
  24968=>"101100111",
  24969=>"001111110",
  24970=>"000100010",
  24971=>"010000001",
  24972=>"001101110",
  24973=>"001010001",
  24974=>"100110001",
  24975=>"110110011",
  24976=>"001111111",
  24977=>"111001000",
  24978=>"010011011",
  24979=>"000000101",
  24980=>"000000111",
  24981=>"101111110",
  24982=>"001011100",
  24983=>"100111010",
  24984=>"110010101",
  24985=>"010000001",
  24986=>"100110011",
  24987=>"111000000",
  24988=>"000010111",
  24989=>"011010010",
  24990=>"011010101",
  24991=>"110100101",
  24992=>"111001010",
  24993=>"101101111",
  24994=>"011110100",
  24995=>"001101110",
  24996=>"001011000",
  24997=>"011111111",
  24998=>"000101000",
  24999=>"111001110",
  25000=>"101001000",
  25001=>"001000110",
  25002=>"100111111",
  25003=>"011111010",
  25004=>"110000101",
  25005=>"000001100",
  25006=>"010000111",
  25007=>"111010111",
  25008=>"001110000",
  25009=>"010101001",
  25010=>"111111010",
  25011=>"101011001",
  25012=>"001110111",
  25013=>"110101011",
  25014=>"100111100",
  25015=>"100011100",
  25016=>"111111011",
  25017=>"111001111",
  25018=>"101011101",
  25019=>"011010011",
  25020=>"000010001",
  25021=>"000111111",
  25022=>"111011001",
  25023=>"000111001",
  25024=>"001001101",
  25025=>"111000010",
  25026=>"110010110",
  25027=>"000111001",
  25028=>"001011000",
  25029=>"000101001",
  25030=>"011101110",
  25031=>"101001000",
  25032=>"011111110",
  25033=>"111111011",
  25034=>"100000111",
  25035=>"001100000",
  25036=>"101010010",
  25037=>"111000100",
  25038=>"010001101",
  25039=>"000110010",
  25040=>"111110011",
  25041=>"111001001",
  25042=>"000011001",
  25043=>"010101010",
  25044=>"011100100",
  25045=>"011000001",
  25046=>"000111110",
  25047=>"100000001",
  25048=>"111001101",
  25049=>"010110001",
  25050=>"101111100",
  25051=>"111000110",
  25052=>"101100101",
  25053=>"000100100",
  25054=>"000011111",
  25055=>"110000101",
  25056=>"000000011",
  25057=>"100011000",
  25058=>"010011001",
  25059=>"111111111",
  25060=>"001000101",
  25061=>"111011000",
  25062=>"011110100",
  25063=>"100000001",
  25064=>"101100100",
  25065=>"010101000",
  25066=>"110000001",
  25067=>"110000000",
  25068=>"111101111",
  25069=>"101101000",
  25070=>"110111111",
  25071=>"010000010",
  25072=>"000011111",
  25073=>"011100000",
  25074=>"000001010",
  25075=>"001100100",
  25076=>"001111001",
  25077=>"110010001",
  25078=>"001011001",
  25079=>"001110000",
  25080=>"000011001",
  25081=>"001101001",
  25082=>"011000011",
  25083=>"001111111",
  25084=>"101000110",
  25085=>"110001011",
  25086=>"011011100",
  25087=>"111001001",
  25088=>"001001010",
  25089=>"001011111",
  25090=>"110001011",
  25091=>"000010111",
  25092=>"100000001",
  25093=>"111000011",
  25094=>"001001101",
  25095=>"100001001",
  25096=>"100100011",
  25097=>"101101101",
  25098=>"111010110",
  25099=>"101100110",
  25100=>"000000100",
  25101=>"111001010",
  25102=>"010100011",
  25103=>"110000001",
  25104=>"111010111",
  25105=>"110000010",
  25106=>"110000100",
  25107=>"110000101",
  25108=>"001100001",
  25109=>"111100110",
  25110=>"111010001",
  25111=>"000000001",
  25112=>"011100011",
  25113=>"010011010",
  25114=>"001111011",
  25115=>"000000100",
  25116=>"001111110",
  25117=>"110000101",
  25118=>"000011110",
  25119=>"110101111",
  25120=>"001001001",
  25121=>"110011111",
  25122=>"000010000",
  25123=>"101001000",
  25124=>"101111111",
  25125=>"000101001",
  25126=>"010000011",
  25127=>"110110001",
  25128=>"000111001",
  25129=>"100011110",
  25130=>"001101000",
  25131=>"100110011",
  25132=>"110111110",
  25133=>"010010010",
  25134=>"110001001",
  25135=>"100110100",
  25136=>"101110011",
  25137=>"001100000",
  25138=>"100100000",
  25139=>"101111111",
  25140=>"111100111",
  25141=>"111110010",
  25142=>"010001100",
  25143=>"011001001",
  25144=>"010110110",
  25145=>"001011001",
  25146=>"100001110",
  25147=>"101010111",
  25148=>"001110111",
  25149=>"100010010",
  25150=>"011101010",
  25151=>"010001111",
  25152=>"101011001",
  25153=>"111101110",
  25154=>"101111001",
  25155=>"101110010",
  25156=>"101101111",
  25157=>"011001001",
  25158=>"001111101",
  25159=>"100101010",
  25160=>"000111101",
  25161=>"100010010",
  25162=>"000111010",
  25163=>"001100101",
  25164=>"111010011",
  25165=>"100100010",
  25166=>"101010110",
  25167=>"001100111",
  25168=>"101111011",
  25169=>"001110001",
  25170=>"010110011",
  25171=>"000001001",
  25172=>"100110110",
  25173=>"110100100",
  25174=>"001000100",
  25175=>"010001001",
  25176=>"100010011",
  25177=>"001010100",
  25178=>"011101100",
  25179=>"110011000",
  25180=>"011011101",
  25181=>"001100101",
  25182=>"011001110",
  25183=>"001101101",
  25184=>"001111000",
  25185=>"101000000",
  25186=>"001011000",
  25187=>"011100111",
  25188=>"000010100",
  25189=>"010001000",
  25190=>"011001011",
  25191=>"001001001",
  25192=>"100001000",
  25193=>"011011100",
  25194=>"100011100",
  25195=>"110100110",
  25196=>"101100011",
  25197=>"111000011",
  25198=>"101101111",
  25199=>"100001111",
  25200=>"000001111",
  25201=>"010101101",
  25202=>"001000100",
  25203=>"000000001",
  25204=>"000010100",
  25205=>"000010010",
  25206=>"001001000",
  25207=>"001010101",
  25208=>"010101110",
  25209=>"011110001",
  25210=>"111111011",
  25211=>"111001011",
  25212=>"100100010",
  25213=>"101011110",
  25214=>"110111111",
  25215=>"010101001",
  25216=>"111010110",
  25217=>"111100101",
  25218=>"010110111",
  25219=>"111011010",
  25220=>"111110101",
  25221=>"011000000",
  25222=>"101011000",
  25223=>"010000001",
  25224=>"111011000",
  25225=>"111101011",
  25226=>"101100011",
  25227=>"010100010",
  25228=>"000111000",
  25229=>"101000111",
  25230=>"001001000",
  25231=>"000100101",
  25232=>"001000110",
  25233=>"110110011",
  25234=>"100010001",
  25235=>"111000011",
  25236=>"010101101",
  25237=>"001001101",
  25238=>"111101110",
  25239=>"101110001",
  25240=>"001000010",
  25241=>"001000001",
  25242=>"110110000",
  25243=>"100101101",
  25244=>"100001000",
  25245=>"101010111",
  25246=>"000001110",
  25247=>"000101011",
  25248=>"011100000",
  25249=>"011000000",
  25250=>"011000001",
  25251=>"010011010",
  25252=>"010010010",
  25253=>"001101111",
  25254=>"100101111",
  25255=>"110100101",
  25256=>"110001110",
  25257=>"001101010",
  25258=>"111000001",
  25259=>"001100101",
  25260=>"111111010",
  25261=>"011010101",
  25262=>"111111101",
  25263=>"100111101",
  25264=>"111111110",
  25265=>"011100100",
  25266=>"001011000",
  25267=>"110110011",
  25268=>"001111000",
  25269=>"111001101",
  25270=>"001001101",
  25271=>"011101110",
  25272=>"000100110",
  25273=>"000101110",
  25274=>"110011100",
  25275=>"100111000",
  25276=>"001101100",
  25277=>"101111100",
  25278=>"110011001",
  25279=>"111110000",
  25280=>"001011000",
  25281=>"100100100",
  25282=>"001110101",
  25283=>"000000010",
  25284=>"101001100",
  25285=>"010100000",
  25286=>"110100100",
  25287=>"001001111",
  25288=>"111101011",
  25289=>"001101011",
  25290=>"010011100",
  25291=>"101110011",
  25292=>"010101101",
  25293=>"001110011",
  25294=>"110100010",
  25295=>"110001110",
  25296=>"001011101",
  25297=>"100101111",
  25298=>"000010000",
  25299=>"000100001",
  25300=>"110010111",
  25301=>"000011010",
  25302=>"101010100",
  25303=>"000010000",
  25304=>"111010100",
  25305=>"110110101",
  25306=>"110000100",
  25307=>"010101111",
  25308=>"011011010",
  25309=>"100100101",
  25310=>"001001110",
  25311=>"000011011",
  25312=>"101001100",
  25313=>"100000011",
  25314=>"011100111",
  25315=>"001000101",
  25316=>"111111011",
  25317=>"101101001",
  25318=>"111001111",
  25319=>"110000101",
  25320=>"001001110",
  25321=>"000001100",
  25322=>"101100101",
  25323=>"110101010",
  25324=>"000010001",
  25325=>"010111001",
  25326=>"101111111",
  25327=>"100101101",
  25328=>"011111000",
  25329=>"011101100",
  25330=>"110000000",
  25331=>"101100110",
  25332=>"010010011",
  25333=>"101011010",
  25334=>"000101101",
  25335=>"110011101",
  25336=>"100111011",
  25337=>"001000101",
  25338=>"111101100",
  25339=>"110000000",
  25340=>"000000010",
  25341=>"111100111",
  25342=>"010110111",
  25343=>"001101110",
  25344=>"100101100",
  25345=>"110001000",
  25346=>"110010001",
  25347=>"010001010",
  25348=>"000000110",
  25349=>"110001011",
  25350=>"101000111",
  25351=>"001010111",
  25352=>"111100110",
  25353=>"001010001",
  25354=>"111000010",
  25355=>"111010011",
  25356=>"111101111",
  25357=>"111011100",
  25358=>"100111100",
  25359=>"100111100",
  25360=>"111100101",
  25361=>"000110110",
  25362=>"000101100",
  25363=>"100111000",
  25364=>"110100110",
  25365=>"000001111",
  25366=>"010110011",
  25367=>"010010001",
  25368=>"111110110",
  25369=>"010001000",
  25370=>"111111010",
  25371=>"001000111",
  25372=>"101110101",
  25373=>"001000110",
  25374=>"111100101",
  25375=>"110100001",
  25376=>"111000011",
  25377=>"100111110",
  25378=>"110011000",
  25379=>"100000001",
  25380=>"111010000",
  25381=>"010011100",
  25382=>"111100111",
  25383=>"111001011",
  25384=>"111001001",
  25385=>"001110100",
  25386=>"000000001",
  25387=>"010010010",
  25388=>"101111010",
  25389=>"111001110",
  25390=>"001100010",
  25391=>"000100011",
  25392=>"010111100",
  25393=>"011100011",
  25394=>"111001111",
  25395=>"001100010",
  25396=>"001011001",
  25397=>"010110010",
  25398=>"100100001",
  25399=>"010111001",
  25400=>"100000100",
  25401=>"101000101",
  25402=>"100100010",
  25403=>"000111101",
  25404=>"110111010",
  25405=>"100000110",
  25406=>"001000100",
  25407=>"100111011",
  25408=>"100001110",
  25409=>"111110111",
  25410=>"001000000",
  25411=>"001101100",
  25412=>"101101111",
  25413=>"110011010",
  25414=>"100101101",
  25415=>"000111101",
  25416=>"011110000",
  25417=>"000010111",
  25418=>"001000111",
  25419=>"000110001",
  25420=>"100110100",
  25421=>"011000010",
  25422=>"000000001",
  25423=>"010011001",
  25424=>"111010110",
  25425=>"011011011",
  25426=>"101111000",
  25427=>"111000000",
  25428=>"011111001",
  25429=>"000101110",
  25430=>"000110101",
  25431=>"100111111",
  25432=>"011101000",
  25433=>"110100010",
  25434=>"111001101",
  25435=>"010000010",
  25436=>"111111101",
  25437=>"111101010",
  25438=>"000110010",
  25439=>"010001110",
  25440=>"001000000",
  25441=>"011100000",
  25442=>"001001111",
  25443=>"110101100",
  25444=>"111001011",
  25445=>"111100110",
  25446=>"101111110",
  25447=>"100001111",
  25448=>"101011001",
  25449=>"111111001",
  25450=>"101111000",
  25451=>"110110100",
  25452=>"000011101",
  25453=>"111110101",
  25454=>"111011001",
  25455=>"101101011",
  25456=>"110110101",
  25457=>"110111100",
  25458=>"111001000",
  25459=>"100001010",
  25460=>"101010110",
  25461=>"001011010",
  25462=>"110000010",
  25463=>"000100110",
  25464=>"010000110",
  25465=>"100111000",
  25466=>"011100100",
  25467=>"111111101",
  25468=>"011001001",
  25469=>"101010111",
  25470=>"111010101",
  25471=>"110111010",
  25472=>"001100101",
  25473=>"000001101",
  25474=>"000011010",
  25475=>"110000111",
  25476=>"111100100",
  25477=>"110010000",
  25478=>"100000000",
  25479=>"100101110",
  25480=>"110100110",
  25481=>"000010000",
  25482=>"010011001",
  25483=>"000011000",
  25484=>"100110110",
  25485=>"010010101",
  25486=>"010110110",
  25487=>"010111111",
  25488=>"110110001",
  25489=>"010011001",
  25490=>"000110001",
  25491=>"110100001",
  25492=>"001001001",
  25493=>"000100100",
  25494=>"000110011",
  25495=>"010010101",
  25496=>"001011101",
  25497=>"001001101",
  25498=>"010010010",
  25499=>"110101110",
  25500=>"001010000",
  25501=>"001100000",
  25502=>"011001101",
  25503=>"010101011",
  25504=>"010111001",
  25505=>"111110110",
  25506=>"101010011",
  25507=>"100101011",
  25508=>"110100100",
  25509=>"010001110",
  25510=>"010010001",
  25511=>"000111101",
  25512=>"000001010",
  25513=>"111001000",
  25514=>"011111011",
  25515=>"111110101",
  25516=>"110110111",
  25517=>"101101010",
  25518=>"000101111",
  25519=>"111011111",
  25520=>"001110101",
  25521=>"001111011",
  25522=>"111011000",
  25523=>"000111000",
  25524=>"001111110",
  25525=>"110110100",
  25526=>"010010011",
  25527=>"100000100",
  25528=>"011011101",
  25529=>"011101001",
  25530=>"010001001",
  25531=>"100000011",
  25532=>"111001111",
  25533=>"010101000",
  25534=>"111111110",
  25535=>"110001011",
  25536=>"110000000",
  25537=>"001011011",
  25538=>"101001010",
  25539=>"100010100",
  25540=>"000010110",
  25541=>"111010111",
  25542=>"111011001",
  25543=>"000100111",
  25544=>"010100100",
  25545=>"011111011",
  25546=>"000110001",
  25547=>"101011000",
  25548=>"110100110",
  25549=>"100000101",
  25550=>"100110101",
  25551=>"101101011",
  25552=>"111101111",
  25553=>"101110100",
  25554=>"101011001",
  25555=>"101110000",
  25556=>"000101100",
  25557=>"111010101",
  25558=>"101100111",
  25559=>"111111101",
  25560=>"101001001",
  25561=>"001110110",
  25562=>"101011001",
  25563=>"010000011",
  25564=>"011111111",
  25565=>"100110110",
  25566=>"111000110",
  25567=>"011000000",
  25568=>"011100000",
  25569=>"011101011",
  25570=>"100000111",
  25571=>"001000000",
  25572=>"101110001",
  25573=>"000001100",
  25574=>"000000001",
  25575=>"000100010",
  25576=>"100001110",
  25577=>"101101011",
  25578=>"101110110",
  25579=>"000011110",
  25580=>"100100001",
  25581=>"101011000",
  25582=>"001000111",
  25583=>"000101111",
  25584=>"010110001",
  25585=>"000001010",
  25586=>"000001111",
  25587=>"010010011",
  25588=>"101101100",
  25589=>"010101101",
  25590=>"111011111",
  25591=>"111001011",
  25592=>"000000110",
  25593=>"011001000",
  25594=>"010111001",
  25595=>"101010001",
  25596=>"000101000",
  25597=>"000010001",
  25598=>"000010110",
  25599=>"011001110",
  25600=>"100101000",
  25601=>"010010010",
  25602=>"110001101",
  25603=>"001111101",
  25604=>"100110110",
  25605=>"000101100",
  25606=>"111001110",
  25607=>"001011100",
  25608=>"100101101",
  25609=>"110000110",
  25610=>"111110001",
  25611=>"110010110",
  25612=>"110000100",
  25613=>"100011001",
  25614=>"011111100",
  25615=>"011010100",
  25616=>"110111100",
  25617=>"101001100",
  25618=>"100101111",
  25619=>"001100010",
  25620=>"110000100",
  25621=>"001011011",
  25622=>"010100011",
  25623=>"110011011",
  25624=>"000010100",
  25625=>"111001100",
  25626=>"010101010",
  25627=>"110101101",
  25628=>"100111110",
  25629=>"110111110",
  25630=>"110110100",
  25631=>"110110110",
  25632=>"111001000",
  25633=>"100100111",
  25634=>"100000101",
  25635=>"011000011",
  25636=>"110001101",
  25637=>"011010001",
  25638=>"001000001",
  25639=>"101110111",
  25640=>"000010100",
  25641=>"011111101",
  25642=>"001011111",
  25643=>"100001110",
  25644=>"010110011",
  25645=>"000111010",
  25646=>"011101010",
  25647=>"101010110",
  25648=>"111110011",
  25649=>"000001000",
  25650=>"101000110",
  25651=>"000000000",
  25652=>"001000100",
  25653=>"001100001",
  25654=>"000001010",
  25655=>"111100110",
  25656=>"000111101",
  25657=>"101110101",
  25658=>"100000100",
  25659=>"100100011",
  25660=>"001000100",
  25661=>"000011100",
  25662=>"000100101",
  25663=>"101110101",
  25664=>"100111000",
  25665=>"001001110",
  25666=>"110111000",
  25667=>"000110010",
  25668=>"100010011",
  25669=>"011010001",
  25670=>"100000100",
  25671=>"000001100",
  25672=>"111111010",
  25673=>"100010101",
  25674=>"001100000",
  25675=>"111110101",
  25676=>"010000000",
  25677=>"101011110",
  25678=>"110100110",
  25679=>"111000011",
  25680=>"000000110",
  25681=>"101110011",
  25682=>"101100111",
  25683=>"111000000",
  25684=>"101000000",
  25685=>"101010111",
  25686=>"100101100",
  25687=>"010100111",
  25688=>"011010110",
  25689=>"111010010",
  25690=>"101110111",
  25691=>"000010111",
  25692=>"001001010",
  25693=>"011101011",
  25694=>"010100101",
  25695=>"100001001",
  25696=>"101010000",
  25697=>"100000110",
  25698=>"010100010",
  25699=>"000011001",
  25700=>"100001111",
  25701=>"101101000",
  25702=>"111010110",
  25703=>"000000111",
  25704=>"000000011",
  25705=>"100100101",
  25706=>"111110001",
  25707=>"110010010",
  25708=>"110111001",
  25709=>"010011011",
  25710=>"011110000",
  25711=>"101001000",
  25712=>"111010010",
  25713=>"011100000",
  25714=>"100111110",
  25715=>"110011100",
  25716=>"100110100",
  25717=>"011011101",
  25718=>"010001101",
  25719=>"001110011",
  25720=>"001100011",
  25721=>"001111100",
  25722=>"111111011",
  25723=>"111101100",
  25724=>"001100110",
  25725=>"010111000",
  25726=>"000001000",
  25727=>"000001100",
  25728=>"100010111",
  25729=>"101010011",
  25730=>"000000000",
  25731=>"001010011",
  25732=>"010000010",
  25733=>"011001100",
  25734=>"110111000",
  25735=>"000011100",
  25736=>"000001011",
  25737=>"100111101",
  25738=>"011000000",
  25739=>"100110101",
  25740=>"100110100",
  25741=>"101001001",
  25742=>"110100111",
  25743=>"011000001",
  25744=>"101111010",
  25745=>"110001001",
  25746=>"001001000",
  25747=>"111011101",
  25748=>"111101110",
  25749=>"000000011",
  25750=>"000010001",
  25751=>"000110101",
  25752=>"010000011",
  25753=>"100000101",
  25754=>"111000111",
  25755=>"001111011",
  25756=>"101001101",
  25757=>"000110100",
  25758=>"111110101",
  25759=>"111101001",
  25760=>"101000100",
  25761=>"110111011",
  25762=>"110011111",
  25763=>"100100011",
  25764=>"101111111",
  25765=>"110111111",
  25766=>"110011101",
  25767=>"010100110",
  25768=>"011011000",
  25769=>"000001001",
  25770=>"001100011",
  25771=>"011111000",
  25772=>"011010100",
  25773=>"111011000",
  25774=>"101111011",
  25775=>"111011101",
  25776=>"011010010",
  25777=>"111111101",
  25778=>"000101001",
  25779=>"010010001",
  25780=>"101101000",
  25781=>"101111111",
  25782=>"011001101",
  25783=>"100110011",
  25784=>"110000010",
  25785=>"010110101",
  25786=>"011010000",
  25787=>"111000101",
  25788=>"111000010",
  25789=>"010100001",
  25790=>"110101000",
  25791=>"111111101",
  25792=>"110110110",
  25793=>"011101101",
  25794=>"010100010",
  25795=>"100010000",
  25796=>"101101000",
  25797=>"000101000",
  25798=>"101110011",
  25799=>"000010011",
  25800=>"010110011",
  25801=>"101011011",
  25802=>"011101111",
  25803=>"010001011",
  25804=>"010111010",
  25805=>"001101111",
  25806=>"011110111",
  25807=>"101000110",
  25808=>"000100100",
  25809=>"010010111",
  25810=>"000001110",
  25811=>"111101110",
  25812=>"000100100",
  25813=>"111110101",
  25814=>"101010101",
  25815=>"100001101",
  25816=>"110110111",
  25817=>"010010110",
  25818=>"011111000",
  25819=>"111010000",
  25820=>"000000101",
  25821=>"001101001",
  25822=>"001010111",
  25823=>"010110101",
  25824=>"111100110",
  25825=>"010010100",
  25826=>"100100110",
  25827=>"000100101",
  25828=>"100010110",
  25829=>"001001010",
  25830=>"100111110",
  25831=>"111111110",
  25832=>"111010010",
  25833=>"011110110",
  25834=>"101100001",
  25835=>"001100110",
  25836=>"101101100",
  25837=>"110110100",
  25838=>"001000110",
  25839=>"000000010",
  25840=>"011111101",
  25841=>"111101100",
  25842=>"011101111",
  25843=>"111110100",
  25844=>"011001101",
  25845=>"001101110",
  25846=>"111110010",
  25847=>"011110001",
  25848=>"000001001",
  25849=>"111100000",
  25850=>"001001100",
  25851=>"000001000",
  25852=>"000100101",
  25853=>"111011000",
  25854=>"101010110",
  25855=>"100011101",
  25856=>"000101101",
  25857=>"101001100",
  25858=>"101000001",
  25859=>"010010011",
  25860=>"001110010",
  25861=>"110000000",
  25862=>"011000111",
  25863=>"111001000",
  25864=>"010011101",
  25865=>"010100110",
  25866=>"000000100",
  25867=>"000010000",
  25868=>"010000111",
  25869=>"110110110",
  25870=>"101100110",
  25871=>"000110010",
  25872=>"010101010",
  25873=>"001100100",
  25874=>"111100011",
  25875=>"010000000",
  25876=>"100010010",
  25877=>"011101001",
  25878=>"001000111",
  25879=>"101000110",
  25880=>"111000011",
  25881=>"001010101",
  25882=>"011011101",
  25883=>"000010110",
  25884=>"001111011",
  25885=>"111001101",
  25886=>"101001100",
  25887=>"100101110",
  25888=>"100011111",
  25889=>"110000010",
  25890=>"111011000",
  25891=>"100001111",
  25892=>"110110111",
  25893=>"110010101",
  25894=>"100000011",
  25895=>"000011100",
  25896=>"100011111",
  25897=>"111101110",
  25898=>"111011101",
  25899=>"000110100",
  25900=>"100001101",
  25901=>"110111000",
  25902=>"001001001",
  25903=>"111001010",
  25904=>"111100111",
  25905=>"101011011",
  25906=>"001001100",
  25907=>"000000110",
  25908=>"100100010",
  25909=>"010010001",
  25910=>"101000011",
  25911=>"100001111",
  25912=>"001000010",
  25913=>"110111000",
  25914=>"001000000",
  25915=>"011000111",
  25916=>"001001110",
  25917=>"110011011",
  25918=>"000010110",
  25919=>"111101000",
  25920=>"001100101",
  25921=>"101010010",
  25922=>"100101110",
  25923=>"000011001",
  25924=>"100010111",
  25925=>"001000000",
  25926=>"000010000",
  25927=>"001011001",
  25928=>"110011000",
  25929=>"000101010",
  25930=>"101110000",
  25931=>"000010110",
  25932=>"000011000",
  25933=>"101010110",
  25934=>"000001100",
  25935=>"100000010",
  25936=>"011010111",
  25937=>"111001011",
  25938=>"000101111",
  25939=>"011101000",
  25940=>"100100000",
  25941=>"100110001",
  25942=>"110100000",
  25943=>"110111000",
  25944=>"001111111",
  25945=>"001001011",
  25946=>"011101000",
  25947=>"110001111",
  25948=>"111001001",
  25949=>"101111010",
  25950=>"011010100",
  25951=>"000101111",
  25952=>"011010100",
  25953=>"011011001",
  25954=>"101011011",
  25955=>"000010011",
  25956=>"100101001",
  25957=>"010011010",
  25958=>"111101101",
  25959=>"000010010",
  25960=>"011110101",
  25961=>"000000110",
  25962=>"111011111",
  25963=>"100100010",
  25964=>"110101000",
  25965=>"101010000",
  25966=>"110100100",
  25967=>"010010100",
  25968=>"111000110",
  25969=>"000100101",
  25970=>"000110011",
  25971=>"010111111",
  25972=>"000111111",
  25973=>"010001110",
  25974=>"111001000",
  25975=>"001100010",
  25976=>"110101101",
  25977=>"011000011",
  25978=>"011000001",
  25979=>"000101100",
  25980=>"100000011",
  25981=>"111110101",
  25982=>"000111011",
  25983=>"010000110",
  25984=>"110000111",
  25985=>"000111010",
  25986=>"111010000",
  25987=>"111000011",
  25988=>"001011000",
  25989=>"110001010",
  25990=>"000010000",
  25991=>"001010011",
  25992=>"000100100",
  25993=>"000010000",
  25994=>"101011001",
  25995=>"011011010",
  25996=>"011000001",
  25997=>"111111010",
  25998=>"001110010",
  25999=>"000010010",
  26000=>"000100011",
  26001=>"010101111",
  26002=>"110010100",
  26003=>"001100100",
  26004=>"011111110",
  26005=>"001110000",
  26006=>"111100110",
  26007=>"011010000",
  26008=>"101010101",
  26009=>"011000001",
  26010=>"001001110",
  26011=>"000100001",
  26012=>"100011000",
  26013=>"111111000",
  26014=>"110010011",
  26015=>"111000011",
  26016=>"001010100",
  26017=>"111011001",
  26018=>"111011000",
  26019=>"100000000",
  26020=>"110010100",
  26021=>"000100010",
  26022=>"000110001",
  26023=>"111011010",
  26024=>"111010011",
  26025=>"110001101",
  26026=>"101111111",
  26027=>"000000001",
  26028=>"010101000",
  26029=>"110011111",
  26030=>"000110000",
  26031=>"000111011",
  26032=>"000001001",
  26033=>"001101111",
  26034=>"011010110",
  26035=>"011011001",
  26036=>"011001100",
  26037=>"010110101",
  26038=>"101011001",
  26039=>"111101000",
  26040=>"000000110",
  26041=>"100100000",
  26042=>"000100000",
  26043=>"110100100",
  26044=>"110110001",
  26045=>"110111010",
  26046=>"101011111",
  26047=>"000101110",
  26048=>"001010000",
  26049=>"011111011",
  26050=>"100010100",
  26051=>"000100010",
  26052=>"010000110",
  26053=>"111000011",
  26054=>"100010011",
  26055=>"110101000",
  26056=>"101100011",
  26057=>"100011100",
  26058=>"101011011",
  26059=>"010001001",
  26060=>"010001111",
  26061=>"001110100",
  26062=>"001110001",
  26063=>"101110010",
  26064=>"110110001",
  26065=>"011000100",
  26066=>"000001010",
  26067=>"000111111",
  26068=>"011101100",
  26069=>"000000011",
  26070=>"111001001",
  26071=>"110101101",
  26072=>"000100100",
  26073=>"100010000",
  26074=>"111010111",
  26075=>"011001000",
  26076=>"100010001",
  26077=>"101110100",
  26078=>"110111000",
  26079=>"110111010",
  26080=>"001101101",
  26081=>"010111101",
  26082=>"101011100",
  26083=>"001001100",
  26084=>"101001000",
  26085=>"001111100",
  26086=>"001011010",
  26087=>"001111000",
  26088=>"111001111",
  26089=>"111100111",
  26090=>"010001011",
  26091=>"000110010",
  26092=>"101001011",
  26093=>"010000010",
  26094=>"001001100",
  26095=>"100101111",
  26096=>"001000011",
  26097=>"100111100",
  26098=>"010011001",
  26099=>"001011010",
  26100=>"101000111",
  26101=>"000111101",
  26102=>"100110001",
  26103=>"111001011",
  26104=>"000111000",
  26105=>"101110000",
  26106=>"111110101",
  26107=>"100001101",
  26108=>"000101011",
  26109=>"000000110",
  26110=>"000100101",
  26111=>"110101001",
  26112=>"000011001",
  26113=>"000000110",
  26114=>"111011110",
  26115=>"000000000",
  26116=>"111101100",
  26117=>"010110100",
  26118=>"011000001",
  26119=>"111111101",
  26120=>"100101001",
  26121=>"010011000",
  26122=>"111100100",
  26123=>"010000001",
  26124=>"001000010",
  26125=>"001010011",
  26126=>"000000110",
  26127=>"001011010",
  26128=>"100000011",
  26129=>"111001111",
  26130=>"100011111",
  26131=>"110010011",
  26132=>"100110000",
  26133=>"110001011",
  26134=>"010100101",
  26135=>"011001010",
  26136=>"110010111",
  26137=>"101010111",
  26138=>"101110011",
  26139=>"001101010",
  26140=>"110111111",
  26141=>"100001010",
  26142=>"101111000",
  26143=>"010001110",
  26144=>"101000000",
  26145=>"010100011",
  26146=>"000001010",
  26147=>"100001001",
  26148=>"010011011",
  26149=>"111111100",
  26150=>"100111010",
  26151=>"011001000",
  26152=>"110001001",
  26153=>"001110111",
  26154=>"111101001",
  26155=>"100000011",
  26156=>"011100111",
  26157=>"000000010",
  26158=>"100101111",
  26159=>"101101011",
  26160=>"010001111",
  26161=>"101010100",
  26162=>"000000110",
  26163=>"010001000",
  26164=>"001111001",
  26165=>"110010010",
  26166=>"010010110",
  26167=>"001001001",
  26168=>"011010100",
  26169=>"010111001",
  26170=>"011000010",
  26171=>"101111010",
  26172=>"011011110",
  26173=>"010100100",
  26174=>"111011001",
  26175=>"110010000",
  26176=>"110010110",
  26177=>"001100001",
  26178=>"001101011",
  26179=>"101110100",
  26180=>"101100001",
  26181=>"011100101",
  26182=>"101001011",
  26183=>"001100101",
  26184=>"011111110",
  26185=>"000001101",
  26186=>"111000010",
  26187=>"111111111",
  26188=>"101110011",
  26189=>"110101110",
  26190=>"111101000",
  26191=>"000001110",
  26192=>"000101010",
  26193=>"101111111",
  26194=>"010000001",
  26195=>"101101101",
  26196=>"101101001",
  26197=>"100110011",
  26198=>"111111011",
  26199=>"111100010",
  26200=>"001101001",
  26201=>"000100110",
  26202=>"001100010",
  26203=>"000101000",
  26204=>"000011101",
  26205=>"000001010",
  26206=>"100010101",
  26207=>"110101100",
  26208=>"100010100",
  26209=>"101001010",
  26210=>"001110000",
  26211=>"100110001",
  26212=>"000000001",
  26213=>"010100011",
  26214=>"001110011",
  26215=>"110101111",
  26216=>"010100110",
  26217=>"010100100",
  26218=>"101111100",
  26219=>"111011010",
  26220=>"001111111",
  26221=>"001010001",
  26222=>"011000001",
  26223=>"011000011",
  26224=>"100100011",
  26225=>"010000100",
  26226=>"010010100",
  26227=>"101100111",
  26228=>"000110001",
  26229=>"011001101",
  26230=>"101010111",
  26231=>"000100000",
  26232=>"111101111",
  26233=>"011101101",
  26234=>"011101100",
  26235=>"001110011",
  26236=>"110010010",
  26237=>"010010001",
  26238=>"100111011",
  26239=>"001000000",
  26240=>"111011000",
  26241=>"001010100",
  26242=>"011010100",
  26243=>"111011111",
  26244=>"111100111",
  26245=>"010000001",
  26246=>"101001001",
  26247=>"100111010",
  26248=>"000011110",
  26249=>"000001000",
  26250=>"011101011",
  26251=>"110010001",
  26252=>"110101011",
  26253=>"001100001",
  26254=>"101000000",
  26255=>"000001111",
  26256=>"000101110",
  26257=>"010111011",
  26258=>"101101111",
  26259=>"111110011",
  26260=>"010010111",
  26261=>"001111000",
  26262=>"011111100",
  26263=>"000101100",
  26264=>"010010100",
  26265=>"100110111",
  26266=>"001110001",
  26267=>"100001110",
  26268=>"011000001",
  26269=>"110000001",
  26270=>"010101011",
  26271=>"101000111",
  26272=>"100110011",
  26273=>"000000010",
  26274=>"101111000",
  26275=>"010110011",
  26276=>"111101100",
  26277=>"010110000",
  26278=>"000011000",
  26279=>"000011000",
  26280=>"000001011",
  26281=>"011000110",
  26282=>"000100001",
  26283=>"110111000",
  26284=>"001011100",
  26285=>"011000110",
  26286=>"101111011",
  26287=>"000010010",
  26288=>"110111101",
  26289=>"111010000",
  26290=>"111110111",
  26291=>"011010101",
  26292=>"110101101",
  26293=>"101101100",
  26294=>"100000011",
  26295=>"010001001",
  26296=>"010110001",
  26297=>"001010100",
  26298=>"110111111",
  26299=>"000001010",
  26300=>"100001101",
  26301=>"011100010",
  26302=>"011000010",
  26303=>"100111010",
  26304=>"100011010",
  26305=>"110100111",
  26306=>"110101001",
  26307=>"001001010",
  26308=>"100110100",
  26309=>"011111111",
  26310=>"110000011",
  26311=>"001111110",
  26312=>"100000110",
  26313=>"001000000",
  26314=>"111110011",
  26315=>"000001000",
  26316=>"001000011",
  26317=>"010111001",
  26318=>"110010001",
  26319=>"000010001",
  26320=>"000010001",
  26321=>"010101111",
  26322=>"101000011",
  26323=>"110000100",
  26324=>"101101010",
  26325=>"000000100",
  26326=>"111110110",
  26327=>"111111110",
  26328=>"001100001",
  26329=>"100101010",
  26330=>"111000101",
  26331=>"000011010",
  26332=>"111111110",
  26333=>"111011010",
  26334=>"111110100",
  26335=>"111011110",
  26336=>"111111110",
  26337=>"100100000",
  26338=>"100001101",
  26339=>"000001100",
  26340=>"010010010",
  26341=>"000110100",
  26342=>"011000110",
  26343=>"000110001",
  26344=>"101100000",
  26345=>"101000011",
  26346=>"000011111",
  26347=>"110100101",
  26348=>"000010100",
  26349=>"001110010",
  26350=>"101101010",
  26351=>"000001001",
  26352=>"001100101",
  26353=>"101101110",
  26354=>"011100001",
  26355=>"001001001",
  26356=>"100010010",
  26357=>"111101101",
  26358=>"111000100",
  26359=>"110100100",
  26360=>"100111100",
  26361=>"000011011",
  26362=>"011110101",
  26363=>"110010010",
  26364=>"001111110",
  26365=>"110000111",
  26366=>"111101100",
  26367=>"010000100",
  26368=>"111001001",
  26369=>"011010110",
  26370=>"101110010",
  26371=>"010011010",
  26372=>"000000110",
  26373=>"101000001",
  26374=>"101101011",
  26375=>"100110011",
  26376=>"100101101",
  26377=>"101111110",
  26378=>"110010011",
  26379=>"100010101",
  26380=>"010010110",
  26381=>"100100101",
  26382=>"011001010",
  26383=>"001101101",
  26384=>"011111100",
  26385=>"100000001",
  26386=>"011100010",
  26387=>"111111111",
  26388=>"101111010",
  26389=>"011111000",
  26390=>"111010000",
  26391=>"011011011",
  26392=>"000110000",
  26393=>"010000111",
  26394=>"111011111",
  26395=>"110010101",
  26396=>"100110001",
  26397=>"111010001",
  26398=>"001110000",
  26399=>"111011101",
  26400=>"101111011",
  26401=>"101001111",
  26402=>"011101011",
  26403=>"000100101",
  26404=>"101111001",
  26405=>"001011010",
  26406=>"010101111",
  26407=>"011000110",
  26408=>"100101010",
  26409=>"011011001",
  26410=>"111111101",
  26411=>"110111000",
  26412=>"011001101",
  26413=>"000010100",
  26414=>"001111000",
  26415=>"111001011",
  26416=>"100100010",
  26417=>"000001100",
  26418=>"101001001",
  26419=>"000001101",
  26420=>"111101101",
  26421=>"100001111",
  26422=>"101000100",
  26423=>"110011100",
  26424=>"110001000",
  26425=>"100001011",
  26426=>"010101011",
  26427=>"101001100",
  26428=>"011010010",
  26429=>"100101110",
  26430=>"101000000",
  26431=>"110110001",
  26432=>"001101110",
  26433=>"101100110",
  26434=>"100010010",
  26435=>"110011111",
  26436=>"110100101",
  26437=>"101001101",
  26438=>"110101011",
  26439=>"111100010",
  26440=>"011110010",
  26441=>"100001100",
  26442=>"001000010",
  26443=>"100000111",
  26444=>"000001110",
  26445=>"000011000",
  26446=>"010100000",
  26447=>"000101001",
  26448=>"010010100",
  26449=>"010110010",
  26450=>"000101011",
  26451=>"000011001",
  26452=>"110001101",
  26453=>"101111000",
  26454=>"100110101",
  26455=>"000001110",
  26456=>"001111111",
  26457=>"001000111",
  26458=>"101110110",
  26459=>"101010101",
  26460=>"011111100",
  26461=>"111010001",
  26462=>"101000001",
  26463=>"000001101",
  26464=>"100110001",
  26465=>"111111111",
  26466=>"100100101",
  26467=>"100100001",
  26468=>"011111001",
  26469=>"101101101",
  26470=>"110011011",
  26471=>"010110111",
  26472=>"110001110",
  26473=>"110000111",
  26474=>"001010010",
  26475=>"100100011",
  26476=>"000001000",
  26477=>"001000010",
  26478=>"001010000",
  26479=>"000101011",
  26480=>"010000001",
  26481=>"110000101",
  26482=>"000111110",
  26483=>"001011101",
  26484=>"000000000",
  26485=>"000111111",
  26486=>"110101110",
  26487=>"001000111",
  26488=>"101100010",
  26489=>"111000111",
  26490=>"000100010",
  26491=>"100101001",
  26492=>"000010000",
  26493=>"111001000",
  26494=>"100101011",
  26495=>"101011101",
  26496=>"001001100",
  26497=>"100110111",
  26498=>"000100000",
  26499=>"110011110",
  26500=>"110110111",
  26501=>"011111001",
  26502=>"110100100",
  26503=>"100001011",
  26504=>"110101010",
  26505=>"110100101",
  26506=>"000010010",
  26507=>"000110000",
  26508=>"011111001",
  26509=>"101111111",
  26510=>"001110100",
  26511=>"100010101",
  26512=>"111011011",
  26513=>"000001001",
  26514=>"000000000",
  26515=>"001011001",
  26516=>"100010111",
  26517=>"111011111",
  26518=>"000110110",
  26519=>"100011011",
  26520=>"110000000",
  26521=>"000011011",
  26522=>"111111111",
  26523=>"100010100",
  26524=>"111110000",
  26525=>"001001100",
  26526=>"101001000",
  26527=>"101010110",
  26528=>"000001000",
  26529=>"001111010",
  26530=>"001111011",
  26531=>"010010111",
  26532=>"010010000",
  26533=>"010001111",
  26534=>"000110110",
  26535=>"010100001",
  26536=>"001111001",
  26537=>"011011010",
  26538=>"100111100",
  26539=>"011100100",
  26540=>"000011111",
  26541=>"000101101",
  26542=>"101000111",
  26543=>"001011000",
  26544=>"000111011",
  26545=>"101011001",
  26546=>"011101101",
  26547=>"000100001",
  26548=>"100000010",
  26549=>"100000010",
  26550=>"100111110",
  26551=>"011101010",
  26552=>"111111000",
  26553=>"100101011",
  26554=>"011010101",
  26555=>"111101010",
  26556=>"000111100",
  26557=>"111110111",
  26558=>"001010010",
  26559=>"100010011",
  26560=>"110011111",
  26561=>"010000100",
  26562=>"111110110",
  26563=>"101111100",
  26564=>"111101101",
  26565=>"110010010",
  26566=>"000000010",
  26567=>"000000000",
  26568=>"100101000",
  26569=>"000000011",
  26570=>"000111110",
  26571=>"001011111",
  26572=>"110010111",
  26573=>"011000011",
  26574=>"011111001",
  26575=>"000010000",
  26576=>"101101001",
  26577=>"011000111",
  26578=>"110110010",
  26579=>"000010001",
  26580=>"110000011",
  26581=>"101011000",
  26582=>"110100011",
  26583=>"011001100",
  26584=>"011100011",
  26585=>"011110010",
  26586=>"011111100",
  26587=>"000100000",
  26588=>"111111111",
  26589=>"100000011",
  26590=>"110000100",
  26591=>"111110011",
  26592=>"111110010",
  26593=>"000111000",
  26594=>"001100001",
  26595=>"111100001",
  26596=>"000000000",
  26597=>"011001000",
  26598=>"100001010",
  26599=>"010110011",
  26600=>"000101010",
  26601=>"010011011",
  26602=>"010000001",
  26603=>"111111010",
  26604=>"011111000",
  26605=>"100010111",
  26606=>"101110010",
  26607=>"001001011",
  26608=>"111011100",
  26609=>"000110000",
  26610=>"110010010",
  26611=>"101101101",
  26612=>"001010000",
  26613=>"010110100",
  26614=>"100000000",
  26615=>"011110101",
  26616=>"110100001",
  26617=>"110010001",
  26618=>"001000010",
  26619=>"110011000",
  26620=>"010010100",
  26621=>"010010000",
  26622=>"000111000",
  26623=>"011000010",
  26624=>"100111110",
  26625=>"011100101",
  26626=>"100101111",
  26627=>"100111101",
  26628=>"100010101",
  26629=>"110101100",
  26630=>"001111011",
  26631=>"011111001",
  26632=>"001111000",
  26633=>"001011001",
  26634=>"100000001",
  26635=>"110010000",
  26636=>"111111000",
  26637=>"100111000",
  26638=>"011001001",
  26639=>"001101010",
  26640=>"100100010",
  26641=>"111100001",
  26642=>"111000010",
  26643=>"110010011",
  26644=>"101000001",
  26645=>"111001001",
  26646=>"100001100",
  26647=>"011111001",
  26648=>"101001000",
  26649=>"101000000",
  26650=>"001100010",
  26651=>"000111111",
  26652=>"000010100",
  26653=>"111001111",
  26654=>"001101110",
  26655=>"100000100",
  26656=>"101000010",
  26657=>"110100111",
  26658=>"000110100",
  26659=>"001110101",
  26660=>"101100100",
  26661=>"111011001",
  26662=>"100010110",
  26663=>"001001111",
  26664=>"111110010",
  26665=>"101001000",
  26666=>"101010111",
  26667=>"100011010",
  26668=>"000111111",
  26669=>"001000011",
  26670=>"100010000",
  26671=>"001100101",
  26672=>"111000000",
  26673=>"011000000",
  26674=>"110111101",
  26675=>"000111001",
  26676=>"110111010",
  26677=>"100110011",
  26678=>"010111100",
  26679=>"110100011",
  26680=>"011001101",
  26681=>"110010111",
  26682=>"010110100",
  26683=>"000001110",
  26684=>"101010000",
  26685=>"101010110",
  26686=>"101000011",
  26687=>"000011011",
  26688=>"110100010",
  26689=>"101001100",
  26690=>"110011100",
  26691=>"000011000",
  26692=>"011010000",
  26693=>"100110101",
  26694=>"110000100",
  26695=>"100110101",
  26696=>"100000110",
  26697=>"110111011",
  26698=>"101100011",
  26699=>"000001001",
  26700=>"111101110",
  26701=>"110111010",
  26702=>"111100100",
  26703=>"111000011",
  26704=>"110000111",
  26705=>"000100011",
  26706=>"110001111",
  26707=>"011111110",
  26708=>"010000110",
  26709=>"000111001",
  26710=>"110110111",
  26711=>"101110100",
  26712=>"011111111",
  26713=>"001011101",
  26714=>"100111001",
  26715=>"111110100",
  26716=>"000010011",
  26717=>"000101110",
  26718=>"000011111",
  26719=>"010000111",
  26720=>"100100011",
  26721=>"111101001",
  26722=>"100100111",
  26723=>"111001100",
  26724=>"011011101",
  26725=>"100100110",
  26726=>"010111010",
  26727=>"001011010",
  26728=>"111111100",
  26729=>"110001110",
  26730=>"000110101",
  26731=>"001101010",
  26732=>"011000000",
  26733=>"101101001",
  26734=>"010001011",
  26735=>"101100000",
  26736=>"110000001",
  26737=>"001001000",
  26738=>"101101000",
  26739=>"110000001",
  26740=>"111001010",
  26741=>"101110110",
  26742=>"110110010",
  26743=>"111101001",
  26744=>"011001101",
  26745=>"100000101",
  26746=>"110000111",
  26747=>"000001000",
  26748=>"100101010",
  26749=>"100101000",
  26750=>"000000000",
  26751=>"111101111",
  26752=>"000011101",
  26753=>"000100101",
  26754=>"101000110",
  26755=>"000010001",
  26756=>"110001101",
  26757=>"101100100",
  26758=>"110101000",
  26759=>"000000111",
  26760=>"011011001",
  26761=>"010101100",
  26762=>"000011110",
  26763=>"000111000",
  26764=>"000010001",
  26765=>"000101111",
  26766=>"010011001",
  26767=>"011000100",
  26768=>"100100100",
  26769=>"100001110",
  26770=>"101100100",
  26771=>"111100000",
  26772=>"101010000",
  26773=>"000100100",
  26774=>"011111010",
  26775=>"010100110",
  26776=>"101111010",
  26777=>"100100111",
  26778=>"000000111",
  26779=>"001100001",
  26780=>"001000101",
  26781=>"000000111",
  26782=>"011010100",
  26783=>"010111001",
  26784=>"110001010",
  26785=>"100101001",
  26786=>"100101001",
  26787=>"111100101",
  26788=>"111100111",
  26789=>"101111110",
  26790=>"110011110",
  26791=>"010101110",
  26792=>"111000111",
  26793=>"110110011",
  26794=>"011000110",
  26795=>"101001001",
  26796=>"001111110",
  26797=>"100101011",
  26798=>"010011010",
  26799=>"110110110",
  26800=>"011111100",
  26801=>"000010100",
  26802=>"101101001",
  26803=>"001010000",
  26804=>"111100001",
  26805=>"000101100",
  26806=>"000000100",
  26807=>"111010111",
  26808=>"010000011",
  26809=>"101011010",
  26810=>"010001011",
  26811=>"111010111",
  26812=>"101110001",
  26813=>"001111000",
  26814=>"011110000",
  26815=>"111100001",
  26816=>"110011111",
  26817=>"110110011",
  26818=>"100111100",
  26819=>"010110101",
  26820=>"110000011",
  26821=>"101111111",
  26822=>"000001101",
  26823=>"101111000",
  26824=>"010000110",
  26825=>"001101001",
  26826=>"111010000",
  26827=>"111110111",
  26828=>"010010010",
  26829=>"111111100",
  26830=>"101000111",
  26831=>"010111001",
  26832=>"111111000",
  26833=>"001100000",
  26834=>"000100010",
  26835=>"010001101",
  26836=>"110010100",
  26837=>"100001001",
  26838=>"011011110",
  26839=>"011100011",
  26840=>"000101000",
  26841=>"011010001",
  26842=>"010000101",
  26843=>"100111011",
  26844=>"110001110",
  26845=>"111111001",
  26846=>"111110110",
  26847=>"100001001",
  26848=>"010101011",
  26849=>"011101110",
  26850=>"010000100",
  26851=>"000000001",
  26852=>"010111100",
  26853=>"000000011",
  26854=>"100010010",
  26855=>"010101000",
  26856=>"011010100",
  26857=>"110000100",
  26858=>"111111001",
  26859=>"000101111",
  26860=>"101000011",
  26861=>"100110111",
  26862=>"001000001",
  26863=>"111000000",
  26864=>"110010100",
  26865=>"110010011",
  26866=>"001000001",
  26867=>"010101010",
  26868=>"001100100",
  26869=>"100110010",
  26870=>"101011001",
  26871=>"000110000",
  26872=>"100101110",
  26873=>"100011110",
  26874=>"001010011",
  26875=>"000011110",
  26876=>"111001111",
  26877=>"000011101",
  26878=>"111101111",
  26879=>"000001001",
  26880=>"110111101",
  26881=>"100100000",
  26882=>"101010010",
  26883=>"010110101",
  26884=>"000111001",
  26885=>"000011110",
  26886=>"010111011",
  26887=>"100100001",
  26888=>"100100100",
  26889=>"001100100",
  26890=>"100100110",
  26891=>"101101100",
  26892=>"111010100",
  26893=>"000111111",
  26894=>"001111001",
  26895=>"111111110",
  26896=>"110011000",
  26897=>"001100011",
  26898=>"010111110",
  26899=>"000101000",
  26900=>"100001001",
  26901=>"111011010",
  26902=>"011000010",
  26903=>"001101011",
  26904=>"001111111",
  26905=>"000000010",
  26906=>"000111101",
  26907=>"110111011",
  26908=>"001100010",
  26909=>"010101100",
  26910=>"011000011",
  26911=>"100101010",
  26912=>"101001001",
  26913=>"010101000",
  26914=>"101000100",
  26915=>"110100100",
  26916=>"110110100",
  26917=>"111000111",
  26918=>"011001101",
  26919=>"000110110",
  26920=>"100000100",
  26921=>"001100010",
  26922=>"111111001",
  26923=>"000011100",
  26924=>"111001110",
  26925=>"000001001",
  26926=>"000100010",
  26927=>"010010110",
  26928=>"101000001",
  26929=>"001001100",
  26930=>"100100111",
  26931=>"110111110",
  26932=>"011111010",
  26933=>"000111000",
  26934=>"000111000",
  26935=>"000101011",
  26936=>"001000001",
  26937=>"010000110",
  26938=>"000101011",
  26939=>"011111010",
  26940=>"001000101",
  26941=>"011001010",
  26942=>"000101001",
  26943=>"010101100",
  26944=>"000100000",
  26945=>"010011011",
  26946=>"000001001",
  26947=>"010000000",
  26948=>"001011100",
  26949=>"010000001",
  26950=>"010101100",
  26951=>"010111001",
  26952=>"000110101",
  26953=>"001011011",
  26954=>"011010110",
  26955=>"111001001",
  26956=>"100011011",
  26957=>"110100010",
  26958=>"001110011",
  26959=>"000110011",
  26960=>"100110010",
  26961=>"101010001",
  26962=>"000001000",
  26963=>"000000010",
  26964=>"100000011",
  26965=>"011101000",
  26966=>"100010110",
  26967=>"000110101",
  26968=>"000100101",
  26969=>"101110000",
  26970=>"011100110",
  26971=>"110010101",
  26972=>"000101100",
  26973=>"100100110",
  26974=>"111100011",
  26975=>"000011000",
  26976=>"110010000",
  26977=>"000011010",
  26978=>"010001101",
  26979=>"100101001",
  26980=>"011100010",
  26981=>"011101110",
  26982=>"111110111",
  26983=>"110001000",
  26984=>"001011011",
  26985=>"101100010",
  26986=>"111001101",
  26987=>"101100111",
  26988=>"010101101",
  26989=>"011000100",
  26990=>"000000001",
  26991=>"001010011",
  26992=>"100111000",
  26993=>"101100010",
  26994=>"010100101",
  26995=>"010101101",
  26996=>"110000101",
  26997=>"100011011",
  26998=>"010010100",
  26999=>"100010001",
  27000=>"011110100",
  27001=>"100101101",
  27002=>"000010010",
  27003=>"000100100",
  27004=>"010100111",
  27005=>"110010011",
  27006=>"101011110",
  27007=>"001000110",
  27008=>"110101100",
  27009=>"011110011",
  27010=>"010011110",
  27011=>"101000011",
  27012=>"110110111",
  27013=>"111101100",
  27014=>"000111010",
  27015=>"011101000",
  27016=>"010010000",
  27017=>"100010100",
  27018=>"011011010",
  27019=>"011111100",
  27020=>"000100010",
  27021=>"100111101",
  27022=>"010111001",
  27023=>"111010001",
  27024=>"001010101",
  27025=>"000001001",
  27026=>"111001110",
  27027=>"001010111",
  27028=>"101101010",
  27029=>"101101101",
  27030=>"010001000",
  27031=>"000110110",
  27032=>"011110100",
  27033=>"011100000",
  27034=>"010100100",
  27035=>"110000010",
  27036=>"101111001",
  27037=>"001101001",
  27038=>"101001011",
  27039=>"111110011",
  27040=>"011101111",
  27041=>"010100100",
  27042=>"111001010",
  27043=>"000001101",
  27044=>"011011011",
  27045=>"010001000",
  27046=>"010101011",
  27047=>"110101111",
  27048=>"011101001",
  27049=>"111001001",
  27050=>"100101110",
  27051=>"110010000",
  27052=>"110110010",
  27053=>"100110000",
  27054=>"100010001",
  27055=>"110100001",
  27056=>"101010110",
  27057=>"111110011",
  27058=>"000111010",
  27059=>"000111010",
  27060=>"100000011",
  27061=>"011001011",
  27062=>"000100000",
  27063=>"110010001",
  27064=>"001111111",
  27065=>"000001001",
  27066=>"000000101",
  27067=>"011010111",
  27068=>"110001100",
  27069=>"000011111",
  27070=>"100011000",
  27071=>"010010110",
  27072=>"000000010",
  27073=>"000010000",
  27074=>"011101101",
  27075=>"010011100",
  27076=>"110010010",
  27077=>"101010101",
  27078=>"011000000",
  27079=>"101100100",
  27080=>"010000101",
  27081=>"001100010",
  27082=>"100000100",
  27083=>"111100001",
  27084=>"000111100",
  27085=>"000101010",
  27086=>"000000101",
  27087=>"001110100",
  27088=>"100101000",
  27089=>"001010100",
  27090=>"111001010",
  27091=>"101100001",
  27092=>"001010010",
  27093=>"000110110",
  27094=>"101110011",
  27095=>"011100101",
  27096=>"011000011",
  27097=>"010001011",
  27098=>"100110010",
  27099=>"101011100",
  27100=>"001110001",
  27101=>"110001110",
  27102=>"000111111",
  27103=>"000111001",
  27104=>"101011001",
  27105=>"011110110",
  27106=>"101111000",
  27107=>"001111110",
  27108=>"000010100",
  27109=>"101010011",
  27110=>"100100000",
  27111=>"111000000",
  27112=>"010111111",
  27113=>"110001001",
  27114=>"100101100",
  27115=>"010001101",
  27116=>"111100011",
  27117=>"011011010",
  27118=>"001000010",
  27119=>"000101100",
  27120=>"111011110",
  27121=>"111111010",
  27122=>"001000011",
  27123=>"110101000",
  27124=>"100001101",
  27125=>"011111101",
  27126=>"111100011",
  27127=>"100001001",
  27128=>"111001110",
  27129=>"111100001",
  27130=>"100000101",
  27131=>"101101000",
  27132=>"100011000",
  27133=>"110011000",
  27134=>"101110000",
  27135=>"011011001",
  27136=>"100111011",
  27137=>"001100110",
  27138=>"111110100",
  27139=>"000001000",
  27140=>"000111111",
  27141=>"110110011",
  27142=>"111110010",
  27143=>"101000111",
  27144=>"111000000",
  27145=>"011010010",
  27146=>"010110010",
  27147=>"010000000",
  27148=>"011001011",
  27149=>"100111111",
  27150=>"111100000",
  27151=>"001100100",
  27152=>"011110010",
  27153=>"000110010",
  27154=>"011101000",
  27155=>"111100100",
  27156=>"000001011",
  27157=>"100000110",
  27158=>"101010101",
  27159=>"001100101",
  27160=>"000111000",
  27161=>"001111010",
  27162=>"110010000",
  27163=>"101101001",
  27164=>"100100101",
  27165=>"111011000",
  27166=>"111011000",
  27167=>"000011010",
  27168=>"000000000",
  27169=>"010110101",
  27170=>"000001110",
  27171=>"011101010",
  27172=>"111101010",
  27173=>"110011000",
  27174=>"101011101",
  27175=>"100111001",
  27176=>"011000100",
  27177=>"011011010",
  27178=>"111101101",
  27179=>"100101010",
  27180=>"110110001",
  27181=>"101110000",
  27182=>"000101010",
  27183=>"000010000",
  27184=>"100000110",
  27185=>"101111001",
  27186=>"010000010",
  27187=>"100011011",
  27188=>"001100101",
  27189=>"001000101",
  27190=>"000011110",
  27191=>"010000001",
  27192=>"011110100",
  27193=>"000101010",
  27194=>"011001001",
  27195=>"101101000",
  27196=>"011011010",
  27197=>"101000100",
  27198=>"011001100",
  27199=>"111110100",
  27200=>"110100000",
  27201=>"101001100",
  27202=>"100010101",
  27203=>"011110101",
  27204=>"111000000",
  27205=>"101110001",
  27206=>"011001000",
  27207=>"000101101",
  27208=>"100001011",
  27209=>"001101001",
  27210=>"011010110",
  27211=>"011010100",
  27212=>"000110111",
  27213=>"001000100",
  27214=>"000011111",
  27215=>"101011011",
  27216=>"000100110",
  27217=>"011110101",
  27218=>"110011010",
  27219=>"010100101",
  27220=>"101111101",
  27221=>"100100101",
  27222=>"001011101",
  27223=>"110111000",
  27224=>"100001111",
  27225=>"100101000",
  27226=>"001101010",
  27227=>"000001100",
  27228=>"001010011",
  27229=>"001100001",
  27230=>"001110011",
  27231=>"011001001",
  27232=>"111001001",
  27233=>"110100011",
  27234=>"111101111",
  27235=>"010010100",
  27236=>"010010100",
  27237=>"111101011",
  27238=>"110110010",
  27239=>"000010101",
  27240=>"000100111",
  27241=>"001000100",
  27242=>"100101011",
  27243=>"001111000",
  27244=>"000010111",
  27245=>"001011001",
  27246=>"111011000",
  27247=>"001001010",
  27248=>"100000011",
  27249=>"000011100",
  27250=>"011011000",
  27251=>"101000100",
  27252=>"100100100",
  27253=>"010110000",
  27254=>"100101111",
  27255=>"111111110",
  27256=>"111100010",
  27257=>"110111111",
  27258=>"110010101",
  27259=>"101110011",
  27260=>"100100001",
  27261=>"011010001",
  27262=>"110110000",
  27263=>"110000101",
  27264=>"111111011",
  27265=>"001011000",
  27266=>"110001001",
  27267=>"100001001",
  27268=>"110010010",
  27269=>"101100001",
  27270=>"101110001",
  27271=>"100000110",
  27272=>"110000000",
  27273=>"101100100",
  27274=>"100110011",
  27275=>"000000111",
  27276=>"011101000",
  27277=>"100100010",
  27278=>"100110101",
  27279=>"010010000",
  27280=>"011001101",
  27281=>"001010000",
  27282=>"011111011",
  27283=>"101111111",
  27284=>"000110010",
  27285=>"000001100",
  27286=>"100010011",
  27287=>"111100111",
  27288=>"101011010",
  27289=>"000101001",
  27290=>"001100010",
  27291=>"010010111",
  27292=>"100111001",
  27293=>"000011011",
  27294=>"011001010",
  27295=>"000000010",
  27296=>"001110010",
  27297=>"110100101",
  27298=>"010101001",
  27299=>"000101001",
  27300=>"010010101",
  27301=>"000110110",
  27302=>"110101110",
  27303=>"011000001",
  27304=>"001101000",
  27305=>"010000100",
  27306=>"110000000",
  27307=>"011010110",
  27308=>"101011011",
  27309=>"110001110",
  27310=>"111000010",
  27311=>"110000101",
  27312=>"000001110",
  27313=>"001000101",
  27314=>"010101100",
  27315=>"110000000",
  27316=>"010000011",
  27317=>"111001111",
  27318=>"100100000",
  27319=>"111011000",
  27320=>"110001001",
  27321=>"101111110",
  27322=>"100011011",
  27323=>"100011001",
  27324=>"100100010",
  27325=>"000000101",
  27326=>"001000000",
  27327=>"000111001",
  27328=>"111100101",
  27329=>"101100110",
  27330=>"000100000",
  27331=>"011011011",
  27332=>"110000101",
  27333=>"110001100",
  27334=>"010100101",
  27335=>"001000001",
  27336=>"100100000",
  27337=>"101001101",
  27338=>"110101001",
  27339=>"100010011",
  27340=>"011110110",
  27341=>"011100010",
  27342=>"001011011",
  27343=>"100011101",
  27344=>"011000100",
  27345=>"100000101",
  27346=>"111101000",
  27347=>"001101111",
  27348=>"110000011",
  27349=>"001010111",
  27350=>"011110011",
  27351=>"000001000",
  27352=>"001010101",
  27353=>"111000010",
  27354=>"001110011",
  27355=>"100111111",
  27356=>"101101101",
  27357=>"000011001",
  27358=>"100001000",
  27359=>"011111101",
  27360=>"101000011",
  27361=>"001110000",
  27362=>"111110110",
  27363=>"000001010",
  27364=>"000010000",
  27365=>"011100000",
  27366=>"001100000",
  27367=>"101010010",
  27368=>"001100101",
  27369=>"000000011",
  27370=>"001101100",
  27371=>"000000011",
  27372=>"001010100",
  27373=>"000110100",
  27374=>"010100111",
  27375=>"000000100",
  27376=>"001001010",
  27377=>"000100100",
  27378=>"001010111",
  27379=>"110010010",
  27380=>"001010101",
  27381=>"101011010",
  27382=>"000001101",
  27383=>"010010100",
  27384=>"110111100",
  27385=>"001110000",
  27386=>"111010111",
  27387=>"001011001",
  27388=>"001011011",
  27389=>"011100000",
  27390=>"101101100",
  27391=>"010010110",
  27392=>"100111001",
  27393=>"110111001",
  27394=>"000111010",
  27395=>"000000001",
  27396=>"010110001",
  27397=>"010110101",
  27398=>"010010110",
  27399=>"100101000",
  27400=>"011010010",
  27401=>"111100010",
  27402=>"101100010",
  27403=>"000000011",
  27404=>"001010010",
  27405=>"011111110",
  27406=>"011110111",
  27407=>"110100110",
  27408=>"001011100",
  27409=>"111100111",
  27410=>"111000001",
  27411=>"101001100",
  27412=>"100100000",
  27413=>"011010101",
  27414=>"010010101",
  27415=>"111101000",
  27416=>"000000101",
  27417=>"100110110",
  27418=>"000000001",
  27419=>"011010010",
  27420=>"110000101",
  27421=>"110100010",
  27422=>"010111010",
  27423=>"000011111",
  27424=>"001101001",
  27425=>"110111100",
  27426=>"110000011",
  27427=>"101000001",
  27428=>"001110001",
  27429=>"110011011",
  27430=>"010011111",
  27431=>"001001010",
  27432=>"010010010",
  27433=>"111101011",
  27434=>"000000001",
  27435=>"011100100",
  27436=>"001001010",
  27437=>"011001110",
  27438=>"001100000",
  27439=>"100101111",
  27440=>"011001010",
  27441=>"000110000",
  27442=>"011100001",
  27443=>"100110100",
  27444=>"000100110",
  27445=>"001110100",
  27446=>"000000111",
  27447=>"001110100",
  27448=>"001011001",
  27449=>"010000110",
  27450=>"110011110",
  27451=>"001001110",
  27452=>"011000011",
  27453=>"001110010",
  27454=>"110110000",
  27455=>"000110010",
  27456=>"110001001",
  27457=>"101101001",
  27458=>"110010101",
  27459=>"100100110",
  27460=>"111000010",
  27461=>"111011010",
  27462=>"100011110",
  27463=>"111001010",
  27464=>"010101010",
  27465=>"010000000",
  27466=>"101101111",
  27467=>"000110110",
  27468=>"110011001",
  27469=>"000001010",
  27470=>"111001110",
  27471=>"010101001",
  27472=>"101110100",
  27473=>"100101110",
  27474=>"111010001",
  27475=>"011000001",
  27476=>"101010110",
  27477=>"101110101",
  27478=>"001100101",
  27479=>"111110001",
  27480=>"100001111",
  27481=>"111110001",
  27482=>"111111000",
  27483=>"100001100",
  27484=>"100001010",
  27485=>"000000100",
  27486=>"110101010",
  27487=>"011001010",
  27488=>"001101000",
  27489=>"100110011",
  27490=>"000000011",
  27491=>"001011000",
  27492=>"011011111",
  27493=>"111111001",
  27494=>"000011000",
  27495=>"100011111",
  27496=>"000000010",
  27497=>"010101001",
  27498=>"111001000",
  27499=>"011101001",
  27500=>"111110110",
  27501=>"111110011",
  27502=>"000001000",
  27503=>"110100110",
  27504=>"101000011",
  27505=>"110111101",
  27506=>"000001101",
  27507=>"010010111",
  27508=>"000110000",
  27509=>"111111000",
  27510=>"010111010",
  27511=>"001011111",
  27512=>"011110000",
  27513=>"000010101",
  27514=>"011011010",
  27515=>"010010111",
  27516=>"000000010",
  27517=>"101111100",
  27518=>"110011011",
  27519=>"011001010",
  27520=>"001000010",
  27521=>"111000001",
  27522=>"001011101",
  27523=>"010011001",
  27524=>"101100000",
  27525=>"000011011",
  27526=>"101101010",
  27527=>"101111001",
  27528=>"110001110",
  27529=>"001100110",
  27530=>"100010111",
  27531=>"100110110",
  27532=>"001010011",
  27533=>"111101101",
  27534=>"111100000",
  27535=>"011110111",
  27536=>"000111001",
  27537=>"000110001",
  27538=>"101101000",
  27539=>"010110000",
  27540=>"010110110",
  27541=>"111100000",
  27542=>"100001001",
  27543=>"110111001",
  27544=>"000100011",
  27545=>"100000110",
  27546=>"100110011",
  27547=>"010001101",
  27548=>"111010011",
  27549=>"110000110",
  27550=>"111001100",
  27551=>"010101111",
  27552=>"111010111",
  27553=>"100001110",
  27554=>"100101110",
  27555=>"101001001",
  27556=>"010101111",
  27557=>"100000111",
  27558=>"001000110",
  27559=>"011001100",
  27560=>"011010000",
  27561=>"100000111",
  27562=>"011001111",
  27563=>"001011011",
  27564=>"001100100",
  27565=>"001010010",
  27566=>"101011000",
  27567=>"100110000",
  27568=>"001010101",
  27569=>"101010001",
  27570=>"100001110",
  27571=>"111000001",
  27572=>"111111001",
  27573=>"001001110",
  27574=>"111011101",
  27575=>"110101010",
  27576=>"001101011",
  27577=>"000100010",
  27578=>"010111000",
  27579=>"110010111",
  27580=>"101110100",
  27581=>"101110011",
  27582=>"011000001",
  27583=>"111000000",
  27584=>"000111101",
  27585=>"110110001",
  27586=>"001011000",
  27587=>"110010111",
  27588=>"100000011",
  27589=>"011010100",
  27590=>"101110001",
  27591=>"101011011",
  27592=>"000000011",
  27593=>"111100001",
  27594=>"110100111",
  27595=>"101011000",
  27596=>"111001011",
  27597=>"000010000",
  27598=>"101111000",
  27599=>"110001111",
  27600=>"111100110",
  27601=>"100001111",
  27602=>"001100001",
  27603=>"100110101",
  27604=>"100000101",
  27605=>"110000000",
  27606=>"101001111",
  27607=>"101100100",
  27608=>"000000111",
  27609=>"101010100",
  27610=>"010010001",
  27611=>"001110001",
  27612=>"101100001",
  27613=>"100110110",
  27614=>"011001010",
  27615=>"111100101",
  27616=>"110001100",
  27617=>"101101001",
  27618=>"011011000",
  27619=>"010001000",
  27620=>"110110111",
  27621=>"010010111",
  27622=>"010100001",
  27623=>"011000101",
  27624=>"000111001",
  27625=>"001011001",
  27626=>"100001110",
  27627=>"000101001",
  27628=>"101011110",
  27629=>"011100001",
  27630=>"100100111",
  27631=>"111010000",
  27632=>"000100100",
  27633=>"100001111",
  27634=>"011101100",
  27635=>"101011010",
  27636=>"010101011",
  27637=>"111010001",
  27638=>"110110110",
  27639=>"000010101",
  27640=>"001000110",
  27641=>"010000001",
  27642=>"010101101",
  27643=>"000011001",
  27644=>"101100001",
  27645=>"000011000",
  27646=>"001010011",
  27647=>"100110000",
  27648=>"101100101",
  27649=>"000111010",
  27650=>"100010010",
  27651=>"111000100",
  27652=>"010100001",
  27653=>"111001001",
  27654=>"101100001",
  27655=>"001101000",
  27656=>"000000100",
  27657=>"100011101",
  27658=>"110010011",
  27659=>"111000000",
  27660=>"101111111",
  27661=>"110101011",
  27662=>"100100001",
  27663=>"010100011",
  27664=>"111100011",
  27665=>"111101011",
  27666=>"101010001",
  27667=>"100000000",
  27668=>"100101000",
  27669=>"100001000",
  27670=>"111001000",
  27671=>"000101011",
  27672=>"110010010",
  27673=>"011001100",
  27674=>"110001100",
  27675=>"000000001",
  27676=>"110010001",
  27677=>"010010010",
  27678=>"000111101",
  27679=>"110000110",
  27680=>"010010001",
  27681=>"011111101",
  27682=>"001010101",
  27683=>"000000110",
  27684=>"100101001",
  27685=>"100010100",
  27686=>"010111100",
  27687=>"011010000",
  27688=>"011001111",
  27689=>"101011111",
  27690=>"011011010",
  27691=>"001011000",
  27692=>"111111010",
  27693=>"100000100",
  27694=>"001100010",
  27695=>"000011100",
  27696=>"100010100",
  27697=>"111100111",
  27698=>"000000000",
  27699=>"011110110",
  27700=>"100011010",
  27701=>"001100011",
  27702=>"110001000",
  27703=>"001010000",
  27704=>"001011010",
  27705=>"101001111",
  27706=>"000010010",
  27707=>"001001101",
  27708=>"110001101",
  27709=>"000111010",
  27710=>"100101011",
  27711=>"110010100",
  27712=>"000001000",
  27713=>"011101101",
  27714=>"011001000",
  27715=>"110100011",
  27716=>"110001111",
  27717=>"001011101",
  27718=>"011011110",
  27719=>"011001010",
  27720=>"111110101",
  27721=>"010101110",
  27722=>"101010010",
  27723=>"000011111",
  27724=>"001000000",
  27725=>"100101100",
  27726=>"110110110",
  27727=>"111011010",
  27728=>"111101101",
  27729=>"000111101",
  27730=>"010010001",
  27731=>"001101011",
  27732=>"010100010",
  27733=>"110010111",
  27734=>"001010100",
  27735=>"000001101",
  27736=>"111111010",
  27737=>"000001010",
  27738=>"011011100",
  27739=>"011100000",
  27740=>"010000101",
  27741=>"100001011",
  27742=>"101001000",
  27743=>"101001011",
  27744=>"111100001",
  27745=>"100111000",
  27746=>"001111011",
  27747=>"011100000",
  27748=>"101000110",
  27749=>"100010101",
  27750=>"011011001",
  27751=>"101010000",
  27752=>"011010010",
  27753=>"111000011",
  27754=>"100110100",
  27755=>"100110110",
  27756=>"001000110",
  27757=>"110110110",
  27758=>"000101000",
  27759=>"101000010",
  27760=>"000100111",
  27761=>"111001010",
  27762=>"110000001",
  27763=>"011101110",
  27764=>"111111011",
  27765=>"011011011",
  27766=>"100000100",
  27767=>"111010011",
  27768=>"100101011",
  27769=>"111011100",
  27770=>"100100100",
  27771=>"101111110",
  27772=>"111111010",
  27773=>"110010000",
  27774=>"101111111",
  27775=>"100111100",
  27776=>"010000101",
  27777=>"000110001",
  27778=>"100011010",
  27779=>"001110101",
  27780=>"110011100",
  27781=>"101101111",
  27782=>"011100111",
  27783=>"011111000",
  27784=>"111100110",
  27785=>"111001011",
  27786=>"011101100",
  27787=>"011111011",
  27788=>"101101011",
  27789=>"011110111",
  27790=>"110000111",
  27791=>"001011110",
  27792=>"111010110",
  27793=>"010001001",
  27794=>"111101001",
  27795=>"000011101",
  27796=>"000100100",
  27797=>"111100110",
  27798=>"001000000",
  27799=>"100111101",
  27800=>"000011110",
  27801=>"000010101",
  27802=>"000001010",
  27803=>"111011001",
  27804=>"001000001",
  27805=>"100010110",
  27806=>"010111011",
  27807=>"001101010",
  27808=>"001010001",
  27809=>"100010001",
  27810=>"011100101",
  27811=>"110101111",
  27812=>"001010101",
  27813=>"101110110",
  27814=>"101011001",
  27815=>"011111111",
  27816=>"111000011",
  27817=>"011111001",
  27818=>"100101001",
  27819=>"010011011",
  27820=>"011000100",
  27821=>"110101110",
  27822=>"101010111",
  27823=>"000010001",
  27824=>"111100101",
  27825=>"101011111",
  27826=>"000010110",
  27827=>"010000010",
  27828=>"001101000",
  27829=>"000111010",
  27830=>"110000010",
  27831=>"000111011",
  27832=>"001000100",
  27833=>"100100011",
  27834=>"000001001",
  27835=>"111001010",
  27836=>"111001011",
  27837=>"100010011",
  27838=>"000000110",
  27839=>"101110010",
  27840=>"000111100",
  27841=>"111101101",
  27842=>"100111100",
  27843=>"100010000",
  27844=>"010110100",
  27845=>"000000000",
  27846=>"011110101",
  27847=>"111011100",
  27848=>"001110110",
  27849=>"000011100",
  27850=>"111010011",
  27851=>"100000000",
  27852=>"000101010",
  27853=>"001101010",
  27854=>"010111010",
  27855=>"000101011",
  27856=>"110001111",
  27857=>"001101000",
  27858=>"100100001",
  27859=>"101110011",
  27860=>"011001111",
  27861=>"000010111",
  27862=>"001101011",
  27863=>"100000100",
  27864=>"100000010",
  27865=>"111111001",
  27866=>"011101000",
  27867=>"000110111",
  27868=>"001000011",
  27869=>"100101111",
  27870=>"110100111",
  27871=>"111111101",
  27872=>"001001101",
  27873=>"110100111",
  27874=>"111111011",
  27875=>"101100110",
  27876=>"011100111",
  27877=>"000000110",
  27878=>"010111111",
  27879=>"101000100",
  27880=>"011100001",
  27881=>"111101110",
  27882=>"011000100",
  27883=>"101001101",
  27884=>"101010101",
  27885=>"111100101",
  27886=>"110111001",
  27887=>"111101001",
  27888=>"011111101",
  27889=>"101101101",
  27890=>"101100010",
  27891=>"001100101",
  27892=>"010110000",
  27893=>"001000110",
  27894=>"010110001",
  27895=>"001001010",
  27896=>"011111011",
  27897=>"111100010",
  27898=>"101011010",
  27899=>"000001001",
  27900=>"111101101",
  27901=>"000001100",
  27902=>"110100101",
  27903=>"010001011",
  27904=>"011111110",
  27905=>"011001101",
  27906=>"001110101",
  27907=>"100001111",
  27908=>"101110001",
  27909=>"010110110",
  27910=>"010000110",
  27911=>"100001100",
  27912=>"010110100",
  27913=>"010111010",
  27914=>"111000001",
  27915=>"001001101",
  27916=>"000001000",
  27917=>"000011110",
  27918=>"100000000",
  27919=>"100000101",
  27920=>"110010000",
  27921=>"011110110",
  27922=>"011110000",
  27923=>"101011011",
  27924=>"101111111",
  27925=>"110011110",
  27926=>"010010000",
  27927=>"110110001",
  27928=>"101000000",
  27929=>"000100111",
  27930=>"101111110",
  27931=>"011111110",
  27932=>"001110101",
  27933=>"101101100",
  27934=>"000101010",
  27935=>"010011010",
  27936=>"101001100",
  27937=>"001011001",
  27938=>"101011000",
  27939=>"001110011",
  27940=>"110000001",
  27941=>"001000101",
  27942=>"111100111",
  27943=>"011111111",
  27944=>"100000001",
  27945=>"000110100",
  27946=>"101000000",
  27947=>"011010000",
  27948=>"101101110",
  27949=>"000111001",
  27950=>"101101101",
  27951=>"101001111",
  27952=>"001011101",
  27953=>"000010010",
  27954=>"011110011",
  27955=>"100100011",
  27956=>"010110100",
  27957=>"010110001",
  27958=>"111010101",
  27959=>"111110010",
  27960=>"101010111",
  27961=>"110111000",
  27962=>"101110010",
  27963=>"101101000",
  27964=>"101111101",
  27965=>"101100010",
  27966=>"101010010",
  27967=>"101101111",
  27968=>"101010010",
  27969=>"000000000",
  27970=>"000011011",
  27971=>"100010111",
  27972=>"001101101",
  27973=>"000010000",
  27974=>"001110100",
  27975=>"110100010",
  27976=>"011110001",
  27977=>"101101000",
  27978=>"111011000",
  27979=>"010111011",
  27980=>"011100110",
  27981=>"000100101",
  27982=>"000110011",
  27983=>"011100001",
  27984=>"110001001",
  27985=>"110011111",
  27986=>"010010011",
  27987=>"100000000",
  27988=>"001001000",
  27989=>"011101011",
  27990=>"100111111",
  27991=>"101010110",
  27992=>"000000001",
  27993=>"110000010",
  27994=>"101010111",
  27995=>"110110001",
  27996=>"001100001",
  27997=>"111101001",
  27998=>"011110001",
  27999=>"000000100",
  28000=>"001010101",
  28001=>"111011100",
  28002=>"000011010",
  28003=>"110001111",
  28004=>"010100000",
  28005=>"111111011",
  28006=>"111001001",
  28007=>"001000010",
  28008=>"011010011",
  28009=>"000100101",
  28010=>"010000101",
  28011=>"101010000",
  28012=>"011010111",
  28013=>"000001010",
  28014=>"100100001",
  28015=>"000011001",
  28016=>"101011011",
  28017=>"011000110",
  28018=>"011010000",
  28019=>"010010011",
  28020=>"000001000",
  28021=>"101111111",
  28022=>"011000000",
  28023=>"111011101",
  28024=>"000111111",
  28025=>"010010111",
  28026=>"100101011",
  28027=>"111000001",
  28028=>"101110011",
  28029=>"010001001",
  28030=>"101110010",
  28031=>"000011100",
  28032=>"100111011",
  28033=>"111110001",
  28034=>"011111101",
  28035=>"011111100",
  28036=>"110111001",
  28037=>"001110000",
  28038=>"100010001",
  28039=>"100011000",
  28040=>"010100110",
  28041=>"110111000",
  28042=>"001000000",
  28043=>"111010111",
  28044=>"000000001",
  28045=>"001000000",
  28046=>"101000110",
  28047=>"110110110",
  28048=>"101101110",
  28049=>"111000100",
  28050=>"000101111",
  28051=>"011111000",
  28052=>"010011100",
  28053=>"110000010",
  28054=>"000011010",
  28055=>"100100000",
  28056=>"110101000",
  28057=>"111001001",
  28058=>"010000100",
  28059=>"101100110",
  28060=>"101111111",
  28061=>"111111110",
  28062=>"000111011",
  28063=>"010100000",
  28064=>"110101111",
  28065=>"111101111",
  28066=>"010011101",
  28067=>"011001111",
  28068=>"011010100",
  28069=>"000110111",
  28070=>"001011011",
  28071=>"101110011",
  28072=>"100011000",
  28073=>"100001010",
  28074=>"010111100",
  28075=>"101011110",
  28076=>"000110001",
  28077=>"111110001",
  28078=>"101110101",
  28079=>"000111010",
  28080=>"011000101",
  28081=>"100110010",
  28082=>"000111010",
  28083=>"101111101",
  28084=>"100000110",
  28085=>"100111000",
  28086=>"101100100",
  28087=>"010101010",
  28088=>"001100011",
  28089=>"100011011",
  28090=>"000101011",
  28091=>"111011011",
  28092=>"111011011",
  28093=>"001010001",
  28094=>"101110000",
  28095=>"000110100",
  28096=>"010010001",
  28097=>"001111110",
  28098=>"001000110",
  28099=>"011000010",
  28100=>"110111110",
  28101=>"100100110",
  28102=>"000101011",
  28103=>"101111011",
  28104=>"001101101",
  28105=>"101110001",
  28106=>"111100011",
  28107=>"110000101",
  28108=>"111110011",
  28109=>"000011101",
  28110=>"101101110",
  28111=>"010001111",
  28112=>"100011110",
  28113=>"011010101",
  28114=>"111110101",
  28115=>"111111110",
  28116=>"001111010",
  28117=>"110110010",
  28118=>"000101010",
  28119=>"100011101",
  28120=>"111111100",
  28121=>"101000001",
  28122=>"010101001",
  28123=>"010100111",
  28124=>"010100100",
  28125=>"010111000",
  28126=>"011111111",
  28127=>"000111110",
  28128=>"011000100",
  28129=>"001010000",
  28130=>"100000000",
  28131=>"000100010",
  28132=>"100010111",
  28133=>"111111110",
  28134=>"000100111",
  28135=>"010100110",
  28136=>"010000111",
  28137=>"010010111",
  28138=>"001111011",
  28139=>"010101101",
  28140=>"101111011",
  28141=>"110011111",
  28142=>"010101110",
  28143=>"111111000",
  28144=>"100011111",
  28145=>"011010001",
  28146=>"110000010",
  28147=>"001101110",
  28148=>"110110010",
  28149=>"101001100",
  28150=>"110000111",
  28151=>"000111111",
  28152=>"111001111",
  28153=>"001100100",
  28154=>"010100010",
  28155=>"001101000",
  28156=>"001100100",
  28157=>"011111111",
  28158=>"111111111",
  28159=>"111111110",
  28160=>"010110011",
  28161=>"111110110",
  28162=>"101011111",
  28163=>"101100001",
  28164=>"100100001",
  28165=>"011100011",
  28166=>"011100001",
  28167=>"011001000",
  28168=>"010001010",
  28169=>"000001100",
  28170=>"100110010",
  28171=>"011001111",
  28172=>"100101101",
  28173=>"100101010",
  28174=>"110111100",
  28175=>"011101010",
  28176=>"110101110",
  28177=>"000001100",
  28178=>"000000000",
  28179=>"000000110",
  28180=>"110110101",
  28181=>"110100111",
  28182=>"001110011",
  28183=>"010001101",
  28184=>"101100001",
  28185=>"001001110",
  28186=>"010101110",
  28187=>"000000111",
  28188=>"011101100",
  28189=>"100010010",
  28190=>"001011100",
  28191=>"000010111",
  28192=>"100011010",
  28193=>"011000100",
  28194=>"000100011",
  28195=>"110000110",
  28196=>"011111101",
  28197=>"110001000",
  28198=>"100011100",
  28199=>"001011010",
  28200=>"100110011",
  28201=>"001010101",
  28202=>"000111001",
  28203=>"000011010",
  28204=>"110011101",
  28205=>"110101110",
  28206=>"100110010",
  28207=>"111001111",
  28208=>"100000000",
  28209=>"010011000",
  28210=>"101101110",
  28211=>"001000001",
  28212=>"100000001",
  28213=>"010011001",
  28214=>"100011101",
  28215=>"011101001",
  28216=>"011011011",
  28217=>"110110111",
  28218=>"000011111",
  28219=>"011000000",
  28220=>"101100110",
  28221=>"100110100",
  28222=>"001011011",
  28223=>"111100101",
  28224=>"011000000",
  28225=>"000011010",
  28226=>"100011010",
  28227=>"000000011",
  28228=>"001001110",
  28229=>"010000010",
  28230=>"000100001",
  28231=>"000101000",
  28232=>"100100011",
  28233=>"111001010",
  28234=>"010000001",
  28235=>"011101100",
  28236=>"111101111",
  28237=>"000100100",
  28238=>"010000110",
  28239=>"110011101",
  28240=>"101100001",
  28241=>"101101000",
  28242=>"100100101",
  28243=>"000000101",
  28244=>"110000000",
  28245=>"001100111",
  28246=>"001011100",
  28247=>"011011001",
  28248=>"110000010",
  28249=>"011110010",
  28250=>"001000000",
  28251=>"110101010",
  28252=>"011001010",
  28253=>"100001100",
  28254=>"000001000",
  28255=>"010001011",
  28256=>"101001001",
  28257=>"000000001",
  28258=>"110110111",
  28259=>"101010010",
  28260=>"111011101",
  28261=>"110000010",
  28262=>"110110101",
  28263=>"001001010",
  28264=>"100100000",
  28265=>"100100011",
  28266=>"010010001",
  28267=>"100000001",
  28268=>"100101011",
  28269=>"010000000",
  28270=>"110101111",
  28271=>"100011111",
  28272=>"010110001",
  28273=>"000001110",
  28274=>"011001011",
  28275=>"100011101",
  28276=>"011111101",
  28277=>"111110011",
  28278=>"000011000",
  28279=>"111001110",
  28280=>"111100010",
  28281=>"100100010",
  28282=>"100010110",
  28283=>"000111011",
  28284=>"110100110",
  28285=>"010010111",
  28286=>"111111001",
  28287=>"100011110",
  28288=>"000110111",
  28289=>"010001100",
  28290=>"101010001",
  28291=>"011010001",
  28292=>"001100010",
  28293=>"001111011",
  28294=>"001001100",
  28295=>"110101000",
  28296=>"101101001",
  28297=>"010110101",
  28298=>"010111100",
  28299=>"010001010",
  28300=>"000001100",
  28301=>"010110110",
  28302=>"101110100",
  28303=>"100100011",
  28304=>"100001001",
  28305=>"110101111",
  28306=>"111101101",
  28307=>"001000001",
  28308=>"011010111",
  28309=>"100010111",
  28310=>"111100000",
  28311=>"111011111",
  28312=>"000101001",
  28313=>"000110110",
  28314=>"100011010",
  28315=>"010001101",
  28316=>"001110010",
  28317=>"011001111",
  28318=>"111110110",
  28319=>"100000000",
  28320=>"011100101",
  28321=>"101010001",
  28322=>"000011010",
  28323=>"000011001",
  28324=>"110010111",
  28325=>"111101011",
  28326=>"011101110",
  28327=>"010000111",
  28328=>"111101101",
  28329=>"001001110",
  28330=>"010000101",
  28331=>"101011010",
  28332=>"000011111",
  28333=>"101010000",
  28334=>"110010100",
  28335=>"101011110",
  28336=>"000000001",
  28337=>"011001010",
  28338=>"011010101",
  28339=>"111000100",
  28340=>"101110101",
  28341=>"001101011",
  28342=>"101100010",
  28343=>"101000110",
  28344=>"010110111",
  28345=>"000011001",
  28346=>"010101111",
  28347=>"001000110",
  28348=>"101101101",
  28349=>"100011100",
  28350=>"001101110",
  28351=>"100100011",
  28352=>"111010011",
  28353=>"110010111",
  28354=>"100101111",
  28355=>"001010011",
  28356=>"001100110",
  28357=>"100111011",
  28358=>"110110011",
  28359=>"000001110",
  28360=>"000001011",
  28361=>"111010100",
  28362=>"000110010",
  28363=>"110010101",
  28364=>"001001110",
  28365=>"011011011",
  28366=>"011110011",
  28367=>"110110001",
  28368=>"001000001",
  28369=>"111110100",
  28370=>"010011011",
  28371=>"011001110",
  28372=>"010110100",
  28373=>"100100100",
  28374=>"011100111",
  28375=>"110011000",
  28376=>"011011111",
  28377=>"100111101",
  28378=>"111101000",
  28379=>"111011100",
  28380=>"101001101",
  28381=>"000000101",
  28382=>"000100010",
  28383=>"000011100",
  28384=>"110010111",
  28385=>"000110001",
  28386=>"000001011",
  28387=>"011110100",
  28388=>"000111010",
  28389=>"010010001",
  28390=>"101111001",
  28391=>"000101001",
  28392=>"100110010",
  28393=>"110010101",
  28394=>"000010011",
  28395=>"111001101",
  28396=>"111100101",
  28397=>"000001000",
  28398=>"010100011",
  28399=>"011111000",
  28400=>"001001110",
  28401=>"010110010",
  28402=>"011101110",
  28403=>"101001010",
  28404=>"101000010",
  28405=>"111100100",
  28406=>"000010111",
  28407=>"111111111",
  28408=>"011001100",
  28409=>"010110100",
  28410=>"001001010",
  28411=>"011000000",
  28412=>"101101011",
  28413=>"001111010",
  28414=>"000110010",
  28415=>"110001101",
  28416=>"100011101",
  28417=>"101011011",
  28418=>"000010101",
  28419=>"010011100",
  28420=>"101011110",
  28421=>"101010110",
  28422=>"100010110",
  28423=>"010100011",
  28424=>"101101100",
  28425=>"100111000",
  28426=>"010011110",
  28427=>"111110011",
  28428=>"100010010",
  28429=>"111011000",
  28430=>"011001000",
  28431=>"101000100",
  28432=>"001001001",
  28433=>"101011000",
  28434=>"110111001",
  28435=>"111110100",
  28436=>"100001001",
  28437=>"100001010",
  28438=>"011110100",
  28439=>"111010110",
  28440=>"111001001",
  28441=>"010110001",
  28442=>"010110000",
  28443=>"010000100",
  28444=>"110011101",
  28445=>"010001011",
  28446=>"011101110",
  28447=>"001010001",
  28448=>"100001101",
  28449=>"101000101",
  28450=>"000101101",
  28451=>"010000010",
  28452=>"000111010",
  28453=>"111001101",
  28454=>"000101111",
  28455=>"000001010",
  28456=>"000010010",
  28457=>"100101101",
  28458=>"101101010",
  28459=>"011000101",
  28460=>"101101000",
  28461=>"000011110",
  28462=>"111101001",
  28463=>"101110011",
  28464=>"101001101",
  28465=>"111101011",
  28466=>"101001011",
  28467=>"011110111",
  28468=>"110000110",
  28469=>"000111100",
  28470=>"101010010",
  28471=>"100101100",
  28472=>"101110111",
  28473=>"100101011",
  28474=>"111110011",
  28475=>"111100110",
  28476=>"111110000",
  28477=>"010110111",
  28478=>"110011010",
  28479=>"000100111",
  28480=>"110000110",
  28481=>"101101110",
  28482=>"111010100",
  28483=>"100100000",
  28484=>"111111101",
  28485=>"000110100",
  28486=>"011001001",
  28487=>"010000001",
  28488=>"111111001",
  28489=>"101101010",
  28490=>"111100111",
  28491=>"101100001",
  28492=>"011000000",
  28493=>"100000100",
  28494=>"011111111",
  28495=>"100010010",
  28496=>"101100001",
  28497=>"001101001",
  28498=>"110000100",
  28499=>"110000110",
  28500=>"011101110",
  28501=>"010101111",
  28502=>"000010010",
  28503=>"011111010",
  28504=>"001001110",
  28505=>"111000101",
  28506=>"111100111",
  28507=>"101111111",
  28508=>"111100100",
  28509=>"001011101",
  28510=>"111100001",
  28511=>"111100001",
  28512=>"111001001",
  28513=>"110111000",
  28514=>"010010101",
  28515=>"101001000",
  28516=>"110000101",
  28517=>"100111011",
  28518=>"011110111",
  28519=>"111110100",
  28520=>"000111110",
  28521=>"110011010",
  28522=>"001101110",
  28523=>"011011011",
  28524=>"100100110",
  28525=>"001010101",
  28526=>"000100100",
  28527=>"100001110",
  28528=>"110100111",
  28529=>"100011110",
  28530=>"000111100",
  28531=>"000001000",
  28532=>"100101110",
  28533=>"000010000",
  28534=>"100111100",
  28535=>"110101110",
  28536=>"010101111",
  28537=>"000111110",
  28538=>"100111000",
  28539=>"101001000",
  28540=>"101010101",
  28541=>"011011101",
  28542=>"001000111",
  28543=>"100110011",
  28544=>"100001011",
  28545=>"101000001",
  28546=>"000001011",
  28547=>"001110111",
  28548=>"110111101",
  28549=>"000111001",
  28550=>"101010000",
  28551=>"011101010",
  28552=>"111110001",
  28553=>"010110000",
  28554=>"111111101",
  28555=>"111011111",
  28556=>"111100110",
  28557=>"001000001",
  28558=>"000100110",
  28559=>"011111001",
  28560=>"101100011",
  28561=>"001001100",
  28562=>"001000011",
  28563=>"100000010",
  28564=>"001111000",
  28565=>"101101110",
  28566=>"011110001",
  28567=>"101111100",
  28568=>"000110101",
  28569=>"101001011",
  28570=>"000001000",
  28571=>"110101011",
  28572=>"001010111",
  28573=>"101001111",
  28574=>"011110011",
  28575=>"101000001",
  28576=>"101001000",
  28577=>"111101111",
  28578=>"001101100",
  28579=>"111101001",
  28580=>"100101101",
  28581=>"111101111",
  28582=>"110100110",
  28583=>"001010010",
  28584=>"010111011",
  28585=>"000011001",
  28586=>"011100100",
  28587=>"111111011",
  28588=>"100000111",
  28589=>"100111011",
  28590=>"001010001",
  28591=>"000101100",
  28592=>"001011010",
  28593=>"000010110",
  28594=>"100100000",
  28595=>"001010111",
  28596=>"001111000",
  28597=>"010111011",
  28598=>"011110111",
  28599=>"110101010",
  28600=>"010001111",
  28601=>"010100101",
  28602=>"111011100",
  28603=>"000000011",
  28604=>"100100001",
  28605=>"001001100",
  28606=>"000001010",
  28607=>"101010110",
  28608=>"011111111",
  28609=>"010101000",
  28610=>"010010110",
  28611=>"111010110",
  28612=>"000011100",
  28613=>"010110101",
  28614=>"011011100",
  28615=>"110111110",
  28616=>"010101011",
  28617=>"111011001",
  28618=>"101001000",
  28619=>"001111110",
  28620=>"100011001",
  28621=>"001101101",
  28622=>"011111101",
  28623=>"110100110",
  28624=>"100000010",
  28625=>"000110110",
  28626=>"000110011",
  28627=>"110101111",
  28628=>"111110111",
  28629=>"100001000",
  28630=>"000101010",
  28631=>"110101010",
  28632=>"001000100",
  28633=>"111101001",
  28634=>"100000010",
  28635=>"101111101",
  28636=>"101010010",
  28637=>"010111101",
  28638=>"111000000",
  28639=>"100001100",
  28640=>"101100001",
  28641=>"101100001",
  28642=>"101110000",
  28643=>"110111100",
  28644=>"100100111",
  28645=>"100010000",
  28646=>"010100001",
  28647=>"111110011",
  28648=>"100111101",
  28649=>"010001110",
  28650=>"110001000",
  28651=>"111010101",
  28652=>"000111100",
  28653=>"111111100",
  28654=>"001100101",
  28655=>"111111011",
  28656=>"011001010",
  28657=>"101011110",
  28658=>"111110010",
  28659=>"111010110",
  28660=>"100011011",
  28661=>"111110001",
  28662=>"111110011",
  28663=>"111101001",
  28664=>"111000111",
  28665=>"100110000",
  28666=>"010000001",
  28667=>"001101000",
  28668=>"100110010",
  28669=>"001110010",
  28670=>"001101111",
  28671=>"000000110",
  28672=>"111000010",
  28673=>"000100101",
  28674=>"000111001",
  28675=>"010010010",
  28676=>"000110011",
  28677=>"111001000",
  28678=>"001100110",
  28679=>"011100111",
  28680=>"110100111",
  28681=>"101101010",
  28682=>"011011001",
  28683=>"001001110",
  28684=>"001011110",
  28685=>"101111111",
  28686=>"010010100",
  28687=>"011001101",
  28688=>"100111110",
  28689=>"110001001",
  28690=>"101111010",
  28691=>"100000100",
  28692=>"111000001",
  28693=>"010100101",
  28694=>"000101111",
  28695=>"011001010",
  28696=>"100101100",
  28697=>"010011100",
  28698=>"000000011",
  28699=>"001001010",
  28700=>"010010101",
  28701=>"110100001",
  28702=>"000100011",
  28703=>"001110011",
  28704=>"010000000",
  28705=>"101000011",
  28706=>"101001000",
  28707=>"001110100",
  28708=>"111000100",
  28709=>"110111011",
  28710=>"000100001",
  28711=>"011010110",
  28712=>"011110101",
  28713=>"111011001",
  28714=>"110011001",
  28715=>"001111100",
  28716=>"011101110",
  28717=>"011010010",
  28718=>"011001100",
  28719=>"100000011",
  28720=>"100110101",
  28721=>"111001100",
  28722=>"101111010",
  28723=>"110111011",
  28724=>"001000000",
  28725=>"111111001",
  28726=>"110000101",
  28727=>"001111011",
  28728=>"110010011",
  28729=>"101011110",
  28730=>"010101010",
  28731=>"000000011",
  28732=>"111001010",
  28733=>"110110010",
  28734=>"100100001",
  28735=>"010000111",
  28736=>"111010111",
  28737=>"110110101",
  28738=>"010100001",
  28739=>"100011000",
  28740=>"011101000",
  28741=>"111001001",
  28742=>"011100111",
  28743=>"010100001",
  28744=>"100010010",
  28745=>"100001000",
  28746=>"111111101",
  28747=>"001001011",
  28748=>"000110101",
  28749=>"100111001",
  28750=>"001100001",
  28751=>"011101011",
  28752=>"111001001",
  28753=>"011110110",
  28754=>"111001111",
  28755=>"010101010",
  28756=>"100000100",
  28757=>"111011011",
  28758=>"011101010",
  28759=>"000010100",
  28760=>"101100011",
  28761=>"111101000",
  28762=>"100000011",
  28763=>"000101010",
  28764=>"111000100",
  28765=>"010100101",
  28766=>"100010010",
  28767=>"100110100",
  28768=>"111000110",
  28769=>"001100011",
  28770=>"011111011",
  28771=>"011011011",
  28772=>"000010000",
  28773=>"000011011",
  28774=>"110101010",
  28775=>"010011110",
  28776=>"111001011",
  28777=>"010110111",
  28778=>"100110110",
  28779=>"001100000",
  28780=>"101000110",
  28781=>"010101010",
  28782=>"001010100",
  28783=>"000001110",
  28784=>"110011101",
  28785=>"111110101",
  28786=>"110010101",
  28787=>"000011100",
  28788=>"101010100",
  28789=>"110110100",
  28790=>"010100110",
  28791=>"101011010",
  28792=>"000100110",
  28793=>"110111000",
  28794=>"001100001",
  28795=>"101110001",
  28796=>"001000110",
  28797=>"001000010",
  28798=>"000000100",
  28799=>"001101011",
  28800=>"111111000",
  28801=>"100110011",
  28802=>"111010111",
  28803=>"101110001",
  28804=>"000011100",
  28805=>"110100110",
  28806=>"110000001",
  28807=>"000000010",
  28808=>"011100011",
  28809=>"111100111",
  28810=>"011110001",
  28811=>"100111000",
  28812=>"010101100",
  28813=>"101001001",
  28814=>"001100010",
  28815=>"011001001",
  28816=>"001100110",
  28817=>"000111001",
  28818=>"111011011",
  28819=>"100101100",
  28820=>"110000001",
  28821=>"010010101",
  28822=>"011010000",
  28823=>"111010111",
  28824=>"000100011",
  28825=>"001000011",
  28826=>"011011100",
  28827=>"010000001",
  28828=>"000111100",
  28829=>"000100110",
  28830=>"010101100",
  28831=>"001010000",
  28832=>"000100000",
  28833=>"010101101",
  28834=>"101010101",
  28835=>"000000011",
  28836=>"110101000",
  28837=>"010000011",
  28838=>"111010100",
  28839=>"101101101",
  28840=>"001111100",
  28841=>"010000110",
  28842=>"010001011",
  28843=>"011011100",
  28844=>"101010100",
  28845=>"100101110",
  28846=>"110001101",
  28847=>"000110000",
  28848=>"010000101",
  28849=>"111001100",
  28850=>"010111101",
  28851=>"001011100",
  28852=>"111010001",
  28853=>"100110000",
  28854=>"001100010",
  28855=>"011001001",
  28856=>"101000100",
  28857=>"110000101",
  28858=>"011010110",
  28859=>"101010111",
  28860=>"101000001",
  28861=>"111111100",
  28862=>"000110011",
  28863=>"000001110",
  28864=>"001111100",
  28865=>"000010111",
  28866=>"111110001",
  28867=>"000000000",
  28868=>"100111100",
  28869=>"010011111",
  28870=>"010100110",
  28871=>"001110000",
  28872=>"001010010",
  28873=>"011011001",
  28874=>"001001101",
  28875=>"101100010",
  28876=>"101001010",
  28877=>"111100001",
  28878=>"010110111",
  28879=>"000011000",
  28880=>"101000011",
  28881=>"001111111",
  28882=>"000100000",
  28883=>"110110110",
  28884=>"100101000",
  28885=>"001111101",
  28886=>"100010011",
  28887=>"101101011",
  28888=>"100100100",
  28889=>"010110011",
  28890=>"001011110",
  28891=>"001011110",
  28892=>"000000000",
  28893=>"010011100",
  28894=>"110100100",
  28895=>"101100001",
  28896=>"000011101",
  28897=>"001100001",
  28898=>"010101011",
  28899=>"110001001",
  28900=>"001100100",
  28901=>"000111000",
  28902=>"111100111",
  28903=>"001000000",
  28904=>"011001001",
  28905=>"001100110",
  28906=>"110100111",
  28907=>"111101011",
  28908=>"010110010",
  28909=>"100000111",
  28910=>"110010000",
  28911=>"100100110",
  28912=>"001001001",
  28913=>"011000010",
  28914=>"000000110",
  28915=>"011001001",
  28916=>"010001100",
  28917=>"000110100",
  28918=>"010100000",
  28919=>"011010011",
  28920=>"110101010",
  28921=>"110110100",
  28922=>"111011000",
  28923=>"010001001",
  28924=>"001111101",
  28925=>"010010000",
  28926=>"000110100",
  28927=>"110110001",
  28928=>"001101110",
  28929=>"100110000",
  28930=>"000101101",
  28931=>"001111110",
  28932=>"110101000",
  28933=>"100011001",
  28934=>"011100110",
  28935=>"110100101",
  28936=>"001000101",
  28937=>"110110110",
  28938=>"110001001",
  28939=>"110000010",
  28940=>"011010010",
  28941=>"000001001",
  28942=>"011101111",
  28943=>"000110001",
  28944=>"100001011",
  28945=>"111110011",
  28946=>"110110010",
  28947=>"000100001",
  28948=>"101111000",
  28949=>"111011001",
  28950=>"111101101",
  28951=>"110100000",
  28952=>"101011000",
  28953=>"101111111",
  28954=>"100110101",
  28955=>"101100010",
  28956=>"010100000",
  28957=>"001010100",
  28958=>"110011110",
  28959=>"011000010",
  28960=>"000010000",
  28961=>"011001111",
  28962=>"111111111",
  28963=>"010001111",
  28964=>"000001111",
  28965=>"000111000",
  28966=>"110100001",
  28967=>"011110001",
  28968=>"100101001",
  28969=>"000100110",
  28970=>"110100000",
  28971=>"100110011",
  28972=>"111100111",
  28973=>"111000000",
  28974=>"101111001",
  28975=>"100100010",
  28976=>"111011011",
  28977=>"101010111",
  28978=>"100010111",
  28979=>"111111000",
  28980=>"111111111",
  28981=>"011001001",
  28982=>"110101010",
  28983=>"101100110",
  28984=>"100011000",
  28985=>"011110001",
  28986=>"010001101",
  28987=>"011110110",
  28988=>"100001101",
  28989=>"001000101",
  28990=>"110100111",
  28991=>"110110110",
  28992=>"101000011",
  28993=>"110100110",
  28994=>"100010011",
  28995=>"101100010",
  28996=>"001010000",
  28997=>"010110110",
  28998=>"101100011",
  28999=>"011001000",
  29000=>"111000111",
  29001=>"101000000",
  29002=>"101111101",
  29003=>"000000110",
  29004=>"101111011",
  29005=>"011110011",
  29006=>"011000111",
  29007=>"000100010",
  29008=>"100111101",
  29009=>"110110010",
  29010=>"001010000",
  29011=>"111111011",
  29012=>"001101011",
  29013=>"000111000",
  29014=>"001101110",
  29015=>"101100111",
  29016=>"010101111",
  29017=>"101010100",
  29018=>"010010011",
  29019=>"000000000",
  29020=>"011001101",
  29021=>"000001011",
  29022=>"100011101",
  29023=>"011110011",
  29024=>"011011010",
  29025=>"100000000",
  29026=>"000001001",
  29027=>"011110110",
  29028=>"010000010",
  29029=>"111111110",
  29030=>"100000000",
  29031=>"001011100",
  29032=>"011110110",
  29033=>"001000111",
  29034=>"011000010",
  29035=>"111111101",
  29036=>"011000100",
  29037=>"101101001",
  29038=>"101000111",
  29039=>"000011011",
  29040=>"011010000",
  29041=>"011010011",
  29042=>"000010011",
  29043=>"001010101",
  29044=>"000110101",
  29045=>"000101010",
  29046=>"101101011",
  29047=>"101111101",
  29048=>"101101000",
  29049=>"101011000",
  29050=>"011000111",
  29051=>"111010100",
  29052=>"100101101",
  29053=>"010111100",
  29054=>"101101100",
  29055=>"111101001",
  29056=>"110000000",
  29057=>"011010000",
  29058=>"111010100",
  29059=>"010010100",
  29060=>"001110011",
  29061=>"010010001",
  29062=>"010100101",
  29063=>"101000011",
  29064=>"010000110",
  29065=>"110101000",
  29066=>"011111101",
  29067=>"101011101",
  29068=>"000010011",
  29069=>"011101000",
  29070=>"111111111",
  29071=>"001010110",
  29072=>"001001101",
  29073=>"001000101",
  29074=>"111000011",
  29075=>"000010001",
  29076=>"111111110",
  29077=>"000100110",
  29078=>"011001010",
  29079=>"111010000",
  29080=>"001000100",
  29081=>"111001101",
  29082=>"110010100",
  29083=>"001011001",
  29084=>"110111111",
  29085=>"010000101",
  29086=>"110111101",
  29087=>"100111111",
  29088=>"101111101",
  29089=>"100111101",
  29090=>"111000001",
  29091=>"011010001",
  29092=>"011010001",
  29093=>"100110010",
  29094=>"111100000",
  29095=>"010011010",
  29096=>"011111001",
  29097=>"010010011",
  29098=>"000101011",
  29099=>"011010110",
  29100=>"011011000",
  29101=>"001110101",
  29102=>"110001111",
  29103=>"101101111",
  29104=>"001011011",
  29105=>"111010111",
  29106=>"000011111",
  29107=>"001110000",
  29108=>"001010100",
  29109=>"110001001",
  29110=>"100111110",
  29111=>"010001000",
  29112=>"011010100",
  29113=>"011111101",
  29114=>"011011101",
  29115=>"101101011",
  29116=>"000101000",
  29117=>"011101110",
  29118=>"000011010",
  29119=>"001111010",
  29120=>"110010010",
  29121=>"001100000",
  29122=>"010010010",
  29123=>"011111100",
  29124=>"100010011",
  29125=>"101111110",
  29126=>"001000000",
  29127=>"100101110",
  29128=>"101011010",
  29129=>"110110000",
  29130=>"101111011",
  29131=>"100111000",
  29132=>"110011011",
  29133=>"110111010",
  29134=>"010010110",
  29135=>"000101011",
  29136=>"010000110",
  29137=>"111111000",
  29138=>"010100000",
  29139=>"101100011",
  29140=>"111100100",
  29141=>"110100110",
  29142=>"011011010",
  29143=>"100110011",
  29144=>"010101111",
  29145=>"000000111",
  29146=>"101011000",
  29147=>"000001011",
  29148=>"111000101",
  29149=>"110101000",
  29150=>"111000101",
  29151=>"000010100",
  29152=>"110000101",
  29153=>"010100110",
  29154=>"100111011",
  29155=>"111001110",
  29156=>"010111000",
  29157=>"101111001",
  29158=>"110111010",
  29159=>"101100010",
  29160=>"111101111",
  29161=>"011111100",
  29162=>"100101101",
  29163=>"000010110",
  29164=>"100100100",
  29165=>"100011010",
  29166=>"110110011",
  29167=>"111111011",
  29168=>"011011011",
  29169=>"011010000",
  29170=>"110111011",
  29171=>"011111000",
  29172=>"011011101",
  29173=>"001110100",
  29174=>"111000010",
  29175=>"100111101",
  29176=>"100000010",
  29177=>"011101011",
  29178=>"011010111",
  29179=>"110100110",
  29180=>"010001010",
  29181=>"101101011",
  29182=>"100101011",
  29183=>"111011000",
  29184=>"101000011",
  29185=>"000111101",
  29186=>"110001101",
  29187=>"111100110",
  29188=>"000111100",
  29189=>"111010111",
  29190=>"000101100",
  29191=>"101101110",
  29192=>"011100000",
  29193=>"001001000",
  29194=>"100011111",
  29195=>"001101000",
  29196=>"011011110",
  29197=>"100010010",
  29198=>"010100111",
  29199=>"000101011",
  29200=>"111111011",
  29201=>"101100100",
  29202=>"010000011",
  29203=>"011010000",
  29204=>"110100011",
  29205=>"111001111",
  29206=>"101100010",
  29207=>"010010110",
  29208=>"000111100",
  29209=>"011111100",
  29210=>"001011000",
  29211=>"110110110",
  29212=>"100000101",
  29213=>"111111011",
  29214=>"001101111",
  29215=>"110100011",
  29216=>"000010101",
  29217=>"111100110",
  29218=>"001001000",
  29219=>"101010010",
  29220=>"011000110",
  29221=>"100100101",
  29222=>"111110101",
  29223=>"000010110",
  29224=>"000101100",
  29225=>"100010010",
  29226=>"010011000",
  29227=>"111100010",
  29228=>"101100010",
  29229=>"101000111",
  29230=>"010011110",
  29231=>"111010111",
  29232=>"100100001",
  29233=>"110110111",
  29234=>"110111110",
  29235=>"100000000",
  29236=>"110001101",
  29237=>"100011010",
  29238=>"001100100",
  29239=>"000101111",
  29240=>"101011101",
  29241=>"101101000",
  29242=>"100101011",
  29243=>"110010000",
  29244=>"010011100",
  29245=>"100110110",
  29246=>"010011100",
  29247=>"101001000",
  29248=>"111111110",
  29249=>"010110111",
  29250=>"001101111",
  29251=>"011100010",
  29252=>"111111101",
  29253=>"011000001",
  29254=>"010000010",
  29255=>"010011000",
  29256=>"110100110",
  29257=>"110111001",
  29258=>"010100011",
  29259=>"011010111",
  29260=>"101100100",
  29261=>"001000101",
  29262=>"010110111",
  29263=>"010101101",
  29264=>"111110001",
  29265=>"101100101",
  29266=>"111000101",
  29267=>"111001001",
  29268=>"001101111",
  29269=>"100100110",
  29270=>"000001010",
  29271=>"010001001",
  29272=>"010010010",
  29273=>"011010011",
  29274=>"000100110",
  29275=>"010000001",
  29276=>"000100001",
  29277=>"101011110",
  29278=>"111001011",
  29279=>"111111010",
  29280=>"010011110",
  29281=>"110101101",
  29282=>"010001010",
  29283=>"010001101",
  29284=>"111111110",
  29285=>"000010000",
  29286=>"100100110",
  29287=>"100010111",
  29288=>"110001100",
  29289=>"100001100",
  29290=>"111010000",
  29291=>"000100000",
  29292=>"110010110",
  29293=>"100000100",
  29294=>"000011111",
  29295=>"101001001",
  29296=>"000001101",
  29297=>"100101001",
  29298=>"101101101",
  29299=>"110111111",
  29300=>"111111110",
  29301=>"111110000",
  29302=>"001110001",
  29303=>"101111011",
  29304=>"000000011",
  29305=>"010010110",
  29306=>"000100100",
  29307=>"010111001",
  29308=>"000000110",
  29309=>"110000000",
  29310=>"111110010",
  29311=>"111001100",
  29312=>"010010010",
  29313=>"100011011",
  29314=>"110100010",
  29315=>"010011110",
  29316=>"000000000",
  29317=>"101010110",
  29318=>"100010001",
  29319=>"001100000",
  29320=>"010101111",
  29321=>"000101010",
  29322=>"011001101",
  29323=>"100111000",
  29324=>"100001100",
  29325=>"111111110",
  29326=>"010111011",
  29327=>"000101110",
  29328=>"000101111",
  29329=>"111011110",
  29330=>"000000110",
  29331=>"001010110",
  29332=>"100100001",
  29333=>"111001000",
  29334=>"010101001",
  29335=>"100011000",
  29336=>"011011011",
  29337=>"100110110",
  29338=>"000001001",
  29339=>"010111000",
  29340=>"011101100",
  29341=>"011000110",
  29342=>"010110000",
  29343=>"110111111",
  29344=>"001101111",
  29345=>"100010111",
  29346=>"001111000",
  29347=>"110001000",
  29348=>"111111101",
  29349=>"000011000",
  29350=>"111001111",
  29351=>"011011111",
  29352=>"110001011",
  29353=>"010110010",
  29354=>"001000001",
  29355=>"001100101",
  29356=>"100000001",
  29357=>"111000011",
  29358=>"110100001",
  29359=>"100110111",
  29360=>"000000101",
  29361=>"010101100",
  29362=>"001001001",
  29363=>"100010010",
  29364=>"101011100",
  29365=>"000100011",
  29366=>"001110011",
  29367=>"000111100",
  29368=>"000001100",
  29369=>"111100111",
  29370=>"111000110",
  29371=>"000010001",
  29372=>"100000000",
  29373=>"111011001",
  29374=>"111010110",
  29375=>"000001101",
  29376=>"000011010",
  29377=>"100100011",
  29378=>"110110010",
  29379=>"000001010",
  29380=>"110011110",
  29381=>"011010110",
  29382=>"110100001",
  29383=>"000000101",
  29384=>"010100110",
  29385=>"011011110",
  29386=>"100001111",
  29387=>"111101111",
  29388=>"100100111",
  29389=>"001000011",
  29390=>"011100100",
  29391=>"010010111",
  29392=>"100111111",
  29393=>"100101000",
  29394=>"100110011",
  29395=>"000000000",
  29396=>"101000100",
  29397=>"100000100",
  29398=>"101010110",
  29399=>"001010001",
  29400=>"000000111",
  29401=>"001001111",
  29402=>"110110000",
  29403=>"100010000",
  29404=>"011110100",
  29405=>"000100010",
  29406=>"111011101",
  29407=>"010010010",
  29408=>"000010000",
  29409=>"110111001",
  29410=>"010011001",
  29411=>"111101100",
  29412=>"100110010",
  29413=>"000111111",
  29414=>"000001101",
  29415=>"001101001",
  29416=>"101101101",
  29417=>"110110101",
  29418=>"001110011",
  29419=>"011001110",
  29420=>"011001010",
  29421=>"000111000",
  29422=>"111000101",
  29423=>"000000100",
  29424=>"100111010",
  29425=>"101000011",
  29426=>"100000000",
  29427=>"111000111",
  29428=>"101101010",
  29429=>"111000010",
  29430=>"101010111",
  29431=>"000111001",
  29432=>"011011110",
  29433=>"111010011",
  29434=>"010111110",
  29435=>"100111010",
  29436=>"110101111",
  29437=>"111000111",
  29438=>"010000111",
  29439=>"000111100",
  29440=>"101010000",
  29441=>"010110010",
  29442=>"111000100",
  29443=>"101110001",
  29444=>"110111110",
  29445=>"100011101",
  29446=>"010100111",
  29447=>"000001011",
  29448=>"011011000",
  29449=>"111100110",
  29450=>"100111100",
  29451=>"110011100",
  29452=>"011101101",
  29453=>"101110101",
  29454=>"110101101",
  29455=>"100011110",
  29456=>"100101010",
  29457=>"111000010",
  29458=>"011100000",
  29459=>"001110001",
  29460=>"110100100",
  29461=>"010111001",
  29462=>"100000100",
  29463=>"000111010",
  29464=>"011010101",
  29465=>"110111110",
  29466=>"000001011",
  29467=>"001000111",
  29468=>"110111010",
  29469=>"101111010",
  29470=>"011100000",
  29471=>"110111101",
  29472=>"100100001",
  29473=>"000010011",
  29474=>"001100001",
  29475=>"010101011",
  29476=>"011011100",
  29477=>"101111111",
  29478=>"110101011",
  29479=>"101000001",
  29480=>"101000001",
  29481=>"000100100",
  29482=>"100010001",
  29483=>"010110010",
  29484=>"010010110",
  29485=>"011000011",
  29486=>"010111010",
  29487=>"001111001",
  29488=>"101110111",
  29489=>"100100100",
  29490=>"001010011",
  29491=>"000110011",
  29492=>"000011011",
  29493=>"100100110",
  29494=>"100100111",
  29495=>"000100010",
  29496=>"111111100",
  29497=>"111111101",
  29498=>"011011110",
  29499=>"001101011",
  29500=>"110111100",
  29501=>"000100010",
  29502=>"011001010",
  29503=>"001011010",
  29504=>"001111111",
  29505=>"111001100",
  29506=>"111100111",
  29507=>"111011101",
  29508=>"110110111",
  29509=>"011111001",
  29510=>"101001101",
  29511=>"000110000",
  29512=>"111101110",
  29513=>"001000010",
  29514=>"011111000",
  29515=>"000010010",
  29516=>"101001110",
  29517=>"010010100",
  29518=>"001010101",
  29519=>"011000010",
  29520=>"010011101",
  29521=>"111000011",
  29522=>"011100001",
  29523=>"111010000",
  29524=>"100010000",
  29525=>"000100101",
  29526=>"010010110",
  29527=>"010011101",
  29528=>"000111001",
  29529=>"001001100",
  29530=>"111011111",
  29531=>"000110001",
  29532=>"000110100",
  29533=>"111110010",
  29534=>"110000011",
  29535=>"100101111",
  29536=>"101010110",
  29537=>"000011011",
  29538=>"001010101",
  29539=>"101000110",
  29540=>"001101111",
  29541=>"010000100",
  29542=>"100010011",
  29543=>"011100111",
  29544=>"101001011",
  29545=>"100101011",
  29546=>"111000001",
  29547=>"110101100",
  29548=>"010001101",
  29549=>"110000100",
  29550=>"011110011",
  29551=>"101011000",
  29552=>"111110111",
  29553=>"111000101",
  29554=>"001101111",
  29555=>"011111100",
  29556=>"010111010",
  29557=>"000011111",
  29558=>"101111110",
  29559=>"000110000",
  29560=>"010001011",
  29561=>"010010100",
  29562=>"011110101",
  29563=>"000001000",
  29564=>"011110011",
  29565=>"110110100",
  29566=>"001110000",
  29567=>"011111011",
  29568=>"010111101",
  29569=>"101000001",
  29570=>"001001010",
  29571=>"110000111",
  29572=>"000000111",
  29573=>"011000011",
  29574=>"011110011",
  29575=>"001110011",
  29576=>"110010010",
  29577=>"010000010",
  29578=>"110111111",
  29579=>"010001101",
  29580=>"101111100",
  29581=>"001010001",
  29582=>"110000000",
  29583=>"011110111",
  29584=>"101100011",
  29585=>"001110111",
  29586=>"001101110",
  29587=>"111111001",
  29588=>"111011010",
  29589=>"010000000",
  29590=>"010001001",
  29591=>"110001101",
  29592=>"000000100",
  29593=>"111111000",
  29594=>"010101001",
  29595=>"000110001",
  29596=>"101010100",
  29597=>"001110110",
  29598=>"010010010",
  29599=>"001110000",
  29600=>"111100011",
  29601=>"111000010",
  29602=>"111011111",
  29603=>"001011100",
  29604=>"001101001",
  29605=>"000100100",
  29606=>"000010010",
  29607=>"110011110",
  29608=>"101111000",
  29609=>"010010110",
  29610=>"000001101",
  29611=>"101111001",
  29612=>"001001111",
  29613=>"011011101",
  29614=>"011000101",
  29615=>"101000001",
  29616=>"110011101",
  29617=>"001011011",
  29618=>"001100100",
  29619=>"001101010",
  29620=>"011100001",
  29621=>"011111111",
  29622=>"010010100",
  29623=>"001101001",
  29624=>"001010010",
  29625=>"011010001",
  29626=>"111100111",
  29627=>"101010011",
  29628=>"101100011",
  29629=>"001011010",
  29630=>"000100100",
  29631=>"101100001",
  29632=>"000001000",
  29633=>"000011111",
  29634=>"110100111",
  29635=>"100011101",
  29636=>"110010000",
  29637=>"110111111",
  29638=>"101100011",
  29639=>"100101101",
  29640=>"001001000",
  29641=>"011110111",
  29642=>"100101000",
  29643=>"110111100",
  29644=>"010011011",
  29645=>"110011101",
  29646=>"100101011",
  29647=>"111010100",
  29648=>"011111100",
  29649=>"010001110",
  29650=>"001110001",
  29651=>"110111111",
  29652=>"001010100",
  29653=>"111100101",
  29654=>"110101110",
  29655=>"100101111",
  29656=>"011001001",
  29657=>"010010000",
  29658=>"100001011",
  29659=>"101000001",
  29660=>"011110010",
  29661=>"010111010",
  29662=>"011010010",
  29663=>"011010010",
  29664=>"101111010",
  29665=>"010001010",
  29666=>"100100101",
  29667=>"011001000",
  29668=>"100000000",
  29669=>"000011011",
  29670=>"110101010",
  29671=>"010101000",
  29672=>"010111001",
  29673=>"111101101",
  29674=>"100111010",
  29675=>"011101001",
  29676=>"010100101",
  29677=>"001010011",
  29678=>"101000001",
  29679=>"001101001",
  29680=>"000100000",
  29681=>"100100011",
  29682=>"101001000",
  29683=>"001111100",
  29684=>"011011101",
  29685=>"100010001",
  29686=>"010011110",
  29687=>"110000101",
  29688=>"111110101",
  29689=>"111100110",
  29690=>"000001111",
  29691=>"000010101",
  29692=>"010000011",
  29693=>"101100111",
  29694=>"010011001",
  29695=>"011001001",
  29696=>"111111000",
  29697=>"000110010",
  29698=>"010110000",
  29699=>"100111111",
  29700=>"100010010",
  29701=>"111111111",
  29702=>"111111010",
  29703=>"101010101",
  29704=>"000100110",
  29705=>"001101001",
  29706=>"111111111",
  29707=>"111110000",
  29708=>"101101010",
  29709=>"100001110",
  29710=>"101101100",
  29711=>"111011101",
  29712=>"011001110",
  29713=>"011000010",
  29714=>"100101011",
  29715=>"101110001",
  29716=>"100101000",
  29717=>"000100001",
  29718=>"100001000",
  29719=>"111101110",
  29720=>"110001011",
  29721=>"110011001",
  29722=>"010101111",
  29723=>"011100100",
  29724=>"110001101",
  29725=>"011010001",
  29726=>"111100100",
  29727=>"011010000",
  29728=>"011001000",
  29729=>"101001111",
  29730=>"110011001",
  29731=>"111100000",
  29732=>"100011101",
  29733=>"101001111",
  29734=>"101010000",
  29735=>"111101001",
  29736=>"100111001",
  29737=>"111001000",
  29738=>"001110000",
  29739=>"011001001",
  29740=>"011011110",
  29741=>"010010111",
  29742=>"010101010",
  29743=>"100100110",
  29744=>"100100101",
  29745=>"101101010",
  29746=>"001000110",
  29747=>"111111110",
  29748=>"101001010",
  29749=>"100101101",
  29750=>"111011111",
  29751=>"100101000",
  29752=>"100100000",
  29753=>"111010111",
  29754=>"111111000",
  29755=>"110011010",
  29756=>"010110001",
  29757=>"011111010",
  29758=>"010011111",
  29759=>"111100000",
  29760=>"010010010",
  29761=>"111110000",
  29762=>"001011111",
  29763=>"000011010",
  29764=>"000000001",
  29765=>"000100000",
  29766=>"000010011",
  29767=>"101111011",
  29768=>"101010001",
  29769=>"110101100",
  29770=>"011101000",
  29771=>"010100110",
  29772=>"100000101",
  29773=>"101001110",
  29774=>"101001000",
  29775=>"110100001",
  29776=>"011111111",
  29777=>"111100111",
  29778=>"010101101",
  29779=>"000101001",
  29780=>"010101100",
  29781=>"100111010",
  29782=>"010010011",
  29783=>"111101001",
  29784=>"000001001",
  29785=>"011011011",
  29786=>"111000110",
  29787=>"000001011",
  29788=>"111010101",
  29789=>"000000100",
  29790=>"010100100",
  29791=>"010000011",
  29792=>"001000110",
  29793=>"110101101",
  29794=>"010011101",
  29795=>"101110001",
  29796=>"110001001",
  29797=>"000000110",
  29798=>"000011011",
  29799=>"001000001",
  29800=>"110001111",
  29801=>"100000010",
  29802=>"111111001",
  29803=>"100001111",
  29804=>"100000100",
  29805=>"011000011",
  29806=>"010100110",
  29807=>"111000010",
  29808=>"101110111",
  29809=>"101000001",
  29810=>"100011000",
  29811=>"010111011",
  29812=>"001111101",
  29813=>"111100111",
  29814=>"111111000",
  29815=>"101001100",
  29816=>"111010001",
  29817=>"010001000",
  29818=>"011110011",
  29819=>"111101111",
  29820=>"100000101",
  29821=>"110011000",
  29822=>"000001010",
  29823=>"111011010",
  29824=>"111111000",
  29825=>"000111111",
  29826=>"111011111",
  29827=>"101001100",
  29828=>"111111111",
  29829=>"010001110",
  29830=>"001000100",
  29831=>"000100110",
  29832=>"001100110",
  29833=>"001110011",
  29834=>"101110110",
  29835=>"010000011",
  29836=>"110111100",
  29837=>"011100101",
  29838=>"001100101",
  29839=>"110011111",
  29840=>"111011110",
  29841=>"011111000",
  29842=>"110011111",
  29843=>"011110110",
  29844=>"000101101",
  29845=>"000010101",
  29846=>"111010111",
  29847=>"001000000",
  29848=>"111010000",
  29849=>"100111001",
  29850=>"000100100",
  29851=>"010101011",
  29852=>"111101110",
  29853=>"111011010",
  29854=>"011011001",
  29855=>"100001111",
  29856=>"001000111",
  29857=>"111010111",
  29858=>"110011111",
  29859=>"000010010",
  29860=>"010011110",
  29861=>"000010010",
  29862=>"001100011",
  29863=>"111100100",
  29864=>"111010011",
  29865=>"101000101",
  29866=>"110100110",
  29867=>"110111110",
  29868=>"100100001",
  29869=>"101010010",
  29870=>"001100100",
  29871=>"111110000",
  29872=>"110000110",
  29873=>"111100110",
  29874=>"111101100",
  29875=>"100110100",
  29876=>"010111111",
  29877=>"111000110",
  29878=>"001011101",
  29879=>"101011000",
  29880=>"111100000",
  29881=>"110000100",
  29882=>"111001000",
  29883=>"000010100",
  29884=>"011111111",
  29885=>"011001000",
  29886=>"011000001",
  29887=>"000011100",
  29888=>"010001011",
  29889=>"110110000",
  29890=>"101000111",
  29891=>"010001100",
  29892=>"101101010",
  29893=>"001011000",
  29894=>"111110100",
  29895=>"111101101",
  29896=>"001000010",
  29897=>"100100111",
  29898=>"110101111",
  29899=>"100011000",
  29900=>"001000100",
  29901=>"110111111",
  29902=>"111100101",
  29903=>"000011001",
  29904=>"111001110",
  29905=>"000011100",
  29906=>"011000010",
  29907=>"100100001",
  29908=>"111101101",
  29909=>"100000100",
  29910=>"010100100",
  29911=>"001011011",
  29912=>"011100111",
  29913=>"100011010",
  29914=>"100110000",
  29915=>"100011100",
  29916=>"110011010",
  29917=>"111100100",
  29918=>"010101111",
  29919=>"011111101",
  29920=>"111101001",
  29921=>"101100111",
  29922=>"110111111",
  29923=>"111110110",
  29924=>"000110111",
  29925=>"001010110",
  29926=>"001110100",
  29927=>"010010110",
  29928=>"011011101",
  29929=>"010101100",
  29930=>"011000110",
  29931=>"101000100",
  29932=>"100110110",
  29933=>"100001100",
  29934=>"101111001",
  29935=>"110110010",
  29936=>"000001101",
  29937=>"101111011",
  29938=>"001111011",
  29939=>"000111001",
  29940=>"100110101",
  29941=>"000001000",
  29942=>"110001001",
  29943=>"111001001",
  29944=>"111001010",
  29945=>"011111100",
  29946=>"100111100",
  29947=>"110001001",
  29948=>"000100010",
  29949=>"010001001",
  29950=>"111111110",
  29951=>"000000111",
  29952=>"101100000",
  29953=>"111001011",
  29954=>"101111011",
  29955=>"101001010",
  29956=>"101010111",
  29957=>"100010010",
  29958=>"101011100",
  29959=>"010000010",
  29960=>"110000000",
  29961=>"110000000",
  29962=>"110010001",
  29963=>"111101111",
  29964=>"101010000",
  29965=>"100101101",
  29966=>"011110011",
  29967=>"111000100",
  29968=>"010011111",
  29969=>"000011000",
  29970=>"100111001",
  29971=>"000000111",
  29972=>"111100101",
  29973=>"111111110",
  29974=>"101111001",
  29975=>"100011010",
  29976=>"101100101",
  29977=>"101011110",
  29978=>"000101111",
  29979=>"100110111",
  29980=>"100000000",
  29981=>"010111011",
  29982=>"100110110",
  29983=>"100100011",
  29984=>"101111010",
  29985=>"101000111",
  29986=>"001111010",
  29987=>"100000001",
  29988=>"111001001",
  29989=>"001111010",
  29990=>"010010111",
  29991=>"111010010",
  29992=>"011101001",
  29993=>"010110111",
  29994=>"000111000",
  29995=>"110110000",
  29996=>"010111000",
  29997=>"001101010",
  29998=>"111110111",
  29999=>"001100010",
  30000=>"011101010",
  30001=>"110110110",
  30002=>"001000010",
  30003=>"100000000",
  30004=>"000010011",
  30005=>"101111111",
  30006=>"101110101",
  30007=>"111001111",
  30008=>"111011110",
  30009=>"111111101",
  30010=>"111011100",
  30011=>"010001000",
  30012=>"100001010",
  30013=>"100000110",
  30014=>"100001011",
  30015=>"111111001",
  30016=>"101010101",
  30017=>"101100101",
  30018=>"111100100",
  30019=>"110110011",
  30020=>"001101101",
  30021=>"000110000",
  30022=>"001111111",
  30023=>"111100010",
  30024=>"011011000",
  30025=>"011111101",
  30026=>"010011101",
  30027=>"111111010",
  30028=>"111001111",
  30029=>"011010010",
  30030=>"100111001",
  30031=>"101011011",
  30032=>"111011100",
  30033=>"000001110",
  30034=>"100010000",
  30035=>"100111000",
  30036=>"000101110",
  30037=>"111000111",
  30038=>"011110100",
  30039=>"010100001",
  30040=>"001001000",
  30041=>"000001111",
  30042=>"001011101",
  30043=>"010011110",
  30044=>"110010011",
  30045=>"011101001",
  30046=>"111110110",
  30047=>"110111111",
  30048=>"101100011",
  30049=>"011101111",
  30050=>"111011100",
  30051=>"111000100",
  30052=>"110110110",
  30053=>"110111111",
  30054=>"010010010",
  30055=>"111111111",
  30056=>"000111111",
  30057=>"111001000",
  30058=>"111101010",
  30059=>"110010101",
  30060=>"111101111",
  30061=>"111111000",
  30062=>"110000000",
  30063=>"111000000",
  30064=>"110010000",
  30065=>"101100010",
  30066=>"001010011",
  30067=>"011111111",
  30068=>"111010000",
  30069=>"000100010",
  30070=>"111001010",
  30071=>"010110001",
  30072=>"001100010",
  30073=>"000110000",
  30074=>"000001010",
  30075=>"001011010",
  30076=>"010100000",
  30077=>"000100110",
  30078=>"100000101",
  30079=>"100111000",
  30080=>"101111100",
  30081=>"011011110",
  30082=>"100000111",
  30083=>"100101111",
  30084=>"001101011",
  30085=>"000001111",
  30086=>"111100100",
  30087=>"111001010",
  30088=>"000100010",
  30089=>"100101010",
  30090=>"111111011",
  30091=>"001101000",
  30092=>"101111111",
  30093=>"111000100",
  30094=>"011111000",
  30095=>"110110110",
  30096=>"001101000",
  30097=>"111110000",
  30098=>"110100010",
  30099=>"000111011",
  30100=>"001101100",
  30101=>"101101000",
  30102=>"101010110",
  30103=>"000000011",
  30104=>"011010011",
  30105=>"110100101",
  30106=>"010000011",
  30107=>"101001111",
  30108=>"010111001",
  30109=>"101101110",
  30110=>"100110011",
  30111=>"110011010",
  30112=>"111100110",
  30113=>"110110111",
  30114=>"101110110",
  30115=>"110001100",
  30116=>"010101110",
  30117=>"110111000",
  30118=>"110111111",
  30119=>"001101011",
  30120=>"100000000",
  30121=>"101110111",
  30122=>"101000000",
  30123=>"101011001",
  30124=>"000000010",
  30125=>"111100100",
  30126=>"111011001",
  30127=>"001110010",
  30128=>"010100100",
  30129=>"010001111",
  30130=>"101000100",
  30131=>"101011111",
  30132=>"110111010",
  30133=>"101101011",
  30134=>"000000001",
  30135=>"001100101",
  30136=>"100101011",
  30137=>"001001011",
  30138=>"111001001",
  30139=>"000011010",
  30140=>"001100111",
  30141=>"011111001",
  30142=>"100100111",
  30143=>"110000000",
  30144=>"111011110",
  30145=>"010010101",
  30146=>"010000110",
  30147=>"010111000",
  30148=>"110111100",
  30149=>"000011110",
  30150=>"110000010",
  30151=>"111110100",
  30152=>"100100110",
  30153=>"100101000",
  30154=>"111100001",
  30155=>"100110101",
  30156=>"001011010",
  30157=>"011001101",
  30158=>"010110100",
  30159=>"011101111",
  30160=>"111100000",
  30161=>"100000001",
  30162=>"001101000",
  30163=>"000000110",
  30164=>"110010101",
  30165=>"011001000",
  30166=>"000001110",
  30167=>"111011111",
  30168=>"011001011",
  30169=>"010011111",
  30170=>"000101101",
  30171=>"101011011",
  30172=>"110010000",
  30173=>"101010101",
  30174=>"100011101",
  30175=>"001010100",
  30176=>"011011100",
  30177=>"010110110",
  30178=>"010101000",
  30179=>"101000100",
  30180=>"110000011",
  30181=>"101110000",
  30182=>"111111111",
  30183=>"111111011",
  30184=>"111111001",
  30185=>"000111011",
  30186=>"011110101",
  30187=>"110110111",
  30188=>"111000001",
  30189=>"000001101",
  30190=>"011101011",
  30191=>"111101111",
  30192=>"101010111",
  30193=>"001001100",
  30194=>"111110011",
  30195=>"110001010",
  30196=>"101010011",
  30197=>"111111101",
  30198=>"100001111",
  30199=>"000011011",
  30200=>"011111000",
  30201=>"010110001",
  30202=>"111100000",
  30203=>"100110011",
  30204=>"101000101",
  30205=>"000101011",
  30206=>"000111011",
  30207=>"010010001",
  30208=>"011110111",
  30209=>"010000100",
  30210=>"110010111",
  30211=>"100111100",
  30212=>"010100011",
  30213=>"110100100",
  30214=>"111111010",
  30215=>"101011100",
  30216=>"100011010",
  30217=>"100000100",
  30218=>"100001000",
  30219=>"110010010",
  30220=>"001000101",
  30221=>"001100101",
  30222=>"110110111",
  30223=>"001010000",
  30224=>"001101101",
  30225=>"010100111",
  30226=>"111110100",
  30227=>"000111011",
  30228=>"000001011",
  30229=>"110011011",
  30230=>"000110100",
  30231=>"001011010",
  30232=>"000111001",
  30233=>"000011001",
  30234=>"101000010",
  30235=>"001010111",
  30236=>"111100101",
  30237=>"111111101",
  30238=>"011011111",
  30239=>"101111101",
  30240=>"101101110",
  30241=>"101001111",
  30242=>"111101000",
  30243=>"011111101",
  30244=>"000111111",
  30245=>"110001111",
  30246=>"001001100",
  30247=>"101110001",
  30248=>"101110111",
  30249=>"010000011",
  30250=>"101011000",
  30251=>"010000000",
  30252=>"110101000",
  30253=>"001101011",
  30254=>"100000001",
  30255=>"101111111",
  30256=>"100011100",
  30257=>"110110011",
  30258=>"011010101",
  30259=>"100111111",
  30260=>"110100000",
  30261=>"111000001",
  30262=>"000010101",
  30263=>"001010110",
  30264=>"110100010",
  30265=>"110101110",
  30266=>"000111011",
  30267=>"101000110",
  30268=>"011101011",
  30269=>"101110010",
  30270=>"001001100",
  30271=>"011101011",
  30272=>"110100000",
  30273=>"111100110",
  30274=>"100111001",
  30275=>"101001100",
  30276=>"001001101",
  30277=>"100110101",
  30278=>"110000011",
  30279=>"011110001",
  30280=>"010100101",
  30281=>"010011001",
  30282=>"010001010",
  30283=>"101001100",
  30284=>"100100101",
  30285=>"101110100",
  30286=>"000111000",
  30287=>"010010000",
  30288=>"001001101",
  30289=>"111110010",
  30290=>"001011010",
  30291=>"011100000",
  30292=>"001111111",
  30293=>"000000101",
  30294=>"111101111",
  30295=>"100001000",
  30296=>"111010100",
  30297=>"000010110",
  30298=>"100010110",
  30299=>"011111110",
  30300=>"111111111",
  30301=>"111110001",
  30302=>"001101010",
  30303=>"100000100",
  30304=>"111101110",
  30305=>"011100100",
  30306=>"110111110",
  30307=>"010011011",
  30308=>"101001100",
  30309=>"100110111",
  30310=>"111101001",
  30311=>"110110001",
  30312=>"010000111",
  30313=>"111101000",
  30314=>"101000000",
  30315=>"111101000",
  30316=>"101010001",
  30317=>"010111000",
  30318=>"110110100",
  30319=>"011011001",
  30320=>"110000011",
  30321=>"110111011",
  30322=>"011101111",
  30323=>"111000100",
  30324=>"101101101",
  30325=>"110010110",
  30326=>"110101000",
  30327=>"101001010",
  30328=>"110110110",
  30329=>"101010011",
  30330=>"010011011",
  30331=>"010011000",
  30332=>"111111111",
  30333=>"001100001",
  30334=>"110111000",
  30335=>"110000001",
  30336=>"011111100",
  30337=>"100010010",
  30338=>"000101101",
  30339=>"011110111",
  30340=>"100000010",
  30341=>"101101110",
  30342=>"100000001",
  30343=>"101110000",
  30344=>"101011110",
  30345=>"110100100",
  30346=>"111000000",
  30347=>"001100100",
  30348=>"100111111",
  30349=>"101001011",
  30350=>"010001011",
  30351=>"111000010",
  30352=>"101001011",
  30353=>"110010001",
  30354=>"111000100",
  30355=>"010001101",
  30356=>"101111011",
  30357=>"011000001",
  30358=>"010110100",
  30359=>"101011001",
  30360=>"100000001",
  30361=>"111101000",
  30362=>"101010010",
  30363=>"111110110",
  30364=>"111011101",
  30365=>"001001110",
  30366=>"110111011",
  30367=>"001111010",
  30368=>"111100011",
  30369=>"001111101",
  30370=>"110000111",
  30371=>"001101111",
  30372=>"000111111",
  30373=>"101001101",
  30374=>"111101101",
  30375=>"011110111",
  30376=>"101001011",
  30377=>"110111100",
  30378=>"111110010",
  30379=>"111101001",
  30380=>"011010111",
  30381=>"111110100",
  30382=>"011001001",
  30383=>"101111001",
  30384=>"111111100",
  30385=>"011010010",
  30386=>"111010010",
  30387=>"100111001",
  30388=>"000101010",
  30389=>"100010000",
  30390=>"101110011",
  30391=>"000110001",
  30392=>"011110101",
  30393=>"001010010",
  30394=>"001011001",
  30395=>"111111100",
  30396=>"111001001",
  30397=>"011011110",
  30398=>"111000111",
  30399=>"000111000",
  30400=>"100101011",
  30401=>"011011010",
  30402=>"000010110",
  30403=>"010111101",
  30404=>"101010000",
  30405=>"111110111",
  30406=>"110001011",
  30407=>"111000010",
  30408=>"011111111",
  30409=>"100101000",
  30410=>"111110001",
  30411=>"111110101",
  30412=>"000000011",
  30413=>"010011011",
  30414=>"010000100",
  30415=>"100010111",
  30416=>"001101010",
  30417=>"011101011",
  30418=>"001000111",
  30419=>"111001001",
  30420=>"101000100",
  30421=>"100000011",
  30422=>"001001100",
  30423=>"101011111",
  30424=>"011101110",
  30425=>"001110011",
  30426=>"011111101",
  30427=>"010000111",
  30428=>"111001000",
  30429=>"011010110",
  30430=>"100000100",
  30431=>"011000110",
  30432=>"011000000",
  30433=>"111001011",
  30434=>"000010001",
  30435=>"010000111",
  30436=>"000011010",
  30437=>"011100010",
  30438=>"000101010",
  30439=>"100001110",
  30440=>"100101000",
  30441=>"101111100",
  30442=>"110001110",
  30443=>"001001100",
  30444=>"110000000",
  30445=>"010111100",
  30446=>"110111110",
  30447=>"111110100",
  30448=>"001010101",
  30449=>"000110000",
  30450=>"111001000",
  30451=>"111100100",
  30452=>"000110001",
  30453=>"000000111",
  30454=>"111101101",
  30455=>"110110111",
  30456=>"110101110",
  30457=>"011100011",
  30458=>"100100111",
  30459=>"111111111",
  30460=>"100101010",
  30461=>"100100001",
  30462=>"011011100",
  30463=>"011010010",
  30464=>"110011001",
  30465=>"110000101",
  30466=>"000001000",
  30467=>"011111010",
  30468=>"110001100",
  30469=>"101101100",
  30470=>"101000000",
  30471=>"101100011",
  30472=>"000000001",
  30473=>"111010101",
  30474=>"010000000",
  30475=>"111110100",
  30476=>"101110100",
  30477=>"100011010",
  30478=>"101000010",
  30479=>"000000010",
  30480=>"101111000",
  30481=>"111011011",
  30482=>"010111001",
  30483=>"011100000",
  30484=>"000001000",
  30485=>"101010100",
  30486=>"011101010",
  30487=>"010000000",
  30488=>"111100111",
  30489=>"111111001",
  30490=>"001111110",
  30491=>"000000001",
  30492=>"010001100",
  30493=>"101111100",
  30494=>"111111100",
  30495=>"000010111",
  30496=>"101101110",
  30497=>"011100000",
  30498=>"000011101",
  30499=>"110000010",
  30500=>"000110000",
  30501=>"111100000",
  30502=>"100001111",
  30503=>"101010110",
  30504=>"101011001",
  30505=>"111111100",
  30506=>"110111100",
  30507=>"011011011",
  30508=>"100111001",
  30509=>"001101100",
  30510=>"011010000",
  30511=>"100100111",
  30512=>"111100001",
  30513=>"101101010",
  30514=>"111011111",
  30515=>"101100101",
  30516=>"111010100",
  30517=>"010101111",
  30518=>"111110110",
  30519=>"111000000",
  30520=>"101010011",
  30521=>"000100111",
  30522=>"001111001",
  30523=>"110110111",
  30524=>"011101011",
  30525=>"111101001",
  30526=>"111100111",
  30527=>"001000100",
  30528=>"111100000",
  30529=>"000001100",
  30530=>"001000111",
  30531=>"110101010",
  30532=>"000111001",
  30533=>"001001100",
  30534=>"001100100",
  30535=>"100111001",
  30536=>"111011010",
  30537=>"011010011",
  30538=>"000101000",
  30539=>"101110001",
  30540=>"000011001",
  30541=>"100011111",
  30542=>"101000111",
  30543=>"101100111",
  30544=>"111010000",
  30545=>"100110110",
  30546=>"110110000",
  30547=>"111000000",
  30548=>"111110110",
  30549=>"001101100",
  30550=>"011111011",
  30551=>"100010011",
  30552=>"000011000",
  30553=>"100000100",
  30554=>"100000100",
  30555=>"111110101",
  30556=>"100110011",
  30557=>"001110000",
  30558=>"101110100",
  30559=>"111010011",
  30560=>"110101100",
  30561=>"101011110",
  30562=>"001001111",
  30563=>"100000110",
  30564=>"010000110",
  30565=>"110110111",
  30566=>"011010010",
  30567=>"000111110",
  30568=>"110111110",
  30569=>"000011110",
  30570=>"100011000",
  30571=>"001110100",
  30572=>"111110111",
  30573=>"111001001",
  30574=>"101100111",
  30575=>"100010011",
  30576=>"011000111",
  30577=>"110100111",
  30578=>"100011101",
  30579=>"100100001",
  30580=>"110001001",
  30581=>"111001111",
  30582=>"001001110",
  30583=>"001101011",
  30584=>"110101110",
  30585=>"011000110",
  30586=>"101101100",
  30587=>"001001010",
  30588=>"111011001",
  30589=>"011111010",
  30590=>"000100111",
  30591=>"011010110",
  30592=>"110010101",
  30593=>"110111001",
  30594=>"110110001",
  30595=>"101110010",
  30596=>"111011101",
  30597=>"111110100",
  30598=>"111101000",
  30599=>"100011110",
  30600=>"101000111",
  30601=>"011011111",
  30602=>"000001000",
  30603=>"111101001",
  30604=>"101000110",
  30605=>"000110010",
  30606=>"000100001",
  30607=>"010100111",
  30608=>"100000001",
  30609=>"100010100",
  30610=>"111000110",
  30611=>"101000111",
  30612=>"000110000",
  30613=>"101100110",
  30614=>"001101111",
  30615=>"111011011",
  30616=>"101101001",
  30617=>"101110100",
  30618=>"000010100",
  30619=>"111010100",
  30620=>"010000000",
  30621=>"110000100",
  30622=>"101111100",
  30623=>"111010010",
  30624=>"101111100",
  30625=>"011111111",
  30626=>"010000000",
  30627=>"111111001",
  30628=>"111111000",
  30629=>"011000000",
  30630=>"101000111",
  30631=>"101011001",
  30632=>"100011000",
  30633=>"111110011",
  30634=>"111101101",
  30635=>"011010010",
  30636=>"010111001",
  30637=>"111011100",
  30638=>"101001011",
  30639=>"000011100",
  30640=>"111110101",
  30641=>"100010101",
  30642=>"000011110",
  30643=>"100010100",
  30644=>"101101111",
  30645=>"010100001",
  30646=>"101110011",
  30647=>"110000101",
  30648=>"101000011",
  30649=>"101011010",
  30650=>"001010011",
  30651=>"111101011",
  30652=>"000111110",
  30653=>"110001100",
  30654=>"000101110",
  30655=>"100111111",
  30656=>"010100110",
  30657=>"010011111",
  30658=>"010011001",
  30659=>"010110000",
  30660=>"000010100",
  30661=>"000101010",
  30662=>"001101001",
  30663=>"001101000",
  30664=>"111001101",
  30665=>"011101011",
  30666=>"001101100",
  30667=>"101001011",
  30668=>"000001111",
  30669=>"111111110",
  30670=>"000100011",
  30671=>"010111101",
  30672=>"100101000",
  30673=>"011000101",
  30674=>"111010100",
  30675=>"111011110",
  30676=>"101110010",
  30677=>"100001001",
  30678=>"000011111",
  30679=>"001000110",
  30680=>"000000111",
  30681=>"010000010",
  30682=>"111111111",
  30683=>"100000111",
  30684=>"000010100",
  30685=>"001011100",
  30686=>"111010001",
  30687=>"111011111",
  30688=>"101100100",
  30689=>"001101101",
  30690=>"010101011",
  30691=>"100110110",
  30692=>"111111000",
  30693=>"111001011",
  30694=>"110110101",
  30695=>"110011010",
  30696=>"111011011",
  30697=>"110010110",
  30698=>"101110001",
  30699=>"111010001",
  30700=>"101101011",
  30701=>"110010000",
  30702=>"000011101",
  30703=>"011100010",
  30704=>"101000011",
  30705=>"110110000",
  30706=>"101001110",
  30707=>"000000011",
  30708=>"100001101",
  30709=>"111111001",
  30710=>"001000000",
  30711=>"110000011",
  30712=>"001111111",
  30713=>"111010000",
  30714=>"001100111",
  30715=>"010100100",
  30716=>"011000010",
  30717=>"011001110",
  30718=>"001101001",
  30719=>"111001010",
  30720=>"111101001",
  30721=>"001011100",
  30722=>"111010011",
  30723=>"010000000",
  30724=>"111110001",
  30725=>"100110001",
  30726=>"000000011",
  30727=>"110111001",
  30728=>"011011000",
  30729=>"100011100",
  30730=>"010101011",
  30731=>"101010000",
  30732=>"111001111",
  30733=>"111110010",
  30734=>"110001011",
  30735=>"111111010",
  30736=>"001000001",
  30737=>"001100001",
  30738=>"011000000",
  30739=>"101111111",
  30740=>"111101101",
  30741=>"110001001",
  30742=>"101101110",
  30743=>"000100001",
  30744=>"111000111",
  30745=>"011000010",
  30746=>"000101101",
  30747=>"100001000",
  30748=>"100101000",
  30749=>"100011100",
  30750=>"000100010",
  30751=>"100000010",
  30752=>"011001011",
  30753=>"000010000",
  30754=>"010111110",
  30755=>"010001000",
  30756=>"000101100",
  30757=>"011110000",
  30758=>"111001111",
  30759=>"101101001",
  30760=>"111001100",
  30761=>"111111110",
  30762=>"000100000",
  30763=>"100000000",
  30764=>"101100001",
  30765=>"111011010",
  30766=>"010010110",
  30767=>"111011110",
  30768=>"011010111",
  30769=>"010010001",
  30770=>"100001100",
  30771=>"100101101",
  30772=>"110000101",
  30773=>"111000110",
  30774=>"000010111",
  30775=>"101011101",
  30776=>"100010000",
  30777=>"010100010",
  30778=>"110111111",
  30779=>"110000110",
  30780=>"100010010",
  30781=>"100001010",
  30782=>"110011101",
  30783=>"101011001",
  30784=>"010101111",
  30785=>"101100110",
  30786=>"001001101",
  30787=>"111000111",
  30788=>"000000100",
  30789=>"111000111",
  30790=>"011110010",
  30791=>"110001101",
  30792=>"101001000",
  30793=>"001111100",
  30794=>"110001011",
  30795=>"100110110",
  30796=>"010001010",
  30797=>"001001001",
  30798=>"110000000",
  30799=>"100010000",
  30800=>"100010110",
  30801=>"010010001",
  30802=>"100000001",
  30803=>"100001000",
  30804=>"101011000",
  30805=>"001010110",
  30806=>"000000000",
  30807=>"011111110",
  30808=>"011100111",
  30809=>"001010110",
  30810=>"000010010",
  30811=>"000000001",
  30812=>"000001011",
  30813=>"001111010",
  30814=>"011110001",
  30815=>"010000011",
  30816=>"010001100",
  30817=>"100110111",
  30818=>"111100101",
  30819=>"011001110",
  30820=>"110111111",
  30821=>"111111001",
  30822=>"110001000",
  30823=>"111110010",
  30824=>"101100100",
  30825=>"010010010",
  30826=>"110110001",
  30827=>"110101010",
  30828=>"011001010",
  30829=>"001001100",
  30830=>"011000010",
  30831=>"010111000",
  30832=>"010000000",
  30833=>"000111010",
  30834=>"001000001",
  30835=>"011101110",
  30836=>"101101011",
  30837=>"010000001",
  30838=>"010000110",
  30839=>"100100011",
  30840=>"000100100",
  30841=>"001011001",
  30842=>"010100110",
  30843=>"000101011",
  30844=>"010011111",
  30845=>"100011110",
  30846=>"010010110",
  30847=>"100011111",
  30848=>"010001011",
  30849=>"000001011",
  30850=>"111001000",
  30851=>"100001110",
  30852=>"101000110",
  30853=>"100111010",
  30854=>"101011110",
  30855=>"001011100",
  30856=>"111001001",
  30857=>"011001101",
  30858=>"010011011",
  30859=>"011000110",
  30860=>"111000000",
  30861=>"001111000",
  30862=>"100001100",
  30863=>"001111011",
  30864=>"010110110",
  30865=>"000011100",
  30866=>"011101011",
  30867=>"000110011",
  30868=>"101111000",
  30869=>"111101011",
  30870=>"000001000",
  30871=>"110001000",
  30872=>"101100011",
  30873=>"101101000",
  30874=>"111010110",
  30875=>"110011101",
  30876=>"000101100",
  30877=>"100100101",
  30878=>"111111100",
  30879=>"111000101",
  30880=>"011100000",
  30881=>"111011010",
  30882=>"010100110",
  30883=>"110101110",
  30884=>"111011100",
  30885=>"001011010",
  30886=>"101101110",
  30887=>"101001101",
  30888=>"001111011",
  30889=>"100100111",
  30890=>"110111111",
  30891=>"000110001",
  30892=>"001100110",
  30893=>"010101010",
  30894=>"000110011",
  30895=>"110100010",
  30896=>"100011001",
  30897=>"011111111",
  30898=>"111111101",
  30899=>"001100001",
  30900=>"111110010",
  30901=>"010100101",
  30902=>"111100000",
  30903=>"001001100",
  30904=>"010011110",
  30905=>"110100011",
  30906=>"010101011",
  30907=>"001110000",
  30908=>"010010100",
  30909=>"110100111",
  30910=>"101100001",
  30911=>"101001011",
  30912=>"100101101",
  30913=>"001011100",
  30914=>"110010011",
  30915=>"010111111",
  30916=>"111000010",
  30917=>"100010001",
  30918=>"111010111",
  30919=>"011101111",
  30920=>"110010110",
  30921=>"101110101",
  30922=>"111000011",
  30923=>"110010111",
  30924=>"111101111",
  30925=>"111101011",
  30926=>"110010001",
  30927=>"011000100",
  30928=>"100001000",
  30929=>"111001001",
  30930=>"000000000",
  30931=>"001010001",
  30932=>"111110101",
  30933=>"111011101",
  30934=>"100000000",
  30935=>"010111111",
  30936=>"101011000",
  30937=>"111111110",
  30938=>"101001000",
  30939=>"111011001",
  30940=>"100001111",
  30941=>"100101111",
  30942=>"000011001",
  30943=>"011010010",
  30944=>"110101010",
  30945=>"010001111",
  30946=>"010000101",
  30947=>"000000011",
  30948=>"110100100",
  30949=>"010000000",
  30950=>"010011110",
  30951=>"011001000",
  30952=>"110101100",
  30953=>"110000101",
  30954=>"001000011",
  30955=>"110001010",
  30956=>"010010000",
  30957=>"100100001",
  30958=>"110100111",
  30959=>"110100001",
  30960=>"000001111",
  30961=>"011000101",
  30962=>"101000010",
  30963=>"001010100",
  30964=>"010011111",
  30965=>"100010110",
  30966=>"101111100",
  30967=>"110010000",
  30968=>"111110110",
  30969=>"010101000",
  30970=>"100000001",
  30971=>"100101111",
  30972=>"110100010",
  30973=>"101101101",
  30974=>"011010100",
  30975=>"111010100",
  30976=>"100000100",
  30977=>"001111101",
  30978=>"111001100",
  30979=>"101011111",
  30980=>"111110000",
  30981=>"000110101",
  30982=>"001001001",
  30983=>"010011001",
  30984=>"101110001",
  30985=>"011111111",
  30986=>"000110001",
  30987=>"010100100",
  30988=>"100111001",
  30989=>"110101101",
  30990=>"101100101",
  30991=>"011000111",
  30992=>"000000110",
  30993=>"111011000",
  30994=>"000000011",
  30995=>"001011110",
  30996=>"101010001",
  30997=>"000010111",
  30998=>"101001110",
  30999=>"100111110",
  31000=>"100111000",
  31001=>"110000111",
  31002=>"000010100",
  31003=>"001010010",
  31004=>"000101010",
  31005=>"111000010",
  31006=>"101101101",
  31007=>"000010110",
  31008=>"010111100",
  31009=>"110111110",
  31010=>"100110111",
  31011=>"011111111",
  31012=>"000000001",
  31013=>"100001000",
  31014=>"110101001",
  31015=>"110011111",
  31016=>"100100111",
  31017=>"110010001",
  31018=>"000110000",
  31019=>"110101111",
  31020=>"010010011",
  31021=>"111110010",
  31022=>"010110100",
  31023=>"000011010",
  31024=>"101000000",
  31025=>"010100011",
  31026=>"010110101",
  31027=>"000011100",
  31028=>"001110100",
  31029=>"100001111",
  31030=>"111111001",
  31031=>"111010101",
  31032=>"101011001",
  31033=>"111010100",
  31034=>"100100001",
  31035=>"100000000",
  31036=>"100110011",
  31037=>"111110001",
  31038=>"010101011",
  31039=>"011011101",
  31040=>"101000011",
  31041=>"000001000",
  31042=>"101001010",
  31043=>"001000110",
  31044=>"011000001",
  31045=>"111010001",
  31046=>"111011010",
  31047=>"011110010",
  31048=>"101000101",
  31049=>"000101001",
  31050=>"001110000",
  31051=>"000110000",
  31052=>"100101111",
  31053=>"100010001",
  31054=>"100101101",
  31055=>"001101011",
  31056=>"011100001",
  31057=>"101110110",
  31058=>"111011110",
  31059=>"111011010",
  31060=>"000101000",
  31061=>"110010111",
  31062=>"100100100",
  31063=>"010110011",
  31064=>"001111001",
  31065=>"010000110",
  31066=>"100011011",
  31067=>"100100010",
  31068=>"100101000",
  31069=>"110001011",
  31070=>"000110101",
  31071=>"110010001",
  31072=>"111100100",
  31073=>"001100110",
  31074=>"101100011",
  31075=>"100100111",
  31076=>"111011000",
  31077=>"111111011",
  31078=>"000010111",
  31079=>"101100100",
  31080=>"000001010",
  31081=>"011000001",
  31082=>"100001111",
  31083=>"111011110",
  31084=>"101011110",
  31085=>"010001101",
  31086=>"111111011",
  31087=>"010001001",
  31088=>"001000101",
  31089=>"011011101",
  31090=>"100001111",
  31091=>"111110010",
  31092=>"101010111",
  31093=>"010100001",
  31094=>"110110111",
  31095=>"101100000",
  31096=>"110101110",
  31097=>"011111001",
  31098=>"000011011",
  31099=>"001111101",
  31100=>"101101001",
  31101=>"100110010",
  31102=>"100110100",
  31103=>"011001001",
  31104=>"001000111",
  31105=>"011110111",
  31106=>"101111010",
  31107=>"000001010",
  31108=>"010000111",
  31109=>"100110011",
  31110=>"001111010",
  31111=>"111010010",
  31112=>"010010110",
  31113=>"000100001",
  31114=>"000001001",
  31115=>"101000110",
  31116=>"010001010",
  31117=>"000000000",
  31118=>"011000111",
  31119=>"101001110",
  31120=>"000100100",
  31121=>"010001101",
  31122=>"111011010",
  31123=>"001010011",
  31124=>"101011011",
  31125=>"111101010",
  31126=>"001110010",
  31127=>"101010011",
  31128=>"001010010",
  31129=>"111100111",
  31130=>"001101111",
  31131=>"000101000",
  31132=>"010000100",
  31133=>"100111101",
  31134=>"010000101",
  31135=>"110011111",
  31136=>"110010011",
  31137=>"111111011",
  31138=>"111000101",
  31139=>"011010011",
  31140=>"111110001",
  31141=>"100100110",
  31142=>"111111000",
  31143=>"011001011",
  31144=>"000101111",
  31145=>"101110111",
  31146=>"000011000",
  31147=>"100100111",
  31148=>"010000100",
  31149=>"010110001",
  31150=>"101000011",
  31151=>"100011111",
  31152=>"111011011",
  31153=>"101010000",
  31154=>"101010001",
  31155=>"011100110",
  31156=>"101111100",
  31157=>"110101101",
  31158=>"101110011",
  31159=>"101011100",
  31160=>"011000100",
  31161=>"010011100",
  31162=>"010100000",
  31163=>"010110001",
  31164=>"001111111",
  31165=>"100011011",
  31166=>"100110000",
  31167=>"000011000",
  31168=>"001101000",
  31169=>"111101100",
  31170=>"101110011",
  31171=>"100001001",
  31172=>"000111010",
  31173=>"001001000",
  31174=>"000001001",
  31175=>"010110000",
  31176=>"011010110",
  31177=>"100001101",
  31178=>"010010011",
  31179=>"010111100",
  31180=>"100010110",
  31181=>"001010010",
  31182=>"100110101",
  31183=>"000010100",
  31184=>"111000100",
  31185=>"001110111",
  31186=>"100110010",
  31187=>"000010010",
  31188=>"110110100",
  31189=>"101101111",
  31190=>"010000111",
  31191=>"001110110",
  31192=>"110011101",
  31193=>"001001111",
  31194=>"110111100",
  31195=>"100001101",
  31196=>"011001110",
  31197=>"000011110",
  31198=>"000100000",
  31199=>"100010010",
  31200=>"110100110",
  31201=>"001110100",
  31202=>"011000011",
  31203=>"001100111",
  31204=>"000011010",
  31205=>"110011000",
  31206=>"001100000",
  31207=>"111000111",
  31208=>"010001011",
  31209=>"011100111",
  31210=>"101101101",
  31211=>"000110011",
  31212=>"000110100",
  31213=>"110111001",
  31214=>"000001101",
  31215=>"111101001",
  31216=>"011011100",
  31217=>"111001100",
  31218=>"111101111",
  31219=>"111000000",
  31220=>"111001111",
  31221=>"111001101",
  31222=>"001110001",
  31223=>"100100101",
  31224=>"000001000",
  31225=>"101101000",
  31226=>"000011011",
  31227=>"100011111",
  31228=>"010110001",
  31229=>"011100001",
  31230=>"010001010",
  31231=>"010001111",
  31232=>"001110101",
  31233=>"010010111",
  31234=>"101010010",
  31235=>"000111010",
  31236=>"001101100",
  31237=>"000111110",
  31238=>"000000110",
  31239=>"100001100",
  31240=>"101000101",
  31241=>"111011000",
  31242=>"100010011",
  31243=>"011101010",
  31244=>"000000000",
  31245=>"110011010",
  31246=>"100001100",
  31247=>"110001101",
  31248=>"110001111",
  31249=>"010101110",
  31250=>"111101100",
  31251=>"111111111",
  31252=>"101010101",
  31253=>"010000001",
  31254=>"001011101",
  31255=>"101010101",
  31256=>"011111111",
  31257=>"001100111",
  31258=>"110110010",
  31259=>"000111111",
  31260=>"011110111",
  31261=>"100110101",
  31262=>"100011011",
  31263=>"000001101",
  31264=>"110111001",
  31265=>"011011110",
  31266=>"101000010",
  31267=>"001100010",
  31268=>"100010001",
  31269=>"111000001",
  31270=>"010100001",
  31271=>"101100011",
  31272=>"000000000",
  31273=>"011111111",
  31274=>"011110101",
  31275=>"011111010",
  31276=>"011100010",
  31277=>"011101110",
  31278=>"011010111",
  31279=>"111101011",
  31280=>"000000101",
  31281=>"000011111",
  31282=>"001110000",
  31283=>"100011101",
  31284=>"010101110",
  31285=>"110111000",
  31286=>"101001100",
  31287=>"000010000",
  31288=>"101001100",
  31289=>"011101111",
  31290=>"000011110",
  31291=>"101010000",
  31292=>"111010111",
  31293=>"001010011",
  31294=>"111011111",
  31295=>"100011111",
  31296=>"010001100",
  31297=>"000011101",
  31298=>"110010011",
  31299=>"010100011",
  31300=>"001111111",
  31301=>"100000101",
  31302=>"011011111",
  31303=>"101001000",
  31304=>"100101111",
  31305=>"000000101",
  31306=>"111110001",
  31307=>"101000010",
  31308=>"011000001",
  31309=>"011011001",
  31310=>"001000011",
  31311=>"010100000",
  31312=>"101010010",
  31313=>"010000100",
  31314=>"000100010",
  31315=>"101010101",
  31316=>"010010010",
  31317=>"010101010",
  31318=>"100011011",
  31319=>"001100010",
  31320=>"010100000",
  31321=>"010101111",
  31322=>"110101111",
  31323=>"011101110",
  31324=>"010111100",
  31325=>"101111011",
  31326=>"111000110",
  31327=>"111110000",
  31328=>"000010110",
  31329=>"011011111",
  31330=>"101100000",
  31331=>"111011011",
  31332=>"100110101",
  31333=>"011001110",
  31334=>"001000101",
  31335=>"111111101",
  31336=>"001100000",
  31337=>"000000111",
  31338=>"101001110",
  31339=>"111011000",
  31340=>"111110011",
  31341=>"000101100",
  31342=>"001110101",
  31343=>"110101000",
  31344=>"101010111",
  31345=>"100110100",
  31346=>"101110101",
  31347=>"110100110",
  31348=>"001110110",
  31349=>"001101011",
  31350=>"110001000",
  31351=>"111101111",
  31352=>"010001010",
  31353=>"100111100",
  31354=>"101010101",
  31355=>"100100010",
  31356=>"110011010",
  31357=>"111010111",
  31358=>"010100011",
  31359=>"101010100",
  31360=>"000111100",
  31361=>"110101101",
  31362=>"011101011",
  31363=>"001101101",
  31364=>"101111111",
  31365=>"111010001",
  31366=>"100110111",
  31367=>"100000100",
  31368=>"101100110",
  31369=>"011111111",
  31370=>"001110010",
  31371=>"010000001",
  31372=>"001011101",
  31373=>"100000000",
  31374=>"001110001",
  31375=>"100111101",
  31376=>"001010000",
  31377=>"111000111",
  31378=>"001011001",
  31379=>"101001000",
  31380=>"010111111",
  31381=>"101111101",
  31382=>"110000110",
  31383=>"001001000",
  31384=>"100111111",
  31385=>"111010001",
  31386=>"100000011",
  31387=>"110010100",
  31388=>"100010010",
  31389=>"000100100",
  31390=>"011011101",
  31391=>"110000011",
  31392=>"111101010",
  31393=>"110111100",
  31394=>"000000110",
  31395=>"110100101",
  31396=>"010100100",
  31397=>"010101000",
  31398=>"011101101",
  31399=>"010100011",
  31400=>"010010110",
  31401=>"010111110",
  31402=>"010010000",
  31403=>"101010100",
  31404=>"010001001",
  31405=>"111100101",
  31406=>"100110100",
  31407=>"000101110",
  31408=>"101111001",
  31409=>"001000010",
  31410=>"111111100",
  31411=>"101010101",
  31412=>"010011001",
  31413=>"000010100",
  31414=>"101101100",
  31415=>"101110010",
  31416=>"110010100",
  31417=>"101100001",
  31418=>"111010101",
  31419=>"010000000",
  31420=>"010001001",
  31421=>"111011010",
  31422=>"111010000",
  31423=>"110100001",
  31424=>"111110111",
  31425=>"001110111",
  31426=>"000110000",
  31427=>"111001000",
  31428=>"110101000",
  31429=>"001101001",
  31430=>"010101001",
  31431=>"001101111",
  31432=>"010010010",
  31433=>"001100001",
  31434=>"011110000",
  31435=>"100111001",
  31436=>"000101100",
  31437=>"100101110",
  31438=>"101011111",
  31439=>"011101000",
  31440=>"110110111",
  31441=>"100010000",
  31442=>"010100010",
  31443=>"001000010",
  31444=>"010110100",
  31445=>"001101111",
  31446=>"101000100",
  31447=>"110100111",
  31448=>"000100111",
  31449=>"000001000",
  31450=>"000000110",
  31451=>"110101101",
  31452=>"000111001",
  31453=>"010010111",
  31454=>"000100111",
  31455=>"110011101",
  31456=>"101110110",
  31457=>"111011101",
  31458=>"010000111",
  31459=>"010100001",
  31460=>"111100000",
  31461=>"000000110",
  31462=>"000011000",
  31463=>"000001010",
  31464=>"101111111",
  31465=>"110011110",
  31466=>"011110010",
  31467=>"001001010",
  31468=>"000111011",
  31469=>"101011111",
  31470=>"111011100",
  31471=>"100001010",
  31472=>"110011011",
  31473=>"110110011",
  31474=>"000000101",
  31475=>"000000011",
  31476=>"001011000",
  31477=>"001010011",
  31478=>"011110011",
  31479=>"001011110",
  31480=>"001000010",
  31481=>"010101101",
  31482=>"111100000",
  31483=>"001101010",
  31484=>"011111010",
  31485=>"000110110",
  31486=>"110110101",
  31487=>"010110101",
  31488=>"111111000",
  31489=>"101101011",
  31490=>"110001101",
  31491=>"000111110",
  31492=>"000110110",
  31493=>"010011000",
  31494=>"010111110",
  31495=>"100111100",
  31496=>"010101101",
  31497=>"100000101",
  31498=>"000111101",
  31499=>"111111001",
  31500=>"001110011",
  31501=>"100000111",
  31502=>"010101101",
  31503=>"000000110",
  31504=>"110000001",
  31505=>"011000001",
  31506=>"011101001",
  31507=>"001110111",
  31508=>"100110011",
  31509=>"111000001",
  31510=>"101101011",
  31511=>"110000101",
  31512=>"100000110",
  31513=>"000000101",
  31514=>"101100101",
  31515=>"010000111",
  31516=>"010000100",
  31517=>"101100010",
  31518=>"101111110",
  31519=>"000001011",
  31520=>"011001110",
  31521=>"110111100",
  31522=>"011010011",
  31523=>"000111110",
  31524=>"110100001",
  31525=>"101000110",
  31526=>"100001110",
  31527=>"110101010",
  31528=>"001111101",
  31529=>"111011101",
  31530=>"101010001",
  31531=>"001111011",
  31532=>"001101101",
  31533=>"011000111",
  31534=>"000000110",
  31535=>"101001001",
  31536=>"110011010",
  31537=>"110000000",
  31538=>"100110100",
  31539=>"000001111",
  31540=>"100010010",
  31541=>"000110110",
  31542=>"000000110",
  31543=>"010100001",
  31544=>"011011110",
  31545=>"001011000",
  31546=>"110011011",
  31547=>"011101010",
  31548=>"101001110",
  31549=>"100010011",
  31550=>"110000000",
  31551=>"101000001",
  31552=>"100000100",
  31553=>"111011110",
  31554=>"100000001",
  31555=>"000101000",
  31556=>"110100100",
  31557=>"000101110",
  31558=>"010001111",
  31559=>"001111001",
  31560=>"001011110",
  31561=>"101001110",
  31562=>"100011000",
  31563=>"110110001",
  31564=>"010000011",
  31565=>"111000110",
  31566=>"111000000",
  31567=>"010011101",
  31568=>"100110100",
  31569=>"111010111",
  31570=>"100001010",
  31571=>"001101101",
  31572=>"110110010",
  31573=>"011100001",
  31574=>"000100000",
  31575=>"010110101",
  31576=>"000001000",
  31577=>"001111101",
  31578=>"111011110",
  31579=>"111011101",
  31580=>"101100001",
  31581=>"011110110",
  31582=>"011101001",
  31583=>"000011010",
  31584=>"000011111",
  31585=>"001000010",
  31586=>"101111011",
  31587=>"111010011",
  31588=>"010110101",
  31589=>"111011100",
  31590=>"101100000",
  31591=>"000001001",
  31592=>"100011101",
  31593=>"011111000",
  31594=>"010001000",
  31595=>"011111011",
  31596=>"011101010",
  31597=>"011000100",
  31598=>"001101001",
  31599=>"001000010",
  31600=>"000100010",
  31601=>"111011110",
  31602=>"100010110",
  31603=>"001100111",
  31604=>"100011111",
  31605=>"111111011",
  31606=>"100111100",
  31607=>"110010110",
  31608=>"111101000",
  31609=>"010101000",
  31610=>"101111000",
  31611=>"000011000",
  31612=>"011110101",
  31613=>"001101001",
  31614=>"100100010",
  31615=>"100011110",
  31616=>"101111001",
  31617=>"001000100",
  31618=>"101101001",
  31619=>"011010101",
  31620=>"111100110",
  31621=>"100001011",
  31622=>"101101011",
  31623=>"011001001",
  31624=>"010111011",
  31625=>"110100111",
  31626=>"010101001",
  31627=>"100111100",
  31628=>"011110001",
  31629=>"110010110",
  31630=>"010011000",
  31631=>"101110001",
  31632=>"000111001",
  31633=>"001001110",
  31634=>"001101011",
  31635=>"101011011",
  31636=>"011100101",
  31637=>"000011001",
  31638=>"101010100",
  31639=>"101101101",
  31640=>"011111001",
  31641=>"011100111",
  31642=>"011000101",
  31643=>"111110010",
  31644=>"100001010",
  31645=>"010011110",
  31646=>"010101101",
  31647=>"111001111",
  31648=>"011110110",
  31649=>"010011110",
  31650=>"111000100",
  31651=>"010111001",
  31652=>"010000110",
  31653=>"101010001",
  31654=>"010100110",
  31655=>"101011101",
  31656=>"011000010",
  31657=>"111000110",
  31658=>"011101110",
  31659=>"011110111",
  31660=>"100100110",
  31661=>"110000101",
  31662=>"110011101",
  31663=>"101111010",
  31664=>"110011111",
  31665=>"110011010",
  31666=>"111011101",
  31667=>"000000101",
  31668=>"111110111",
  31669=>"011001000",
  31670=>"111010110",
  31671=>"111111000",
  31672=>"000101011",
  31673=>"010111100",
  31674=>"110010001",
  31675=>"100010101",
  31676=>"111101100",
  31677=>"011110110",
  31678=>"100101110",
  31679=>"101011100",
  31680=>"000111000",
  31681=>"000110000",
  31682=>"001110100",
  31683=>"101100101",
  31684=>"000110100",
  31685=>"011001011",
  31686=>"111101111",
  31687=>"111001011",
  31688=>"110111000",
  31689=>"011100101",
  31690=>"111000110",
  31691=>"100111001",
  31692=>"110110111",
  31693=>"001011111",
  31694=>"011011011",
  31695=>"011111110",
  31696=>"011100100",
  31697=>"000001001",
  31698=>"010110101",
  31699=>"001010010",
  31700=>"000010000",
  31701=>"010111100",
  31702=>"011110101",
  31703=>"100010100",
  31704=>"011000011",
  31705=>"110011111",
  31706=>"001100000",
  31707=>"100000110",
  31708=>"110010110",
  31709=>"100000001",
  31710=>"000000101",
  31711=>"011100010",
  31712=>"001100101",
  31713=>"011110110",
  31714=>"000010101",
  31715=>"011000010",
  31716=>"001110111",
  31717=>"000010111",
  31718=>"001110000",
  31719=>"110011110",
  31720=>"000111010",
  31721=>"010011011",
  31722=>"101000100",
  31723=>"001001110",
  31724=>"100111011",
  31725=>"010000000",
  31726=>"111011101",
  31727=>"101110111",
  31728=>"111001011",
  31729=>"100010010",
  31730=>"110100100",
  31731=>"111100011",
  31732=>"101101110",
  31733=>"010010100",
  31734=>"001000111",
  31735=>"000011111",
  31736=>"101100010",
  31737=>"001100010",
  31738=>"001001101",
  31739=>"110100001",
  31740=>"000100001",
  31741=>"100110000",
  31742=>"000110111",
  31743=>"010101100",
  31744=>"000010111",
  31745=>"111101011",
  31746=>"010101010",
  31747=>"110101001",
  31748=>"010000000",
  31749=>"100110100",
  31750=>"101000111",
  31751=>"001001000",
  31752=>"100111001",
  31753=>"001000000",
  31754=>"110100001",
  31755=>"111100101",
  31756=>"100110111",
  31757=>"000110101",
  31758=>"001011010",
  31759=>"110101101",
  31760=>"010101110",
  31761=>"010111101",
  31762=>"010110100",
  31763=>"101000111",
  31764=>"000011111",
  31765=>"010101000",
  31766=>"000010001",
  31767=>"010111000",
  31768=>"101001101",
  31769=>"011110001",
  31770=>"101011000",
  31771=>"111000110",
  31772=>"001000000",
  31773=>"100111110",
  31774=>"010101100",
  31775=>"001001110",
  31776=>"000101100",
  31777=>"001001110",
  31778=>"101011010",
  31779=>"010100001",
  31780=>"100000010",
  31781=>"110011100",
  31782=>"100000010",
  31783=>"110110011",
  31784=>"011111011",
  31785=>"101010001",
  31786=>"100100001",
  31787=>"101111100",
  31788=>"110101001",
  31789=>"111100000",
  31790=>"000001100",
  31791=>"000000010",
  31792=>"011110100",
  31793=>"100011010",
  31794=>"011010010",
  31795=>"001001101",
  31796=>"011111000",
  31797=>"101000001",
  31798=>"011111110",
  31799=>"100100001",
  31800=>"000100001",
  31801=>"110011100",
  31802=>"011000110",
  31803=>"100011101",
  31804=>"011000010",
  31805=>"100010000",
  31806=>"010101010",
  31807=>"100011010",
  31808=>"111010101",
  31809=>"111010110",
  31810=>"010111001",
  31811=>"111010100",
  31812=>"011100111",
  31813=>"000100111",
  31814=>"010110011",
  31815=>"111111010",
  31816=>"001011111",
  31817=>"100110111",
  31818=>"101101111",
  31819=>"010001001",
  31820=>"110011000",
  31821=>"011011001",
  31822=>"100001100",
  31823=>"111100110",
  31824=>"000110001",
  31825=>"010100010",
  31826=>"010001010",
  31827=>"010000011",
  31828=>"001100000",
  31829=>"000101110",
  31830=>"101101100",
  31831=>"001101101",
  31832=>"001100101",
  31833=>"110111100",
  31834=>"001000001",
  31835=>"000000011",
  31836=>"010001110",
  31837=>"001011000",
  31838=>"110100001",
  31839=>"111100101",
  31840=>"101000111",
  31841=>"111100011",
  31842=>"001000110",
  31843=>"001101000",
  31844=>"101011011",
  31845=>"111000100",
  31846=>"001100000",
  31847=>"111011111",
  31848=>"000010000",
  31849=>"011011001",
  31850=>"110100001",
  31851=>"011111101",
  31852=>"001001011",
  31853=>"101110101",
  31854=>"000110110",
  31855=>"010001001",
  31856=>"110001010",
  31857=>"110100111",
  31858=>"001011111",
  31859=>"110111100",
  31860=>"011101001",
  31861=>"011010101",
  31862=>"101000111",
  31863=>"000010001",
  31864=>"011011111",
  31865=>"111110010",
  31866=>"111110101",
  31867=>"010010011",
  31868=>"111111000",
  31869=>"011110011",
  31870=>"101111110",
  31871=>"001001110",
  31872=>"111110100",
  31873=>"010101110",
  31874=>"001011111",
  31875=>"010100000",
  31876=>"100101000",
  31877=>"111010110",
  31878=>"111101000",
  31879=>"001001000",
  31880=>"011010011",
  31881=>"011001010",
  31882=>"110100101",
  31883=>"011000110",
  31884=>"011000100",
  31885=>"110110011",
  31886=>"101011001",
  31887=>"101000110",
  31888=>"001101100",
  31889=>"101011011",
  31890=>"101100001",
  31891=>"001100100",
  31892=>"010110001",
  31893=>"001100110",
  31894=>"100001000",
  31895=>"001001101",
  31896=>"001110111",
  31897=>"011011100",
  31898=>"001101001",
  31899=>"111010110",
  31900=>"010111001",
  31901=>"010000100",
  31902=>"110000001",
  31903=>"101000000",
  31904=>"110010101",
  31905=>"011010011",
  31906=>"000000001",
  31907=>"110001111",
  31908=>"110110111",
  31909=>"001100010",
  31910=>"111110111",
  31911=>"011001101",
  31912=>"011101111",
  31913=>"001010001",
  31914=>"010100101",
  31915=>"010110010",
  31916=>"010010011",
  31917=>"111111001",
  31918=>"100010110",
  31919=>"101011110",
  31920=>"101110000",
  31921=>"010001101",
  31922=>"100110111",
  31923=>"000000100",
  31924=>"011000100",
  31925=>"110000011",
  31926=>"111010110",
  31927=>"111101110",
  31928=>"100101000",
  31929=>"110101110",
  31930=>"110010000",
  31931=>"100101001",
  31932=>"000010000",
  31933=>"110011111",
  31934=>"111011011",
  31935=>"001101000",
  31936=>"011111110",
  31937=>"000110111",
  31938=>"111110010",
  31939=>"101011001",
  31940=>"101011010",
  31941=>"000011001",
  31942=>"011010001",
  31943=>"111101101",
  31944=>"100110100",
  31945=>"111111100",
  31946=>"001110000",
  31947=>"100110111",
  31948=>"000101000",
  31949=>"110000100",
  31950=>"000010001",
  31951=>"100101110",
  31952=>"010010000",
  31953=>"100101110",
  31954=>"000101010",
  31955=>"011011001",
  31956=>"111101000",
  31957=>"110111111",
  31958=>"101100000",
  31959=>"000000011",
  31960=>"101110000",
  31961=>"110110000",
  31962=>"000111011",
  31963=>"011111010",
  31964=>"101000010",
  31965=>"010101110",
  31966=>"001001101",
  31967=>"110111101",
  31968=>"101100111",
  31969=>"011001000",
  31970=>"101111101",
  31971=>"011110010",
  31972=>"101100110",
  31973=>"110111110",
  31974=>"010011110",
  31975=>"111101111",
  31976=>"100110011",
  31977=>"101111111",
  31978=>"110011111",
  31979=>"000011100",
  31980=>"110100110",
  31981=>"110000011",
  31982=>"011011101",
  31983=>"101001011",
  31984=>"100001000",
  31985=>"100000011",
  31986=>"101010000",
  31987=>"001000000",
  31988=>"101111110",
  31989=>"111011111",
  31990=>"011000000",
  31991=>"101100001",
  31992=>"001010111",
  31993=>"110010110",
  31994=>"100010000",
  31995=>"001011111",
  31996=>"010001000",
  31997=>"110110011",
  31998=>"100001111",
  31999=>"100000100",
  32000=>"010111011",
  32001=>"110100110",
  32002=>"001101010",
  32003=>"000100100",
  32004=>"100100011",
  32005=>"000111010",
  32006=>"011001000",
  32007=>"000011101",
  32008=>"010001011",
  32009=>"011001101",
  32010=>"111001111",
  32011=>"000001101",
  32012=>"100000100",
  32013=>"001001101",
  32014=>"010101110",
  32015=>"001011100",
  32016=>"101110110",
  32017=>"111001110",
  32018=>"011001001",
  32019=>"000111010",
  32020=>"000110000",
  32021=>"011000111",
  32022=>"111100110",
  32023=>"001110000",
  32024=>"001010011",
  32025=>"000100110",
  32026=>"001111010",
  32027=>"100001110",
  32028=>"011000001",
  32029=>"110100100",
  32030=>"010010010",
  32031=>"010000001",
  32032=>"011101001",
  32033=>"000110111",
  32034=>"001111010",
  32035=>"000000100",
  32036=>"100110010",
  32037=>"000111100",
  32038=>"000010111",
  32039=>"110100100",
  32040=>"001110101",
  32041=>"110110110",
  32042=>"001100110",
  32043=>"010000000",
  32044=>"100111101",
  32045=>"000101100",
  32046=>"011001001",
  32047=>"110100100",
  32048=>"111001110",
  32049=>"000000000",
  32050=>"111000111",
  32051=>"000000111",
  32052=>"100111110",
  32053=>"111010011",
  32054=>"110111100",
  32055=>"111000010",
  32056=>"011011100",
  32057=>"101101001",
  32058=>"111011011",
  32059=>"011011011",
  32060=>"010001000",
  32061=>"111001100",
  32062=>"111111110",
  32063=>"010111100",
  32064=>"001101000",
  32065=>"001010001",
  32066=>"111010000",
  32067=>"010001011",
  32068=>"010011110",
  32069=>"001100010",
  32070=>"011101111",
  32071=>"011010011",
  32072=>"111011000",
  32073=>"111101100",
  32074=>"001000111",
  32075=>"011111000",
  32076=>"000101101",
  32077=>"111101001",
  32078=>"000000001",
  32079=>"110011011",
  32080=>"001010101",
  32081=>"010000101",
  32082=>"111111011",
  32083=>"100011010",
  32084=>"101000010",
  32085=>"001001000",
  32086=>"000110001",
  32087=>"100001110",
  32088=>"010011000",
  32089=>"000001001",
  32090=>"100101100",
  32091=>"111100110",
  32092=>"101101011",
  32093=>"111110100",
  32094=>"010010001",
  32095=>"110001111",
  32096=>"110010001",
  32097=>"011101010",
  32098=>"010011110",
  32099=>"001010000",
  32100=>"001000001",
  32101=>"101011100",
  32102=>"110110010",
  32103=>"010101000",
  32104=>"110101001",
  32105=>"101011000",
  32106=>"110111001",
  32107=>"000011100",
  32108=>"101101100",
  32109=>"001010010",
  32110=>"010110010",
  32111=>"011011100",
  32112=>"001101101",
  32113=>"101100000",
  32114=>"100000001",
  32115=>"110100010",
  32116=>"100001001",
  32117=>"010101001",
  32118=>"010100100",
  32119=>"000011101",
  32120=>"000011011",
  32121=>"110111110",
  32122=>"110010000",
  32123=>"101111110",
  32124=>"000110010",
  32125=>"111011110",
  32126=>"111101010",
  32127=>"100111111",
  32128=>"101100101",
  32129=>"000100110",
  32130=>"000101110",
  32131=>"011110111",
  32132=>"011111111",
  32133=>"000111101",
  32134=>"101101101",
  32135=>"110101011",
  32136=>"101100101",
  32137=>"001010001",
  32138=>"111010111",
  32139=>"111111000",
  32140=>"011001100",
  32141=>"011001010",
  32142=>"101101011",
  32143=>"101011111",
  32144=>"010110101",
  32145=>"010011000",
  32146=>"100011100",
  32147=>"100010011",
  32148=>"000001100",
  32149=>"010011111",
  32150=>"011101111",
  32151=>"110100010",
  32152=>"001110011",
  32153=>"101011001",
  32154=>"011110110",
  32155=>"110111001",
  32156=>"100101100",
  32157=>"011010100",
  32158=>"011100100",
  32159=>"010010000",
  32160=>"101000001",
  32161=>"100001000",
  32162=>"011000000",
  32163=>"000001001",
  32164=>"110100111",
  32165=>"010000011",
  32166=>"011000001",
  32167=>"110000100",
  32168=>"110001110",
  32169=>"011101111",
  32170=>"111110100",
  32171=>"010010110",
  32172=>"111101010",
  32173=>"000000110",
  32174=>"010110111",
  32175=>"111001011",
  32176=>"111100101",
  32177=>"011111111",
  32178=>"111001110",
  32179=>"001001011",
  32180=>"000011110",
  32181=>"101010001",
  32182=>"101110110",
  32183=>"101010010",
  32184=>"001100000",
  32185=>"000000000",
  32186=>"101110101",
  32187=>"010000011",
  32188=>"010101011",
  32189=>"100111110",
  32190=>"100010110",
  32191=>"000110000",
  32192=>"010101111",
  32193=>"010101010",
  32194=>"101110101",
  32195=>"110011101",
  32196=>"001100000",
  32197=>"110110101",
  32198=>"111000101",
  32199=>"000000001",
  32200=>"001001010",
  32201=>"110011110",
  32202=>"011011010",
  32203=>"000011111",
  32204=>"011100101",
  32205=>"101110011",
  32206=>"001011111",
  32207=>"000111000",
  32208=>"110101110",
  32209=>"101100001",
  32210=>"110000010",
  32211=>"010001100",
  32212=>"010101001",
  32213=>"110010000",
  32214=>"100101010",
  32215=>"010001110",
  32216=>"000011011",
  32217=>"001110111",
  32218=>"010110101",
  32219=>"110001000",
  32220=>"000010000",
  32221=>"111011101",
  32222=>"110011111",
  32223=>"000001111",
  32224=>"110000001",
  32225=>"111111100",
  32226=>"110110111",
  32227=>"010111110",
  32228=>"110010101",
  32229=>"111001011",
  32230=>"010111001",
  32231=>"001010011",
  32232=>"010010011",
  32233=>"100110101",
  32234=>"110110110",
  32235=>"010000001",
  32236=>"101001110",
  32237=>"100100111",
  32238=>"000010000",
  32239=>"111100010",
  32240=>"100100011",
  32241=>"100011111",
  32242=>"111001011",
  32243=>"010001011",
  32244=>"001110011",
  32245=>"011110110",
  32246=>"011111001",
  32247=>"011010111",
  32248=>"111110010",
  32249=>"000001001",
  32250=>"010100001",
  32251=>"001011100",
  32252=>"010011000",
  32253=>"011000010",
  32254=>"000011111",
  32255=>"010111101",
  32256=>"110100000",
  32257=>"001000001",
  32258=>"101111101",
  32259=>"110101111",
  32260=>"101101100",
  32261=>"000001110",
  32262=>"110100111",
  32263=>"011011110",
  32264=>"101001110",
  32265=>"101000011",
  32266=>"100010011",
  32267=>"010000110",
  32268=>"111100100",
  32269=>"010111110",
  32270=>"101100101",
  32271=>"001000001",
  32272=>"110101010",
  32273=>"110110100",
  32274=>"110101011",
  32275=>"100011011",
  32276=>"011000111",
  32277=>"100001110",
  32278=>"000111100",
  32279=>"111111110",
  32280=>"110110100",
  32281=>"110010000",
  32282=>"101001000",
  32283=>"110110001",
  32284=>"101100001",
  32285=>"011111100",
  32286=>"111011110",
  32287=>"001001110",
  32288=>"010001110",
  32289=>"110101000",
  32290=>"100101011",
  32291=>"011011110",
  32292=>"101001110",
  32293=>"101001011",
  32294=>"000111101",
  32295=>"111100110",
  32296=>"000010101",
  32297=>"111011011",
  32298=>"010000111",
  32299=>"000100101",
  32300=>"100010010",
  32301=>"000111011",
  32302=>"011011100",
  32303=>"011011101",
  32304=>"111011001",
  32305=>"110101111",
  32306=>"010111011",
  32307=>"000100000",
  32308=>"001101000",
  32309=>"011100110",
  32310=>"100000100",
  32311=>"011110011",
  32312=>"010100000",
  32313=>"010110101",
  32314=>"011101111",
  32315=>"100110000",
  32316=>"000010110",
  32317=>"010110100",
  32318=>"000011111",
  32319=>"011110001",
  32320=>"010000010",
  32321=>"000111101",
  32322=>"100000000",
  32323=>"101010101",
  32324=>"100101101",
  32325=>"011111010",
  32326=>"010000001",
  32327=>"111011000",
  32328=>"010010101",
  32329=>"110101010",
  32330=>"101011010",
  32331=>"100100000",
  32332=>"000100001",
  32333=>"101100100",
  32334=>"101111110",
  32335=>"000001000",
  32336=>"010101010",
  32337=>"100001100",
  32338=>"101111011",
  32339=>"010010001",
  32340=>"111010110",
  32341=>"101000100",
  32342=>"001000110",
  32343=>"001100110",
  32344=>"101001000",
  32345=>"101111100",
  32346=>"010000011",
  32347=>"010001011",
  32348=>"010100101",
  32349=>"000100000",
  32350=>"100011100",
  32351=>"001100111",
  32352=>"001011000",
  32353=>"001100101",
  32354=>"111110010",
  32355=>"110110110",
  32356=>"001110000",
  32357=>"101110010",
  32358=>"001100111",
  32359=>"011000111",
  32360=>"010110000",
  32361=>"011000100",
  32362=>"111111101",
  32363=>"100100101",
  32364=>"110011100",
  32365=>"100010010",
  32366=>"100000111",
  32367=>"100100101",
  32368=>"101101001",
  32369=>"001000101",
  32370=>"110111001",
  32371=>"010011011",
  32372=>"110101111",
  32373=>"000101010",
  32374=>"111101101",
  32375=>"101111101",
  32376=>"000001010",
  32377=>"011101000",
  32378=>"001011000",
  32379=>"111101001",
  32380=>"010010001",
  32381=>"011011100",
  32382=>"110010101",
  32383=>"100011101",
  32384=>"011110100",
  32385=>"010111111",
  32386=>"010111111",
  32387=>"011000110",
  32388=>"000000011",
  32389=>"101110100",
  32390=>"101011110",
  32391=>"010011000",
  32392=>"111010101",
  32393=>"100010111",
  32394=>"011000000",
  32395=>"010001100",
  32396=>"001101111",
  32397=>"011001101",
  32398=>"010010010",
  32399=>"011111010",
  32400=>"011011110",
  32401=>"110110111",
  32402=>"101000000",
  32403=>"111011111",
  32404=>"110000101",
  32405=>"111111000",
  32406=>"100101101",
  32407=>"101010101",
  32408=>"011011101",
  32409=>"101001101",
  32410=>"000110110",
  32411=>"100111100",
  32412=>"111010110",
  32413=>"100100000",
  32414=>"111110011",
  32415=>"101001000",
  32416=>"000100011",
  32417=>"010011011",
  32418=>"011000110",
  32419=>"111000010",
  32420=>"101000011",
  32421=>"010001101",
  32422=>"101010000",
  32423=>"000001011",
  32424=>"111010010",
  32425=>"000000100",
  32426=>"011110111",
  32427=>"111001001",
  32428=>"010110000",
  32429=>"100001000",
  32430=>"100010000",
  32431=>"101010100",
  32432=>"111001011",
  32433=>"100010000",
  32434=>"100111110",
  32435=>"101000001",
  32436=>"010111111",
  32437=>"001111011",
  32438=>"100000000",
  32439=>"101000110",
  32440=>"111010101",
  32441=>"101100111",
  32442=>"011101001",
  32443=>"111100101",
  32444=>"100101111",
  32445=>"011011100",
  32446=>"111000111",
  32447=>"001000000",
  32448=>"110111110",
  32449=>"000010011",
  32450=>"000111100",
  32451=>"110000000",
  32452=>"000100110",
  32453=>"110111010",
  32454=>"001010111",
  32455=>"111110111",
  32456=>"000010110",
  32457=>"111101101",
  32458=>"011111100",
  32459=>"111001011",
  32460=>"011101001",
  32461=>"010110011",
  32462=>"000000110",
  32463=>"100101011",
  32464=>"101001100",
  32465=>"100111011",
  32466=>"111110010",
  32467=>"100111111",
  32468=>"101000011",
  32469=>"011001011",
  32470=>"000100100",
  32471=>"111110110",
  32472=>"001011111",
  32473=>"110011001",
  32474=>"001001000",
  32475=>"010010111",
  32476=>"010000101",
  32477=>"000000001",
  32478=>"100000010",
  32479=>"100111111",
  32480=>"000110000",
  32481=>"000000011",
  32482=>"101011001",
  32483=>"101101101",
  32484=>"011101101",
  32485=>"000100100",
  32486=>"000001100",
  32487=>"001010000",
  32488=>"100001001",
  32489=>"110111100",
  32490=>"101011101",
  32491=>"010000100",
  32492=>"010001101",
  32493=>"000000000",
  32494=>"000101000",
  32495=>"001010100",
  32496=>"101110100",
  32497=>"000010111",
  32498=>"110111100",
  32499=>"111011100",
  32500=>"001100111",
  32501=>"100000011",
  32502=>"100001000",
  32503=>"111001011",
  32504=>"010101011",
  32505=>"101100101",
  32506=>"100011110",
  32507=>"110001100",
  32508=>"100100111",
  32509=>"011110011",
  32510=>"101111101",
  32511=>"101010010",
  32512=>"010110110",
  32513=>"110100100",
  32514=>"001110110",
  32515=>"001110110",
  32516=>"100000001",
  32517=>"111100001",
  32518=>"001000001",
  32519=>"111011000",
  32520=>"100001000",
  32521=>"001011100",
  32522=>"001101100",
  32523=>"101101000",
  32524=>"001011011",
  32525=>"111011011",
  32526=>"100011111",
  32527=>"000101010",
  32528=>"010001011",
  32529=>"010001001",
  32530=>"101001001",
  32531=>"011010001",
  32532=>"010110101",
  32533=>"000000111",
  32534=>"110101110",
  32535=>"101001111",
  32536=>"111101101",
  32537=>"101100101",
  32538=>"000101111",
  32539=>"111011110",
  32540=>"111100100",
  32541=>"001010111",
  32542=>"101001111",
  32543=>"100000101",
  32544=>"010000000",
  32545=>"001011111",
  32546=>"000101001",
  32547=>"111011100",
  32548=>"101111010",
  32549=>"111101100",
  32550=>"001001011",
  32551=>"101001101",
  32552=>"110000110",
  32553=>"000100100",
  32554=>"010111011",
  32555=>"001101001",
  32556=>"000100000",
  32557=>"001110000",
  32558=>"101110000",
  32559=>"111100001",
  32560=>"001110111",
  32561=>"010000001",
  32562=>"000100110",
  32563=>"001011100",
  32564=>"000010001",
  32565=>"111110010",
  32566=>"000110011",
  32567=>"010101000",
  32568=>"110101011",
  32569=>"010101111",
  32570=>"001000011",
  32571=>"011000110",
  32572=>"010100010",
  32573=>"100110001",
  32574=>"111011100",
  32575=>"011101110",
  32576=>"101001011",
  32577=>"111110010",
  32578=>"101100110",
  32579=>"111111111",
  32580=>"000110001",
  32581=>"111001011",
  32582=>"001110101",
  32583=>"111111011",
  32584=>"010000111",
  32585=>"111001111",
  32586=>"111101100",
  32587=>"111111100",
  32588=>"111111011",
  32589=>"111101001",
  32590=>"111000010",
  32591=>"000000001",
  32592=>"111111101",
  32593=>"000000011",
  32594=>"001001111",
  32595=>"110001001",
  32596=>"101100001",
  32597=>"001011000",
  32598=>"011010011",
  32599=>"001101010",
  32600=>"011100001",
  32601=>"001011110",
  32602=>"010100100",
  32603=>"010110000",
  32604=>"101000111",
  32605=>"010000000",
  32606=>"110000010",
  32607=>"000000010",
  32608=>"011110000",
  32609=>"000011101",
  32610=>"011000000",
  32611=>"101011011",
  32612=>"111110100",
  32613=>"110101011",
  32614=>"101000100",
  32615=>"111000000",
  32616=>"111000011",
  32617=>"100010001",
  32618=>"000011000",
  32619=>"100101000",
  32620=>"000100000",
  32621=>"001011011",
  32622=>"011111111",
  32623=>"110100101",
  32624=>"011110011",
  32625=>"110000000",
  32626=>"011111010",
  32627=>"101011000",
  32628=>"001001101",
  32629=>"110010101",
  32630=>"110001110",
  32631=>"001010010",
  32632=>"011100010",
  32633=>"010001000",
  32634=>"011101011",
  32635=>"010010111",
  32636=>"110111111",
  32637=>"100001010",
  32638=>"111001111",
  32639=>"000110010",
  32640=>"111111110",
  32641=>"111101100",
  32642=>"111000100",
  32643=>"100101010",
  32644=>"001010011",
  32645=>"001011001",
  32646=>"010100110",
  32647=>"011010001",
  32648=>"101111111",
  32649=>"011101100",
  32650=>"011001010",
  32651=>"111010100",
  32652=>"100101001",
  32653=>"100110101",
  32654=>"010100001",
  32655=>"001100111",
  32656=>"100100001",
  32657=>"111000111",
  32658=>"100110100",
  32659=>"100001101",
  32660=>"101011001",
  32661=>"011001000",
  32662=>"111111010",
  32663=>"100101101",
  32664=>"011000101",
  32665=>"110001111",
  32666=>"110101110",
  32667=>"010100001",
  32668=>"001111101",
  32669=>"011111100",
  32670=>"100111011",
  32671=>"010100110",
  32672=>"000000111",
  32673=>"110001011",
  32674=>"010100100",
  32675=>"010001101",
  32676=>"101100101",
  32677=>"100100101",
  32678=>"101001100",
  32679=>"100101111",
  32680=>"101000111",
  32681=>"111001000",
  32682=>"111011100",
  32683=>"011010001",
  32684=>"010100110",
  32685=>"010111111",
  32686=>"100111010",
  32687=>"111100001",
  32688=>"100110101",
  32689=>"101111011",
  32690=>"000110001",
  32691=>"100110001",
  32692=>"000010101",
  32693=>"111010111",
  32694=>"011110101",
  32695=>"100100000",
  32696=>"100011011",
  32697=>"011010001",
  32698=>"000100111",
  32699=>"110100000",
  32700=>"011101001",
  32701=>"100100100",
  32702=>"010010010",
  32703=>"101101111",
  32704=>"011000011",
  32705=>"111100100",
  32706=>"010000001",
  32707=>"011111111",
  32708=>"101001011",
  32709=>"110001111",
  32710=>"110111011",
  32711=>"001101110",
  32712=>"110010010",
  32713=>"001011000",
  32714=>"111110011",
  32715=>"000000110",
  32716=>"101001101",
  32717=>"110101000",
  32718=>"001010111",
  32719=>"110101100",
  32720=>"100000011",
  32721=>"010100000",
  32722=>"110011110",
  32723=>"001010101",
  32724=>"110110000",
  32725=>"001000010",
  32726=>"001110001",
  32727=>"100101110",
  32728=>"100001001",
  32729=>"100001010",
  32730=>"101011001",
  32731=>"101111100",
  32732=>"101101010",
  32733=>"100110011",
  32734=>"000010100",
  32735=>"100100010",
  32736=>"010010001",
  32737=>"011000000",
  32738=>"110101011",
  32739=>"001101110",
  32740=>"001010011",
  32741=>"000001101",
  32742=>"101110000",
  32743=>"110110001",
  32744=>"100010111",
  32745=>"010001000",
  32746=>"010100100",
  32747=>"111111100",
  32748=>"100101010",
  32749=>"111010001",
  32750=>"100000111",
  32751=>"000000001",
  32752=>"000110100",
  32753=>"111110010",
  32754=>"001000010",
  32755=>"110001110",
  32756=>"101000111",
  32757=>"010000000",
  32758=>"010100011",
  32759=>"100001111",
  32760=>"000100011",
  32761=>"010100110",
  32762=>"010001100",
  32763=>"001100000",
  32764=>"111111111",
  32765=>"100000010",
  32766=>"001010011",
  32767=>"010010010",
  32768=>"011101011",
  32769=>"100111111",
  32770=>"110100111",
  32771=>"011010111",
  32772=>"101011000",
  32773=>"000000110",
  32774=>"101101001",
  32775=>"101111001",
  32776=>"111000100",
  32777=>"111110100",
  32778=>"111100010",
  32779=>"010111101",
  32780=>"111101111",
  32781=>"100001010",
  32782=>"011011000",
  32783=>"100010110",
  32784=>"100001001",
  32785=>"101100110",
  32786=>"011111000",
  32787=>"010000101",
  32788=>"000000100",
  32789=>"011001010",
  32790=>"101001011",
  32791=>"100011001",
  32792=>"001000011",
  32793=>"010111011",
  32794=>"101110000",
  32795=>"100111000",
  32796=>"111011101",
  32797=>"010111110",
  32798=>"111110001",
  32799=>"111101110",
  32800=>"111111100",
  32801=>"001011111",
  32802=>"001100100",
  32803=>"111110101",
  32804=>"000110110",
  32805=>"110010100",
  32806=>"100010010",
  32807=>"100010001",
  32808=>"110101100",
  32809=>"001101001",
  32810=>"110111110",
  32811=>"110000101",
  32812=>"110000110",
  32813=>"101111101",
  32814=>"010010000",
  32815=>"001001001",
  32816=>"111111000",
  32817=>"010000111",
  32818=>"111000000",
  32819=>"110100010",
  32820=>"000010001",
  32821=>"011000011",
  32822=>"010100100",
  32823=>"000000111",
  32824=>"100011010",
  32825=>"111101110",
  32826=>"010011101",
  32827=>"110111101",
  32828=>"000111000",
  32829=>"101100110",
  32830=>"101010100",
  32831=>"100111010",
  32832=>"100101110",
  32833=>"011101011",
  32834=>"000000101",
  32835=>"001101000",
  32836=>"011001010",
  32837=>"111101010",
  32838=>"100010000",
  32839=>"010010000",
  32840=>"111101011",
  32841=>"111100111",
  32842=>"010001101",
  32843=>"100001000",
  32844=>"110100001",
  32845=>"010010000",
  32846=>"011011010",
  32847=>"010001001",
  32848=>"001110011",
  32849=>"101000110",
  32850=>"100100011",
  32851=>"001100100",
  32852=>"110000001",
  32853=>"100110000",
  32854=>"010010011",
  32855=>"001110101",
  32856=>"111101110",
  32857=>"100000000",
  32858=>"111101111",
  32859=>"101000010",
  32860=>"000110101",
  32861=>"010111001",
  32862=>"111010010",
  32863=>"100101110",
  32864=>"000111001",
  32865=>"101100001",
  32866=>"011100100",
  32867=>"000101001",
  32868=>"101000100",
  32869=>"011011011",
  32870=>"000010111",
  32871=>"111110010",
  32872=>"110101111",
  32873=>"010011000",
  32874=>"000011100",
  32875=>"110000001",
  32876=>"010001101",
  32877=>"011010111",
  32878=>"001100000",
  32879=>"010110000",
  32880=>"111111010",
  32881=>"011000001",
  32882=>"000111011",
  32883=>"111011100",
  32884=>"001111000",
  32885=>"000101100",
  32886=>"110101101",
  32887=>"001110110",
  32888=>"000111101",
  32889=>"010101110",
  32890=>"110011100",
  32891=>"000111111",
  32892=>"010011001",
  32893=>"101010110",
  32894=>"000110000",
  32895=>"111101100",
  32896=>"011001111",
  32897=>"000011111",
  32898=>"011011000",
  32899=>"111000100",
  32900=>"111000100",
  32901=>"111001000",
  32902=>"000001100",
  32903=>"000110100",
  32904=>"110100110",
  32905=>"100101010",
  32906=>"010010010",
  32907=>"100100011",
  32908=>"010111001",
  32909=>"110010000",
  32910=>"111101001",
  32911=>"101111011",
  32912=>"101111011",
  32913=>"111111001",
  32914=>"010111100",
  32915=>"010111100",
  32916=>"111001010",
  32917=>"101100100",
  32918=>"111001001",
  32919=>"110001010",
  32920=>"110010100",
  32921=>"000100100",
  32922=>"000100101",
  32923=>"100100101",
  32924=>"100000111",
  32925=>"100101000",
  32926=>"010001001",
  32927=>"011011000",
  32928=>"100110111",
  32929=>"011001101",
  32930=>"011001011",
  32931=>"011000000",
  32932=>"111100010",
  32933=>"101100110",
  32934=>"110011000",
  32935=>"000000100",
  32936=>"001100001",
  32937=>"101010001",
  32938=>"101010001",
  32939=>"101000011",
  32940=>"001011111",
  32941=>"111110111",
  32942=>"001011100",
  32943=>"000100111",
  32944=>"100000000",
  32945=>"000100110",
  32946=>"110111111",
  32947=>"000101010",
  32948=>"000000001",
  32949=>"100011101",
  32950=>"000101010",
  32951=>"000010001",
  32952=>"010010001",
  32953=>"010010010",
  32954=>"000101110",
  32955=>"010100000",
  32956=>"010110000",
  32957=>"010100011",
  32958=>"000110011",
  32959=>"110110110",
  32960=>"111000011",
  32961=>"011000100",
  32962=>"101110000",
  32963=>"001101001",
  32964=>"111011010",
  32965=>"010011001",
  32966=>"000110001",
  32967=>"101111101",
  32968=>"001010101",
  32969=>"100110110",
  32970=>"110001010",
  32971=>"100111000",
  32972=>"000111010",
  32973=>"100101111",
  32974=>"011110011",
  32975=>"101011111",
  32976=>"010101111",
  32977=>"111000010",
  32978=>"001111101",
  32979=>"110000110",
  32980=>"001001011",
  32981=>"110110010",
  32982=>"000100001",
  32983=>"000010001",
  32984=>"100110110",
  32985=>"011110000",
  32986=>"111010101",
  32987=>"111000111",
  32988=>"111100111",
  32989=>"110010010",
  32990=>"001100110",
  32991=>"010100100",
  32992=>"111011000",
  32993=>"000111010",
  32994=>"000111000",
  32995=>"010000010",
  32996=>"000111100",
  32997=>"101110001",
  32998=>"000001000",
  32999=>"100111110",
  33000=>"010101000",
  33001=>"100011000",
  33002=>"000111000",
  33003=>"101111111",
  33004=>"000010110",
  33005=>"100100000",
  33006=>"100110101",
  33007=>"001000001",
  33008=>"111111100",
  33009=>"111101101",
  33010=>"110101100",
  33011=>"110000001",
  33012=>"011000011",
  33013=>"111000001",
  33014=>"011000011",
  33015=>"111010001",
  33016=>"100000011",
  33017=>"100000000",
  33018=>"010001111",
  33019=>"010010101",
  33020=>"000011001",
  33021=>"100010001",
  33022=>"010100110",
  33023=>"010110000",
  33024=>"110101100",
  33025=>"000100001",
  33026=>"010001111",
  33027=>"101110000",
  33028=>"101001100",
  33029=>"000000100",
  33030=>"000001001",
  33031=>"111001110",
  33032=>"101101000",
  33033=>"110010111",
  33034=>"111111100",
  33035=>"101111010",
  33036=>"000010100",
  33037=>"101110010",
  33038=>"100111110",
  33039=>"000100010",
  33040=>"001101010",
  33041=>"110110011",
  33042=>"100011011",
  33043=>"101111100",
  33044=>"001111111",
  33045=>"100111001",
  33046=>"000010100",
  33047=>"110001011",
  33048=>"100000101",
  33049=>"101001111",
  33050=>"010010110",
  33051=>"011110001",
  33052=>"100010101",
  33053=>"111100010",
  33054=>"001001010",
  33055=>"000010110",
  33056=>"000010110",
  33057=>"011111011",
  33058=>"001011110",
  33059=>"010010000",
  33060=>"111101010",
  33061=>"100111010",
  33062=>"110011011",
  33063=>"101011000",
  33064=>"100010001",
  33065=>"011000011",
  33066=>"011110111",
  33067=>"011110111",
  33068=>"000010010",
  33069=>"110010010",
  33070=>"011100100",
  33071=>"101110011",
  33072=>"010100110",
  33073=>"110011010",
  33074=>"100101110",
  33075=>"111001110",
  33076=>"101110100",
  33077=>"100101011",
  33078=>"111101101",
  33079=>"111101101",
  33080=>"001000101",
  33081=>"101000001",
  33082=>"111111100",
  33083=>"110001011",
  33084=>"111000110",
  33085=>"011100111",
  33086=>"110000010",
  33087=>"110001001",
  33088=>"110001110",
  33089=>"010100000",
  33090=>"011100000",
  33091=>"011111011",
  33092=>"011110101",
  33093=>"100011101",
  33094=>"010110000",
  33095=>"101000011",
  33096=>"110001100",
  33097=>"110001110",
  33098=>"001000011",
  33099=>"111000110",
  33100=>"101110001",
  33101=>"100001010",
  33102=>"010001110",
  33103=>"000010110",
  33104=>"110010011",
  33105=>"000110110",
  33106=>"110111101",
  33107=>"100111011",
  33108=>"101001110",
  33109=>"101101100",
  33110=>"000101100",
  33111=>"101011100",
  33112=>"111100101",
  33113=>"101001000",
  33114=>"100001111",
  33115=>"101100111",
  33116=>"000100000",
  33117=>"011010110",
  33118=>"011110100",
  33119=>"000111101",
  33120=>"110010001",
  33121=>"011110011",
  33122=>"101001100",
  33123=>"010010001",
  33124=>"011001101",
  33125=>"000000111",
  33126=>"010010111",
  33127=>"000000010",
  33128=>"010100011",
  33129=>"100100001",
  33130=>"101111001",
  33131=>"000111000",
  33132=>"011101000",
  33133=>"111111010",
  33134=>"000011110",
  33135=>"111110000",
  33136=>"000010101",
  33137=>"110110001",
  33138=>"100010111",
  33139=>"100001001",
  33140=>"101110101",
  33141=>"101100001",
  33142=>"011001000",
  33143=>"010101010",
  33144=>"110011101",
  33145=>"111011001",
  33146=>"011010101",
  33147=>"011100011",
  33148=>"111000010",
  33149=>"111111011",
  33150=>"011000111",
  33151=>"110111000",
  33152=>"111001110",
  33153=>"100011110",
  33154=>"001101111",
  33155=>"100101111",
  33156=>"001101110",
  33157=>"100111100",
  33158=>"100111111",
  33159=>"010100111",
  33160=>"010101100",
  33161=>"101101111",
  33162=>"011111011",
  33163=>"000000001",
  33164=>"100110101",
  33165=>"011110111",
  33166=>"100100111",
  33167=>"001110111",
  33168=>"011101111",
  33169=>"101101110",
  33170=>"011110100",
  33171=>"101100101",
  33172=>"010010101",
  33173=>"010100001",
  33174=>"110010001",
  33175=>"111000101",
  33176=>"000101010",
  33177=>"010000111",
  33178=>"100010111",
  33179=>"011111000",
  33180=>"101111010",
  33181=>"011111000",
  33182=>"011111111",
  33183=>"111010111",
  33184=>"110111111",
  33185=>"110001101",
  33186=>"111011110",
  33187=>"110110010",
  33188=>"000001000",
  33189=>"010100111",
  33190=>"001100001",
  33191=>"000111111",
  33192=>"111111010",
  33193=>"101110011",
  33194=>"000000111",
  33195=>"000000111",
  33196=>"101110101",
  33197=>"010100100",
  33198=>"111000000",
  33199=>"000010010",
  33200=>"011010110",
  33201=>"111101100",
  33202=>"110101101",
  33203=>"011110000",
  33204=>"111010111",
  33205=>"100111001",
  33206=>"100111100",
  33207=>"000000001",
  33208=>"100001010",
  33209=>"100001110",
  33210=>"011010111",
  33211=>"011000110",
  33212=>"010010001",
  33213=>"011100010",
  33214=>"110000100",
  33215=>"110001111",
  33216=>"110010011",
  33217=>"110100000",
  33218=>"001101111",
  33219=>"010110000",
  33220=>"000000101",
  33221=>"000000011",
  33222=>"000011100",
  33223=>"111100010",
  33224=>"101111001",
  33225=>"101010001",
  33226=>"010100000",
  33227=>"110011101",
  33228=>"001010000",
  33229=>"010011010",
  33230=>"111000001",
  33231=>"000111110",
  33232=>"110001001",
  33233=>"001111000",
  33234=>"111011010",
  33235=>"111101001",
  33236=>"110010000",
  33237=>"011000101",
  33238=>"100111111",
  33239=>"110001011",
  33240=>"110011100",
  33241=>"101010101",
  33242=>"000010101",
  33243=>"110010110",
  33244=>"100110100",
  33245=>"011110001",
  33246=>"000101000",
  33247=>"001010111",
  33248=>"111111110",
  33249=>"101110100",
  33250=>"010111110",
  33251=>"101010011",
  33252=>"101001010",
  33253=>"001000101",
  33254=>"010101110",
  33255=>"010111011",
  33256=>"010011000",
  33257=>"010111000",
  33258=>"001001000",
  33259=>"110000111",
  33260=>"110111100",
  33261=>"101100100",
  33262=>"110100000",
  33263=>"001011000",
  33264=>"101000110",
  33265=>"010010010",
  33266=>"111110110",
  33267=>"011111010",
  33268=>"111101000",
  33269=>"001010010",
  33270=>"111101010",
  33271=>"000010000",
  33272=>"000011001",
  33273=>"111110110",
  33274=>"110010000",
  33275=>"111110101",
  33276=>"000001111",
  33277=>"011101100",
  33278=>"011010101",
  33279=>"101111111",
  33280=>"011100111",
  33281=>"001110110",
  33282=>"111111100",
  33283=>"110000010",
  33284=>"000101110",
  33285=>"101000111",
  33286=>"100011110",
  33287=>"111001000",
  33288=>"011000000",
  33289=>"100111110",
  33290=>"101101110",
  33291=>"000011010",
  33292=>"000101110",
  33293=>"100101111",
  33294=>"101100110",
  33295=>"110101000",
  33296=>"101010000",
  33297=>"111000001",
  33298=>"000110011",
  33299=>"011001100",
  33300=>"011000010",
  33301=>"011101000",
  33302=>"001101010",
  33303=>"101000010",
  33304=>"000000100",
  33305=>"100011001",
  33306=>"000101000",
  33307=>"110000001",
  33308=>"001110010",
  33309=>"111111000",
  33310=>"110101110",
  33311=>"011101011",
  33312=>"111000100",
  33313=>"100110011",
  33314=>"010011111",
  33315=>"101010101",
  33316=>"000010110",
  33317=>"010111101",
  33318=>"110010001",
  33319=>"001101111",
  33320=>"010011001",
  33321=>"011001111",
  33322=>"111101010",
  33323=>"110011101",
  33324=>"011001000",
  33325=>"010010011",
  33326=>"101000001",
  33327=>"101001001",
  33328=>"010111111",
  33329=>"011111111",
  33330=>"010110101",
  33331=>"110000011",
  33332=>"010011100",
  33333=>"000010111",
  33334=>"100101000",
  33335=>"010111001",
  33336=>"010101100",
  33337=>"110110000",
  33338=>"001010010",
  33339=>"010010000",
  33340=>"101001101",
  33341=>"010011110",
  33342=>"001101111",
  33343=>"010110001",
  33344=>"010111100",
  33345=>"001001010",
  33346=>"111011001",
  33347=>"110110111",
  33348=>"001001011",
  33349=>"011010000",
  33350=>"100100100",
  33351=>"011101000",
  33352=>"110110100",
  33353=>"100111111",
  33354=>"110111010",
  33355=>"111110111",
  33356=>"101110110",
  33357=>"101110110",
  33358=>"011001101",
  33359=>"000100110",
  33360=>"111101111",
  33361=>"000110001",
  33362=>"101001011",
  33363=>"100010010",
  33364=>"000110000",
  33365=>"010100100",
  33366=>"100010100",
  33367=>"100000000",
  33368=>"101110000",
  33369=>"011110010",
  33370=>"110101101",
  33371=>"010101100",
  33372=>"001111010",
  33373=>"110101100",
  33374=>"000001110",
  33375=>"010010010",
  33376=>"101010001",
  33377=>"001001110",
  33378=>"100110110",
  33379=>"001011001",
  33380=>"110000010",
  33381=>"110001101",
  33382=>"101111101",
  33383=>"100001010",
  33384=>"000111110",
  33385=>"001000001",
  33386=>"110101001",
  33387=>"100000011",
  33388=>"101010110",
  33389=>"010110010",
  33390=>"111110010",
  33391=>"011010110",
  33392=>"010111111",
  33393=>"011010000",
  33394=>"011011001",
  33395=>"101100010",
  33396=>"011111000",
  33397=>"101000100",
  33398=>"110000100",
  33399=>"000111101",
  33400=>"011011110",
  33401=>"001000101",
  33402=>"001100111",
  33403=>"101000011",
  33404=>"010011001",
  33405=>"110001010",
  33406=>"011110100",
  33407=>"100001111",
  33408=>"111001001",
  33409=>"000010101",
  33410=>"011110101",
  33411=>"010100101",
  33412=>"000011111",
  33413=>"110110101",
  33414=>"111101101",
  33415=>"010101100",
  33416=>"000010011",
  33417=>"000000110",
  33418=>"111111111",
  33419=>"000100000",
  33420=>"010001100",
  33421=>"000111101",
  33422=>"010001000",
  33423=>"100010010",
  33424=>"111101101",
  33425=>"111001110",
  33426=>"101111010",
  33427=>"001111001",
  33428=>"000100111",
  33429=>"110100010",
  33430=>"111001111",
  33431=>"100101101",
  33432=>"011100100",
  33433=>"100101100",
  33434=>"110000111",
  33435=>"011011100",
  33436=>"100001011",
  33437=>"110010000",
  33438=>"010010011",
  33439=>"010010110",
  33440=>"110110111",
  33441=>"101010100",
  33442=>"110101110",
  33443=>"111111000",
  33444=>"010110101",
  33445=>"111000001",
  33446=>"011110001",
  33447=>"000011011",
  33448=>"011011011",
  33449=>"111101001",
  33450=>"110110101",
  33451=>"111000011",
  33452=>"010110100",
  33453=>"011001111",
  33454=>"001010000",
  33455=>"100111001",
  33456=>"001100100",
  33457=>"000010100",
  33458=>"010111100",
  33459=>"101011000",
  33460=>"001111110",
  33461=>"011010000",
  33462=>"100100110",
  33463=>"101110001",
  33464=>"101110110",
  33465=>"111010000",
  33466=>"100000101",
  33467=>"001111110",
  33468=>"101101000",
  33469=>"111101000",
  33470=>"100100000",
  33471=>"111100101",
  33472=>"011000101",
  33473=>"000100111",
  33474=>"101011111",
  33475=>"000111010",
  33476=>"110101110",
  33477=>"010100001",
  33478=>"101000011",
  33479=>"001000110",
  33480=>"110011010",
  33481=>"001010101",
  33482=>"000111111",
  33483=>"100001000",
  33484=>"000111110",
  33485=>"111111111",
  33486=>"100111001",
  33487=>"011001111",
  33488=>"001110000",
  33489=>"001110000",
  33490=>"100001011",
  33491=>"111101111",
  33492=>"011000011",
  33493=>"001010100",
  33494=>"100101011",
  33495=>"010110100",
  33496=>"100011001",
  33497=>"101100111",
  33498=>"101000110",
  33499=>"010101111",
  33500=>"100010010",
  33501=>"010100010",
  33502=>"100101000",
  33503=>"111110011",
  33504=>"011000010",
  33505=>"001110011",
  33506=>"111111110",
  33507=>"011101001",
  33508=>"101110110",
  33509=>"011111110",
  33510=>"011111111",
  33511=>"011101100",
  33512=>"100000111",
  33513=>"101100101",
  33514=>"000000010",
  33515=>"101001001",
  33516=>"101111011",
  33517=>"011101010",
  33518=>"010111011",
  33519=>"000101010",
  33520=>"011110010",
  33521=>"010110111",
  33522=>"011100010",
  33523=>"110011111",
  33524=>"000000010",
  33525=>"111011001",
  33526=>"001100010",
  33527=>"111111010",
  33528=>"001110011",
  33529=>"110101100",
  33530=>"100000111",
  33531=>"110110100",
  33532=>"010011000",
  33533=>"000111101",
  33534=>"110110011",
  33535=>"110010101",
  33536=>"010010100",
  33537=>"000100011",
  33538=>"001000010",
  33539=>"101000010",
  33540=>"111011000",
  33541=>"111010110",
  33542=>"111101100",
  33543=>"100111010",
  33544=>"001011010",
  33545=>"010101101",
  33546=>"000110110",
  33547=>"100100100",
  33548=>"010101010",
  33549=>"111111111",
  33550=>"010010011",
  33551=>"101111101",
  33552=>"100001001",
  33553=>"101110110",
  33554=>"001110110",
  33555=>"011110011",
  33556=>"010010101",
  33557=>"101100110",
  33558=>"101100001",
  33559=>"011010000",
  33560=>"110100000",
  33561=>"000000011",
  33562=>"010101011",
  33563=>"111110001",
  33564=>"111100110",
  33565=>"001000001",
  33566=>"110010010",
  33567=>"000110100",
  33568=>"000010111",
  33569=>"101011101",
  33570=>"111010100",
  33571=>"100011011",
  33572=>"001011010",
  33573=>"110110000",
  33574=>"101101101",
  33575=>"000011010",
  33576=>"111001101",
  33577=>"000000110",
  33578=>"011001111",
  33579=>"010011000",
  33580=>"111111111",
  33581=>"011111001",
  33582=>"010110101",
  33583=>"111110000",
  33584=>"110110001",
  33585=>"111010100",
  33586=>"010000011",
  33587=>"011110000",
  33588=>"101000001",
  33589=>"110011100",
  33590=>"100010111",
  33591=>"010001000",
  33592=>"001001000",
  33593=>"001010101",
  33594=>"110111100",
  33595=>"000110111",
  33596=>"100000010",
  33597=>"001001001",
  33598=>"011000100",
  33599=>"101110111",
  33600=>"110011110",
  33601=>"100000100",
  33602=>"000001011",
  33603=>"001111000",
  33604=>"110100101",
  33605=>"000111011",
  33606=>"100000000",
  33607=>"110001110",
  33608=>"111010101",
  33609=>"001101000",
  33610=>"001101101",
  33611=>"110011101",
  33612=>"110001101",
  33613=>"101110101",
  33614=>"100011110",
  33615=>"110110100",
  33616=>"000010100",
  33617=>"000000000",
  33618=>"100001011",
  33619=>"111011010",
  33620=>"110100100",
  33621=>"001000000",
  33622=>"000111111",
  33623=>"001011010",
  33624=>"111111100",
  33625=>"010101100",
  33626=>"110101000",
  33627=>"110101011",
  33628=>"110011100",
  33629=>"000111011",
  33630=>"100011101",
  33631=>"001000001",
  33632=>"010000010",
  33633=>"111101000",
  33634=>"111101000",
  33635=>"000010010",
  33636=>"000001010",
  33637=>"000110000",
  33638=>"001010111",
  33639=>"101011001",
  33640=>"101101000",
  33641=>"111111101",
  33642=>"111110010",
  33643=>"101111010",
  33644=>"101010011",
  33645=>"001001010",
  33646=>"000100110",
  33647=>"000110000",
  33648=>"000011011",
  33649=>"001000000",
  33650=>"110000010",
  33651=>"101011001",
  33652=>"000011110",
  33653=>"100000011",
  33654=>"111111111",
  33655=>"110111110",
  33656=>"110111110",
  33657=>"001110101",
  33658=>"000001101",
  33659=>"011100110",
  33660=>"000100101",
  33661=>"110100110",
  33662=>"101110000",
  33663=>"001010011",
  33664=>"100101010",
  33665=>"110100111",
  33666=>"101011000",
  33667=>"110011011",
  33668=>"111010011",
  33669=>"111001010",
  33670=>"011100001",
  33671=>"110101111",
  33672=>"011101010",
  33673=>"110110010",
  33674=>"011010011",
  33675=>"100000110",
  33676=>"111011011",
  33677=>"010101100",
  33678=>"001100110",
  33679=>"000001100",
  33680=>"100010010",
  33681=>"000101100",
  33682=>"100100001",
  33683=>"101010010",
  33684=>"000001100",
  33685=>"101101111",
  33686=>"010110001",
  33687=>"111011001",
  33688=>"010000000",
  33689=>"110010001",
  33690=>"110010100",
  33691=>"010011101",
  33692=>"101011101",
  33693=>"001111001",
  33694=>"101000110",
  33695=>"111011011",
  33696=>"100000001",
  33697=>"011101110",
  33698=>"110001110",
  33699=>"010111101",
  33700=>"101110111",
  33701=>"111110010",
  33702=>"001110101",
  33703=>"110001000",
  33704=>"101001000",
  33705=>"001010100",
  33706=>"001010011",
  33707=>"111000100",
  33708=>"000001011",
  33709=>"101111101",
  33710=>"101001110",
  33711=>"100011100",
  33712=>"001000100",
  33713=>"110110001",
  33714=>"011111001",
  33715=>"111101000",
  33716=>"100000111",
  33717=>"101111001",
  33718=>"001100001",
  33719=>"010010110",
  33720=>"110011000",
  33721=>"010011100",
  33722=>"011000010",
  33723=>"000101101",
  33724=>"000001100",
  33725=>"111111101",
  33726=>"101001001",
  33727=>"000100111",
  33728=>"111100110",
  33729=>"000100000",
  33730=>"100000011",
  33731=>"111110110",
  33732=>"000111101",
  33733=>"011000011",
  33734=>"110101101",
  33735=>"101101110",
  33736=>"001100101",
  33737=>"100110010",
  33738=>"000111010",
  33739=>"011110011",
  33740=>"100001101",
  33741=>"100001111",
  33742=>"100101111",
  33743=>"001111000",
  33744=>"100010100",
  33745=>"011101000",
  33746=>"010100000",
  33747=>"000000010",
  33748=>"101011100",
  33749=>"111111101",
  33750=>"011010100",
  33751=>"110100100",
  33752=>"001010111",
  33753=>"110001101",
  33754=>"100001000",
  33755=>"100101111",
  33756=>"101110100",
  33757=>"111100101",
  33758=>"110111011",
  33759=>"000111011",
  33760=>"101001010",
  33761=>"001000111",
  33762=>"011111011",
  33763=>"000010001",
  33764=>"000100010",
  33765=>"100110010",
  33766=>"111011011",
  33767=>"111010001",
  33768=>"111010100",
  33769=>"010011011",
  33770=>"001111100",
  33771=>"101101011",
  33772=>"000101110",
  33773=>"111101001",
  33774=>"111010000",
  33775=>"100010101",
  33776=>"000100010",
  33777=>"010010001",
  33778=>"001100111",
  33779=>"000100010",
  33780=>"100111111",
  33781=>"010000011",
  33782=>"010010000",
  33783=>"110000001",
  33784=>"000011001",
  33785=>"001010011",
  33786=>"000111110",
  33787=>"000101101",
  33788=>"101110111",
  33789=>"101111101",
  33790=>"101001010",
  33791=>"010111011",
  33792=>"100000010",
  33793=>"110101101",
  33794=>"111111111",
  33795=>"100010101",
  33796=>"000000111",
  33797=>"000001011",
  33798=>"110001110",
  33799=>"000101011",
  33800=>"001100110",
  33801=>"110001111",
  33802=>"000101000",
  33803=>"101111100",
  33804=>"100001000",
  33805=>"010111010",
  33806=>"010011110",
  33807=>"001000010",
  33808=>"111000000",
  33809=>"111111011",
  33810=>"100001001",
  33811=>"100000100",
  33812=>"001010001",
  33813=>"110110000",
  33814=>"110101001",
  33815=>"101000111",
  33816=>"110111000",
  33817=>"000000100",
  33818=>"111000001",
  33819=>"000001110",
  33820=>"111000101",
  33821=>"101011001",
  33822=>"010100101",
  33823=>"100011011",
  33824=>"011000000",
  33825=>"101010000",
  33826=>"100110000",
  33827=>"101010010",
  33828=>"001010000",
  33829=>"011110100",
  33830=>"000010000",
  33831=>"001101111",
  33832=>"011000000",
  33833=>"001001111",
  33834=>"111100110",
  33835=>"100010001",
  33836=>"101001010",
  33837=>"100000000",
  33838=>"011110100",
  33839=>"011101010",
  33840=>"001010110",
  33841=>"101100100",
  33842=>"010001100",
  33843=>"111110101",
  33844=>"110010011",
  33845=>"101111011",
  33846=>"011000000",
  33847=>"010000000",
  33848=>"111111000",
  33849=>"100111100",
  33850=>"010000100",
  33851=>"010000111",
  33852=>"100111001",
  33853=>"101101010",
  33854=>"111010111",
  33855=>"111101111",
  33856=>"100110010",
  33857=>"000011110",
  33858=>"110101111",
  33859=>"011111001",
  33860=>"000100100",
  33861=>"100101010",
  33862=>"100010011",
  33863=>"111010111",
  33864=>"010100100",
  33865=>"100011000",
  33866=>"001000010",
  33867=>"000111001",
  33868=>"001000001",
  33869=>"100011111",
  33870=>"011101100",
  33871=>"001001011",
  33872=>"001000001",
  33873=>"000000101",
  33874=>"111010111",
  33875=>"110101001",
  33876=>"110100000",
  33877=>"100110101",
  33878=>"111011101",
  33879=>"000001010",
  33880=>"011111101",
  33881=>"011011110",
  33882=>"110011100",
  33883=>"001101010",
  33884=>"011101110",
  33885=>"000101001",
  33886=>"010001110",
  33887=>"011101010",
  33888=>"011101111",
  33889=>"010010000",
  33890=>"110100100",
  33891=>"111100100",
  33892=>"010000010",
  33893=>"010110111",
  33894=>"101101101",
  33895=>"010100000",
  33896=>"011001110",
  33897=>"111011110",
  33898=>"110010010",
  33899=>"111100000",
  33900=>"000010101",
  33901=>"110101010",
  33902=>"011001111",
  33903=>"000000010",
  33904=>"110000001",
  33905=>"010011000",
  33906=>"000100001",
  33907=>"000110001",
  33908=>"011011000",
  33909=>"100000010",
  33910=>"110110011",
  33911=>"010101101",
  33912=>"000000100",
  33913=>"010100111",
  33914=>"110101111",
  33915=>"100010001",
  33916=>"001101011",
  33917=>"000110000",
  33918=>"100111100",
  33919=>"100010011",
  33920=>"110000000",
  33921=>"101111101",
  33922=>"001110001",
  33923=>"100000100",
  33924=>"101011011",
  33925=>"111100010",
  33926=>"100111000",
  33927=>"001001111",
  33928=>"010111101",
  33929=>"111101001",
  33930=>"010100000",
  33931=>"100011100",
  33932=>"001000000",
  33933=>"011110101",
  33934=>"010010001",
  33935=>"010101011",
  33936=>"110101011",
  33937=>"110110101",
  33938=>"010001010",
  33939=>"000101000",
  33940=>"101011100",
  33941=>"101111110",
  33942=>"101001000",
  33943=>"001000010",
  33944=>"111111001",
  33945=>"000010011",
  33946=>"011110000",
  33947=>"101110001",
  33948=>"111010001",
  33949=>"101000011",
  33950=>"001111000",
  33951=>"111000010",
  33952=>"001000100",
  33953=>"010000110",
  33954=>"010100011",
  33955=>"010001001",
  33956=>"001110111",
  33957=>"000001110",
  33958=>"001111001",
  33959=>"000010001",
  33960=>"100000101",
  33961=>"100101100",
  33962=>"111110110",
  33963=>"100100100",
  33964=>"001111010",
  33965=>"110000111",
  33966=>"110111101",
  33967=>"100101011",
  33968=>"000100000",
  33969=>"000000011",
  33970=>"000000100",
  33971=>"100010100",
  33972=>"111000000",
  33973=>"011000000",
  33974=>"000111011",
  33975=>"111010110",
  33976=>"100010111",
  33977=>"010100000",
  33978=>"100110000",
  33979=>"010111101",
  33980=>"010001010",
  33981=>"110110110",
  33982=>"010110000",
  33983=>"100100100",
  33984=>"110000001",
  33985=>"110001111",
  33986=>"101001010",
  33987=>"111010011",
  33988=>"011011111",
  33989=>"011000110",
  33990=>"101011110",
  33991=>"110000001",
  33992=>"101110111",
  33993=>"111111110",
  33994=>"011101000",
  33995=>"001001110",
  33996=>"010000111",
  33997=>"001100011",
  33998=>"011101111",
  33999=>"001110010",
  34000=>"010000100",
  34001=>"001101111",
  34002=>"101110001",
  34003=>"011001001",
  34004=>"100000001",
  34005=>"111011000",
  34006=>"001011001",
  34007=>"100110001",
  34008=>"001011100",
  34009=>"111000001",
  34010=>"111010001",
  34011=>"101111101",
  34012=>"011110000",
  34013=>"000011101",
  34014=>"010101101",
  34015=>"111011010",
  34016=>"110001000",
  34017=>"001101100",
  34018=>"110001111",
  34019=>"111110011",
  34020=>"010101010",
  34021=>"010010011",
  34022=>"010000101",
  34023=>"011011001",
  34024=>"111101000",
  34025=>"010011100",
  34026=>"010001101",
  34027=>"000000010",
  34028=>"110101100",
  34029=>"101101001",
  34030=>"100111111",
  34031=>"111110111",
  34032=>"110000000",
  34033=>"101101110",
  34034=>"110000101",
  34035=>"110010100",
  34036=>"100001011",
  34037=>"111000000",
  34038=>"111011100",
  34039=>"110010101",
  34040=>"000000110",
  34041=>"001111010",
  34042=>"011000100",
  34043=>"010101000",
  34044=>"001111101",
  34045=>"011000001",
  34046=>"100101000",
  34047=>"001010011",
  34048=>"100110001",
  34049=>"101011010",
  34050=>"001000000",
  34051=>"100001110",
  34052=>"000011001",
  34053=>"001000001",
  34054=>"111010001",
  34055=>"101111001",
  34056=>"101110001",
  34057=>"111000010",
  34058=>"111000101",
  34059=>"100001010",
  34060=>"111011000",
  34061=>"001100000",
  34062=>"111001111",
  34063=>"001001110",
  34064=>"010101001",
  34065=>"111000100",
  34066=>"100010011",
  34067=>"110000011",
  34068=>"001011110",
  34069=>"111001011",
  34070=>"010010111",
  34071=>"001011010",
  34072=>"100101000",
  34073=>"001111010",
  34074=>"010111000",
  34075=>"101010010",
  34076=>"010000110",
  34077=>"110101011",
  34078=>"111111000",
  34079=>"010010100",
  34080=>"001000001",
  34081=>"000110111",
  34082=>"010000000",
  34083=>"000000101",
  34084=>"010000100",
  34085=>"111001101",
  34086=>"101001011",
  34087=>"110000001",
  34088=>"111010001",
  34089=>"111000011",
  34090=>"101010101",
  34091=>"011111110",
  34092=>"110110110",
  34093=>"001000101",
  34094=>"001100101",
  34095=>"011111010",
  34096=>"001000000",
  34097=>"101110001",
  34098=>"110101001",
  34099=>"100101001",
  34100=>"110001101",
  34101=>"010100100",
  34102=>"101111010",
  34103=>"100101001",
  34104=>"100100101",
  34105=>"110011001",
  34106=>"010001100",
  34107=>"111001100",
  34108=>"100000101",
  34109=>"110011100",
  34110=>"011101011",
  34111=>"011101111",
  34112=>"010001010",
  34113=>"111110001",
  34114=>"011000111",
  34115=>"111110101",
  34116=>"111110111",
  34117=>"000111110",
  34118=>"010011101",
  34119=>"101110010",
  34120=>"000000001",
  34121=>"001001000",
  34122=>"010111110",
  34123=>"100000011",
  34124=>"110100000",
  34125=>"111011001",
  34126=>"000100101",
  34127=>"011100100",
  34128=>"101000001",
  34129=>"110100111",
  34130=>"010011110",
  34131=>"010001011",
  34132=>"010010100",
  34133=>"011100100",
  34134=>"111010001",
  34135=>"011011110",
  34136=>"111111011",
  34137=>"111100010",
  34138=>"001001100",
  34139=>"010111001",
  34140=>"100010011",
  34141=>"110000011",
  34142=>"110010011",
  34143=>"001111001",
  34144=>"010100001",
  34145=>"011011011",
  34146=>"011111011",
  34147=>"010111010",
  34148=>"111100001",
  34149=>"011110100",
  34150=>"001000000",
  34151=>"010000010",
  34152=>"011010111",
  34153=>"001010011",
  34154=>"101000010",
  34155=>"110101101",
  34156=>"100001001",
  34157=>"110001100",
  34158=>"011001100",
  34159=>"011011100",
  34160=>"011100001",
  34161=>"100001010",
  34162=>"100110100",
  34163=>"111100000",
  34164=>"001110110",
  34165=>"110111111",
  34166=>"101110101",
  34167=>"101010011",
  34168=>"000100101",
  34169=>"110000101",
  34170=>"011110111",
  34171=>"100101011",
  34172=>"000101111",
  34173=>"000111001",
  34174=>"101000011",
  34175=>"000101101",
  34176=>"100001111",
  34177=>"100010101",
  34178=>"001111000",
  34179=>"100100001",
  34180=>"101110111",
  34181=>"010011010",
  34182=>"101100010",
  34183=>"111011101",
  34184=>"111110000",
  34185=>"110100010",
  34186=>"011001110",
  34187=>"000010000",
  34188=>"110100111",
  34189=>"000100000",
  34190=>"100001101",
  34191=>"010101111",
  34192=>"111001111",
  34193=>"101101100",
  34194=>"110101101",
  34195=>"011001111",
  34196=>"101001111",
  34197=>"110111100",
  34198=>"010000001",
  34199=>"100100011",
  34200=>"011100111",
  34201=>"110001001",
  34202=>"110010000",
  34203=>"000111001",
  34204=>"100101111",
  34205=>"010001010",
  34206=>"101011000",
  34207=>"111010101",
  34208=>"100100010",
  34209=>"100011110",
  34210=>"101001000",
  34211=>"101101010",
  34212=>"001100000",
  34213=>"001000110",
  34214=>"111110000",
  34215=>"000010000",
  34216=>"111110100",
  34217=>"101011110",
  34218=>"001000011",
  34219=>"000000011",
  34220=>"011000001",
  34221=>"100001110",
  34222=>"110111111",
  34223=>"100101110",
  34224=>"111110001",
  34225=>"111110111",
  34226=>"011101000",
  34227=>"111011001",
  34228=>"101111011",
  34229=>"110111110",
  34230=>"010110000",
  34231=>"000111001",
  34232=>"011110100",
  34233=>"011101000",
  34234=>"010011110",
  34235=>"101101010",
  34236=>"011001010",
  34237=>"110001011",
  34238=>"010001001",
  34239=>"001000011",
  34240=>"000010000",
  34241=>"010011110",
  34242=>"000001010",
  34243=>"100000100",
  34244=>"110001100",
  34245=>"100111011",
  34246=>"101111110",
  34247=>"101001010",
  34248=>"001011110",
  34249=>"110100101",
  34250=>"110111010",
  34251=>"001000111",
  34252=>"001000011",
  34253=>"100010111",
  34254=>"001000000",
  34255=>"000000110",
  34256=>"000011011",
  34257=>"000011101",
  34258=>"100110100",
  34259=>"010111000",
  34260=>"000101001",
  34261=>"100101111",
  34262=>"101000001",
  34263=>"111011110",
  34264=>"101001110",
  34265=>"001100101",
  34266=>"010111100",
  34267=>"010100110",
  34268=>"100101101",
  34269=>"100000100",
  34270=>"010100110",
  34271=>"001100001",
  34272=>"101101010",
  34273=>"001000110",
  34274=>"111100101",
  34275=>"101100010",
  34276=>"111001110",
  34277=>"001011011",
  34278=>"110010110",
  34279=>"100100101",
  34280=>"100100111",
  34281=>"011000001",
  34282=>"110011101",
  34283=>"100010000",
  34284=>"110111010",
  34285=>"001110011",
  34286=>"000000011",
  34287=>"001111000",
  34288=>"110010111",
  34289=>"001001101",
  34290=>"100100100",
  34291=>"001000001",
  34292=>"000000111",
  34293=>"101111111",
  34294=>"001101011",
  34295=>"011101000",
  34296=>"101011011",
  34297=>"010100011",
  34298=>"000001001",
  34299=>"110100101",
  34300=>"001111011",
  34301=>"111011110",
  34302=>"101110100",
  34303=>"011100111",
  34304=>"000010010",
  34305=>"101010101",
  34306=>"101001001",
  34307=>"010101001",
  34308=>"000100111",
  34309=>"100100000",
  34310=>"111010100",
  34311=>"111111100",
  34312=>"000101001",
  34313=>"000101100",
  34314=>"101000100",
  34315=>"001001100",
  34316=>"110000101",
  34317=>"110000111",
  34318=>"001000011",
  34319=>"011000010",
  34320=>"100111100",
  34321=>"101011110",
  34322=>"110011000",
  34323=>"001101011",
  34324=>"000110001",
  34325=>"010110100",
  34326=>"100100001",
  34327=>"011011001",
  34328=>"111011111",
  34329=>"110101000",
  34330=>"001011111",
  34331=>"101101011",
  34332=>"010001100",
  34333=>"100101100",
  34334=>"100000011",
  34335=>"100000011",
  34336=>"010001011",
  34337=>"110011011",
  34338=>"000100001",
  34339=>"011100010",
  34340=>"111011000",
  34341=>"101010100",
  34342=>"111111011",
  34343=>"000010000",
  34344=>"100100101",
  34345=>"011010100",
  34346=>"110010001",
  34347=>"100100101",
  34348=>"001001110",
  34349=>"001010000",
  34350=>"110001100",
  34351=>"110000011",
  34352=>"100001111",
  34353=>"011001111",
  34354=>"001011100",
  34355=>"001111110",
  34356=>"010001110",
  34357=>"111010001",
  34358=>"100100111",
  34359=>"111101101",
  34360=>"111010111",
  34361=>"110110110",
  34362=>"000010111",
  34363=>"101100000",
  34364=>"000001001",
  34365=>"010110001",
  34366=>"010111100",
  34367=>"010001001",
  34368=>"011101011",
  34369=>"100100100",
  34370=>"111100001",
  34371=>"001010101",
  34372=>"000010001",
  34373=>"101101011",
  34374=>"000000111",
  34375=>"000111001",
  34376=>"001010010",
  34377=>"010010011",
  34378=>"101010101",
  34379=>"001000000",
  34380=>"011101100",
  34381=>"001010111",
  34382=>"100011001",
  34383=>"101100101",
  34384=>"011100000",
  34385=>"111110000",
  34386=>"100100011",
  34387=>"111111101",
  34388=>"111011101",
  34389=>"001000001",
  34390=>"111010101",
  34391=>"010110111",
  34392=>"110011000",
  34393=>"000010101",
  34394=>"010100010",
  34395=>"000000000",
  34396=>"000010000",
  34397=>"100100000",
  34398=>"010011100",
  34399=>"111111111",
  34400=>"000100011",
  34401=>"111000010",
  34402=>"000101010",
  34403=>"010001001",
  34404=>"111011011",
  34405=>"000001101",
  34406=>"101001100",
  34407=>"010010011",
  34408=>"100110101",
  34409=>"101100101",
  34410=>"000111100",
  34411=>"100000110",
  34412=>"011101101",
  34413=>"010100111",
  34414=>"111000111",
  34415=>"010111111",
  34416=>"111111111",
  34417=>"011100111",
  34418=>"010101100",
  34419=>"100011001",
  34420=>"100101001",
  34421=>"001100011",
  34422=>"010110001",
  34423=>"100010000",
  34424=>"111111011",
  34425=>"101101100",
  34426=>"000000000",
  34427=>"011100101",
  34428=>"010000101",
  34429=>"100001101",
  34430=>"010100101",
  34431=>"011110101",
  34432=>"001011110",
  34433=>"111110011",
  34434=>"000110000",
  34435=>"110000001",
  34436=>"101100000",
  34437=>"100010100",
  34438=>"110100110",
  34439=>"010111110",
  34440=>"110011010",
  34441=>"100011110",
  34442=>"111110000",
  34443=>"101101000",
  34444=>"111101011",
  34445=>"000010011",
  34446=>"100110010",
  34447=>"101111000",
  34448=>"001010110",
  34449=>"101011111",
  34450=>"111111001",
  34451=>"011010001",
  34452=>"011001010",
  34453=>"010011011",
  34454=>"111001011",
  34455=>"111100001",
  34456=>"110001000",
  34457=>"100000111",
  34458=>"010111001",
  34459=>"110000110",
  34460=>"100001001",
  34461=>"101010111",
  34462=>"110111000",
  34463=>"000110101",
  34464=>"001001100",
  34465=>"001011000",
  34466=>"000011101",
  34467=>"101011000",
  34468=>"101001011",
  34469=>"101000110",
  34470=>"000010001",
  34471=>"000000111",
  34472=>"010111111",
  34473=>"000001001",
  34474=>"011010001",
  34475=>"010100010",
  34476=>"110110000",
  34477=>"011100100",
  34478=>"110110110",
  34479=>"110111100",
  34480=>"000101001",
  34481=>"010111011",
  34482=>"001101100",
  34483=>"111001011",
  34484=>"111111001",
  34485=>"011100010",
  34486=>"111101001",
  34487=>"000100101",
  34488=>"000101100",
  34489=>"111000001",
  34490=>"101010001",
  34491=>"111000110",
  34492=>"101100001",
  34493=>"111000011",
  34494=>"110000110",
  34495=>"110101100",
  34496=>"110000010",
  34497=>"001010111",
  34498=>"110011001",
  34499=>"111101011",
  34500=>"101101111",
  34501=>"001100100",
  34502=>"110000001",
  34503=>"010000100",
  34504=>"101100000",
  34505=>"111010111",
  34506=>"111010011",
  34507=>"100100011",
  34508=>"100000001",
  34509=>"111110001",
  34510=>"000011000",
  34511=>"110011101",
  34512=>"011000000",
  34513=>"000010100",
  34514=>"110100001",
  34515=>"100001011",
  34516=>"100111101",
  34517=>"011010111",
  34518=>"111111100",
  34519=>"001010011",
  34520=>"100000111",
  34521=>"000111011",
  34522=>"001111001",
  34523=>"000001010",
  34524=>"111011001",
  34525=>"010100010",
  34526=>"001010001",
  34527=>"111000101",
  34528=>"010000000",
  34529=>"110011010",
  34530=>"000001101",
  34531=>"100010110",
  34532=>"110001011",
  34533=>"110001001",
  34534=>"010000011",
  34535=>"000100001",
  34536=>"110110110",
  34537=>"110101100",
  34538=>"101110011",
  34539=>"011101010",
  34540=>"010000000",
  34541=>"110110100",
  34542=>"001110101",
  34543=>"001001001",
  34544=>"100111110",
  34545=>"001000011",
  34546=>"110011101",
  34547=>"011000011",
  34548=>"010111010",
  34549=>"010100110",
  34550=>"000010110",
  34551=>"000101010",
  34552=>"010001010",
  34553=>"111000000",
  34554=>"110000001",
  34555=>"110010010",
  34556=>"000110101",
  34557=>"010001000",
  34558=>"001000110",
  34559=>"010000110",
  34560=>"000101101",
  34561=>"110100011",
  34562=>"100001011",
  34563=>"011000000",
  34564=>"000111000",
  34565=>"010010011",
  34566=>"111110001",
  34567=>"010110111",
  34568=>"111001011",
  34569=>"110111001",
  34570=>"001010000",
  34571=>"000101100",
  34572=>"110010011",
  34573=>"101000000",
  34574=>"011100100",
  34575=>"101111000",
  34576=>"000100110",
  34577=>"100001001",
  34578=>"011101101",
  34579=>"001100101",
  34580=>"000011001",
  34581=>"111100100",
  34582=>"111100010",
  34583=>"001111111",
  34584=>"010101000",
  34585=>"010100110",
  34586=>"111001101",
  34587=>"110011110",
  34588=>"111100101",
  34589=>"110000001",
  34590=>"000101011",
  34591=>"000010000",
  34592=>"111010111",
  34593=>"011010010",
  34594=>"110110100",
  34595=>"001100001",
  34596=>"000110110",
  34597=>"011101100",
  34598=>"000011000",
  34599=>"110111011",
  34600=>"110101101",
  34601=>"110101110",
  34602=>"101100000",
  34603=>"111000101",
  34604=>"100110110",
  34605=>"100010001",
  34606=>"000101000",
  34607=>"100110100",
  34608=>"010000010",
  34609=>"111100010",
  34610=>"101100001",
  34611=>"100100000",
  34612=>"111110111",
  34613=>"100101101",
  34614=>"100111011",
  34615=>"010101101",
  34616=>"010111000",
  34617=>"100110110",
  34618=>"000000001",
  34619=>"011101100",
  34620=>"000011101",
  34621=>"011000001",
  34622=>"100001110",
  34623=>"010100010",
  34624=>"011101011",
  34625=>"110000011",
  34626=>"011000011",
  34627=>"101000011",
  34628=>"100111101",
  34629=>"011111000",
  34630=>"111010010",
  34631=>"010100100",
  34632=>"110111011",
  34633=>"001011000",
  34634=>"000001100",
  34635=>"101110000",
  34636=>"100110111",
  34637=>"010100011",
  34638=>"010100010",
  34639=>"111010010",
  34640=>"001001010",
  34641=>"111110101",
  34642=>"001101101",
  34643=>"011000001",
  34644=>"010001010",
  34645=>"110001100",
  34646=>"101000011",
  34647=>"000111110",
  34648=>"110111010",
  34649=>"010000001",
  34650=>"101000001",
  34651=>"001010001",
  34652=>"011000111",
  34653=>"111111010",
  34654=>"100001100",
  34655=>"001011101",
  34656=>"000000011",
  34657=>"101011001",
  34658=>"001010011",
  34659=>"010110001",
  34660=>"100101001",
  34661=>"111000101",
  34662=>"011010010",
  34663=>"001000010",
  34664=>"011111101",
  34665=>"100110010",
  34666=>"111000000",
  34667=>"011101110",
  34668=>"010011010",
  34669=>"000001001",
  34670=>"111101101",
  34671=>"111000101",
  34672=>"111000010",
  34673=>"001011001",
  34674=>"101101101",
  34675=>"001010011",
  34676=>"010000001",
  34677=>"111010000",
  34678=>"101001111",
  34679=>"000110100",
  34680=>"010101111",
  34681=>"110001110",
  34682=>"101010111",
  34683=>"111010001",
  34684=>"000011000",
  34685=>"001010111",
  34686=>"100000001",
  34687=>"101111110",
  34688=>"001101000",
  34689=>"001000110",
  34690=>"001000011",
  34691=>"000010101",
  34692=>"001100100",
  34693=>"101000100",
  34694=>"011111100",
  34695=>"001111101",
  34696=>"011111111",
  34697=>"010110001",
  34698=>"000100011",
  34699=>"000110001",
  34700=>"110100011",
  34701=>"000010001",
  34702=>"100001100",
  34703=>"100100100",
  34704=>"100100001",
  34705=>"010110001",
  34706=>"011110000",
  34707=>"110110111",
  34708=>"000010010",
  34709=>"101111001",
  34710=>"001110000",
  34711=>"101010100",
  34712=>"010000011",
  34713=>"010100000",
  34714=>"101100111",
  34715=>"100000011",
  34716=>"111111011",
  34717=>"110110011",
  34718=>"100100111",
  34719=>"010101010",
  34720=>"111001001",
  34721=>"110100111",
  34722=>"000101000",
  34723=>"101110101",
  34724=>"011100101",
  34725=>"010100111",
  34726=>"111000100",
  34727=>"011111111",
  34728=>"001100010",
  34729=>"010110111",
  34730=>"111110010",
  34731=>"011110011",
  34732=>"010100001",
  34733=>"011110001",
  34734=>"111011001",
  34735=>"100010011",
  34736=>"001001000",
  34737=>"011010110",
  34738=>"000011111",
  34739=>"101111000",
  34740=>"100001111",
  34741=>"010001100",
  34742=>"010111111",
  34743=>"001110011",
  34744=>"010100000",
  34745=>"111000101",
  34746=>"011101101",
  34747=>"100000110",
  34748=>"111011011",
  34749=>"110111000",
  34750=>"010100010",
  34751=>"100001100",
  34752=>"010011000",
  34753=>"111000001",
  34754=>"111000001",
  34755=>"010111001",
  34756=>"100011101",
  34757=>"000010100",
  34758=>"001100100",
  34759=>"100100110",
  34760=>"000011011",
  34761=>"101000001",
  34762=>"101010101",
  34763=>"000100111",
  34764=>"101000011",
  34765=>"011111111",
  34766=>"100000011",
  34767=>"111110010",
  34768=>"001100101",
  34769=>"111111011",
  34770=>"000000011",
  34771=>"001011110",
  34772=>"000000011",
  34773=>"110101010",
  34774=>"111010000",
  34775=>"001000110",
  34776=>"111001111",
  34777=>"101110110",
  34778=>"111101000",
  34779=>"100111101",
  34780=>"001011100",
  34781=>"010011011",
  34782=>"101011111",
  34783=>"000100101",
  34784=>"110010001",
  34785=>"000001000",
  34786=>"001000000",
  34787=>"111000110",
  34788=>"101110000",
  34789=>"011111110",
  34790=>"100110001",
  34791=>"101010011",
  34792=>"001100111",
  34793=>"101111100",
  34794=>"011101011",
  34795=>"111001001",
  34796=>"010000000",
  34797=>"101000001",
  34798=>"000110100",
  34799=>"010000011",
  34800=>"110100011",
  34801=>"101000000",
  34802=>"110011111",
  34803=>"100100101",
  34804=>"011011101",
  34805=>"001001100",
  34806=>"110011101",
  34807=>"100101000",
  34808=>"101111111",
  34809=>"000111100",
  34810=>"010010001",
  34811=>"100001111",
  34812=>"100111100",
  34813=>"101111111",
  34814=>"001000100",
  34815=>"000001101",
  34816=>"100110001",
  34817=>"001000010",
  34818=>"001111000",
  34819=>"010100110",
  34820=>"000001010",
  34821=>"001010010",
  34822=>"010001110",
  34823=>"010001101",
  34824=>"011010000",
  34825=>"101101101",
  34826=>"101100000",
  34827=>"111000011",
  34828=>"001010000",
  34829=>"101111010",
  34830=>"010100011",
  34831=>"110000010",
  34832=>"010110000",
  34833=>"001001111",
  34834=>"111101011",
  34835=>"010000001",
  34836=>"111101111",
  34837=>"110100011",
  34838=>"100010101",
  34839=>"001000101",
  34840=>"010110110",
  34841=>"110000001",
  34842=>"011110001",
  34843=>"110010101",
  34844=>"100110001",
  34845=>"011011111",
  34846=>"101110100",
  34847=>"110110010",
  34848=>"010010010",
  34849=>"010010101",
  34850=>"110101111",
  34851=>"110001010",
  34852=>"100111111",
  34853=>"110010110",
  34854=>"110000011",
  34855=>"101011100",
  34856=>"011010011",
  34857=>"111100001",
  34858=>"010100010",
  34859=>"110100101",
  34860=>"000000100",
  34861=>"001110101",
  34862=>"101100010",
  34863=>"111010000",
  34864=>"100100001",
  34865=>"100000110",
  34866=>"100011010",
  34867=>"100100001",
  34868=>"110001101",
  34869=>"101001101",
  34870=>"010001100",
  34871=>"000010000",
  34872=>"111101101",
  34873=>"010100011",
  34874=>"100000010",
  34875=>"101000110",
  34876=>"100010000",
  34877=>"110011111",
  34878=>"101001101",
  34879=>"011000111",
  34880=>"100010001",
  34881=>"011100110",
  34882=>"111010001",
  34883=>"011110010",
  34884=>"001110101",
  34885=>"100111000",
  34886=>"101100001",
  34887=>"111110111",
  34888=>"100100111",
  34889=>"100000101",
  34890=>"100111001",
  34891=>"000001011",
  34892=>"011000000",
  34893=>"101101111",
  34894=>"001111000",
  34895=>"001110101",
  34896=>"011100110",
  34897=>"100110010",
  34898=>"111101111",
  34899=>"010111101",
  34900=>"101000011",
  34901=>"100101001",
  34902=>"010010011",
  34903=>"000100000",
  34904=>"100011111",
  34905=>"011100100",
  34906=>"001110110",
  34907=>"011101011",
  34908=>"100010000",
  34909=>"010111111",
  34910=>"000000011",
  34911=>"010100010",
  34912=>"000111001",
  34913=>"111111111",
  34914=>"010100101",
  34915=>"001001000",
  34916=>"001000010",
  34917=>"111101011",
  34918=>"111000111",
  34919=>"100010001",
  34920=>"011111101",
  34921=>"000010010",
  34922=>"111000001",
  34923=>"100111010",
  34924=>"110011100",
  34925=>"110001100",
  34926=>"111100110",
  34927=>"001010111",
  34928=>"101000000",
  34929=>"010011100",
  34930=>"000000010",
  34931=>"010011111",
  34932=>"011101011",
  34933=>"100100010",
  34934=>"010101011",
  34935=>"000010010",
  34936=>"110001000",
  34937=>"111110011",
  34938=>"010011100",
  34939=>"101110011",
  34940=>"010001001",
  34941=>"110110000",
  34942=>"100010110",
  34943=>"111111110",
  34944=>"011010101",
  34945=>"100100011",
  34946=>"010111000",
  34947=>"111001110",
  34948=>"100111011",
  34949=>"111000111",
  34950=>"001011010",
  34951=>"110010110",
  34952=>"010100010",
  34953=>"100010000",
  34954=>"101101100",
  34955=>"010110111",
  34956=>"101000011",
  34957=>"010110011",
  34958=>"100111001",
  34959=>"111110111",
  34960=>"111101001",
  34961=>"001110011",
  34962=>"100100101",
  34963=>"110010100",
  34964=>"101001001",
  34965=>"001000001",
  34966=>"011011011",
  34967=>"010110101",
  34968=>"101110010",
  34969=>"111000001",
  34970=>"000101010",
  34971=>"010101101",
  34972=>"101000111",
  34973=>"110001000",
  34974=>"100101000",
  34975=>"110111011",
  34976=>"100010000",
  34977=>"101101000",
  34978=>"100110100",
  34979=>"010000110",
  34980=>"100011101",
  34981=>"001010100",
  34982=>"001010101",
  34983=>"011011111",
  34984=>"011001011",
  34985=>"011011001",
  34986=>"110011100",
  34987=>"101000110",
  34988=>"111001100",
  34989=>"100110100",
  34990=>"101011110",
  34991=>"011101001",
  34992=>"100001111",
  34993=>"001011110",
  34994=>"010110001",
  34995=>"110111101",
  34996=>"111111100",
  34997=>"000010100",
  34998=>"001101010",
  34999=>"100010100",
  35000=>"000111011",
  35001=>"001100001",
  35002=>"110001010",
  35003=>"111101101",
  35004=>"000011000",
  35005=>"111000101",
  35006=>"011110000",
  35007=>"011111001",
  35008=>"111011001",
  35009=>"010000110",
  35010=>"001000001",
  35011=>"000001011",
  35012=>"111100000",
  35013=>"110110011",
  35014=>"101100010",
  35015=>"110111010",
  35016=>"001110110",
  35017=>"011110001",
  35018=>"110010100",
  35019=>"010110011",
  35020=>"011110010",
  35021=>"101010100",
  35022=>"010010010",
  35023=>"011000110",
  35024=>"011011100",
  35025=>"110111101",
  35026=>"000010110",
  35027=>"011011111",
  35028=>"011101011",
  35029=>"111010111",
  35030=>"111010001",
  35031=>"001111111",
  35032=>"011101100",
  35033=>"100000000",
  35034=>"000000000",
  35035=>"000000001",
  35036=>"110011101",
  35037=>"001000101",
  35038=>"010011011",
  35039=>"101001111",
  35040=>"000000101",
  35041=>"011010000",
  35042=>"110010000",
  35043=>"100101001",
  35044=>"000010110",
  35045=>"100011000",
  35046=>"011001100",
  35047=>"111110001",
  35048=>"111111011",
  35049=>"010100010",
  35050=>"110000100",
  35051=>"100110000",
  35052=>"111101110",
  35053=>"111110011",
  35054=>"110110000",
  35055=>"001101011",
  35056=>"010000001",
  35057=>"001000011",
  35058=>"001100000",
  35059=>"101010100",
  35060=>"100110000",
  35061=>"100100101",
  35062=>"111011010",
  35063=>"011111000",
  35064=>"011010001",
  35065=>"101111100",
  35066=>"100001000",
  35067=>"001111010",
  35068=>"101101011",
  35069=>"000000101",
  35070=>"111100111",
  35071=>"001110100",
  35072=>"100100110",
  35073=>"101111010",
  35074=>"101011001",
  35075=>"000110111",
  35076=>"100001010",
  35077=>"001111101",
  35078=>"001100100",
  35079=>"111010100",
  35080=>"001110101",
  35081=>"001100111",
  35082=>"011011000",
  35083=>"001001000",
  35084=>"111001001",
  35085=>"001101110",
  35086=>"010110110",
  35087=>"001101011",
  35088=>"110100101",
  35089=>"010101001",
  35090=>"101001101",
  35091=>"000010000",
  35092=>"111110101",
  35093=>"111000100",
  35094=>"101011111",
  35095=>"101001111",
  35096=>"001101100",
  35097=>"101001000",
  35098=>"010000100",
  35099=>"100000010",
  35100=>"110110000",
  35101=>"101010001",
  35102=>"100010010",
  35103=>"110010011",
  35104=>"101010110",
  35105=>"010011010",
  35106=>"000110000",
  35107=>"011101100",
  35108=>"001011100",
  35109=>"011101011",
  35110=>"111101011",
  35111=>"010010111",
  35112=>"010011011",
  35113=>"011110100",
  35114=>"010110100",
  35115=>"000001011",
  35116=>"011010100",
  35117=>"001001101",
  35118=>"001001100",
  35119=>"110111011",
  35120=>"111011110",
  35121=>"110010001",
  35122=>"000101101",
  35123=>"000001101",
  35124=>"101111100",
  35125=>"001000010",
  35126=>"111011100",
  35127=>"100010000",
  35128=>"100010011",
  35129=>"001100100",
  35130=>"111110101",
  35131=>"000000001",
  35132=>"101111111",
  35133=>"110101010",
  35134=>"100101101",
  35135=>"111110011",
  35136=>"110011101",
  35137=>"010000011",
  35138=>"000110100",
  35139=>"111110011",
  35140=>"100011101",
  35141=>"011111010",
  35142=>"000101001",
  35143=>"110101110",
  35144=>"101001111",
  35145=>"110001011",
  35146=>"001110101",
  35147=>"010101010",
  35148=>"000000101",
  35149=>"010111111",
  35150=>"001111110",
  35151=>"011110000",
  35152=>"101000100",
  35153=>"011111100",
  35154=>"001011000",
  35155=>"100000000",
  35156=>"100010100",
  35157=>"010101110",
  35158=>"000011001",
  35159=>"000000101",
  35160=>"111100001",
  35161=>"100000101",
  35162=>"000011010",
  35163=>"110000001",
  35164=>"101100000",
  35165=>"111111001",
  35166=>"111011010",
  35167=>"110000001",
  35168=>"100010110",
  35169=>"101101100",
  35170=>"001101010",
  35171=>"110111100",
  35172=>"100010010",
  35173=>"100101101",
  35174=>"100100010",
  35175=>"100000010",
  35176=>"011010110",
  35177=>"000000101",
  35178=>"001010101",
  35179=>"001110001",
  35180=>"011000100",
  35181=>"001011101",
  35182=>"001100001",
  35183=>"010000010",
  35184=>"010101010",
  35185=>"010110111",
  35186=>"111101111",
  35187=>"111001011",
  35188=>"100010001",
  35189=>"110010100",
  35190=>"110011101",
  35191=>"011110011",
  35192=>"010100001",
  35193=>"001011001",
  35194=>"001001000",
  35195=>"011000011",
  35196=>"011000000",
  35197=>"000110110",
  35198=>"111101101",
  35199=>"011101110",
  35200=>"010010011",
  35201=>"111011000",
  35202=>"111101011",
  35203=>"110110010",
  35204=>"010001000",
  35205=>"011001111",
  35206=>"001100001",
  35207=>"111101101",
  35208=>"011010000",
  35209=>"110110010",
  35210=>"111001101",
  35211=>"000010110",
  35212=>"001010100",
  35213=>"110000110",
  35214=>"110101000",
  35215=>"000100010",
  35216=>"101101010",
  35217=>"011000000",
  35218=>"101010111",
  35219=>"110001001",
  35220=>"111010111",
  35221=>"001110111",
  35222=>"110010111",
  35223=>"000000100",
  35224=>"000000100",
  35225=>"101101111",
  35226=>"001101101",
  35227=>"100110011",
  35228=>"001000010",
  35229=>"011101010",
  35230=>"011111111",
  35231=>"011110111",
  35232=>"110010000",
  35233=>"111010011",
  35234=>"010111011",
  35235=>"101101001",
  35236=>"100000100",
  35237=>"011011000",
  35238=>"000010100",
  35239=>"111000110",
  35240=>"111110100",
  35241=>"001001001",
  35242=>"101001000",
  35243=>"001110000",
  35244=>"100000010",
  35245=>"011101010",
  35246=>"100010101",
  35247=>"010111011",
  35248=>"111010011",
  35249=>"111111111",
  35250=>"110000011",
  35251=>"001000100",
  35252=>"010111011",
  35253=>"000110000",
  35254=>"000000111",
  35255=>"011010001",
  35256=>"011111011",
  35257=>"011100010",
  35258=>"111011011",
  35259=>"111111001",
  35260=>"110110011",
  35261=>"100111100",
  35262=>"010000111",
  35263=>"101000110",
  35264=>"110000100",
  35265=>"100101100",
  35266=>"010110110",
  35267=>"001101110",
  35268=>"111111010",
  35269=>"011111110",
  35270=>"011010000",
  35271=>"011110010",
  35272=>"001001010",
  35273=>"110110100",
  35274=>"000110000",
  35275=>"111011110",
  35276=>"110111100",
  35277=>"010101110",
  35278=>"001001000",
  35279=>"000010011",
  35280=>"011111011",
  35281=>"100011001",
  35282=>"000100100",
  35283=>"011110100",
  35284=>"001100011",
  35285=>"000100001",
  35286=>"010000000",
  35287=>"011100000",
  35288=>"000110101",
  35289=>"011101011",
  35290=>"101111000",
  35291=>"010101000",
  35292=>"001000000",
  35293=>"100110110",
  35294=>"111100010",
  35295=>"010000110",
  35296=>"000100101",
  35297=>"010010100",
  35298=>"110110111",
  35299=>"011101011",
  35300=>"011011100",
  35301=>"101110101",
  35302=>"110010000",
  35303=>"110111011",
  35304=>"010101000",
  35305=>"000100010",
  35306=>"000110001",
  35307=>"111100110",
  35308=>"111111111",
  35309=>"010001101",
  35310=>"101001010",
  35311=>"011101011",
  35312=>"110111101",
  35313=>"011101111",
  35314=>"011000011",
  35315=>"100010101",
  35316=>"001010111",
  35317=>"101100011",
  35318=>"101111101",
  35319=>"111100100",
  35320=>"001001010",
  35321=>"100100010",
  35322=>"010110000",
  35323=>"101111101",
  35324=>"101110111",
  35325=>"000010111",
  35326=>"101011110",
  35327=>"100000000",
  35328=>"100100000",
  35329=>"111011111",
  35330=>"110001010",
  35331=>"101011111",
  35332=>"011011100",
  35333=>"101011011",
  35334=>"001110001",
  35335=>"110110101",
  35336=>"011001000",
  35337=>"100110000",
  35338=>"100000100",
  35339=>"010010010",
  35340=>"100111111",
  35341=>"000111000",
  35342=>"000111011",
  35343=>"111111011",
  35344=>"100110100",
  35345=>"100111011",
  35346=>"000000000",
  35347=>"000101100",
  35348=>"011001001",
  35349=>"001101000",
  35350=>"110110000",
  35351=>"101111001",
  35352=>"010101101",
  35353=>"000111000",
  35354=>"001001010",
  35355=>"111111111",
  35356=>"001001010",
  35357=>"101111000",
  35358=>"001011000",
  35359=>"010000101",
  35360=>"111101101",
  35361=>"100111101",
  35362=>"001111111",
  35363=>"000111111",
  35364=>"111100001",
  35365=>"010000001",
  35366=>"110001001",
  35367=>"010101111",
  35368=>"000001010",
  35369=>"100010110",
  35370=>"100000000",
  35371=>"000101101",
  35372=>"111101011",
  35373=>"010100101",
  35374=>"000001101",
  35375=>"000000101",
  35376=>"100101101",
  35377=>"010110001",
  35378=>"010011001",
  35379=>"111010101",
  35380=>"001011001",
  35381=>"111010111",
  35382=>"001001000",
  35383=>"001010111",
  35384=>"100011011",
  35385=>"101000000",
  35386=>"111011110",
  35387=>"110101100",
  35388=>"001000011",
  35389=>"010101001",
  35390=>"001100111",
  35391=>"000101101",
  35392=>"110101110",
  35393=>"101110000",
  35394=>"101000000",
  35395=>"101110111",
  35396=>"110100010",
  35397=>"101101100",
  35398=>"111001101",
  35399=>"010101101",
  35400=>"011010100",
  35401=>"001101000",
  35402=>"100000100",
  35403=>"011001000",
  35404=>"001001011",
  35405=>"110111101",
  35406=>"110100000",
  35407=>"101011000",
  35408=>"100110001",
  35409=>"001001111",
  35410=>"000000110",
  35411=>"100011011",
  35412=>"010101111",
  35413=>"000001000",
  35414=>"100110000",
  35415=>"001111000",
  35416=>"111001000",
  35417=>"110010010",
  35418=>"000100101",
  35419=>"000001011",
  35420=>"010011011",
  35421=>"110100101",
  35422=>"000101010",
  35423=>"100101110",
  35424=>"101010111",
  35425=>"001111000",
  35426=>"110010011",
  35427=>"010111010",
  35428=>"110010000",
  35429=>"101001001",
  35430=>"110001110",
  35431=>"000011101",
  35432=>"101000001",
  35433=>"110100110",
  35434=>"011100111",
  35435=>"001000000",
  35436=>"101000110",
  35437=>"101111111",
  35438=>"000011000",
  35439=>"101010111",
  35440=>"010100011",
  35441=>"001100010",
  35442=>"110000111",
  35443=>"011000010",
  35444=>"110111011",
  35445=>"010000000",
  35446=>"100101111",
  35447=>"101110100",
  35448=>"100011010",
  35449=>"111001110",
  35450=>"001110011",
  35451=>"010100011",
  35452=>"001010101",
  35453=>"110101111",
  35454=>"110100100",
  35455=>"000001001",
  35456=>"001001101",
  35457=>"101001011",
  35458=>"011100000",
  35459=>"001100101",
  35460=>"000011001",
  35461=>"101110110",
  35462=>"110001011",
  35463=>"000110101",
  35464=>"000110001",
  35465=>"111101001",
  35466=>"010001011",
  35467=>"001000011",
  35468=>"100100000",
  35469=>"110011111",
  35470=>"101111100",
  35471=>"111110111",
  35472=>"011011000",
  35473=>"011100011",
  35474=>"010001010",
  35475=>"011111100",
  35476=>"101100100",
  35477=>"111010010",
  35478=>"000100100",
  35479=>"001111001",
  35480=>"110001100",
  35481=>"010100000",
  35482=>"011101000",
  35483=>"010010010",
  35484=>"001111111",
  35485=>"001111001",
  35486=>"010111110",
  35487=>"100111010",
  35488=>"100110101",
  35489=>"010011010",
  35490=>"000100001",
  35491=>"011110011",
  35492=>"000001111",
  35493=>"000111110",
  35494=>"100011010",
  35495=>"110000001",
  35496=>"000110010",
  35497=>"000000010",
  35498=>"001101001",
  35499=>"010110010",
  35500=>"101110111",
  35501=>"001011101",
  35502=>"111010111",
  35503=>"001011011",
  35504=>"000000011",
  35505=>"010011101",
  35506=>"111010111",
  35507=>"101011000",
  35508=>"101100000",
  35509=>"111110010",
  35510=>"000000000",
  35511=>"100100111",
  35512=>"000001000",
  35513=>"011111100",
  35514=>"100010110",
  35515=>"001011001",
  35516=>"000011001",
  35517=>"111101011",
  35518=>"000001011",
  35519=>"111101101",
  35520=>"011010101",
  35521=>"110001000",
  35522=>"101001111",
  35523=>"111001100",
  35524=>"010110011",
  35525=>"010111101",
  35526=>"000100100",
  35527=>"000010001",
  35528=>"110010110",
  35529=>"000001101",
  35530=>"110001010",
  35531=>"110001111",
  35532=>"000000100",
  35533=>"101000001",
  35534=>"010000000",
  35535=>"100001001",
  35536=>"001010110",
  35537=>"110010110",
  35538=>"101011001",
  35539=>"110010010",
  35540=>"010110110",
  35541=>"110011111",
  35542=>"111010001",
  35543=>"101110001",
  35544=>"101100101",
  35545=>"000110100",
  35546=>"100101101",
  35547=>"000010000",
  35548=>"101100011",
  35549=>"001100000",
  35550=>"001100111",
  35551=>"010111010",
  35552=>"111000000",
  35553=>"111110000",
  35554=>"011011000",
  35555=>"111001110",
  35556=>"010011000",
  35557=>"000010010",
  35558=>"111010000",
  35559=>"111011100",
  35560=>"101101110",
  35561=>"100000101",
  35562=>"101101111",
  35563=>"100010101",
  35564=>"100011011",
  35565=>"010001001",
  35566=>"011011001",
  35567=>"010010111",
  35568=>"101001111",
  35569=>"110111001",
  35570=>"100010011",
  35571=>"001011010",
  35572=>"111100110",
  35573=>"001111010",
  35574=>"101110011",
  35575=>"111001110",
  35576=>"000110010",
  35577=>"111110110",
  35578=>"111011010",
  35579=>"101010001",
  35580=>"110110111",
  35581=>"100001001",
  35582=>"100101111",
  35583=>"100011110",
  35584=>"100100110",
  35585=>"111010011",
  35586=>"100001000",
  35587=>"010110101",
  35588=>"000110110",
  35589=>"111110100",
  35590=>"010110110",
  35591=>"011011110",
  35592=>"000010111",
  35593=>"000011011",
  35594=>"100110110",
  35595=>"111101001",
  35596=>"000001010",
  35597=>"010100011",
  35598=>"111101001",
  35599=>"000100000",
  35600=>"110000010",
  35601=>"101100001",
  35602=>"011110111",
  35603=>"000101101",
  35604=>"111010001",
  35605=>"011010110",
  35606=>"011011101",
  35607=>"100000000",
  35608=>"110000000",
  35609=>"101100010",
  35610=>"000001110",
  35611=>"001010110",
  35612=>"111011010",
  35613=>"100111001",
  35614=>"001001111",
  35615=>"000100011",
  35616=>"000001011",
  35617=>"001000101",
  35618=>"100101011",
  35619=>"010110000",
  35620=>"010100100",
  35621=>"101001000",
  35622=>"011011011",
  35623=>"100111100",
  35624=>"101000111",
  35625=>"000100101",
  35626=>"010101110",
  35627=>"110101101",
  35628=>"000011110",
  35629=>"101001010",
  35630=>"101011101",
  35631=>"010100010",
  35632=>"001100011",
  35633=>"110101100",
  35634=>"111001100",
  35635=>"111010100",
  35636=>"001000101",
  35637=>"000000010",
  35638=>"000001001",
  35639=>"001110111",
  35640=>"001101010",
  35641=>"011111101",
  35642=>"000010111",
  35643=>"000100101",
  35644=>"100101101",
  35645=>"101110110",
  35646=>"111010110",
  35647=>"011000011",
  35648=>"000000011",
  35649=>"101101111",
  35650=>"100001011",
  35651=>"101110101",
  35652=>"100111011",
  35653=>"100111011",
  35654=>"100100110",
  35655=>"000100100",
  35656=>"001001011",
  35657=>"111010010",
  35658=>"010011000",
  35659=>"000000101",
  35660=>"111101011",
  35661=>"000101010",
  35662=>"101001100",
  35663=>"011010100",
  35664=>"000000101",
  35665=>"101001101",
  35666=>"000101000",
  35667=>"101010100",
  35668=>"110100011",
  35669=>"100100100",
  35670=>"111001001",
  35671=>"000100011",
  35672=>"101100111",
  35673=>"011110011",
  35674=>"000100100",
  35675=>"000101111",
  35676=>"101000001",
  35677=>"111111111",
  35678=>"000001001",
  35679=>"110011111",
  35680=>"000001011",
  35681=>"011100001",
  35682=>"111011111",
  35683=>"001110011",
  35684=>"001100001",
  35685=>"110001100",
  35686=>"100001110",
  35687=>"000101000",
  35688=>"100100100",
  35689=>"101011110",
  35690=>"010110110",
  35691=>"100100010",
  35692=>"000000100",
  35693=>"101100110",
  35694=>"010100110",
  35695=>"111010101",
  35696=>"000010110",
  35697=>"011110100",
  35698=>"101001001",
  35699=>"011011001",
  35700=>"110101011",
  35701=>"010111011",
  35702=>"010000100",
  35703=>"010001010",
  35704=>"100011101",
  35705=>"110110101",
  35706=>"100111111",
  35707=>"111110001",
  35708=>"101011100",
  35709=>"011101100",
  35710=>"010001111",
  35711=>"111111100",
  35712=>"011111010",
  35713=>"100010001",
  35714=>"000101110",
  35715=>"000010100",
  35716=>"011000110",
  35717=>"101101100",
  35718=>"110101000",
  35719=>"110111100",
  35720=>"100110000",
  35721=>"100100011",
  35722=>"110101111",
  35723=>"111110111",
  35724=>"000001111",
  35725=>"011011011",
  35726=>"011101100",
  35727=>"100101111",
  35728=>"101000000",
  35729=>"110101010",
  35730=>"110100100",
  35731=>"011110111",
  35732=>"011000010",
  35733=>"011111101",
  35734=>"011111110",
  35735=>"000011011",
  35736=>"011010110",
  35737=>"101001111",
  35738=>"100011111",
  35739=>"101000100",
  35740=>"011110010",
  35741=>"010110110",
  35742=>"010000001",
  35743=>"100111100",
  35744=>"000110011",
  35745=>"101110000",
  35746=>"001010011",
  35747=>"001110111",
  35748=>"000111111",
  35749=>"110000000",
  35750=>"011110100",
  35751=>"000110000",
  35752=>"100000100",
  35753=>"100110111",
  35754=>"010010011",
  35755=>"100010000",
  35756=>"000101001",
  35757=>"110101101",
  35758=>"010110100",
  35759=>"000011111",
  35760=>"110000110",
  35761=>"110010100",
  35762=>"100000100",
  35763=>"001011000",
  35764=>"101110110",
  35765=>"000000001",
  35766=>"100010000",
  35767=>"110111110",
  35768=>"000011111",
  35769=>"010110110",
  35770=>"010111001",
  35771=>"100010011",
  35772=>"011111010",
  35773=>"111100100",
  35774=>"010111100",
  35775=>"000001111",
  35776=>"010000010",
  35777=>"101101000",
  35778=>"100001010",
  35779=>"001110010",
  35780=>"010100011",
  35781=>"100100101",
  35782=>"110010111",
  35783=>"010001011",
  35784=>"101100010",
  35785=>"010001001",
  35786=>"100100110",
  35787=>"001001011",
  35788=>"010000111",
  35789=>"100001110",
  35790=>"101010000",
  35791=>"101111000",
  35792=>"001011001",
  35793=>"011011011",
  35794=>"000000111",
  35795=>"110110000",
  35796=>"010000101",
  35797=>"101111011",
  35798=>"010000000",
  35799=>"000110000",
  35800=>"010110100",
  35801=>"100010001",
  35802=>"011000011",
  35803=>"101101001",
  35804=>"010001001",
  35805=>"101011111",
  35806=>"101101101",
  35807=>"111111110",
  35808=>"000011000",
  35809=>"111010010",
  35810=>"001100100",
  35811=>"101110010",
  35812=>"100100100",
  35813=>"101110000",
  35814=>"101110111",
  35815=>"111101000",
  35816=>"010011001",
  35817=>"010000110",
  35818=>"001101110",
  35819=>"001001111",
  35820=>"110100100",
  35821=>"000001101",
  35822=>"111111000",
  35823=>"000110110",
  35824=>"100001101",
  35825=>"000000100",
  35826=>"011101111",
  35827=>"110001111",
  35828=>"000010011",
  35829=>"100010110",
  35830=>"111011111",
  35831=>"101011010",
  35832=>"111000000",
  35833=>"111111100",
  35834=>"010000101",
  35835=>"110111011",
  35836=>"101101110",
  35837=>"011101111",
  35838=>"000011100",
  35839=>"010101101",
  35840=>"111000100",
  35841=>"001001111",
  35842=>"010111010",
  35843=>"010001011",
  35844=>"110100101",
  35845=>"111000011",
  35846=>"001000111",
  35847=>"110010010",
  35848=>"001111011",
  35849=>"001000111",
  35850=>"100010101",
  35851=>"011011011",
  35852=>"110011010",
  35853=>"001000010",
  35854=>"111111100",
  35855=>"001010100",
  35856=>"010111010",
  35857=>"100010100",
  35858=>"000011111",
  35859=>"100100010",
  35860=>"000000110",
  35861=>"100000011",
  35862=>"010110111",
  35863=>"110010000",
  35864=>"100101001",
  35865=>"001110110",
  35866=>"110111111",
  35867=>"100000010",
  35868=>"110101001",
  35869=>"000101100",
  35870=>"100100101",
  35871=>"100110011",
  35872=>"011010010",
  35873=>"001001011",
  35874=>"000100000",
  35875=>"100111010",
  35876=>"111100111",
  35877=>"010001011",
  35878=>"101010011",
  35879=>"010110100",
  35880=>"011110100",
  35881=>"000000110",
  35882=>"111001111",
  35883=>"001100001",
  35884=>"101010011",
  35885=>"110010101",
  35886=>"110001111",
  35887=>"000010110",
  35888=>"001001100",
  35889=>"110001000",
  35890=>"010100001",
  35891=>"101100100",
  35892=>"011111111",
  35893=>"010001011",
  35894=>"110010001",
  35895=>"000101110",
  35896=>"001011101",
  35897=>"011001110",
  35898=>"110001111",
  35899=>"000011001",
  35900=>"111000111",
  35901=>"101100011",
  35902=>"100111001",
  35903=>"011101100",
  35904=>"001010000",
  35905=>"111110101",
  35906=>"010010110",
  35907=>"111110010",
  35908=>"101000110",
  35909=>"110111011",
  35910=>"011100110",
  35911=>"101010101",
  35912=>"000001110",
  35913=>"110001100",
  35914=>"111110110",
  35915=>"010111001",
  35916=>"111001111",
  35917=>"010010001",
  35918=>"001100010",
  35919=>"111010011",
  35920=>"101111111",
  35921=>"100010000",
  35922=>"000000011",
  35923=>"111010001",
  35924=>"101111111",
  35925=>"101000010",
  35926=>"110000001",
  35927=>"000100010",
  35928=>"001101100",
  35929=>"011110101",
  35930=>"101000000",
  35931=>"111110110",
  35932=>"000111010",
  35933=>"100001010",
  35934=>"000111001",
  35935=>"101011100",
  35936=>"011110000",
  35937=>"001100001",
  35938=>"010100100",
  35939=>"001110011",
  35940=>"110010001",
  35941=>"000101000",
  35942=>"001001111",
  35943=>"000000001",
  35944=>"101101100",
  35945=>"101111011",
  35946=>"111100101",
  35947=>"101010000",
  35948=>"000010100",
  35949=>"000101011",
  35950=>"110011000",
  35951=>"001001100",
  35952=>"101100000",
  35953=>"010010111",
  35954=>"010010000",
  35955=>"001100010",
  35956=>"001100001",
  35957=>"111011011",
  35958=>"100010101",
  35959=>"011000111",
  35960=>"001010011",
  35961=>"001110010",
  35962=>"111110000",
  35963=>"000111110",
  35964=>"011010010",
  35965=>"011101011",
  35966=>"110010000",
  35967=>"111011001",
  35968=>"001010011",
  35969=>"001100100",
  35970=>"010011011",
  35971=>"111100001",
  35972=>"111111101",
  35973=>"100111010",
  35974=>"110011011",
  35975=>"010011110",
  35976=>"101100111",
  35977=>"010110101",
  35978=>"101110110",
  35979=>"110001011",
  35980=>"001110000",
  35981=>"000010000",
  35982=>"001000111",
  35983=>"111001111",
  35984=>"011000101",
  35985=>"010011000",
  35986=>"111110010",
  35987=>"010100110",
  35988=>"111111111",
  35989=>"111111110",
  35990=>"110000000",
  35991=>"011110111",
  35992=>"010110110",
  35993=>"011100111",
  35994=>"111101101",
  35995=>"101101101",
  35996=>"010001110",
  35997=>"000101000",
  35998=>"100010001",
  35999=>"011111000",
  36000=>"111001111",
  36001=>"000001110",
  36002=>"010100110",
  36003=>"100100100",
  36004=>"011110010",
  36005=>"111111001",
  36006=>"001011101",
  36007=>"011010010",
  36008=>"100110110",
  36009=>"100111001",
  36010=>"000110100",
  36011=>"011000001",
  36012=>"100110111",
  36013=>"011000000",
  36014=>"011011001",
  36015=>"000010110",
  36016=>"001111101",
  36017=>"101110000",
  36018=>"111101111",
  36019=>"010011111",
  36020=>"111000010",
  36021=>"101000011",
  36022=>"011111001",
  36023=>"001010110",
  36024=>"111000100",
  36025=>"011001001",
  36026=>"101011010",
  36027=>"010110011",
  36028=>"101111011",
  36029=>"010111000",
  36030=>"000101110",
  36031=>"101000010",
  36032=>"001001000",
  36033=>"100010101",
  36034=>"000100111",
  36035=>"111000001",
  36036=>"000000111",
  36037=>"000000100",
  36038=>"011001011",
  36039=>"000101010",
  36040=>"011010001",
  36041=>"000111100",
  36042=>"101000110",
  36043=>"100011011",
  36044=>"011000000",
  36045=>"000000011",
  36046=>"111111010",
  36047=>"001110111",
  36048=>"110010000",
  36049=>"010100000",
  36050=>"000001000",
  36051=>"110110110",
  36052=>"000100000",
  36053=>"010111100",
  36054=>"010100000",
  36055=>"010000101",
  36056=>"101100010",
  36057=>"011000011",
  36058=>"111001001",
  36059=>"000110111",
  36060=>"001100110",
  36061=>"100110010",
  36062=>"101110100",
  36063=>"111000110",
  36064=>"101001001",
  36065=>"111011000",
  36066=>"011001011",
  36067=>"000101110",
  36068=>"100111001",
  36069=>"100101010",
  36070=>"111101000",
  36071=>"111111001",
  36072=>"001110110",
  36073=>"100100110",
  36074=>"010110011",
  36075=>"110010010",
  36076=>"011100100",
  36077=>"111001110",
  36078=>"111011001",
  36079=>"000001000",
  36080=>"100100111",
  36081=>"000110101",
  36082=>"100100000",
  36083=>"100001110",
  36084=>"111101111",
  36085=>"111100101",
  36086=>"001100000",
  36087=>"010011101",
  36088=>"001000010",
  36089=>"011001110",
  36090=>"010110100",
  36091=>"010000000",
  36092=>"010110010",
  36093=>"010001111",
  36094=>"101111001",
  36095=>"001110000",
  36096=>"010111101",
  36097=>"110101100",
  36098=>"010011100",
  36099=>"110100111",
  36100=>"100101010",
  36101=>"100010001",
  36102=>"010010110",
  36103=>"101100110",
  36104=>"100111111",
  36105=>"001110000",
  36106=>"011100101",
  36107=>"000110000",
  36108=>"100001001",
  36109=>"111100111",
  36110=>"110110101",
  36111=>"000110101",
  36112=>"111000100",
  36113=>"100101100",
  36114=>"000100000",
  36115=>"101111011",
  36116=>"001100100",
  36117=>"100100001",
  36118=>"001101001",
  36119=>"100111010",
  36120=>"111101011",
  36121=>"000100000",
  36122=>"110011101",
  36123=>"110111100",
  36124=>"010110001",
  36125=>"101110111",
  36126=>"010001100",
  36127=>"001000011",
  36128=>"010010100",
  36129=>"010001010",
  36130=>"000000011",
  36131=>"101101001",
  36132=>"111101000",
  36133=>"111110001",
  36134=>"010001101",
  36135=>"000010010",
  36136=>"110010011",
  36137=>"010101110",
  36138=>"000000010",
  36139=>"010111010",
  36140=>"001001001",
  36141=>"100011101",
  36142=>"111000011",
  36143=>"101001111",
  36144=>"110011011",
  36145=>"101100000",
  36146=>"000000101",
  36147=>"000000011",
  36148=>"011001001",
  36149=>"110111001",
  36150=>"010001000",
  36151=>"111011000",
  36152=>"000001000",
  36153=>"100100000",
  36154=>"011100111",
  36155=>"000001010",
  36156=>"110000111",
  36157=>"100011100",
  36158=>"000000001",
  36159=>"010010001",
  36160=>"111011010",
  36161=>"010111100",
  36162=>"111001111",
  36163=>"101110000",
  36164=>"100001101",
  36165=>"011100110",
  36166=>"100010100",
  36167=>"010000110",
  36168=>"000010000",
  36169=>"100100000",
  36170=>"101111011",
  36171=>"001010001",
  36172=>"110011011",
  36173=>"110100001",
  36174=>"011011001",
  36175=>"010001111",
  36176=>"010001110",
  36177=>"100000011",
  36178=>"110101100",
  36179=>"011111001",
  36180=>"100001000",
  36181=>"111110101",
  36182=>"010100101",
  36183=>"000101100",
  36184=>"111111011",
  36185=>"100001010",
  36186=>"000010000",
  36187=>"110100101",
  36188=>"100001111",
  36189=>"011000101",
  36190=>"001101000",
  36191=>"000011100",
  36192=>"110100110",
  36193=>"100001000",
  36194=>"000110000",
  36195=>"010010101",
  36196=>"111110001",
  36197=>"010001100",
  36198=>"001001110",
  36199=>"111001000",
  36200=>"001011100",
  36201=>"110111101",
  36202=>"111000110",
  36203=>"011100101",
  36204=>"011000110",
  36205=>"101001111",
  36206=>"100001111",
  36207=>"111101011",
  36208=>"100001100",
  36209=>"101000000",
  36210=>"000000010",
  36211=>"111011100",
  36212=>"001110110",
  36213=>"000011111",
  36214=>"110000000",
  36215=>"100110101",
  36216=>"101001100",
  36217=>"010000011",
  36218=>"100010011",
  36219=>"111100000",
  36220=>"000111010",
  36221=>"101000101",
  36222=>"010010001",
  36223=>"001100101",
  36224=>"011001000",
  36225=>"010000100",
  36226=>"101011001",
  36227=>"000010100",
  36228=>"111000101",
  36229=>"001000101",
  36230=>"000000100",
  36231=>"000100101",
  36232=>"111000000",
  36233=>"011100000",
  36234=>"010100001",
  36235=>"111001010",
  36236=>"000000100",
  36237=>"100111010",
  36238=>"110110110",
  36239=>"110110101",
  36240=>"110101001",
  36241=>"001000111",
  36242=>"100010001",
  36243=>"001101100",
  36244=>"100011110",
  36245=>"111110000",
  36246=>"111111111",
  36247=>"010100111",
  36248=>"001101110",
  36249=>"100111101",
  36250=>"110001011",
  36251=>"100010000",
  36252=>"000000110",
  36253=>"001111001",
  36254=>"100001011",
  36255=>"001101111",
  36256=>"001010011",
  36257=>"101100001",
  36258=>"110001010",
  36259=>"110010001",
  36260=>"000101111",
  36261=>"110011100",
  36262=>"001100111",
  36263=>"011110010",
  36264=>"000101000",
  36265=>"101100100",
  36266=>"011001100",
  36267=>"001000100",
  36268=>"101001100",
  36269=>"110000000",
  36270=>"100101100",
  36271=>"011101111",
  36272=>"001011010",
  36273=>"100010011",
  36274=>"110011110",
  36275=>"000001001",
  36276=>"011011100",
  36277=>"000101011",
  36278=>"100111111",
  36279=>"100101001",
  36280=>"111011010",
  36281=>"110011100",
  36282=>"100010000",
  36283=>"001001100",
  36284=>"100101111",
  36285=>"001110101",
  36286=>"100001010",
  36287=>"111001001",
  36288=>"010111111",
  36289=>"100110011",
  36290=>"010011011",
  36291=>"101110010",
  36292=>"001100100",
  36293=>"100010101",
  36294=>"101001000",
  36295=>"001110000",
  36296=>"001111100",
  36297=>"100111001",
  36298=>"001100101",
  36299=>"010100010",
  36300=>"000000111",
  36301=>"101011000",
  36302=>"011001001",
  36303=>"010011001",
  36304=>"001011000",
  36305=>"001111011",
  36306=>"110101011",
  36307=>"000010110",
  36308=>"111011101",
  36309=>"010000000",
  36310=>"111011111",
  36311=>"111011111",
  36312=>"110000111",
  36313=>"101110110",
  36314=>"101000000",
  36315=>"001111000",
  36316=>"010100101",
  36317=>"001000100",
  36318=>"010000010",
  36319=>"000000001",
  36320=>"100100111",
  36321=>"000111001",
  36322=>"011011100",
  36323=>"111111100",
  36324=>"011100110",
  36325=>"010001111",
  36326=>"011101000",
  36327=>"010110100",
  36328=>"100010011",
  36329=>"011010011",
  36330=>"111100011",
  36331=>"011011100",
  36332=>"110001000",
  36333=>"000111000",
  36334=>"110111100",
  36335=>"010010100",
  36336=>"111111101",
  36337=>"111000011",
  36338=>"110100011",
  36339=>"000011011",
  36340=>"010001000",
  36341=>"110101111",
  36342=>"111110010",
  36343=>"011000001",
  36344=>"010011000",
  36345=>"101100100",
  36346=>"101111011",
  36347=>"110011100",
  36348=>"010101101",
  36349=>"111000010",
  36350=>"011001011",
  36351=>"001010101",
  36352=>"111011011",
  36353=>"101100000",
  36354=>"001101110",
  36355=>"011100101",
  36356=>"101111101",
  36357=>"110011010",
  36358=>"001010011",
  36359=>"011000110",
  36360=>"001000001",
  36361=>"011010001",
  36362=>"001010011",
  36363=>"010101001",
  36364=>"010011110",
  36365=>"100111010",
  36366=>"010101011",
  36367=>"010100010",
  36368=>"100000111",
  36369=>"010100100",
  36370=>"110110110",
  36371=>"111010000",
  36372=>"110011100",
  36373=>"011000011",
  36374=>"111100111",
  36375=>"101011001",
  36376=>"000000111",
  36377=>"101111011",
  36378=>"010100110",
  36379=>"110001001",
  36380=>"111111000",
  36381=>"101000000",
  36382=>"111111001",
  36383=>"100101011",
  36384=>"111001110",
  36385=>"010010001",
  36386=>"010100010",
  36387=>"000001000",
  36388=>"000000111",
  36389=>"111100111",
  36390=>"011101111",
  36391=>"101000010",
  36392=>"001101111",
  36393=>"011111000",
  36394=>"000110111",
  36395=>"100011111",
  36396=>"101110010",
  36397=>"110100110",
  36398=>"010100001",
  36399=>"000101000",
  36400=>"111101001",
  36401=>"101101000",
  36402=>"111110110",
  36403=>"100011010",
  36404=>"110101100",
  36405=>"101110101",
  36406=>"011101101",
  36407=>"100100001",
  36408=>"111100101",
  36409=>"100101010",
  36410=>"011000010",
  36411=>"000010111",
  36412=>"001100010",
  36413=>"110001000",
  36414=>"010000101",
  36415=>"101100100",
  36416=>"001100101",
  36417=>"100001011",
  36418=>"000010100",
  36419=>"100111001",
  36420=>"010100101",
  36421=>"110110110",
  36422=>"010101001",
  36423=>"110111110",
  36424=>"000101010",
  36425=>"100111101",
  36426=>"001001001",
  36427=>"010001101",
  36428=>"111110101",
  36429=>"101000000",
  36430=>"010100000",
  36431=>"001000000",
  36432=>"011111100",
  36433=>"001101101",
  36434=>"010100001",
  36435=>"110100000",
  36436=>"010001110",
  36437=>"011011001",
  36438=>"010011010",
  36439=>"111010101",
  36440=>"110101100",
  36441=>"001111010",
  36442=>"101011001",
  36443=>"111011011",
  36444=>"100001101",
  36445=>"101010100",
  36446=>"100100101",
  36447=>"111101101",
  36448=>"100010110",
  36449=>"010111111",
  36450=>"100110000",
  36451=>"101101001",
  36452=>"101110010",
  36453=>"000011010",
  36454=>"011011110",
  36455=>"100100010",
  36456=>"001101001",
  36457=>"010000100",
  36458=>"101111101",
  36459=>"111100111",
  36460=>"000001110",
  36461=>"000011111",
  36462=>"110101111",
  36463=>"111001000",
  36464=>"111110000",
  36465=>"100010000",
  36466=>"010000110",
  36467=>"110110100",
  36468=>"011011000",
  36469=>"101011000",
  36470=>"001010110",
  36471=>"011011100",
  36472=>"110001001",
  36473=>"101011001",
  36474=>"111010101",
  36475=>"001110101",
  36476=>"000011101",
  36477=>"001010100",
  36478=>"111000011",
  36479=>"000010111",
  36480=>"110000010",
  36481=>"100000111",
  36482=>"110101111",
  36483=>"100100000",
  36484=>"011100100",
  36485=>"011110111",
  36486=>"111010010",
  36487=>"011100110",
  36488=>"110010001",
  36489=>"110100001",
  36490=>"011010100",
  36491=>"101100100",
  36492=>"111110111",
  36493=>"100000100",
  36494=>"101111101",
  36495=>"000001001",
  36496=>"011110011",
  36497=>"110111101",
  36498=>"100001110",
  36499=>"011000011",
  36500=>"001000001",
  36501=>"110001011",
  36502=>"111000101",
  36503=>"001011110",
  36504=>"000000111",
  36505=>"111110110",
  36506=>"100100010",
  36507=>"100111011",
  36508=>"110010110",
  36509=>"001101110",
  36510=>"101110011",
  36511=>"100110000",
  36512=>"101000111",
  36513=>"110001001",
  36514=>"110000010",
  36515=>"101111100",
  36516=>"110111010",
  36517=>"110001101",
  36518=>"111001110",
  36519=>"000111100",
  36520=>"100111001",
  36521=>"110101011",
  36522=>"011100000",
  36523=>"101011111",
  36524=>"011011100",
  36525=>"010001010",
  36526=>"111011101",
  36527=>"011000010",
  36528=>"000100011",
  36529=>"011100000",
  36530=>"010000100",
  36531=>"011000111",
  36532=>"001111001",
  36533=>"110010111",
  36534=>"100000011",
  36535=>"001110100",
  36536=>"010001111",
  36537=>"101101000",
  36538=>"000111000",
  36539=>"110010111",
  36540=>"100001101",
  36541=>"001100101",
  36542=>"001000110",
  36543=>"001100011",
  36544=>"100111110",
  36545=>"110111101",
  36546=>"001001101",
  36547=>"110110000",
  36548=>"010010001",
  36549=>"100001111",
  36550=>"100011011",
  36551=>"101101101",
  36552=>"101000101",
  36553=>"111111111",
  36554=>"000110111",
  36555=>"001011001",
  36556=>"101111011",
  36557=>"100011110",
  36558=>"000000011",
  36559=>"000110101",
  36560=>"100101000",
  36561=>"101100110",
  36562=>"111010110",
  36563=>"111001101",
  36564=>"100001011",
  36565=>"000010000",
  36566=>"000110101",
  36567=>"010001000",
  36568=>"011111001",
  36569=>"100110100",
  36570=>"100110101",
  36571=>"110110011",
  36572=>"010001011",
  36573=>"101110110",
  36574=>"000111000",
  36575=>"001011010",
  36576=>"100001000",
  36577=>"000010111",
  36578=>"000100110",
  36579=>"100101011",
  36580=>"000010111",
  36581=>"000000001",
  36582=>"011000001",
  36583=>"010101010",
  36584=>"010011111",
  36585=>"011011110",
  36586=>"001101001",
  36587=>"111000000",
  36588=>"000010101",
  36589=>"010101110",
  36590=>"000010110",
  36591=>"010010001",
  36592=>"100011111",
  36593=>"000000001",
  36594=>"101101100",
  36595=>"111101100",
  36596=>"111011010",
  36597=>"001001010",
  36598=>"111111111",
  36599=>"011010010",
  36600=>"000001101",
  36601=>"101100111",
  36602=>"000111101",
  36603=>"000010010",
  36604=>"010100000",
  36605=>"011010110",
  36606=>"100001010",
  36607=>"101100100",
  36608=>"011100100",
  36609=>"010011100",
  36610=>"111111001",
  36611=>"001101001",
  36612=>"110110111",
  36613=>"001101100",
  36614=>"011011110",
  36615=>"101110110",
  36616=>"110000011",
  36617=>"000011111",
  36618=>"111001111",
  36619=>"001001011",
  36620=>"111010101",
  36621=>"101100000",
  36622=>"101000011",
  36623=>"110100111",
  36624=>"100000110",
  36625=>"010010010",
  36626=>"110011010",
  36627=>"100101111",
  36628=>"000110111",
  36629=>"000110100",
  36630=>"111100010",
  36631=>"111110010",
  36632=>"110111001",
  36633=>"111001001",
  36634=>"001000100",
  36635=>"011111010",
  36636=>"100010001",
  36637=>"000001110",
  36638=>"011011000",
  36639=>"001001111",
  36640=>"000010011",
  36641=>"011010101",
  36642=>"010111101",
  36643=>"011000001",
  36644=>"100101110",
  36645=>"011100000",
  36646=>"110100110",
  36647=>"100001010",
  36648=>"000111010",
  36649=>"110011101",
  36650=>"111101111",
  36651=>"000100111",
  36652=>"100101100",
  36653=>"000011100",
  36654=>"111110000",
  36655=>"101011001",
  36656=>"010001110",
  36657=>"111001001",
  36658=>"001110011",
  36659=>"000111010",
  36660=>"111100110",
  36661=>"010001010",
  36662=>"000100101",
  36663=>"101010111",
  36664=>"100100000",
  36665=>"000010010",
  36666=>"000000100",
  36667=>"001011110",
  36668=>"011000010",
  36669=>"111110111",
  36670=>"100010100",
  36671=>"010110100",
  36672=>"011011111",
  36673=>"110010001",
  36674=>"100110110",
  36675=>"000000011",
  36676=>"100100000",
  36677=>"000010010",
  36678=>"001000111",
  36679=>"111111011",
  36680=>"010100110",
  36681=>"011000010",
  36682=>"110101011",
  36683=>"000111000",
  36684=>"101101010",
  36685=>"000111001",
  36686=>"011110111",
  36687=>"111101010",
  36688=>"101110111",
  36689=>"100100000",
  36690=>"000011000",
  36691=>"000000111",
  36692=>"000010111",
  36693=>"001101111",
  36694=>"111111101",
  36695=>"010110000",
  36696=>"110001111",
  36697=>"110111001",
  36698=>"101101001",
  36699=>"111111011",
  36700=>"010010001",
  36701=>"001101100",
  36702=>"100011111",
  36703=>"111010100",
  36704=>"000100101",
  36705=>"111100000",
  36706=>"100010111",
  36707=>"000010101",
  36708=>"011101001",
  36709=>"110001111",
  36710=>"101010101",
  36711=>"000101010",
  36712=>"000101100",
  36713=>"000010011",
  36714=>"000110000",
  36715=>"110110011",
  36716=>"111010101",
  36717=>"101110101",
  36718=>"011111010",
  36719=>"011000110",
  36720=>"100101111",
  36721=>"110001010",
  36722=>"111001000",
  36723=>"001010100",
  36724=>"000010100",
  36725=>"010010010",
  36726=>"101111111",
  36727=>"000111111",
  36728=>"000000101",
  36729=>"100011010",
  36730=>"001110011",
  36731=>"111110000",
  36732=>"000010100",
  36733=>"000000001",
  36734=>"011001101",
  36735=>"101110011",
  36736=>"110011011",
  36737=>"100111011",
  36738=>"101010010",
  36739=>"011100011",
  36740=>"111001110",
  36741=>"111111010",
  36742=>"010110111",
  36743=>"110000101",
  36744=>"001110000",
  36745=>"101101100",
  36746=>"110110111",
  36747=>"111000111",
  36748=>"011010001",
  36749=>"101010001",
  36750=>"000000000",
  36751=>"111001110",
  36752=>"011011101",
  36753=>"011001110",
  36754=>"010010001",
  36755=>"000100111",
  36756=>"100001000",
  36757=>"000001111",
  36758=>"101101101",
  36759=>"001000101",
  36760=>"110111010",
  36761=>"000110010",
  36762=>"111110110",
  36763=>"000010011",
  36764=>"001000011",
  36765=>"111100000",
  36766=>"111001101",
  36767=>"111101011",
  36768=>"100001010",
  36769=>"100100100",
  36770=>"110000110",
  36771=>"011100010",
  36772=>"100110010",
  36773=>"011100001",
  36774=>"000101111",
  36775=>"111011011",
  36776=>"000101111",
  36777=>"110101000",
  36778=>"110011001",
  36779=>"101111110",
  36780=>"001010101",
  36781=>"001011001",
  36782=>"111001011",
  36783=>"010010100",
  36784=>"010001010",
  36785=>"001111100",
  36786=>"101010111",
  36787=>"111111011",
  36788=>"001101011",
  36789=>"111000111",
  36790=>"001100110",
  36791=>"100100000",
  36792=>"100001101",
  36793=>"000001100",
  36794=>"000010011",
  36795=>"010000100",
  36796=>"001101011",
  36797=>"111001101",
  36798=>"010110100",
  36799=>"010111110",
  36800=>"010110110",
  36801=>"110011010",
  36802=>"010110011",
  36803=>"110000110",
  36804=>"110001001",
  36805=>"010001011",
  36806=>"010010000",
  36807=>"001010100",
  36808=>"101010100",
  36809=>"000100101",
  36810=>"111101111",
  36811=>"011100111",
  36812=>"001000110",
  36813=>"111111011",
  36814=>"110011010",
  36815=>"001001001",
  36816=>"001101111",
  36817=>"010011101",
  36818=>"100101100",
  36819=>"000110111",
  36820=>"101110111",
  36821=>"111100000",
  36822=>"001000100",
  36823=>"110111100",
  36824=>"101101111",
  36825=>"111011111",
  36826=>"000011000",
  36827=>"011010000",
  36828=>"110110011",
  36829=>"111111011",
  36830=>"101000111",
  36831=>"010000111",
  36832=>"100111010",
  36833=>"110010111",
  36834=>"010010001",
  36835=>"101101011",
  36836=>"101011100",
  36837=>"100111011",
  36838=>"101010010",
  36839=>"011000110",
  36840=>"001101111",
  36841=>"110010010",
  36842=>"001000001",
  36843=>"111100010",
  36844=>"111001000",
  36845=>"110000011",
  36846=>"111101011",
  36847=>"011010001",
  36848=>"110111111",
  36849=>"000010000",
  36850=>"100110110",
  36851=>"100000111",
  36852=>"011011000",
  36853=>"001101101",
  36854=>"010000011",
  36855=>"000011111",
  36856=>"001011101",
  36857=>"100001100",
  36858=>"111100001",
  36859=>"000111111",
  36860=>"011001001",
  36861=>"100100110",
  36862=>"111001110",
  36863=>"011110111",
  36864=>"000001000",
  36865=>"110110000",
  36866=>"011110010",
  36867=>"100110101",
  36868=>"011101101",
  36869=>"101011011",
  36870=>"100101101",
  36871=>"110010000",
  36872=>"000101100",
  36873=>"000010000",
  36874=>"001110011",
  36875=>"010101111",
  36876=>"100011110",
  36877=>"101000101",
  36878=>"101111001",
  36879=>"100111110",
  36880=>"000010011",
  36881=>"011010101",
  36882=>"100001110",
  36883=>"100010000",
  36884=>"110011000",
  36885=>"011010010",
  36886=>"011000110",
  36887=>"010001011",
  36888=>"010011110",
  36889=>"111001000",
  36890=>"001101111",
  36891=>"110010110",
  36892=>"001001001",
  36893=>"100010000",
  36894=>"011111110",
  36895=>"001101000",
  36896=>"110100110",
  36897=>"110010011",
  36898=>"101000110",
  36899=>"111010101",
  36900=>"000111101",
  36901=>"101000001",
  36902=>"010100101",
  36903=>"110100110",
  36904=>"101011001",
  36905=>"001100100",
  36906=>"010100010",
  36907=>"010000100",
  36908=>"111011000",
  36909=>"100101101",
  36910=>"101010001",
  36911=>"101010100",
  36912=>"011100100",
  36913=>"011010011",
  36914=>"100001001",
  36915=>"101110001",
  36916=>"010100010",
  36917=>"000011111",
  36918=>"010100101",
  36919=>"111111010",
  36920=>"000100010",
  36921=>"100000000",
  36922=>"111010000",
  36923=>"001001110",
  36924=>"000110101",
  36925=>"110001111",
  36926=>"100001011",
  36927=>"111101111",
  36928=>"000001110",
  36929=>"001001000",
  36930=>"100110000",
  36931=>"001010001",
  36932=>"100110101",
  36933=>"100110001",
  36934=>"010001000",
  36935=>"111110101",
  36936=>"101111111",
  36937=>"110000101",
  36938=>"110111111",
  36939=>"000000000",
  36940=>"011111001",
  36941=>"110001000",
  36942=>"011010000",
  36943=>"101101110",
  36944=>"100010100",
  36945=>"111111111",
  36946=>"001011111",
  36947=>"011000101",
  36948=>"100011011",
  36949=>"010101101",
  36950=>"000010100",
  36951=>"001001010",
  36952=>"001101000",
  36953=>"110001100",
  36954=>"001001101",
  36955=>"111111001",
  36956=>"111100000",
  36957=>"000101100",
  36958=>"000001000",
  36959=>"001100101",
  36960=>"011111111",
  36961=>"100110001",
  36962=>"111110111",
  36963=>"000111101",
  36964=>"100110110",
  36965=>"110110000",
  36966=>"100001001",
  36967=>"001111101",
  36968=>"011010000",
  36969=>"111001011",
  36970=>"111010110",
  36971=>"100100000",
  36972=>"110101011",
  36973=>"110100010",
  36974=>"001100010",
  36975=>"101111010",
  36976=>"111110011",
  36977=>"011101010",
  36978=>"000110111",
  36979=>"100101010",
  36980=>"111101110",
  36981=>"110000001",
  36982=>"001111010",
  36983=>"100101110",
  36984=>"111101100",
  36985=>"000011001",
  36986=>"011001011",
  36987=>"011101010",
  36988=>"111000101",
  36989=>"010011101",
  36990=>"010000110",
  36991=>"110010010",
  36992=>"100110100",
  36993=>"010000011",
  36994=>"000100000",
  36995=>"011100000",
  36996=>"001010000",
  36997=>"001111001",
  36998=>"010101011",
  36999=>"101001100",
  37000=>"001000011",
  37001=>"110100010",
  37002=>"100100001",
  37003=>"010100011",
  37004=>"010010001",
  37005=>"010111011",
  37006=>"011011000",
  37007=>"111011010",
  37008=>"101000101",
  37009=>"111011000",
  37010=>"000010111",
  37011=>"111101111",
  37012=>"100101111",
  37013=>"111111011",
  37014=>"011010010",
  37015=>"101100001",
  37016=>"100001010",
  37017=>"100111011",
  37018=>"101101111",
  37019=>"000101111",
  37020=>"110011100",
  37021=>"111101000",
  37022=>"011010000",
  37023=>"111001010",
  37024=>"000000001",
  37025=>"000000000",
  37026=>"001110011",
  37027=>"101100011",
  37028=>"101100000",
  37029=>"111101111",
  37030=>"001000110",
  37031=>"000000101",
  37032=>"100010100",
  37033=>"111100000",
  37034=>"000110001",
  37035=>"101011000",
  37036=>"011111101",
  37037=>"101111110",
  37038=>"011101001",
  37039=>"011101010",
  37040=>"000111110",
  37041=>"101000101",
  37042=>"001001101",
  37043=>"011010110",
  37044=>"101100101",
  37045=>"101000011",
  37046=>"101110010",
  37047=>"101110010",
  37048=>"011001000",
  37049=>"001000110",
  37050=>"001010100",
  37051=>"110001011",
  37052=>"110010010",
  37053=>"111101101",
  37054=>"000000000",
  37055=>"111111110",
  37056=>"000111011",
  37057=>"010110011",
  37058=>"000111110",
  37059=>"010001101",
  37060=>"111010110",
  37061=>"011101111",
  37062=>"110110000",
  37063=>"100101100",
  37064=>"011011001",
  37065=>"100110001",
  37066=>"100100001",
  37067=>"111011000",
  37068=>"101001111",
  37069=>"011001000",
  37070=>"100100100",
  37071=>"000110100",
  37072=>"100010100",
  37073=>"101011011",
  37074=>"000100100",
  37075=>"011100101",
  37076=>"100000001",
  37077=>"000000011",
  37078=>"101011111",
  37079=>"100000110",
  37080=>"111110010",
  37081=>"101010010",
  37082=>"001000100",
  37083=>"010010110",
  37084=>"000010110",
  37085=>"011010010",
  37086=>"010110000",
  37087=>"101101101",
  37088=>"100100110",
  37089=>"011001100",
  37090=>"101111100",
  37091=>"010010001",
  37092=>"101101011",
  37093=>"101000111",
  37094=>"100111001",
  37095=>"110100011",
  37096=>"111111111",
  37097=>"111100100",
  37098=>"110101110",
  37099=>"101100001",
  37100=>"110111000",
  37101=>"010111101",
  37102=>"001100101",
  37103=>"001100110",
  37104=>"100110101",
  37105=>"000001000",
  37106=>"010001110",
  37107=>"111110100",
  37108=>"001110000",
  37109=>"110000100",
  37110=>"100110101",
  37111=>"101001101",
  37112=>"001000001",
  37113=>"101010001",
  37114=>"100000001",
  37115=>"001101001",
  37116=>"100110101",
  37117=>"110000111",
  37118=>"111010000",
  37119=>"110100110",
  37120=>"000111000",
  37121=>"111011001",
  37122=>"100101100",
  37123=>"000001101",
  37124=>"001001000",
  37125=>"011100011",
  37126=>"010001011",
  37127=>"111000010",
  37128=>"100000000",
  37129=>"000100000",
  37130=>"101100001",
  37131=>"110100011",
  37132=>"011011010",
  37133=>"010111000",
  37134=>"110101010",
  37135=>"101000010",
  37136=>"000011101",
  37137=>"110111010",
  37138=>"010000010",
  37139=>"100000010",
  37140=>"011101101",
  37141=>"100111101",
  37142=>"101001000",
  37143=>"001101011",
  37144=>"010101100",
  37145=>"011000010",
  37146=>"110010000",
  37147=>"111100111",
  37148=>"111010111",
  37149=>"100100011",
  37150=>"010110111",
  37151=>"110001101",
  37152=>"010111000",
  37153=>"100111011",
  37154=>"000111001",
  37155=>"101101100",
  37156=>"111101101",
  37157=>"101110100",
  37158=>"010000101",
  37159=>"011010111",
  37160=>"101100011",
  37161=>"110001100",
  37162=>"010100111",
  37163=>"110100101",
  37164=>"101011101",
  37165=>"101101111",
  37166=>"111101110",
  37167=>"100111001",
  37168=>"101110100",
  37169=>"000100010",
  37170=>"000001010",
  37171=>"001101100",
  37172=>"111011010",
  37173=>"011000100",
  37174=>"100001000",
  37175=>"110011000",
  37176=>"111001100",
  37177=>"011011110",
  37178=>"100111000",
  37179=>"000001001",
  37180=>"010001111",
  37181=>"110101100",
  37182=>"111011100",
  37183=>"000011010",
  37184=>"011111010",
  37185=>"100001011",
  37186=>"001000111",
  37187=>"011101001",
  37188=>"000001110",
  37189=>"100000101",
  37190=>"100100000",
  37191=>"010101100",
  37192=>"010000110",
  37193=>"101001100",
  37194=>"011111111",
  37195=>"000100001",
  37196=>"010010001",
  37197=>"101001010",
  37198=>"001001001",
  37199=>"001101110",
  37200=>"011011000",
  37201=>"000111011",
  37202=>"101010111",
  37203=>"000110010",
  37204=>"011000001",
  37205=>"111101101",
  37206=>"000110000",
  37207=>"010111010",
  37208=>"000000100",
  37209=>"101100011",
  37210=>"010001010",
  37211=>"010011111",
  37212=>"010010000",
  37213=>"111011011",
  37214=>"000001111",
  37215=>"001011100",
  37216=>"111010001",
  37217=>"101001010",
  37218=>"011000000",
  37219=>"100011101",
  37220=>"001011110",
  37221=>"100011000",
  37222=>"000000100",
  37223=>"000100001",
  37224=>"001010000",
  37225=>"100100111",
  37226=>"101111110",
  37227=>"110110000",
  37228=>"110110101",
  37229=>"011110000",
  37230=>"000100010",
  37231=>"001110001",
  37232=>"011001010",
  37233=>"001110000",
  37234=>"110001110",
  37235=>"001111101",
  37236=>"111001011",
  37237=>"001101011",
  37238=>"000001000",
  37239=>"000110010",
  37240=>"011100100",
  37241=>"011110101",
  37242=>"001101001",
  37243=>"010010001",
  37244=>"000101000",
  37245=>"111101100",
  37246=>"101010100",
  37247=>"010000011",
  37248=>"100010010",
  37249=>"000001000",
  37250=>"001000110",
  37251=>"110011100",
  37252=>"111100111",
  37253=>"111000111",
  37254=>"010110100",
  37255=>"111110100",
  37256=>"001011011",
  37257=>"110010000",
  37258=>"001111100",
  37259=>"000001011",
  37260=>"000011011",
  37261=>"110000000",
  37262=>"101101001",
  37263=>"101011100",
  37264=>"100001110",
  37265=>"010111001",
  37266=>"000000100",
  37267=>"000111101",
  37268=>"010100000",
  37269=>"011110110",
  37270=>"111111011",
  37271=>"100111010",
  37272=>"101100100",
  37273=>"110101111",
  37274=>"101001011",
  37275=>"000011010",
  37276=>"000101011",
  37277=>"001101001",
  37278=>"011110001",
  37279=>"101110110",
  37280=>"110111011",
  37281=>"000001011",
  37282=>"010000100",
  37283=>"111111101",
  37284=>"111101001",
  37285=>"001101010",
  37286=>"111110000",
  37287=>"000001111",
  37288=>"010000011",
  37289=>"001110111",
  37290=>"100011001",
  37291=>"010000010",
  37292=>"110110010",
  37293=>"101111111",
  37294=>"001101011",
  37295=>"100011011",
  37296=>"100110001",
  37297=>"001001100",
  37298=>"001001001",
  37299=>"011011011",
  37300=>"101011110",
  37301=>"101110100",
  37302=>"101011111",
  37303=>"111001010",
  37304=>"010111011",
  37305=>"001100101",
  37306=>"010011000",
  37307=>"001111010",
  37308=>"100011010",
  37309=>"011001110",
  37310=>"101111101",
  37311=>"101110000",
  37312=>"001100000",
  37313=>"110001111",
  37314=>"100010000",
  37315=>"011100100",
  37316=>"010001110",
  37317=>"000001000",
  37318=>"010000000",
  37319=>"110011000",
  37320=>"000111001",
  37321=>"110011000",
  37322=>"010100011",
  37323=>"000100100",
  37324=>"101010001",
  37325=>"010011010",
  37326=>"011010101",
  37327=>"001011111",
  37328=>"001100010",
  37329=>"001011000",
  37330=>"111010101",
  37331=>"000100101",
  37332=>"100111111",
  37333=>"111100100",
  37334=>"101001101",
  37335=>"001100001",
  37336=>"010000001",
  37337=>"100110001",
  37338=>"111110011",
  37339=>"001001000",
  37340=>"110100010",
  37341=>"000010100",
  37342=>"011001000",
  37343=>"011010010",
  37344=>"110000000",
  37345=>"100100110",
  37346=>"101100000",
  37347=>"110011010",
  37348=>"101111001",
  37349=>"011101011",
  37350=>"110000001",
  37351=>"010011100",
  37352=>"010011110",
  37353=>"011010011",
  37354=>"111010101",
  37355=>"100101110",
  37356=>"101101000",
  37357=>"111100010",
  37358=>"111011001",
  37359=>"100010001",
  37360=>"101011110",
  37361=>"001010101",
  37362=>"010010110",
  37363=>"101000001",
  37364=>"011010101",
  37365=>"100101110",
  37366=>"000100000",
  37367=>"111101000",
  37368=>"010010001",
  37369=>"001011011",
  37370=>"101010111",
  37371=>"001111010",
  37372=>"101110010",
  37373=>"001010110",
  37374=>"001111110",
  37375=>"100110100",
  37376=>"011111001",
  37377=>"110110001",
  37378=>"001110101",
  37379=>"100110100",
  37380=>"100010111",
  37381=>"110011010",
  37382=>"011000011",
  37383=>"110000110",
  37384=>"100111011",
  37385=>"110101001",
  37386=>"011001011",
  37387=>"001000100",
  37388=>"001101110",
  37389=>"010001100",
  37390=>"011010100",
  37391=>"000011110",
  37392=>"111101001",
  37393=>"010011011",
  37394=>"110111010",
  37395=>"010011011",
  37396=>"011101011",
  37397=>"110110011",
  37398=>"111001110",
  37399=>"010100110",
  37400=>"001111110",
  37401=>"000100100",
  37402=>"010011000",
  37403=>"001100110",
  37404=>"111011010",
  37405=>"110100000",
  37406=>"111100110",
  37407=>"110101111",
  37408=>"011000001",
  37409=>"001110011",
  37410=>"001100111",
  37411=>"110011100",
  37412=>"011011001",
  37413=>"110001001",
  37414=>"111110010",
  37415=>"111010100",
  37416=>"001001111",
  37417=>"010000101",
  37418=>"101100100",
  37419=>"110101100",
  37420=>"001000001",
  37421=>"101101001",
  37422=>"110110011",
  37423=>"000000101",
  37424=>"001111010",
  37425=>"000001010",
  37426=>"101001001",
  37427=>"000111101",
  37428=>"110100100",
  37429=>"010110010",
  37430=>"001001000",
  37431=>"000010111",
  37432=>"010000111",
  37433=>"100011111",
  37434=>"110101011",
  37435=>"100101110",
  37436=>"001100010",
  37437=>"111101000",
  37438=>"101000101",
  37439=>"110100101",
  37440=>"110101111",
  37441=>"111110110",
  37442=>"110000001",
  37443=>"111000000",
  37444=>"100001111",
  37445=>"000000101",
  37446=>"111000111",
  37447=>"111101111",
  37448=>"111010100",
  37449=>"001111011",
  37450=>"100101000",
  37451=>"111010000",
  37452=>"000101000",
  37453=>"001110010",
  37454=>"010010000",
  37455=>"100111011",
  37456=>"111110100",
  37457=>"111011010",
  37458=>"101111100",
  37459=>"000011010",
  37460=>"101100001",
  37461=>"011101111",
  37462=>"010001001",
  37463=>"011100001",
  37464=>"011011010",
  37465=>"011101001",
  37466=>"000001111",
  37467=>"100001010",
  37468=>"001001011",
  37469=>"110100101",
  37470=>"001001010",
  37471=>"110000010",
  37472=>"010010000",
  37473=>"000010011",
  37474=>"000100110",
  37475=>"001101101",
  37476=>"110000010",
  37477=>"001101110",
  37478=>"111011000",
  37479=>"110001000",
  37480=>"110010010",
  37481=>"100001001",
  37482=>"001000110",
  37483=>"000110101",
  37484=>"100000000",
  37485=>"111010010",
  37486=>"001010111",
  37487=>"101001000",
  37488=>"100101000",
  37489=>"000100110",
  37490=>"001110100",
  37491=>"111111101",
  37492=>"110101000",
  37493=>"110110100",
  37494=>"111001011",
  37495=>"010011110",
  37496=>"011000011",
  37497=>"101101000",
  37498=>"110010001",
  37499=>"010101101",
  37500=>"110101101",
  37501=>"111111110",
  37502=>"101001101",
  37503=>"010110001",
  37504=>"000010101",
  37505=>"010110011",
  37506=>"101101000",
  37507=>"000100000",
  37508=>"001110101",
  37509=>"011100000",
  37510=>"111001011",
  37511=>"100000010",
  37512=>"100010010",
  37513=>"111100101",
  37514=>"010010110",
  37515=>"100111001",
  37516=>"110111010",
  37517=>"000000100",
  37518=>"000111111",
  37519=>"010001101",
  37520=>"000011101",
  37521=>"000100010",
  37522=>"111001000",
  37523=>"010100011",
  37524=>"001011011",
  37525=>"111101110",
  37526=>"001000001",
  37527=>"110001100",
  37528=>"110111000",
  37529=>"001110010",
  37530=>"111000110",
  37531=>"011101110",
  37532=>"001110001",
  37533=>"101000011",
  37534=>"000001001",
  37535=>"111001111",
  37536=>"001100110",
  37537=>"111001001",
  37538=>"100011110",
  37539=>"110000111",
  37540=>"010001101",
  37541=>"010010000",
  37542=>"000010110",
  37543=>"110111101",
  37544=>"111000001",
  37545=>"000000111",
  37546=>"011010110",
  37547=>"010000110",
  37548=>"000100000",
  37549=>"010111001",
  37550=>"111000010",
  37551=>"100001000",
  37552=>"000100101",
  37553=>"100100010",
  37554=>"001011110",
  37555=>"001100101",
  37556=>"011100000",
  37557=>"001000011",
  37558=>"011011000",
  37559=>"000001000",
  37560=>"000110011",
  37561=>"111010100",
  37562=>"101110111",
  37563=>"111100000",
  37564=>"101011001",
  37565=>"010111000",
  37566=>"001111111",
  37567=>"011011000",
  37568=>"000010001",
  37569=>"110111111",
  37570=>"100110011",
  37571=>"101100001",
  37572=>"010011111",
  37573=>"110001011",
  37574=>"100111111",
  37575=>"110111111",
  37576=>"011100100",
  37577=>"110000110",
  37578=>"101111000",
  37579=>"010110000",
  37580=>"001110101",
  37581=>"000000000",
  37582=>"011100100",
  37583=>"101111001",
  37584=>"000001100",
  37585=>"011100010",
  37586=>"111010001",
  37587=>"001101001",
  37588=>"101000110",
  37589=>"100011010",
  37590=>"010100111",
  37591=>"011011101",
  37592=>"011011101",
  37593=>"000100101",
  37594=>"011000110",
  37595=>"100100011",
  37596=>"010100111",
  37597=>"111000001",
  37598=>"100111010",
  37599=>"011000000",
  37600=>"111010100",
  37601=>"000011111",
  37602=>"111101110",
  37603=>"000110011",
  37604=>"011100111",
  37605=>"010100000",
  37606=>"001100111",
  37607=>"111000001",
  37608=>"000000001",
  37609=>"111100110",
  37610=>"110100010",
  37611=>"100000011",
  37612=>"110100101",
  37613=>"000111110",
  37614=>"111001100",
  37615=>"101111000",
  37616=>"111001111",
  37617=>"010000000",
  37618=>"111010000",
  37619=>"010111010",
  37620=>"001100011",
  37621=>"010100011",
  37622=>"001011100",
  37623=>"111110111",
  37624=>"100011100",
  37625=>"110101011",
  37626=>"101101110",
  37627=>"100101100",
  37628=>"111011110",
  37629=>"011110100",
  37630=>"000101010",
  37631=>"011111010",
  37632=>"001011001",
  37633=>"001100100",
  37634=>"110011100",
  37635=>"010000001",
  37636=>"000110101",
  37637=>"101000000",
  37638=>"111011001",
  37639=>"100110001",
  37640=>"000011011",
  37641=>"111110100",
  37642=>"011000100",
  37643=>"101101110",
  37644=>"000101111",
  37645=>"011110101",
  37646=>"011001110",
  37647=>"100101110",
  37648=>"110111011",
  37649=>"111011101",
  37650=>"101110111",
  37651=>"010010000",
  37652=>"111100010",
  37653=>"101101110",
  37654=>"100001110",
  37655=>"110111100",
  37656=>"011110000",
  37657=>"110011001",
  37658=>"000010111",
  37659=>"110111011",
  37660=>"110100011",
  37661=>"100100000",
  37662=>"101110100",
  37663=>"111010011",
  37664=>"100001111",
  37665=>"100000010",
  37666=>"111000110",
  37667=>"100100111",
  37668=>"000010001",
  37669=>"011001010",
  37670=>"001001110",
  37671=>"111001100",
  37672=>"011001100",
  37673=>"101110000",
  37674=>"010011000",
  37675=>"101000000",
  37676=>"001110101",
  37677=>"110010001",
  37678=>"000100000",
  37679=>"011111111",
  37680=>"101101111",
  37681=>"011000010",
  37682=>"001110000",
  37683=>"011100000",
  37684=>"001101100",
  37685=>"100010001",
  37686=>"010011000",
  37687=>"010110111",
  37688=>"101110101",
  37689=>"010110011",
  37690=>"110001101",
  37691=>"011101001",
  37692=>"010010111",
  37693=>"101001110",
  37694=>"110110001",
  37695=>"111001010",
  37696=>"100111100",
  37697=>"000101000",
  37698=>"011001100",
  37699=>"110000000",
  37700=>"111001110",
  37701=>"010100100",
  37702=>"101010011",
  37703=>"000111100",
  37704=>"111101001",
  37705=>"010000100",
  37706=>"010000000",
  37707=>"000010101",
  37708=>"011010000",
  37709=>"100100010",
  37710=>"011011110",
  37711=>"011101010",
  37712=>"110110111",
  37713=>"110110100",
  37714=>"001101011",
  37715=>"111100001",
  37716=>"111000000",
  37717=>"010001001",
  37718=>"111110100",
  37719=>"011000100",
  37720=>"001010100",
  37721=>"000000011",
  37722=>"010111010",
  37723=>"110001110",
  37724=>"010101101",
  37725=>"001110110",
  37726=>"100111001",
  37727=>"000000100",
  37728=>"100101011",
  37729=>"010000000",
  37730=>"010111000",
  37731=>"010001100",
  37732=>"101111000",
  37733=>"111000110",
  37734=>"100000111",
  37735=>"010001101",
  37736=>"001001101",
  37737=>"001011000",
  37738=>"001111100",
  37739=>"111000011",
  37740=>"100101110",
  37741=>"001101001",
  37742=>"001111011",
  37743=>"100011110",
  37744=>"100010101",
  37745=>"110100010",
  37746=>"001011001",
  37747=>"001001011",
  37748=>"110011100",
  37749=>"001010011",
  37750=>"000001101",
  37751=>"110100011",
  37752=>"001010010",
  37753=>"000001101",
  37754=>"000000101",
  37755=>"010001010",
  37756=>"001111000",
  37757=>"001100000",
  37758=>"000101011",
  37759=>"000111101",
  37760=>"010010010",
  37761=>"010000110",
  37762=>"001000101",
  37763=>"000111000",
  37764=>"010001011",
  37765=>"001111010",
  37766=>"110111111",
  37767=>"010101101",
  37768=>"000001001",
  37769=>"010000110",
  37770=>"011100110",
  37771=>"000001110",
  37772=>"101010000",
  37773=>"011011101",
  37774=>"010101011",
  37775=>"001111101",
  37776=>"111010011",
  37777=>"111101111",
  37778=>"100100000",
  37779=>"111110001",
  37780=>"001101111",
  37781=>"011001000",
  37782=>"001111010",
  37783=>"010001001",
  37784=>"100100011",
  37785=>"011110110",
  37786=>"111101110",
  37787=>"111001111",
  37788=>"100010000",
  37789=>"111111111",
  37790=>"010101011",
  37791=>"111110001",
  37792=>"000001000",
  37793=>"111011100",
  37794=>"011111110",
  37795=>"110101011",
  37796=>"001111100",
  37797=>"011011011",
  37798=>"101001011",
  37799=>"001111111",
  37800=>"001100110",
  37801=>"000001000",
  37802=>"110011010",
  37803=>"101010011",
  37804=>"111100000",
  37805=>"101011000",
  37806=>"100101111",
  37807=>"000100101",
  37808=>"000100101",
  37809=>"000100110",
  37810=>"111010111",
  37811=>"011000001",
  37812=>"110001011",
  37813=>"010100100",
  37814=>"000101101",
  37815=>"011111001",
  37816=>"100000110",
  37817=>"001110000",
  37818=>"001100110",
  37819=>"100011101",
  37820=>"001110101",
  37821=>"100100100",
  37822=>"110000011",
  37823=>"000000101",
  37824=>"011100001",
  37825=>"010011111",
  37826=>"101100111",
  37827=>"111010011",
  37828=>"011010000",
  37829=>"111001010",
  37830=>"111011110",
  37831=>"000001101",
  37832=>"000001001",
  37833=>"001010010",
  37834=>"111001000",
  37835=>"001100110",
  37836=>"111111001",
  37837=>"000000001",
  37838=>"000000000",
  37839=>"001111010",
  37840=>"110010111",
  37841=>"011101000",
  37842=>"001011001",
  37843=>"100001111",
  37844=>"011111011",
  37845=>"010011010",
  37846=>"011111110",
  37847=>"101100000",
  37848=>"000110100",
  37849=>"101101000",
  37850=>"000010000",
  37851=>"100001101",
  37852=>"010101000",
  37853=>"111111001",
  37854=>"100100010",
  37855=>"010110001",
  37856=>"111010101",
  37857=>"001100101",
  37858=>"100001011",
  37859=>"110011000",
  37860=>"100011000",
  37861=>"100011000",
  37862=>"100000110",
  37863=>"010001111",
  37864=>"101010110",
  37865=>"000111000",
  37866=>"010010101",
  37867=>"000001000",
  37868=>"111110110",
  37869=>"000110000",
  37870=>"100001111",
  37871=>"010101110",
  37872=>"010001111",
  37873=>"100111101",
  37874=>"100110101",
  37875=>"000000010",
  37876=>"000110101",
  37877=>"000000011",
  37878=>"100011110",
  37879=>"001101100",
  37880=>"011000010",
  37881=>"001000010",
  37882=>"010010011",
  37883=>"001100110",
  37884=>"010001010",
  37885=>"101111101",
  37886=>"000111110",
  37887=>"010010010",
  37888=>"100110010",
  37889=>"111000001",
  37890=>"010111101",
  37891=>"111011001",
  37892=>"101110001",
  37893=>"111001110",
  37894=>"101000111",
  37895=>"111001001",
  37896=>"011011111",
  37897=>"010001010",
  37898=>"001001111",
  37899=>"110000100",
  37900=>"100001110",
  37901=>"111100100",
  37902=>"100011010",
  37903=>"010001011",
  37904=>"101111111",
  37905=>"000100110",
  37906=>"111111011",
  37907=>"111111010",
  37908=>"000001011",
  37909=>"100100101",
  37910=>"010010111",
  37911=>"100001110",
  37912=>"010011100",
  37913=>"000101011",
  37914=>"001101001",
  37915=>"110000010",
  37916=>"101001010",
  37917=>"001100100",
  37918=>"110100010",
  37919=>"111111111",
  37920=>"010000101",
  37921=>"101110001",
  37922=>"000100011",
  37923=>"100010101",
  37924=>"011111101",
  37925=>"011000010",
  37926=>"110100101",
  37927=>"110110011",
  37928=>"000111110",
  37929=>"101001111",
  37930=>"101101111",
  37931=>"010011111",
  37932=>"001111000",
  37933=>"101010111",
  37934=>"000101011",
  37935=>"100110110",
  37936=>"110011100",
  37937=>"010010110",
  37938=>"111010110",
  37939=>"011000100",
  37940=>"000100110",
  37941=>"001111001",
  37942=>"110111000",
  37943=>"110101100",
  37944=>"101100011",
  37945=>"000101011",
  37946=>"101111010",
  37947=>"000010101",
  37948=>"100100100",
  37949=>"110010000",
  37950=>"010010011",
  37951=>"010110011",
  37952=>"000101100",
  37953=>"000000110",
  37954=>"100011001",
  37955=>"010101111",
  37956=>"111101011",
  37957=>"001110101",
  37958=>"000011001",
  37959=>"001011101",
  37960=>"100011011",
  37961=>"011000001",
  37962=>"110101110",
  37963=>"000110001",
  37964=>"111011011",
  37965=>"111011110",
  37966=>"001000000",
  37967=>"101100111",
  37968=>"000000100",
  37969=>"110010001",
  37970=>"111110000",
  37971=>"001000110",
  37972=>"011101111",
  37973=>"011100111",
  37974=>"001001000",
  37975=>"001010111",
  37976=>"000010100",
  37977=>"001000110",
  37978=>"101010110",
  37979=>"000110000",
  37980=>"010011010",
  37981=>"010110111",
  37982=>"000101001",
  37983=>"101100010",
  37984=>"000110111",
  37985=>"111010111",
  37986=>"110101000",
  37987=>"000110101",
  37988=>"101101000",
  37989=>"100010100",
  37990=>"101100011",
  37991=>"000011111",
  37992=>"000110000",
  37993=>"001111011",
  37994=>"011101011",
  37995=>"100000011",
  37996=>"100100010",
  37997=>"010011010",
  37998=>"100010000",
  37999=>"000010001",
  38000=>"110010000",
  38001=>"000110111",
  38002=>"001100011",
  38003=>"111011001",
  38004=>"001101010",
  38005=>"000000101",
  38006=>"000011101",
  38007=>"101010000",
  38008=>"011100000",
  38009=>"101010111",
  38010=>"010010010",
  38011=>"000001011",
  38012=>"110001110",
  38013=>"111111101",
  38014=>"001001000",
  38015=>"011111010",
  38016=>"111000110",
  38017=>"010010010",
  38018=>"010010011",
  38019=>"101110100",
  38020=>"100111001",
  38021=>"000010110",
  38022=>"111110000",
  38023=>"110110001",
  38024=>"111110111",
  38025=>"110010101",
  38026=>"010010011",
  38027=>"010111101",
  38028=>"101000001",
  38029=>"100000101",
  38030=>"100110000",
  38031=>"011001001",
  38032=>"110010101",
  38033=>"111011100",
  38034=>"101000001",
  38035=>"000010111",
  38036=>"000010101",
  38037=>"110111110",
  38038=>"100010100",
  38039=>"011100001",
  38040=>"100110010",
  38041=>"100001011",
  38042=>"011010010",
  38043=>"011011011",
  38044=>"010011011",
  38045=>"001100000",
  38046=>"011011111",
  38047=>"100111101",
  38048=>"110110001",
  38049=>"110111100",
  38050=>"000001010",
  38051=>"010111101",
  38052=>"001001001",
  38053=>"011100001",
  38054=>"111011111",
  38055=>"111111100",
  38056=>"010101101",
  38057=>"101101000",
  38058=>"111100001",
  38059=>"111101001",
  38060=>"010011001",
  38061=>"000001101",
  38062=>"101101001",
  38063=>"001000010",
  38064=>"110111010",
  38065=>"100100010",
  38066=>"000100011",
  38067=>"000000010",
  38068=>"001000011",
  38069=>"000100101",
  38070=>"011111011",
  38071=>"101101100",
  38072=>"001000100",
  38073=>"001101101",
  38074=>"010000000",
  38075=>"001001110",
  38076=>"100000101",
  38077=>"011101010",
  38078=>"011111101",
  38079=>"110111001",
  38080=>"010000101",
  38081=>"100110000",
  38082=>"100010110",
  38083=>"010000001",
  38084=>"000010110",
  38085=>"111111111",
  38086=>"001010100",
  38087=>"000101100",
  38088=>"101100011",
  38089=>"000100011",
  38090=>"111111111",
  38091=>"110101110",
  38092=>"100100100",
  38093=>"001111110",
  38094=>"001110000",
  38095=>"110000001",
  38096=>"010111111",
  38097=>"011100101",
  38098=>"100010100",
  38099=>"001001110",
  38100=>"101010001",
  38101=>"011010101",
  38102=>"001000100",
  38103=>"010001111",
  38104=>"110100001",
  38105=>"010000110",
  38106=>"001000100",
  38107=>"111011000",
  38108=>"010010001",
  38109=>"001100110",
  38110=>"111000000",
  38111=>"000011111",
  38112=>"100100000",
  38113=>"010100010",
  38114=>"110111000",
  38115=>"000010001",
  38116=>"001001011",
  38117=>"000110110",
  38118=>"110101011",
  38119=>"011000111",
  38120=>"111111101",
  38121=>"010000111",
  38122=>"011111111",
  38123=>"100000000",
  38124=>"001111011",
  38125=>"110011110",
  38126=>"010001011",
  38127=>"000100000",
  38128=>"111110101",
  38129=>"110110010",
  38130=>"100110111",
  38131=>"100010001",
  38132=>"011001100",
  38133=>"000001111",
  38134=>"010100110",
  38135=>"111000111",
  38136=>"001111001",
  38137=>"111000010",
  38138=>"111011101",
  38139=>"001100101",
  38140=>"001001111",
  38141=>"001100100",
  38142=>"000100001",
  38143=>"000110011",
  38144=>"011011101",
  38145=>"011010111",
  38146=>"001010000",
  38147=>"110111100",
  38148=>"010100111",
  38149=>"000010110",
  38150=>"001110110",
  38151=>"000110101",
  38152=>"011110001",
  38153=>"101111101",
  38154=>"111010001",
  38155=>"101001010",
  38156=>"000011011",
  38157=>"110110111",
  38158=>"110110010",
  38159=>"000010111",
  38160=>"111010111",
  38161=>"100110101",
  38162=>"111011101",
  38163=>"010110000",
  38164=>"111011001",
  38165=>"100100011",
  38166=>"101001001",
  38167=>"011101001",
  38168=>"010010001",
  38169=>"110000010",
  38170=>"010100110",
  38171=>"111010011",
  38172=>"100001110",
  38173=>"001000100",
  38174=>"111011110",
  38175=>"000110111",
  38176=>"100000001",
  38177=>"101011110",
  38178=>"001001001",
  38179=>"100001100",
  38180=>"111011011",
  38181=>"100101110",
  38182=>"101010100",
  38183=>"101110111",
  38184=>"110011110",
  38185=>"010100110",
  38186=>"110001110",
  38187=>"000110011",
  38188=>"010001111",
  38189=>"010001000",
  38190=>"001000001",
  38191=>"101010100",
  38192=>"110010000",
  38193=>"011111100",
  38194=>"110101110",
  38195=>"000100111",
  38196=>"010101111",
  38197=>"111111100",
  38198=>"011101111",
  38199=>"000011000",
  38200=>"110101100",
  38201=>"010000010",
  38202=>"110110101",
  38203=>"100001010",
  38204=>"101100011",
  38205=>"000101111",
  38206=>"011010000",
  38207=>"001001110",
  38208=>"100000000",
  38209=>"001000001",
  38210=>"100111101",
  38211=>"101001000",
  38212=>"010000111",
  38213=>"000011011",
  38214=>"101100010",
  38215=>"011001100",
  38216=>"110011001",
  38217=>"000101110",
  38218=>"101111011",
  38219=>"011000001",
  38220=>"110011001",
  38221=>"101100111",
  38222=>"011110010",
  38223=>"001011000",
  38224=>"011011101",
  38225=>"101100010",
  38226=>"101010110",
  38227=>"000010111",
  38228=>"101111100",
  38229=>"001001111",
  38230=>"010101011",
  38231=>"000100101",
  38232=>"111100101",
  38233=>"001001110",
  38234=>"111000111",
  38235=>"101100010",
  38236=>"011101111",
  38237=>"001011010",
  38238=>"111111001",
  38239=>"100000111",
  38240=>"010110111",
  38241=>"011011101",
  38242=>"001101010",
  38243=>"001001000",
  38244=>"000010001",
  38245=>"011000011",
  38246=>"000011011",
  38247=>"011101010",
  38248=>"010010001",
  38249=>"000011111",
  38250=>"010000110",
  38251=>"010100000",
  38252=>"110011010",
  38253=>"010100000",
  38254=>"000010101",
  38255=>"111101000",
  38256=>"000111011",
  38257=>"110100111",
  38258=>"100101001",
  38259=>"101100100",
  38260=>"100110111",
  38261=>"001100011",
  38262=>"111100001",
  38263=>"111110001",
  38264=>"111111011",
  38265=>"001110101",
  38266=>"111011100",
  38267=>"010000110",
  38268=>"100110000",
  38269=>"100110001",
  38270=>"100101001",
  38271=>"100000000",
  38272=>"001111001",
  38273=>"101001111",
  38274=>"000100001",
  38275=>"101110111",
  38276=>"001100000",
  38277=>"100010111",
  38278=>"011111101",
  38279=>"111110110",
  38280=>"100000011",
  38281=>"111011111",
  38282=>"110011101",
  38283=>"100101001",
  38284=>"000001111",
  38285=>"110010011",
  38286=>"011001100",
  38287=>"010111010",
  38288=>"010110111",
  38289=>"101100111",
  38290=>"000000001",
  38291=>"001010000",
  38292=>"000000001",
  38293=>"011001100",
  38294=>"110111011",
  38295=>"101110100",
  38296=>"000011100",
  38297=>"001101010",
  38298=>"000111100",
  38299=>"000000100",
  38300=>"110100100",
  38301=>"000000111",
  38302=>"000110000",
  38303=>"101101010",
  38304=>"110110000",
  38305=>"000011000",
  38306=>"100000010",
  38307=>"111001000",
  38308=>"111111100",
  38309=>"100001101",
  38310=>"101000010",
  38311=>"000001111",
  38312=>"111100011",
  38313=>"010010111",
  38314=>"000011101",
  38315=>"101011000",
  38316=>"000011010",
  38317=>"001110010",
  38318=>"100110101",
  38319=>"100110110",
  38320=>"101100101",
  38321=>"110100100",
  38322=>"010010010",
  38323=>"001011000",
  38324=>"011000101",
  38325=>"100011011",
  38326=>"100101111",
  38327=>"101100111",
  38328=>"100110111",
  38329=>"000111010",
  38330=>"001010011",
  38331=>"000000010",
  38332=>"010000000",
  38333=>"001001010",
  38334=>"011100010",
  38335=>"010111010",
  38336=>"100100010",
  38337=>"000010011",
  38338=>"010101110",
  38339=>"011111000",
  38340=>"010011100",
  38341=>"000100110",
  38342=>"111110000",
  38343=>"111100010",
  38344=>"110011100",
  38345=>"100110010",
  38346=>"100011110",
  38347=>"110011111",
  38348=>"000101001",
  38349=>"110101011",
  38350=>"000111100",
  38351=>"111111100",
  38352=>"110101001",
  38353=>"100000110",
  38354=>"100001111",
  38355=>"110101000",
  38356=>"000100111",
  38357=>"001000001",
  38358=>"010111000",
  38359=>"010111111",
  38360=>"011110110",
  38361=>"101000111",
  38362=>"000001111",
  38363=>"010111001",
  38364=>"011001101",
  38365=>"101111111",
  38366=>"011100110",
  38367=>"010000111",
  38368=>"100001110",
  38369=>"100111011",
  38370=>"111100010",
  38371=>"101001000",
  38372=>"000010100",
  38373=>"001110111",
  38374=>"101110000",
  38375=>"110111110",
  38376=>"000100100",
  38377=>"111100001",
  38378=>"010100111",
  38379=>"011100010",
  38380=>"111111101",
  38381=>"110100100",
  38382=>"010110000",
  38383=>"100011111",
  38384=>"001101001",
  38385=>"100001001",
  38386=>"110010001",
  38387=>"011100101",
  38388=>"001011000",
  38389=>"100000101",
  38390=>"011001100",
  38391=>"010111011",
  38392=>"011011100",
  38393=>"100010010",
  38394=>"010010001",
  38395=>"110011100",
  38396=>"010001010",
  38397=>"001000111",
  38398=>"010001111",
  38399=>"001111111",
  38400=>"111110110",
  38401=>"010111101",
  38402=>"110101000",
  38403=>"111100100",
  38404=>"111010000",
  38405=>"010100101",
  38406=>"010001000",
  38407=>"100110111",
  38408=>"001010110",
  38409=>"000110001",
  38410=>"101110001",
  38411=>"000001011",
  38412=>"000000001",
  38413=>"001100100",
  38414=>"111000111",
  38415=>"101100100",
  38416=>"000000000",
  38417=>"011001000",
  38418=>"100110111",
  38419=>"001011001",
  38420=>"110000101",
  38421=>"110000010",
  38422=>"110111001",
  38423=>"001100000",
  38424=>"101111101",
  38425=>"011001111",
  38426=>"100001110",
  38427=>"100010000",
  38428=>"101100101",
  38429=>"010101000",
  38430=>"100010001",
  38431=>"100000110",
  38432=>"011110100",
  38433=>"011011001",
  38434=>"000010111",
  38435=>"111010110",
  38436=>"000100110",
  38437=>"000010101",
  38438=>"011110110",
  38439=>"111110111",
  38440=>"100111011",
  38441=>"001010001",
  38442=>"101100100",
  38443=>"101101010",
  38444=>"100011000",
  38445=>"000011011",
  38446=>"111110000",
  38447=>"100100010",
  38448=>"111101011",
  38449=>"100011100",
  38450=>"011001000",
  38451=>"101001111",
  38452=>"011111011",
  38453=>"010111000",
  38454=>"011010110",
  38455=>"011011011",
  38456=>"000100110",
  38457=>"110101000",
  38458=>"000111000",
  38459=>"000100011",
  38460=>"010000000",
  38461=>"011001111",
  38462=>"101001010",
  38463=>"111001000",
  38464=>"111010001",
  38465=>"000100000",
  38466=>"110100001",
  38467=>"010010100",
  38468=>"010111100",
  38469=>"111010100",
  38470=>"001101111",
  38471=>"001000011",
  38472=>"010001111",
  38473=>"000101100",
  38474=>"111000001",
  38475=>"011010001",
  38476=>"000101000",
  38477=>"100011110",
  38478=>"101111000",
  38479=>"101011000",
  38480=>"101111111",
  38481=>"111111000",
  38482=>"110001100",
  38483=>"110000000",
  38484=>"110000111",
  38485=>"000011111",
  38486=>"000001110",
  38487=>"111111101",
  38488=>"111011110",
  38489=>"001000110",
  38490=>"001001000",
  38491=>"000100101",
  38492=>"001010010",
  38493=>"000011001",
  38494=>"010011111",
  38495=>"000110110",
  38496=>"000101001",
  38497=>"101000110",
  38498=>"011010011",
  38499=>"111011011",
  38500=>"100011110",
  38501=>"100111101",
  38502=>"011110110",
  38503=>"011001111",
  38504=>"001100110",
  38505=>"110011101",
  38506=>"110110111",
  38507=>"000010010",
  38508=>"000101100",
  38509=>"101000010",
  38510=>"110001101",
  38511=>"101010100",
  38512=>"011111011",
  38513=>"001100100",
  38514=>"101100111",
  38515=>"101111101",
  38516=>"010010010",
  38517=>"010001111",
  38518=>"110101110",
  38519=>"101101001",
  38520=>"011100000",
  38521=>"110111011",
  38522=>"101001000",
  38523=>"000010110",
  38524=>"110110100",
  38525=>"001001000",
  38526=>"101100101",
  38527=>"110110001",
  38528=>"111100101",
  38529=>"100100101",
  38530=>"101001000",
  38531=>"001010111",
  38532=>"001110010",
  38533=>"000101110",
  38534=>"110011111",
  38535=>"001110101",
  38536=>"100011010",
  38537=>"111101011",
  38538=>"001001100",
  38539=>"111010001",
  38540=>"000010001",
  38541=>"110010111",
  38542=>"111100010",
  38543=>"000000110",
  38544=>"010110100",
  38545=>"011100011",
  38546=>"001110011",
  38547=>"010010111",
  38548=>"001011001",
  38549=>"100001011",
  38550=>"011110100",
  38551=>"010100100",
  38552=>"111001110",
  38553=>"111100110",
  38554=>"010110110",
  38555=>"011000000",
  38556=>"111001011",
  38557=>"101110001",
  38558=>"011000110",
  38559=>"001101010",
  38560=>"011111010",
  38561=>"110010001",
  38562=>"110000011",
  38563=>"111111011",
  38564=>"100010000",
  38565=>"100000110",
  38566=>"101100011",
  38567=>"100100101",
  38568=>"000001001",
  38569=>"111111001",
  38570=>"101001111",
  38571=>"111110100",
  38572=>"000010001",
  38573=>"011110110",
  38574=>"111000010",
  38575=>"110111001",
  38576=>"010001011",
  38577=>"000100100",
  38578=>"010001110",
  38579=>"011000000",
  38580=>"000010110",
  38581=>"101100010",
  38582=>"111011100",
  38583=>"001000110",
  38584=>"101010110",
  38585=>"011001011",
  38586=>"010100001",
  38587=>"010000010",
  38588=>"001100100",
  38589=>"111010100",
  38590=>"000010101",
  38591=>"011010011",
  38592=>"110111100",
  38593=>"110000100",
  38594=>"000001100",
  38595=>"010011011",
  38596=>"101110000",
  38597=>"001001100",
  38598=>"101011010",
  38599=>"000110110",
  38600=>"111001011",
  38601=>"110001100",
  38602=>"111010011",
  38603=>"000101010",
  38604=>"101001101",
  38605=>"001100000",
  38606=>"111000100",
  38607=>"001100111",
  38608=>"011010000",
  38609=>"101100110",
  38610=>"101101010",
  38611=>"101010010",
  38612=>"101101000",
  38613=>"100011011",
  38614=>"001000010",
  38615=>"001111111",
  38616=>"100000110",
  38617=>"011010111",
  38618=>"000010001",
  38619=>"011001110",
  38620=>"101011010",
  38621=>"010110110",
  38622=>"111111011",
  38623=>"000100011",
  38624=>"110011001",
  38625=>"111110010",
  38626=>"101010000",
  38627=>"110011111",
  38628=>"001001011",
  38629=>"011101000",
  38630=>"000110111",
  38631=>"101010011",
  38632=>"000111111",
  38633=>"000010111",
  38634=>"101100000",
  38635=>"111111010",
  38636=>"001000001",
  38637=>"100101101",
  38638=>"100111111",
  38639=>"000000011",
  38640=>"010000011",
  38641=>"101110101",
  38642=>"101001000",
  38643=>"101110111",
  38644=>"000100011",
  38645=>"000010011",
  38646=>"100100100",
  38647=>"011111110",
  38648=>"111100000",
  38649=>"110011000",
  38650=>"110101111",
  38651=>"110110000",
  38652=>"111001000",
  38653=>"111100101",
  38654=>"111110100",
  38655=>"110010010",
  38656=>"100110011",
  38657=>"111101111",
  38658=>"101001101",
  38659=>"101100010",
  38660=>"100001010",
  38661=>"101000000",
  38662=>"010111001",
  38663=>"011101111",
  38664=>"111111100",
  38665=>"111111001",
  38666=>"100100000",
  38667=>"100011101",
  38668=>"111100011",
  38669=>"110111100",
  38670=>"110000001",
  38671=>"000010011",
  38672=>"101010000",
  38673=>"011011001",
  38674=>"100110110",
  38675=>"011111011",
  38676=>"100111111",
  38677=>"001010111",
  38678=>"001011110",
  38679=>"011110000",
  38680=>"111110101",
  38681=>"110111101",
  38682=>"000001000",
  38683=>"001101101",
  38684=>"101100010",
  38685=>"010110101",
  38686=>"110001101",
  38687=>"111011001",
  38688=>"011100111",
  38689=>"001010001",
  38690=>"001110000",
  38691=>"000111011",
  38692=>"011011111",
  38693=>"110010101",
  38694=>"000100100",
  38695=>"111111000",
  38696=>"000000001",
  38697=>"101000100",
  38698=>"101011011",
  38699=>"111101000",
  38700=>"000011010",
  38701=>"001001001",
  38702=>"100010000",
  38703=>"110100000",
  38704=>"001010000",
  38705=>"100000110",
  38706=>"101100000",
  38707=>"011010001",
  38708=>"101101111",
  38709=>"001000000",
  38710=>"000001000",
  38711=>"001011010",
  38712=>"001010000",
  38713=>"001010001",
  38714=>"001100000",
  38715=>"001010001",
  38716=>"000110011",
  38717=>"100111001",
  38718=>"110101111",
  38719=>"011000001",
  38720=>"011010001",
  38721=>"000011010",
  38722=>"110010010",
  38723=>"001000000",
  38724=>"110001101",
  38725=>"011111110",
  38726=>"010100011",
  38727=>"110001101",
  38728=>"010101110",
  38729=>"000010000",
  38730=>"001000000",
  38731=>"001001001",
  38732=>"110011001",
  38733=>"011100001",
  38734=>"110010011",
  38735=>"111111110",
  38736=>"100010010",
  38737=>"101011100",
  38738=>"100000011",
  38739=>"111001100",
  38740=>"111011001",
  38741=>"011100110",
  38742=>"110101000",
  38743=>"010001001",
  38744=>"001101111",
  38745=>"011100101",
  38746=>"110010101",
  38747=>"111110011",
  38748=>"011110000",
  38749=>"001110011",
  38750=>"110001010",
  38751=>"010010011",
  38752=>"010010111",
  38753=>"011000000",
  38754=>"001111001",
  38755=>"111100110",
  38756=>"001000001",
  38757=>"000101000",
  38758=>"011001110",
  38759=>"011000011",
  38760=>"110011000",
  38761=>"110011000",
  38762=>"111101100",
  38763=>"111011001",
  38764=>"011010010",
  38765=>"111110101",
  38766=>"101110010",
  38767=>"001000101",
  38768=>"000000101",
  38769=>"000110010",
  38770=>"101011110",
  38771=>"010101000",
  38772=>"010010110",
  38773=>"000011000",
  38774=>"101011001",
  38775=>"000010000",
  38776=>"101001011",
  38777=>"100000011",
  38778=>"111010110",
  38779=>"000101001",
  38780=>"001100011",
  38781=>"010101101",
  38782=>"101010110",
  38783=>"111001001",
  38784=>"100111100",
  38785=>"001000000",
  38786=>"011111111",
  38787=>"101010001",
  38788=>"000110101",
  38789=>"100011100",
  38790=>"011010011",
  38791=>"001010000",
  38792=>"100101100",
  38793=>"110100100",
  38794=>"000111010",
  38795=>"001100110",
  38796=>"110110010",
  38797=>"111010011",
  38798=>"010010100",
  38799=>"011001100",
  38800=>"110011110",
  38801=>"111101000",
  38802=>"100000111",
  38803=>"111001000",
  38804=>"101111110",
  38805=>"111110011",
  38806=>"011111111",
  38807=>"010110000",
  38808=>"001010011",
  38809=>"111101111",
  38810=>"100111100",
  38811=>"111110100",
  38812=>"001111101",
  38813=>"001110110",
  38814=>"100100100",
  38815=>"110110010",
  38816=>"110010110",
  38817=>"111010110",
  38818=>"110000001",
  38819=>"110100001",
  38820=>"010111001",
  38821=>"111011111",
  38822=>"100010010",
  38823=>"010000100",
  38824=>"110010111",
  38825=>"100110110",
  38826=>"001001110",
  38827=>"000010101",
  38828=>"111000100",
  38829=>"001100111",
  38830=>"000110010",
  38831=>"000001010",
  38832=>"001011100",
  38833=>"111100111",
  38834=>"011000110",
  38835=>"111010100",
  38836=>"101011101",
  38837=>"000101001",
  38838=>"000111010",
  38839=>"010000010",
  38840=>"001110010",
  38841=>"110100110",
  38842=>"001111000",
  38843=>"101010011",
  38844=>"010110100",
  38845=>"010000011",
  38846=>"101110001",
  38847=>"101010001",
  38848=>"101011111",
  38849=>"101100111",
  38850=>"101110001",
  38851=>"111001011",
  38852=>"010011011",
  38853=>"001101101",
  38854=>"011001000",
  38855=>"110001101",
  38856=>"000001100",
  38857=>"100111111",
  38858=>"011000111",
  38859=>"111110100",
  38860=>"111011110",
  38861=>"000010001",
  38862=>"000001011",
  38863=>"111011111",
  38864=>"000101000",
  38865=>"110111010",
  38866=>"000110111",
  38867=>"011101011",
  38868=>"110111001",
  38869=>"000011100",
  38870=>"010001101",
  38871=>"000000001",
  38872=>"000000010",
  38873=>"101011011",
  38874=>"101010000",
  38875=>"011100000",
  38876=>"001100011",
  38877=>"010011000",
  38878=>"100000000",
  38879=>"000100100",
  38880=>"100111101",
  38881=>"001011001",
  38882=>"010110110",
  38883=>"000101111",
  38884=>"111100100",
  38885=>"100001111",
  38886=>"101111000",
  38887=>"011100100",
  38888=>"111100100",
  38889=>"101000111",
  38890=>"000100110",
  38891=>"100100111",
  38892=>"000100100",
  38893=>"100010101",
  38894=>"100000010",
  38895=>"111100110",
  38896=>"000101111",
  38897=>"011100110",
  38898=>"011000000",
  38899=>"000001010",
  38900=>"111111000",
  38901=>"011100011",
  38902=>"010111111",
  38903=>"111110111",
  38904=>"011011111",
  38905=>"010110110",
  38906=>"111000111",
  38907=>"101110110",
  38908=>"011110110",
  38909=>"101110110",
  38910=>"011000111",
  38911=>"001000101",
  38912=>"010001001",
  38913=>"011000110",
  38914=>"010110011",
  38915=>"011010000",
  38916=>"001100111",
  38917=>"100001010",
  38918=>"100010011",
  38919=>"000100010",
  38920=>"111011000",
  38921=>"010111100",
  38922=>"100101101",
  38923=>"111001011",
  38924=>"000001011",
  38925=>"101001000",
  38926=>"111110001",
  38927=>"000011011",
  38928=>"101101001",
  38929=>"000100110",
  38930=>"000111000",
  38931=>"010010100",
  38932=>"010001001",
  38933=>"111000111",
  38934=>"100000000",
  38935=>"000000110",
  38936=>"101110001",
  38937=>"001001101",
  38938=>"110011010",
  38939=>"101011101",
  38940=>"111101100",
  38941=>"010011100",
  38942=>"001000111",
  38943=>"000101100",
  38944=>"100110000",
  38945=>"110011001",
  38946=>"010101111",
  38947=>"111110001",
  38948=>"000101101",
  38949=>"010001111",
  38950=>"101000101",
  38951=>"101100110",
  38952=>"111010001",
  38953=>"010111010",
  38954=>"110010000",
  38955=>"000111001",
  38956=>"111011100",
  38957=>"110111100",
  38958=>"011110100",
  38959=>"100000101",
  38960=>"010111101",
  38961=>"001101111",
  38962=>"110101011",
  38963=>"101001011",
  38964=>"001101001",
  38965=>"011100000",
  38966=>"111001000",
  38967=>"000001000",
  38968=>"100111110",
  38969=>"010101100",
  38970=>"000001000",
  38971=>"000001111",
  38972=>"001010111",
  38973=>"111100010",
  38974=>"100110011",
  38975=>"100001111",
  38976=>"111000000",
  38977=>"000110010",
  38978=>"011111000",
  38979=>"100001000",
  38980=>"111111100",
  38981=>"110110011",
  38982=>"010111011",
  38983=>"110010011",
  38984=>"111001001",
  38985=>"100110010",
  38986=>"100000100",
  38987=>"001010010",
  38988=>"000000111",
  38989=>"010011101",
  38990=>"111000100",
  38991=>"011100100",
  38992=>"100100101",
  38993=>"010010110",
  38994=>"011001011",
  38995=>"000000110",
  38996=>"110000011",
  38997=>"111101001",
  38998=>"001010010",
  38999=>"000000001",
  39000=>"111100100",
  39001=>"010001100",
  39002=>"101001001",
  39003=>"000001000",
  39004=>"100100010",
  39005=>"001100001",
  39006=>"000000101",
  39007=>"011100101",
  39008=>"011101100",
  39009=>"111011000",
  39010=>"000011011",
  39011=>"000010111",
  39012=>"001010100",
  39013=>"110100011",
  39014=>"111110110",
  39015=>"000101011",
  39016=>"110011111",
  39017=>"111100001",
  39018=>"000000111",
  39019=>"100110101",
  39020=>"011000100",
  39021=>"011001101",
  39022=>"011001111",
  39023=>"100110000",
  39024=>"110001000",
  39025=>"101100010",
  39026=>"000110000",
  39027=>"110010001",
  39028=>"000001000",
  39029=>"011010000",
  39030=>"100010100",
  39031=>"001011000",
  39032=>"000001001",
  39033=>"110110010",
  39034=>"000110011",
  39035=>"001100000",
  39036=>"100110111",
  39037=>"110001011",
  39038=>"100010001",
  39039=>"100001111",
  39040=>"111010110",
  39041=>"110001110",
  39042=>"001001010",
  39043=>"110011101",
  39044=>"000011100",
  39045=>"001101010",
  39046=>"011101111",
  39047=>"100110010",
  39048=>"100111011",
  39049=>"011000011",
  39050=>"100010110",
  39051=>"010111111",
  39052=>"000001000",
  39053=>"111111000",
  39054=>"100010011",
  39055=>"100101101",
  39056=>"010110000",
  39057=>"110000100",
  39058=>"111010100",
  39059=>"011000000",
  39060=>"100101100",
  39061=>"001100010",
  39062=>"000010011",
  39063=>"101111110",
  39064=>"101000011",
  39065=>"100101010",
  39066=>"000010100",
  39067=>"101111001",
  39068=>"001011010",
  39069=>"101000101",
  39070=>"101110000",
  39071=>"110100001",
  39072=>"100100110",
  39073=>"111111100",
  39074=>"000110101",
  39075=>"110101001",
  39076=>"100110101",
  39077=>"010111011",
  39078=>"111110100",
  39079=>"011011011",
  39080=>"100111100",
  39081=>"110011101",
  39082=>"010011000",
  39083=>"011110111",
  39084=>"101011010",
  39085=>"000110101",
  39086=>"100000100",
  39087=>"001110010",
  39088=>"001000011",
  39089=>"010001000",
  39090=>"101111100",
  39091=>"100100011",
  39092=>"101010001",
  39093=>"100001100",
  39094=>"000111010",
  39095=>"110010111",
  39096=>"101000001",
  39097=>"100011000",
  39098=>"000110110",
  39099=>"000101101",
  39100=>"100010011",
  39101=>"001010001",
  39102=>"001001010",
  39103=>"110000010",
  39104=>"100101110",
  39105=>"111111011",
  39106=>"000010011",
  39107=>"010001011",
  39108=>"100111010",
  39109=>"110011010",
  39110=>"000001010",
  39111=>"001101101",
  39112=>"111100011",
  39113=>"101011110",
  39114=>"100100111",
  39115=>"011101000",
  39116=>"110000011",
  39117=>"100011001",
  39118=>"111011111",
  39119=>"111000000",
  39120=>"110000100",
  39121=>"001011110",
  39122=>"110000000",
  39123=>"111001010",
  39124=>"111011010",
  39125=>"110010010",
  39126=>"001110011",
  39127=>"000001111",
  39128=>"111001000",
  39129=>"000110101",
  39130=>"011110000",
  39131=>"011000111",
  39132=>"100011000",
  39133=>"001000000",
  39134=>"010110001",
  39135=>"100110111",
  39136=>"010000001",
  39137=>"000110101",
  39138=>"010110001",
  39139=>"000010101",
  39140=>"110111111",
  39141=>"000100001",
  39142=>"000011000",
  39143=>"110011010",
  39144=>"001110101",
  39145=>"001010000",
  39146=>"100010100",
  39147=>"011111001",
  39148=>"100010001",
  39149=>"000000011",
  39150=>"001000000",
  39151=>"010110001",
  39152=>"000001010",
  39153=>"011000001",
  39154=>"110011011",
  39155=>"111101100",
  39156=>"111111101",
  39157=>"110111101",
  39158=>"110000100",
  39159=>"001010010",
  39160=>"101100110",
  39161=>"110101000",
  39162=>"100110000",
  39163=>"101000111",
  39164=>"000000000",
  39165=>"011000001",
  39166=>"111010111",
  39167=>"010100000",
  39168=>"001111110",
  39169=>"110010010",
  39170=>"100001100",
  39171=>"000000000",
  39172=>"010101111",
  39173=>"010011100",
  39174=>"010101000",
  39175=>"111100010",
  39176=>"001011101",
  39177=>"011101011",
  39178=>"110011111",
  39179=>"110011001",
  39180=>"010100100",
  39181=>"000001001",
  39182=>"100111101",
  39183=>"001001100",
  39184=>"110010000",
  39185=>"001100110",
  39186=>"100001010",
  39187=>"100100100",
  39188=>"000001101",
  39189=>"100011100",
  39190=>"101010010",
  39191=>"100101111",
  39192=>"011110010",
  39193=>"010010010",
  39194=>"011001110",
  39195=>"111011011",
  39196=>"010010101",
  39197=>"001000000",
  39198=>"101110111",
  39199=>"001110001",
  39200=>"001001110",
  39201=>"011010001",
  39202=>"000010110",
  39203=>"111101100",
  39204=>"101110011",
  39205=>"000110001",
  39206=>"111010101",
  39207=>"111100011",
  39208=>"100001000",
  39209=>"010000101",
  39210=>"000111101",
  39211=>"110001100",
  39212=>"111111110",
  39213=>"000001100",
  39214=>"001000001",
  39215=>"101110011",
  39216=>"010001100",
  39217=>"110101111",
  39218=>"010111110",
  39219=>"000001000",
  39220=>"100101101",
  39221=>"000000001",
  39222=>"011011011",
  39223=>"101011111",
  39224=>"001001010",
  39225=>"000010110",
  39226=>"001000111",
  39227=>"100010001",
  39228=>"111100011",
  39229=>"010101000",
  39230=>"100010100",
  39231=>"100101100",
  39232=>"101101111",
  39233=>"001111101",
  39234=>"010111111",
  39235=>"111111100",
  39236=>"011100001",
  39237=>"101001001",
  39238=>"100011110",
  39239=>"100110000",
  39240=>"101110000",
  39241=>"000101010",
  39242=>"110001101",
  39243=>"110000001",
  39244=>"011100011",
  39245=>"100101100",
  39246=>"111110110",
  39247=>"100001100",
  39248=>"001100110",
  39249=>"111011110",
  39250=>"011010000",
  39251=>"000001011",
  39252=>"010101000",
  39253=>"101001000",
  39254=>"111000000",
  39255=>"010101011",
  39256=>"010000011",
  39257=>"000011000",
  39258=>"000110110",
  39259=>"011001100",
  39260=>"011100000",
  39261=>"000011100",
  39262=>"111001101",
  39263=>"100101101",
  39264=>"100010011",
  39265=>"110011001",
  39266=>"110001000",
  39267=>"001100101",
  39268=>"010011001",
  39269=>"001001100",
  39270=>"001100010",
  39271=>"011000000",
  39272=>"111110110",
  39273=>"000111111",
  39274=>"011001111",
  39275=>"011111111",
  39276=>"101111001",
  39277=>"000100001",
  39278=>"100110100",
  39279=>"001111000",
  39280=>"010010000",
  39281=>"101001110",
  39282=>"001001001",
  39283=>"111011010",
  39284=>"100100011",
  39285=>"000000011",
  39286=>"010111101",
  39287=>"111001000",
  39288=>"100011000",
  39289=>"111111010",
  39290=>"100010001",
  39291=>"100001100",
  39292=>"000011010",
  39293=>"110010100",
  39294=>"010011000",
  39295=>"111100011",
  39296=>"000000010",
  39297=>"100011110",
  39298=>"110110001",
  39299=>"100000100",
  39300=>"110011001",
  39301=>"011001100",
  39302=>"000001010",
  39303=>"111001000",
  39304=>"010010001",
  39305=>"101110010",
  39306=>"001010110",
  39307=>"001010110",
  39308=>"010101100",
  39309=>"110011110",
  39310=>"011000000",
  39311=>"100100101",
  39312=>"110001111",
  39313=>"000010011",
  39314=>"001110010",
  39315=>"100110100",
  39316=>"110010001",
  39317=>"001001000",
  39318=>"010000100",
  39319=>"111110111",
  39320=>"100110111",
  39321=>"000001010",
  39322=>"010110101",
  39323=>"011111010",
  39324=>"110000101",
  39325=>"101110000",
  39326=>"001000000",
  39327=>"010111101",
  39328=>"011100101",
  39329=>"000011101",
  39330=>"110111101",
  39331=>"111000011",
  39332=>"000001001",
  39333=>"101110001",
  39334=>"100111001",
  39335=>"101100011",
  39336=>"101111011",
  39337=>"100010000",
  39338=>"000101000",
  39339=>"001111001",
  39340=>"000001010",
  39341=>"101011001",
  39342=>"011000100",
  39343=>"111100001",
  39344=>"100000000",
  39345=>"111100101",
  39346=>"101100110",
  39347=>"111011001",
  39348=>"011100101",
  39349=>"010110110",
  39350=>"000110001",
  39351=>"010111110",
  39352=>"000000100",
  39353=>"111001011",
  39354=>"001010000",
  39355=>"010010110",
  39356=>"011011111",
  39357=>"100111101",
  39358=>"010101011",
  39359=>"000000111",
  39360=>"000100001",
  39361=>"010101101",
  39362=>"101011111",
  39363=>"110011010",
  39364=>"010010000",
  39365=>"010001110",
  39366=>"010001111",
  39367=>"111110000",
  39368=>"011001101",
  39369=>"001100011",
  39370=>"110001101",
  39371=>"010011001",
  39372=>"000110010",
  39373=>"010100010",
  39374=>"001010000",
  39375=>"111101101",
  39376=>"100010111",
  39377=>"010000000",
  39378=>"001000110",
  39379=>"101001011",
  39380=>"001001100",
  39381=>"010111101",
  39382=>"111011101",
  39383=>"100011011",
  39384=>"011001110",
  39385=>"100110010",
  39386=>"010001000",
  39387=>"110111111",
  39388=>"011011101",
  39389=>"011010010",
  39390=>"011010100",
  39391=>"010111101",
  39392=>"101001100",
  39393=>"011111010",
  39394=>"110100101",
  39395=>"100010000",
  39396=>"100001110",
  39397=>"111111010",
  39398=>"010100010",
  39399=>"000100001",
  39400=>"100010110",
  39401=>"000011110",
  39402=>"010000010",
  39403=>"110001101",
  39404=>"010001011",
  39405=>"010111001",
  39406=>"100000111",
  39407=>"111001000",
  39408=>"001111101",
  39409=>"111111010",
  39410=>"101010010",
  39411=>"101101000",
  39412=>"001110000",
  39413=>"001001000",
  39414=>"100100000",
  39415=>"111001100",
  39416=>"001010100",
  39417=>"111010010",
  39418=>"000010111",
  39419=>"010100101",
  39420=>"001100010",
  39421=>"100111010",
  39422=>"110000100",
  39423=>"111110000",
  39424=>"110110111",
  39425=>"001011110",
  39426=>"100000111",
  39427=>"011000010",
  39428=>"100110110",
  39429=>"110110000",
  39430=>"110110100",
  39431=>"100011000",
  39432=>"110101100",
  39433=>"000001001",
  39434=>"110110001",
  39435=>"000110100",
  39436=>"100110010",
  39437=>"011101100",
  39438=>"111001000",
  39439=>"010011110",
  39440=>"110010010",
  39441=>"111010110",
  39442=>"000101001",
  39443=>"100011011",
  39444=>"010100110",
  39445=>"100100001",
  39446=>"010110100",
  39447=>"011110111",
  39448=>"001001101",
  39449=>"000100111",
  39450=>"010011001",
  39451=>"100100000",
  39452=>"111001000",
  39453=>"100001000",
  39454=>"011101000",
  39455=>"001001011",
  39456=>"001111101",
  39457=>"010011000",
  39458=>"000001010",
  39459=>"100000001",
  39460=>"001000011",
  39461=>"001000100",
  39462=>"100001011",
  39463=>"110000101",
  39464=>"011011100",
  39465=>"001011111",
  39466=>"010010100",
  39467=>"000001001",
  39468=>"100000111",
  39469=>"100000101",
  39470=>"100110111",
  39471=>"001000000",
  39472=>"110001110",
  39473=>"111101110",
  39474=>"101001001",
  39475=>"000101000",
  39476=>"000011010",
  39477=>"001101000",
  39478=>"111100110",
  39479=>"101001010",
  39480=>"010001001",
  39481=>"111111000",
  39482=>"001110000",
  39483=>"010011100",
  39484=>"110100001",
  39485=>"110000110",
  39486=>"000001011",
  39487=>"000101010",
  39488=>"111011011",
  39489=>"010110101",
  39490=>"111001111",
  39491=>"111101011",
  39492=>"111001011",
  39493=>"111001010",
  39494=>"101101110",
  39495=>"101001001",
  39496=>"100000011",
  39497=>"011010010",
  39498=>"010100010",
  39499=>"001100000",
  39500=>"110010100",
  39501=>"001011000",
  39502=>"111011111",
  39503=>"101110100",
  39504=>"110011111",
  39505=>"110111011",
  39506=>"101101011",
  39507=>"101101000",
  39508=>"000000011",
  39509=>"000001111",
  39510=>"000011010",
  39511=>"100011011",
  39512=>"010101001",
  39513=>"111001101",
  39514=>"000001000",
  39515=>"000101001",
  39516=>"001111001",
  39517=>"010101010",
  39518=>"000000000",
  39519=>"011011001",
  39520=>"111101011",
  39521=>"001000100",
  39522=>"010110001",
  39523=>"000000100",
  39524=>"000011010",
  39525=>"110101011",
  39526=>"101010111",
  39527=>"101000101",
  39528=>"010000000",
  39529=>"011101110",
  39530=>"101100000",
  39531=>"011001110",
  39532=>"000100101",
  39533=>"110110101",
  39534=>"011011011",
  39535=>"000000101",
  39536=>"010001101",
  39537=>"000100110",
  39538=>"110010101",
  39539=>"001001000",
  39540=>"010100011",
  39541=>"100111111",
  39542=>"110100001",
  39543=>"001101101",
  39544=>"000101110",
  39545=>"110100010",
  39546=>"111001010",
  39547=>"111100110",
  39548=>"110001000",
  39549=>"101110011",
  39550=>"101110000",
  39551=>"100110111",
  39552=>"110110110",
  39553=>"110000100",
  39554=>"111101000",
  39555=>"010001011",
  39556=>"000111000",
  39557=>"010001001",
  39558=>"001111111",
  39559=>"101110111",
  39560=>"011001110",
  39561=>"010011000",
  39562=>"000100000",
  39563=>"010010001",
  39564=>"110011000",
  39565=>"101000110",
  39566=>"001000110",
  39567=>"110011110",
  39568=>"001101101",
  39569=>"001000101",
  39570=>"010010000",
  39571=>"001110010",
  39572=>"000101111",
  39573=>"000110011",
  39574=>"010010001",
  39575=>"110100101",
  39576=>"110111101",
  39577=>"100110100",
  39578=>"111101110",
  39579=>"001010100",
  39580=>"111011010",
  39581=>"111111100",
  39582=>"000001000",
  39583=>"001110010",
  39584=>"100011010",
  39585=>"110110001",
  39586=>"010110100",
  39587=>"000010000",
  39588=>"000001111",
  39589=>"000100001",
  39590=>"000110010",
  39591=>"000001110",
  39592=>"011110110",
  39593=>"011100001",
  39594=>"001111001",
  39595=>"000011011",
  39596=>"000100001",
  39597=>"001010100",
  39598=>"111011000",
  39599=>"010111011",
  39600=>"011100100",
  39601=>"000010000",
  39602=>"000110111",
  39603=>"011001001",
  39604=>"000001101",
  39605=>"011010111",
  39606=>"100110011",
  39607=>"010011110",
  39608=>"010111111",
  39609=>"100000100",
  39610=>"000011010",
  39611=>"101101000",
  39612=>"001110001",
  39613=>"010101000",
  39614=>"110010101",
  39615=>"110110111",
  39616=>"011101010",
  39617=>"101101101",
  39618=>"001111001",
  39619=>"001000000",
  39620=>"000011010",
  39621=>"110001001",
  39622=>"000110010",
  39623=>"011110101",
  39624=>"111111111",
  39625=>"101001000",
  39626=>"100001011",
  39627=>"000011000",
  39628=>"000000101",
  39629=>"111010010",
  39630=>"000001011",
  39631=>"011001011",
  39632=>"101001010",
  39633=>"000110111",
  39634=>"000100110",
  39635=>"001010001",
  39636=>"001110100",
  39637=>"001000100",
  39638=>"101101111",
  39639=>"101000011",
  39640=>"000011000",
  39641=>"111111101",
  39642=>"100100111",
  39643=>"110101110",
  39644=>"101101001",
  39645=>"110001111",
  39646=>"000100110",
  39647=>"011100011",
  39648=>"010001010",
  39649=>"100101111",
  39650=>"111010010",
  39651=>"010110000",
  39652=>"000001110",
  39653=>"110011111",
  39654=>"000101100",
  39655=>"111010100",
  39656=>"010000011",
  39657=>"011111110",
  39658=>"000101001",
  39659=>"111101010",
  39660=>"000111101",
  39661=>"100111011",
  39662=>"010010000",
  39663=>"101001001",
  39664=>"001110011",
  39665=>"100010111",
  39666=>"111000110",
  39667=>"101101111",
  39668=>"000011101",
  39669=>"110101010",
  39670=>"000100101",
  39671=>"111001100",
  39672=>"110010101",
  39673=>"001100011",
  39674=>"111101001",
  39675=>"100011101",
  39676=>"100011011",
  39677=>"101010100",
  39678=>"011101101",
  39679=>"001010010",
  39680=>"010100000",
  39681=>"001101001",
  39682=>"000111110",
  39683=>"000000100",
  39684=>"111011101",
  39685=>"000110010",
  39686=>"001100110",
  39687=>"100000100",
  39688=>"010001001",
  39689=>"000100010",
  39690=>"111100000",
  39691=>"100111011",
  39692=>"001110101",
  39693=>"101111111",
  39694=>"000010011",
  39695=>"101001011",
  39696=>"010100110",
  39697=>"101100100",
  39698=>"101101000",
  39699=>"011111001",
  39700=>"101101010",
  39701=>"111111100",
  39702=>"001011000",
  39703=>"000111101",
  39704=>"011100111",
  39705=>"000011010",
  39706=>"100011110",
  39707=>"011000111",
  39708=>"011000000",
  39709=>"001001110",
  39710=>"100000000",
  39711=>"110010010",
  39712=>"001100110",
  39713=>"111101010",
  39714=>"011110011",
  39715=>"000101010",
  39716=>"001001010",
  39717=>"111011010",
  39718=>"010100011",
  39719=>"010101111",
  39720=>"000001111",
  39721=>"111110011",
  39722=>"101011011",
  39723=>"110110001",
  39724=>"010110010",
  39725=>"000000000",
  39726=>"000100010",
  39727=>"010000111",
  39728=>"000111110",
  39729=>"000101001",
  39730=>"001001001",
  39731=>"111100100",
  39732=>"101110001",
  39733=>"110101101",
  39734=>"010011000",
  39735=>"101101001",
  39736=>"001000001",
  39737=>"111111110",
  39738=>"111101011",
  39739=>"101010010",
  39740=>"110000101",
  39741=>"001010010",
  39742=>"100110111",
  39743=>"001111010",
  39744=>"111101111",
  39745=>"101101111",
  39746=>"010010101",
  39747=>"011000011",
  39748=>"001101011",
  39749=>"111011110",
  39750=>"101101011",
  39751=>"001000101",
  39752=>"011010011",
  39753=>"001101111",
  39754=>"010101101",
  39755=>"101100011",
  39756=>"111100000",
  39757=>"001101001",
  39758=>"110010001",
  39759=>"110010000",
  39760=>"011011010",
  39761=>"110100110",
  39762=>"011100001",
  39763=>"100001011",
  39764=>"010011100",
  39765=>"101101000",
  39766=>"101111010",
  39767=>"111001110",
  39768=>"001101001",
  39769=>"010010100",
  39770=>"110100110",
  39771=>"101010101",
  39772=>"111101110",
  39773=>"001110011",
  39774=>"001001011",
  39775=>"000000000",
  39776=>"111110101",
  39777=>"111011000",
  39778=>"000100000",
  39779=>"010101000",
  39780=>"011011110",
  39781=>"000001001",
  39782=>"010010111",
  39783=>"011111111",
  39784=>"000010111",
  39785=>"001011111",
  39786=>"110011000",
  39787=>"010111101",
  39788=>"010111110",
  39789=>"010101101",
  39790=>"101100010",
  39791=>"010010110",
  39792=>"100011100",
  39793=>"111111010",
  39794=>"110101111",
  39795=>"000111100",
  39796=>"011111000",
  39797=>"001110111",
  39798=>"100001001",
  39799=>"110001100",
  39800=>"010101010",
  39801=>"110000001",
  39802=>"000001010",
  39803=>"100001010",
  39804=>"001000000",
  39805=>"011000001",
  39806=>"001000000",
  39807=>"100100100",
  39808=>"000101110",
  39809=>"010010111",
  39810=>"001000010",
  39811=>"101010001",
  39812=>"000000010",
  39813=>"100001011",
  39814=>"000111010",
  39815=>"101000001",
  39816=>"111111110",
  39817=>"111100011",
  39818=>"001010000",
  39819=>"001001110",
  39820=>"000000010",
  39821=>"110010000",
  39822=>"001110101",
  39823=>"010111100",
  39824=>"110000111",
  39825=>"011000010",
  39826=>"000110000",
  39827=>"001010001",
  39828=>"110011000",
  39829=>"011110011",
  39830=>"010010100",
  39831=>"000111111",
  39832=>"111100111",
  39833=>"111110100",
  39834=>"010001010",
  39835=>"001100101",
  39836=>"000010110",
  39837=>"110011011",
  39838=>"000011110",
  39839=>"000100000",
  39840=>"100101001",
  39841=>"111011001",
  39842=>"110101001",
  39843=>"000100100",
  39844=>"000110010",
  39845=>"000110111",
  39846=>"001000101",
  39847=>"111001101",
  39848=>"010111110",
  39849=>"010110101",
  39850=>"111111011",
  39851=>"001110000",
  39852=>"100001001",
  39853=>"011010001",
  39854=>"000011100",
  39855=>"011111110",
  39856=>"010001101",
  39857=>"011101000",
  39858=>"001111000",
  39859=>"001000011",
  39860=>"000101101",
  39861=>"110011110",
  39862=>"110110100",
  39863=>"000111010",
  39864=>"011100001",
  39865=>"100101001",
  39866=>"111110110",
  39867=>"001101001",
  39868=>"111001011",
  39869=>"001101100",
  39870=>"010000011",
  39871=>"101100100",
  39872=>"100110011",
  39873=>"001110101",
  39874=>"000001001",
  39875=>"111110100",
  39876=>"100110001",
  39877=>"000101011",
  39878=>"110011000",
  39879=>"111110001",
  39880=>"001001000",
  39881=>"100101101",
  39882=>"111111011",
  39883=>"010110101",
  39884=>"110001011",
  39885=>"100000000",
  39886=>"001110010",
  39887=>"001001100",
  39888=>"001010001",
  39889=>"000011111",
  39890=>"010101001",
  39891=>"011001001",
  39892=>"101000000",
  39893=>"001111111",
  39894=>"100000110",
  39895=>"001001111",
  39896=>"110000010",
  39897=>"101101100",
  39898=>"000101011",
  39899=>"001100100",
  39900=>"000001000",
  39901=>"010101011",
  39902=>"110110000",
  39903=>"101000000",
  39904=>"000000101",
  39905=>"001100011",
  39906=>"000111000",
  39907=>"010101010",
  39908=>"111011010",
  39909=>"111000110",
  39910=>"000100101",
  39911=>"100111011",
  39912=>"001001011",
  39913=>"001011100",
  39914=>"100011110",
  39915=>"100111011",
  39916=>"100001111",
  39917=>"100100111",
  39918=>"011101000",
  39919=>"001101000",
  39920=>"100111111",
  39921=>"001010111",
  39922=>"001100000",
  39923=>"101100101",
  39924=>"000001100",
  39925=>"000010001",
  39926=>"111100010",
  39927=>"010001101",
  39928=>"000010000",
  39929=>"110101010",
  39930=>"000101011",
  39931=>"110111010",
  39932=>"100100100",
  39933=>"111110101",
  39934=>"100101101",
  39935=>"001110010",
  39936=>"001100010",
  39937=>"111111100",
  39938=>"100111111",
  39939=>"110101111",
  39940=>"001000101",
  39941=>"100100010",
  39942=>"001111111",
  39943=>"101010110",
  39944=>"111101101",
  39945=>"101100100",
  39946=>"000011110",
  39947=>"101100010",
  39948=>"111000011",
  39949=>"001111111",
  39950=>"100100111",
  39951=>"100001100",
  39952=>"110111001",
  39953=>"000111101",
  39954=>"011001110",
  39955=>"011100111",
  39956=>"000011000",
  39957=>"000101010",
  39958=>"100111000",
  39959=>"000000101",
  39960=>"011010100",
  39961=>"111100101",
  39962=>"100110011",
  39963=>"011011011",
  39964=>"001000011",
  39965=>"111010100",
  39966=>"000111110",
  39967=>"011110100",
  39968=>"010101100",
  39969=>"001100111",
  39970=>"011111010",
  39971=>"001100100",
  39972=>"000111000",
  39973=>"000010110",
  39974=>"010000000",
  39975=>"011010110",
  39976=>"110100111",
  39977=>"001011011",
  39978=>"110011101",
  39979=>"100110010",
  39980=>"010000101",
  39981=>"111001001",
  39982=>"111111111",
  39983=>"010100100",
  39984=>"001110100",
  39985=>"000100011",
  39986=>"110110110",
  39987=>"000001100",
  39988=>"001000000",
  39989=>"111111111",
  39990=>"111010101",
  39991=>"000100011",
  39992=>"001100001",
  39993=>"001001000",
  39994=>"100011100",
  39995=>"011100110",
  39996=>"101000000",
  39997=>"100000010",
  39998=>"101010000",
  39999=>"000011101",
  40000=>"101000110",
  40001=>"011101110",
  40002=>"010100001",
  40003=>"001100001",
  40004=>"100110001",
  40005=>"111011110",
  40006=>"111100010",
  40007=>"101100101",
  40008=>"110111011",
  40009=>"001111101",
  40010=>"110101110",
  40011=>"000000001",
  40012=>"101100000",
  40013=>"010001000",
  40014=>"101100011",
  40015=>"001011000",
  40016=>"000011010",
  40017=>"010010000",
  40018=>"111010011",
  40019=>"011001011",
  40020=>"111100110",
  40021=>"111101101",
  40022=>"111011011",
  40023=>"111101001",
  40024=>"110111101",
  40025=>"000011110",
  40026=>"011011010",
  40027=>"000111100",
  40028=>"100000001",
  40029=>"101111111",
  40030=>"001110100",
  40031=>"101011001",
  40032=>"100111001",
  40033=>"011101110",
  40034=>"011100111",
  40035=>"010011100",
  40036=>"100000101",
  40037=>"010100111",
  40038=>"110110101",
  40039=>"000010111",
  40040=>"001111011",
  40041=>"111000010",
  40042=>"000000010",
  40043=>"110000010",
  40044=>"100111100",
  40045=>"000010011",
  40046=>"001110100",
  40047=>"000111111",
  40048=>"101100100",
  40049=>"011110000",
  40050=>"000011110",
  40051=>"001100010",
  40052=>"111101001",
  40053=>"111110001",
  40054=>"111100110",
  40055=>"100111000",
  40056=>"010111101",
  40057=>"111101011",
  40058=>"000001010",
  40059=>"001001101",
  40060=>"111101001",
  40061=>"001100000",
  40062=>"110000111",
  40063=>"001011110",
  40064=>"100000001",
  40065=>"000010110",
  40066=>"000101100",
  40067=>"101010111",
  40068=>"001101011",
  40069=>"011110001",
  40070=>"100100100",
  40071=>"111011111",
  40072=>"110001001",
  40073=>"000001011",
  40074=>"101001001",
  40075=>"110000011",
  40076=>"001110110",
  40077=>"000001001",
  40078=>"110101111",
  40079=>"010100101",
  40080=>"001010110",
  40081=>"101000111",
  40082=>"000110111",
  40083=>"001000111",
  40084=>"011101011",
  40085=>"001010110",
  40086=>"011110101",
  40087=>"111000000",
  40088=>"001000100",
  40089=>"001001101",
  40090=>"111011101",
  40091=>"010110000",
  40092=>"110110111",
  40093=>"101001101",
  40094=>"111011101",
  40095=>"111111010",
  40096=>"100100101",
  40097=>"000110101",
  40098=>"000100101",
  40099=>"100001000",
  40100=>"100011001",
  40101=>"000111111",
  40102=>"001100000",
  40103=>"010001000",
  40104=>"010010011",
  40105=>"001001001",
  40106=>"111010010",
  40107=>"001011010",
  40108=>"001000100",
  40109=>"000010011",
  40110=>"001010010",
  40111=>"100010101",
  40112=>"000010000",
  40113=>"000011111",
  40114=>"000001000",
  40115=>"001011001",
  40116=>"101001000",
  40117=>"010110000",
  40118=>"011000000",
  40119=>"010111100",
  40120=>"111010011",
  40121=>"101100110",
  40122=>"001001100",
  40123=>"110110011",
  40124=>"011010101",
  40125=>"010001000",
  40126=>"100010111",
  40127=>"010101001",
  40128=>"100000010",
  40129=>"111011001",
  40130=>"001001111",
  40131=>"001011000",
  40132=>"011001001",
  40133=>"001100100",
  40134=>"101011111",
  40135=>"101100111",
  40136=>"001101101",
  40137=>"011101110",
  40138=>"110111100",
  40139=>"110010110",
  40140=>"000100000",
  40141=>"110011111",
  40142=>"011011011",
  40143=>"010101110",
  40144=>"111000101",
  40145=>"011111110",
  40146=>"101001011",
  40147=>"111110001",
  40148=>"011010110",
  40149=>"110100111",
  40150=>"001100011",
  40151=>"110001111",
  40152=>"011000011",
  40153=>"100110100",
  40154=>"000101100",
  40155=>"111111011",
  40156=>"010011001",
  40157=>"000101010",
  40158=>"101001011",
  40159=>"111011111",
  40160=>"011001001",
  40161=>"011000100",
  40162=>"110000011",
  40163=>"001000101",
  40164=>"000000100",
  40165=>"101010110",
  40166=>"010010101",
  40167=>"011011011",
  40168=>"000100111",
  40169=>"001111011",
  40170=>"011011101",
  40171=>"000111111",
  40172=>"010010010",
  40173=>"101110000",
  40174=>"101101001",
  40175=>"111010011",
  40176=>"111111101",
  40177=>"011110000",
  40178=>"001000111",
  40179=>"011101011",
  40180=>"001111000",
  40181=>"111111001",
  40182=>"100000000",
  40183=>"010111111",
  40184=>"010011000",
  40185=>"010001110",
  40186=>"101000111",
  40187=>"100000111",
  40188=>"100010101",
  40189=>"011001110",
  40190=>"011110011",
  40191=>"000001000",
  40192=>"101011100",
  40193=>"011001011",
  40194=>"001000000",
  40195=>"010111010",
  40196=>"000110000",
  40197=>"000100101",
  40198=>"010010111",
  40199=>"100101000",
  40200=>"101111001",
  40201=>"000001011",
  40202=>"100001111",
  40203=>"000100100",
  40204=>"001010110",
  40205=>"001110100",
  40206=>"110110011",
  40207=>"010100110",
  40208=>"101010100",
  40209=>"000011111",
  40210=>"110100100",
  40211=>"000010001",
  40212=>"111100001",
  40213=>"001001111",
  40214=>"010110110",
  40215=>"010100110",
  40216=>"101110110",
  40217=>"011010001",
  40218=>"000100011",
  40219=>"001101010",
  40220=>"101111110",
  40221=>"111111100",
  40222=>"010110000",
  40223=>"010101000",
  40224=>"100011110",
  40225=>"101100101",
  40226=>"000101000",
  40227=>"000000000",
  40228=>"101010110",
  40229=>"010101011",
  40230=>"000000111",
  40231=>"010110001",
  40232=>"101000000",
  40233=>"000001000",
  40234=>"101011001",
  40235=>"101111011",
  40236=>"001101000",
  40237=>"111100110",
  40238=>"001001100",
  40239=>"100010011",
  40240=>"011010111",
  40241=>"000010111",
  40242=>"100010000",
  40243=>"000100100",
  40244=>"001101100",
  40245=>"001001001",
  40246=>"101111110",
  40247=>"101111111",
  40248=>"111011001",
  40249=>"001101011",
  40250=>"101101000",
  40251=>"011111010",
  40252=>"001101100",
  40253=>"111000010",
  40254=>"100100001",
  40255=>"011111110",
  40256=>"110101000",
  40257=>"010100100",
  40258=>"010000100",
  40259=>"110001011",
  40260=>"000000111",
  40261=>"111001111",
  40262=>"010001000",
  40263=>"111001110",
  40264=>"000110010",
  40265=>"000110101",
  40266=>"110001000",
  40267=>"011001101",
  40268=>"011001001",
  40269=>"001110101",
  40270=>"100111000",
  40271=>"100011101",
  40272=>"101111110",
  40273=>"001001011",
  40274=>"011000010",
  40275=>"111101101",
  40276=>"011101111",
  40277=>"000001011",
  40278=>"010011010",
  40279=>"000100010",
  40280=>"100111101",
  40281=>"100110001",
  40282=>"011011001",
  40283=>"010101010",
  40284=>"011111101",
  40285=>"001111011",
  40286=>"001111011",
  40287=>"011101011",
  40288=>"101000011",
  40289=>"101101101",
  40290=>"111110111",
  40291=>"000101001",
  40292=>"101101000",
  40293=>"010101010",
  40294=>"000010000",
  40295=>"111110000",
  40296=>"000011001",
  40297=>"011000001",
  40298=>"000101010",
  40299=>"000001100",
  40300=>"011011000",
  40301=>"110000100",
  40302=>"010000110",
  40303=>"111010000",
  40304=>"000110101",
  40305=>"011110101",
  40306=>"100111101",
  40307=>"101100011",
  40308=>"011110001",
  40309=>"110010110",
  40310=>"000011000",
  40311=>"010101111",
  40312=>"000010001",
  40313=>"110010111",
  40314=>"110010010",
  40315=>"010011000",
  40316=>"001101100",
  40317=>"011011111",
  40318=>"111100000",
  40319=>"100011101",
  40320=>"000001000",
  40321=>"010010111",
  40322=>"111110011",
  40323=>"101111100",
  40324=>"000010001",
  40325=>"110010110",
  40326=>"111110101",
  40327=>"010101111",
  40328=>"010100011",
  40329=>"001100000",
  40330=>"000000000",
  40331=>"101100101",
  40332=>"011110000",
  40333=>"001011111",
  40334=>"011111010",
  40335=>"111111111",
  40336=>"000100101",
  40337=>"101011111",
  40338=>"010000101",
  40339=>"111101101",
  40340=>"011000000",
  40341=>"101111001",
  40342=>"001000111",
  40343=>"001111111",
  40344=>"010011011",
  40345=>"101000010",
  40346=>"111010011",
  40347=>"100110110",
  40348=>"011110100",
  40349=>"000111000",
  40350=>"100001011",
  40351=>"111001110",
  40352=>"000000001",
  40353=>"101100110",
  40354=>"110111111",
  40355=>"001001010",
  40356=>"101100011",
  40357=>"000000001",
  40358=>"000101010",
  40359=>"000010101",
  40360=>"010100101",
  40361=>"011011110",
  40362=>"101000101",
  40363=>"000111010",
  40364=>"010100001",
  40365=>"010001011",
  40366=>"010010011",
  40367=>"010010100",
  40368=>"011001101",
  40369=>"000110100",
  40370=>"000100110",
  40371=>"010100000",
  40372=>"111100110",
  40373=>"010011000",
  40374=>"101001011",
  40375=>"010010000",
  40376=>"001000110",
  40377=>"010010010",
  40378=>"000010111",
  40379=>"011000010",
  40380=>"100010101",
  40381=>"011111110",
  40382=>"001101111",
  40383=>"111110101",
  40384=>"100100110",
  40385=>"001011000",
  40386=>"111101010",
  40387=>"111011011",
  40388=>"101000110",
  40389=>"101010011",
  40390=>"001000000",
  40391=>"101001000",
  40392=>"100100100",
  40393=>"111110001",
  40394=>"100010001",
  40395=>"001110110",
  40396=>"100001100",
  40397=>"101101111",
  40398=>"100010000",
  40399=>"101110011",
  40400=>"011110000",
  40401=>"100101111",
  40402=>"010010000",
  40403=>"101001011",
  40404=>"100111011",
  40405=>"001111100",
  40406=>"101111101",
  40407=>"111001011",
  40408=>"101001010",
  40409=>"010101101",
  40410=>"110111111",
  40411=>"101001100",
  40412=>"101110001",
  40413=>"000110111",
  40414=>"001011111",
  40415=>"110001010",
  40416=>"101001011",
  40417=>"010010101",
  40418=>"001000000",
  40419=>"100011101",
  40420=>"111100100",
  40421=>"001001011",
  40422=>"100100000",
  40423=>"000111100",
  40424=>"000000011",
  40425=>"011001001",
  40426=>"110110110",
  40427=>"100111000",
  40428=>"111101001",
  40429=>"110001010",
  40430=>"111100000",
  40431=>"010000000",
  40432=>"101101111",
  40433=>"001101111",
  40434=>"100000000",
  40435=>"011101001",
  40436=>"100111011",
  40437=>"000101000",
  40438=>"001111101",
  40439=>"010100001",
  40440=>"001101111",
  40441=>"001111000",
  40442=>"110111110",
  40443=>"000101011",
  40444=>"001101010",
  40445=>"110001000",
  40446=>"010110100",
  40447=>"010010101",
  40448=>"101100100",
  40449=>"001100111",
  40450=>"011010010",
  40451=>"111001010",
  40452=>"011101101",
  40453=>"110101101",
  40454=>"111010101",
  40455=>"000110000",
  40456=>"010010001",
  40457=>"011111011",
  40458=>"101011101",
  40459=>"000010010",
  40460=>"100100101",
  40461=>"100001100",
  40462=>"111001010",
  40463=>"100110011",
  40464=>"001000000",
  40465=>"001001100",
  40466=>"000100100",
  40467=>"001100100",
  40468=>"001001000",
  40469=>"000110100",
  40470=>"011001000",
  40471=>"011111001",
  40472=>"010010000",
  40473=>"100001011",
  40474=>"010001011",
  40475=>"110101001",
  40476=>"000011110",
  40477=>"101001101",
  40478=>"100000000",
  40479=>"111110100",
  40480=>"100010000",
  40481=>"110001010",
  40482=>"000000110",
  40483=>"111101110",
  40484=>"111110111",
  40485=>"010110001",
  40486=>"111010110",
  40487=>"011111111",
  40488=>"011100000",
  40489=>"010101011",
  40490=>"110110111",
  40491=>"100100100",
  40492=>"001000001",
  40493=>"000111011",
  40494=>"010111001",
  40495=>"001100001",
  40496=>"111010011",
  40497=>"100100101",
  40498=>"100110000",
  40499=>"000000100",
  40500=>"110100001",
  40501=>"001001111",
  40502=>"111101001",
  40503=>"000001100",
  40504=>"000110110",
  40505=>"000000110",
  40506=>"111011000",
  40507=>"110000000",
  40508=>"100111001",
  40509=>"010110110",
  40510=>"110110000",
  40511=>"110011101",
  40512=>"011101100",
  40513=>"010011001",
  40514=>"000111010",
  40515=>"100111111",
  40516=>"000101111",
  40517=>"111000100",
  40518=>"100101110",
  40519=>"001011110",
  40520=>"001101110",
  40521=>"100111001",
  40522=>"111101111",
  40523=>"000101101",
  40524=>"111110010",
  40525=>"110100101",
  40526=>"100010101",
  40527=>"001111000",
  40528=>"111101011",
  40529=>"011100001",
  40530=>"110111010",
  40531=>"111010001",
  40532=>"011000111",
  40533=>"101111011",
  40534=>"011111000",
  40535=>"101010110",
  40536=>"111011010",
  40537=>"010100101",
  40538=>"000110101",
  40539=>"001011110",
  40540=>"001001111",
  40541=>"101110100",
  40542=>"000001100",
  40543=>"110111101",
  40544=>"010000000",
  40545=>"000101101",
  40546=>"001011100",
  40547=>"000000101",
  40548=>"111110010",
  40549=>"111101111",
  40550=>"110100001",
  40551=>"011101100",
  40552=>"000110110",
  40553=>"101010011",
  40554=>"111011011",
  40555=>"101111101",
  40556=>"100001110",
  40557=>"011100100",
  40558=>"001011100",
  40559=>"101000100",
  40560=>"000001100",
  40561=>"000000000",
  40562=>"111000010",
  40563=>"001101101",
  40564=>"011011100",
  40565=>"001000001",
  40566=>"100101011",
  40567=>"000111100",
  40568=>"101100010",
  40569=>"101111111",
  40570=>"111000010",
  40571=>"010011011",
  40572=>"000001110",
  40573=>"001010101",
  40574=>"011010100",
  40575=>"111010100",
  40576=>"101100110",
  40577=>"100011110",
  40578=>"001011011",
  40579=>"000101010",
  40580=>"001000111",
  40581=>"000000010",
  40582=>"111100110",
  40583=>"010000100",
  40584=>"100000110",
  40585=>"001011001",
  40586=>"000100100",
  40587=>"011111101",
  40588=>"011111100",
  40589=>"001011100",
  40590=>"100100001",
  40591=>"000001100",
  40592=>"011101101",
  40593=>"110111101",
  40594=>"010010001",
  40595=>"111001000",
  40596=>"101011100",
  40597=>"011010010",
  40598=>"100111001",
  40599=>"000000010",
  40600=>"111111000",
  40601=>"000000000",
  40602=>"010001111",
  40603=>"111001100",
  40604=>"110101111",
  40605=>"111100110",
  40606=>"011010110",
  40607=>"011000100",
  40608=>"011001100",
  40609=>"111011111",
  40610=>"111111000",
  40611=>"010001000",
  40612=>"010010010",
  40613=>"111101111",
  40614=>"100001011",
  40615=>"001101010",
  40616=>"010110100",
  40617=>"101000000",
  40618=>"010000110",
  40619=>"011001011",
  40620=>"010100011",
  40621=>"000110110",
  40622=>"101101101",
  40623=>"111000000",
  40624=>"100110101",
  40625=>"110001100",
  40626=>"101011010",
  40627=>"010010000",
  40628=>"000000110",
  40629=>"011001110",
  40630=>"010001101",
  40631=>"110011011",
  40632=>"000111110",
  40633=>"001000110",
  40634=>"010001000",
  40635=>"110101010",
  40636=>"101100101",
  40637=>"111001100",
  40638=>"001110000",
  40639=>"100010011",
  40640=>"000011011",
  40641=>"101000001",
  40642=>"100001101",
  40643=>"001101111",
  40644=>"110011001",
  40645=>"011001000",
  40646=>"110111100",
  40647=>"110100110",
  40648=>"010011011",
  40649=>"100011000",
  40650=>"001000111",
  40651=>"110101000",
  40652=>"000001001",
  40653=>"110000011",
  40654=>"101010111",
  40655=>"001010111",
  40656=>"110011010",
  40657=>"011101011",
  40658=>"101101100",
  40659=>"001100101",
  40660=>"101100101",
  40661=>"100010011",
  40662=>"010011001",
  40663=>"000100001",
  40664=>"110010000",
  40665=>"010101011",
  40666=>"100010010",
  40667=>"111100100",
  40668=>"000001000",
  40669=>"100000011",
  40670=>"111001000",
  40671=>"010111101",
  40672=>"101100011",
  40673=>"000000001",
  40674=>"111101111",
  40675=>"010000001",
  40676=>"001111001",
  40677=>"011011001",
  40678=>"100000100",
  40679=>"101011111",
  40680=>"110101100",
  40681=>"111001010",
  40682=>"010001011",
  40683=>"110111011",
  40684=>"000011101",
  40685=>"000100011",
  40686=>"111010011",
  40687=>"111111111",
  40688=>"011100010",
  40689=>"100000110",
  40690=>"000100011",
  40691=>"001100101",
  40692=>"011111001",
  40693=>"111001011",
  40694=>"100101100",
  40695=>"010110111",
  40696=>"111011011",
  40697=>"000111010",
  40698=>"110100000",
  40699=>"011000000",
  40700=>"111111010",
  40701=>"000000010",
  40702=>"101111111",
  40703=>"001010100",
  40704=>"010100000",
  40705=>"010101000",
  40706=>"100100110",
  40707=>"101001011",
  40708=>"100100110",
  40709=>"001001110",
  40710=>"101110110",
  40711=>"000000111",
  40712=>"000111100",
  40713=>"111001000",
  40714=>"010000101",
  40715=>"011101000",
  40716=>"100100000",
  40717=>"011110000",
  40718=>"100100010",
  40719=>"111110010",
  40720=>"001110011",
  40721=>"110110100",
  40722=>"110001001",
  40723=>"001111111",
  40724=>"100110100",
  40725=>"000010000",
  40726=>"000001100",
  40727=>"111001101",
  40728=>"011001100",
  40729=>"111011011",
  40730=>"000001000",
  40731=>"000000110",
  40732=>"110000101",
  40733=>"001000000",
  40734=>"011011111",
  40735=>"101000011",
  40736=>"000000010",
  40737=>"001100000",
  40738=>"100111101",
  40739=>"011101011",
  40740=>"010100010",
  40741=>"010100100",
  40742=>"001011111",
  40743=>"111001011",
  40744=>"101111110",
  40745=>"110110110",
  40746=>"111101011",
  40747=>"111111000",
  40748=>"111100001",
  40749=>"000111000",
  40750=>"100110101",
  40751=>"010111110",
  40752=>"110000111",
  40753=>"100010100",
  40754=>"100110101",
  40755=>"100100100",
  40756=>"000000001",
  40757=>"110110100",
  40758=>"000011011",
  40759=>"000111111",
  40760=>"100111001",
  40761=>"100100110",
  40762=>"011100100",
  40763=>"111010111",
  40764=>"011100110",
  40765=>"111010001",
  40766=>"001001110",
  40767=>"101001101",
  40768=>"011100010",
  40769=>"110111000",
  40770=>"011001010",
  40771=>"010000100",
  40772=>"011000000",
  40773=>"011010001",
  40774=>"100100101",
  40775=>"111110001",
  40776=>"111110100",
  40777=>"000111011",
  40778=>"111110010",
  40779=>"100011110",
  40780=>"000001100",
  40781=>"111011100",
  40782=>"110000001",
  40783=>"101011111",
  40784=>"000101100",
  40785=>"011110110",
  40786=>"111110001",
  40787=>"111000001",
  40788=>"110001000",
  40789=>"001110011",
  40790=>"001001100",
  40791=>"110110011",
  40792=>"111000101",
  40793=>"111101110",
  40794=>"110111010",
  40795=>"010011011",
  40796=>"010010101",
  40797=>"100011101",
  40798=>"100010010",
  40799=>"001100011",
  40800=>"111001101",
  40801=>"100101100",
  40802=>"000001101",
  40803=>"111101111",
  40804=>"010000010",
  40805=>"101010011",
  40806=>"111110011",
  40807=>"101010010",
  40808=>"100011010",
  40809=>"101010100",
  40810=>"011110101",
  40811=>"111011101",
  40812=>"101011111",
  40813=>"010111011",
  40814=>"001101101",
  40815=>"010000110",
  40816=>"000111111",
  40817=>"111110010",
  40818=>"111110011",
  40819=>"011011010",
  40820=>"010000010",
  40821=>"000011011",
  40822=>"100001000",
  40823=>"000101110",
  40824=>"010011010",
  40825=>"111001110",
  40826=>"011101111",
  40827=>"101100010",
  40828=>"101000111",
  40829=>"101101000",
  40830=>"100111110",
  40831=>"110000101",
  40832=>"000001100",
  40833=>"111101000",
  40834=>"111011010",
  40835=>"111111101",
  40836=>"011000111",
  40837=>"011110111",
  40838=>"010011011",
  40839=>"011000010",
  40840=>"111010001",
  40841=>"001111000",
  40842=>"110111111",
  40843=>"110000101",
  40844=>"101101010",
  40845=>"001010010",
  40846=>"010110111",
  40847=>"111110100",
  40848=>"010110000",
  40849=>"011010000",
  40850=>"100001001",
  40851=>"000011001",
  40852=>"111110000",
  40853=>"111111111",
  40854=>"011011001",
  40855=>"110001010",
  40856=>"001101000",
  40857=>"110101111",
  40858=>"011101100",
  40859=>"111001010",
  40860=>"010010000",
  40861=>"001110001",
  40862=>"010011101",
  40863=>"000000110",
  40864=>"101001101",
  40865=>"001100100",
  40866=>"100110011",
  40867=>"111111110",
  40868=>"100000011",
  40869=>"110110001",
  40870=>"001010111",
  40871=>"100111011",
  40872=>"111000101",
  40873=>"001010110",
  40874=>"001111011",
  40875=>"110010101",
  40876=>"011010011",
  40877=>"010010001",
  40878=>"111101010",
  40879=>"101010011",
  40880=>"001000010",
  40881=>"011011100",
  40882=>"000110000",
  40883=>"110100101",
  40884=>"110011000",
  40885=>"111100000",
  40886=>"111000010",
  40887=>"000100010",
  40888=>"010111111",
  40889=>"101001101",
  40890=>"000011000",
  40891=>"011011100",
  40892=>"000010011",
  40893=>"101001110",
  40894=>"111000010",
  40895=>"011001000",
  40896=>"010101101",
  40897=>"010100000",
  40898=>"010110100",
  40899=>"111000100",
  40900=>"100110011",
  40901=>"111001010",
  40902=>"011100000",
  40903=>"111110011",
  40904=>"010100111",
  40905=>"001010111",
  40906=>"000010001",
  40907=>"111010110",
  40908=>"011001101",
  40909=>"000101100",
  40910=>"010101001",
  40911=>"101100001",
  40912=>"000011000",
  40913=>"010111111",
  40914=>"000000000",
  40915=>"110100100",
  40916=>"000010100",
  40917=>"111000110",
  40918=>"001100111",
  40919=>"010101110",
  40920=>"100000011",
  40921=>"010101110",
  40922=>"111101111",
  40923=>"111100110",
  40924=>"010100010",
  40925=>"010001000",
  40926=>"111100101",
  40927=>"111010110",
  40928=>"100011000",
  40929=>"100000100",
  40930=>"011011111",
  40931=>"000100010",
  40932=>"010010010",
  40933=>"111100101",
  40934=>"111010111",
  40935=>"001110000",
  40936=>"001001101",
  40937=>"100011110",
  40938=>"010100001",
  40939=>"101100111",
  40940=>"001110011",
  40941=>"111010011",
  40942=>"001000000",
  40943=>"010011010",
  40944=>"010111011",
  40945=>"011000110",
  40946=>"000011111",
  40947=>"001111000",
  40948=>"010111110",
  40949=>"110100011",
  40950=>"000000111",
  40951=>"010111111",
  40952=>"101011010",
  40953=>"110101001",
  40954=>"010100000",
  40955=>"100001000",
  40956=>"110000000",
  40957=>"000111011",
  40958=>"110000000",
  40959=>"001111100",
  40960=>"011110011",
  40961=>"010010111",
  40962=>"001101111",
  40963=>"010101111",
  40964=>"100110100",
  40965=>"010111011",
  40966=>"001111111",
  40967=>"101001110",
  40968=>"010010110",
  40969=>"000010000",
  40970=>"011000100",
  40971=>"100000110",
  40972=>"011000101",
  40973=>"111011100",
  40974=>"111011010",
  40975=>"110110100",
  40976=>"011110110",
  40977=>"010100011",
  40978=>"101000001",
  40979=>"010100000",
  40980=>"110101000",
  40981=>"100111111",
  40982=>"101101111",
  40983=>"101001000",
  40984=>"010110100",
  40985=>"000100010",
  40986=>"010000111",
  40987=>"111101011",
  40988=>"100111110",
  40989=>"101111110",
  40990=>"011101101",
  40991=>"101111111",
  40992=>"110110000",
  40993=>"010111110",
  40994=>"000011100",
  40995=>"111000001",
  40996=>"011001001",
  40997=>"010001111",
  40998=>"110101001",
  40999=>"011010001",
  41000=>"110001101",
  41001=>"101101100",
  41002=>"011000100",
  41003=>"001000101",
  41004=>"001000111",
  41005=>"100101011",
  41006=>"100100010",
  41007=>"001111010",
  41008=>"101001011",
  41009=>"000111110",
  41010=>"000100011",
  41011=>"011001111",
  41012=>"011000111",
  41013=>"010001100",
  41014=>"000001111",
  41015=>"100110011",
  41016=>"001000010",
  41017=>"010110111",
  41018=>"000010101",
  41019=>"010111010",
  41020=>"110011010",
  41021=>"110001000",
  41022=>"010001110",
  41023=>"010100110",
  41024=>"000110000",
  41025=>"101001111",
  41026=>"000110111",
  41027=>"000110010",
  41028=>"100011111",
  41029=>"000110100",
  41030=>"001110110",
  41031=>"011111111",
  41032=>"101111100",
  41033=>"101001001",
  41034=>"000000011",
  41035=>"000011110",
  41036=>"001111000",
  41037=>"000110011",
  41038=>"000110011",
  41039=>"000011110",
  41040=>"101111011",
  41041=>"010111110",
  41042=>"110111001",
  41043=>"100101000",
  41044=>"001000100",
  41045=>"011101001",
  41046=>"110011011",
  41047=>"001111100",
  41048=>"111001000",
  41049=>"100110111",
  41050=>"000000110",
  41051=>"111010110",
  41052=>"101011010",
  41053=>"010100001",
  41054=>"100110101",
  41055=>"101001101",
  41056=>"101001001",
  41057=>"101011000",
  41058=>"111111110",
  41059=>"110000011",
  41060=>"011101011",
  41061=>"101011000",
  41062=>"110010010",
  41063=>"111001011",
  41064=>"000111000",
  41065=>"001001100",
  41066=>"110010001",
  41067=>"100100010",
  41068=>"000000110",
  41069=>"111000010",
  41070=>"110011101",
  41071=>"101100000",
  41072=>"000000001",
  41073=>"011101110",
  41074=>"010011001",
  41075=>"111111101",
  41076=>"101101011",
  41077=>"111101000",
  41078=>"011000001",
  41079=>"111000000",
  41080=>"000101001",
  41081=>"100010110",
  41082=>"011110001",
  41083=>"011110010",
  41084=>"110111000",
  41085=>"100001000",
  41086=>"001110110",
  41087=>"000000100",
  41088=>"000000011",
  41089=>"000101100",
  41090=>"010010100",
  41091=>"001111011",
  41092=>"100001101",
  41093=>"010001101",
  41094=>"100000101",
  41095=>"011001100",
  41096=>"100101101",
  41097=>"110000101",
  41098=>"100111111",
  41099=>"000010000",
  41100=>"011100011",
  41101=>"011011000",
  41102=>"110111001",
  41103=>"110110110",
  41104=>"001101100",
  41105=>"010110010",
  41106=>"110111110",
  41107=>"011011011",
  41108=>"000010100",
  41109=>"011010100",
  41110=>"001000000",
  41111=>"001100101",
  41112=>"000101011",
  41113=>"000001010",
  41114=>"100100100",
  41115=>"110101100",
  41116=>"000000101",
  41117=>"001101100",
  41118=>"110110001",
  41119=>"010000010",
  41120=>"000111000",
  41121=>"010111001",
  41122=>"111111101",
  41123=>"111110011",
  41124=>"000010011",
  41125=>"000101011",
  41126=>"101111110",
  41127=>"110110011",
  41128=>"100001100",
  41129=>"111011011",
  41130=>"000000011",
  41131=>"001011110",
  41132=>"110110111",
  41133=>"010000011",
  41134=>"010001110",
  41135=>"100010101",
  41136=>"010000001",
  41137=>"111101011",
  41138=>"101000001",
  41139=>"010101011",
  41140=>"000001000",
  41141=>"111101100",
  41142=>"010110110",
  41143=>"111100000",
  41144=>"000000100",
  41145=>"001100000",
  41146=>"101111111",
  41147=>"110111001",
  41148=>"110011111",
  41149=>"111101101",
  41150=>"010010010",
  41151=>"000011011",
  41152=>"111100001",
  41153=>"101111010",
  41154=>"101000011",
  41155=>"100100001",
  41156=>"011100111",
  41157=>"001000001",
  41158=>"100001001",
  41159=>"010111010",
  41160=>"101010010",
  41161=>"000001000",
  41162=>"000001001",
  41163=>"110101111",
  41164=>"110011110",
  41165=>"100101001",
  41166=>"111001101",
  41167=>"111011110",
  41168=>"011000101",
  41169=>"001010101",
  41170=>"000000101",
  41171=>"001110011",
  41172=>"111001101",
  41173=>"011101011",
  41174=>"100111100",
  41175=>"010101001",
  41176=>"001001000",
  41177=>"111110010",
  41178=>"100001011",
  41179=>"000010001",
  41180=>"001000010",
  41181=>"101101100",
  41182=>"101000001",
  41183=>"110110101",
  41184=>"100101110",
  41185=>"001100110",
  41186=>"100111101",
  41187=>"001001111",
  41188=>"000011011",
  41189=>"000110110",
  41190=>"111110100",
  41191=>"000011101",
  41192=>"000010011",
  41193=>"111010111",
  41194=>"011100011",
  41195=>"001110110",
  41196=>"000011001",
  41197=>"000110100",
  41198=>"101111101",
  41199=>"010011001",
  41200=>"001111011",
  41201=>"001000111",
  41202=>"110011101",
  41203=>"000111011",
  41204=>"100000010",
  41205=>"110000000",
  41206=>"000100010",
  41207=>"000000011",
  41208=>"010110000",
  41209=>"110100101",
  41210=>"011011111",
  41211=>"100000111",
  41212=>"001111100",
  41213=>"011010100",
  41214=>"111001111",
  41215=>"111111100",
  41216=>"000100100",
  41217=>"000001010",
  41218=>"010110001",
  41219=>"110100111",
  41220=>"001011110",
  41221=>"110011010",
  41222=>"010000110",
  41223=>"011101100",
  41224=>"100011111",
  41225=>"010100011",
  41226=>"001111111",
  41227=>"100010001",
  41228=>"010110001",
  41229=>"100011100",
  41230=>"011011011",
  41231=>"011001110",
  41232=>"100001100",
  41233=>"000110011",
  41234=>"101111001",
  41235=>"011010010",
  41236=>"100111001",
  41237=>"101101010",
  41238=>"001001100",
  41239=>"000000100",
  41240=>"110100010",
  41241=>"010111001",
  41242=>"111001000",
  41243=>"110100011",
  41244=>"111010101",
  41245=>"010110110",
  41246=>"010001001",
  41247=>"001110000",
  41248=>"000101101",
  41249=>"110101000",
  41250=>"100100100",
  41251=>"000100101",
  41252=>"010000100",
  41253=>"101101100",
  41254=>"000001110",
  41255=>"010011000",
  41256=>"011100000",
  41257=>"011001101",
  41258=>"101000001",
  41259=>"111111110",
  41260=>"110100011",
  41261=>"101101011",
  41262=>"100011011",
  41263=>"100101010",
  41264=>"011101000",
  41265=>"000011101",
  41266=>"001111111",
  41267=>"101100100",
  41268=>"000110001",
  41269=>"010110010",
  41270=>"010010110",
  41271=>"010111011",
  41272=>"100001001",
  41273=>"110000000",
  41274=>"010101011",
  41275=>"000011010",
  41276=>"100110110",
  41277=>"000101101",
  41278=>"001100010",
  41279=>"111001111",
  41280=>"111101110",
  41281=>"100110001",
  41282=>"000111111",
  41283=>"111010110",
  41284=>"101100010",
  41285=>"100011110",
  41286=>"001010100",
  41287=>"101110010",
  41288=>"110000100",
  41289=>"111101101",
  41290=>"101001011",
  41291=>"100000000",
  41292=>"101011001",
  41293=>"001110101",
  41294=>"110110111",
  41295=>"001111010",
  41296=>"111111001",
  41297=>"101100001",
  41298=>"001001110",
  41299=>"011011010",
  41300=>"000111110",
  41301=>"000010110",
  41302=>"110111111",
  41303=>"110010110",
  41304=>"000001100",
  41305=>"000101100",
  41306=>"111011011",
  41307=>"010011100",
  41308=>"100000001",
  41309=>"001000101",
  41310=>"111110010",
  41311=>"010001010",
  41312=>"101101001",
  41313=>"110011011",
  41314=>"101100011",
  41315=>"101010111",
  41316=>"110101110",
  41317=>"110100110",
  41318=>"011011101",
  41319=>"111011111",
  41320=>"100110000",
  41321=>"001001000",
  41322=>"000010100",
  41323=>"111110010",
  41324=>"010010001",
  41325=>"101111111",
  41326=>"000001001",
  41327=>"100111111",
  41328=>"111110111",
  41329=>"111111100",
  41330=>"100010001",
  41331=>"001111010",
  41332=>"100101010",
  41333=>"011000110",
  41334=>"110101110",
  41335=>"001110100",
  41336=>"100001000",
  41337=>"001011111",
  41338=>"001111000",
  41339=>"000111111",
  41340=>"110100110",
  41341=>"000010111",
  41342=>"011000100",
  41343=>"010110000",
  41344=>"101011011",
  41345=>"111111011",
  41346=>"011011110",
  41347=>"110110011",
  41348=>"011000111",
  41349=>"110000011",
  41350=>"110011001",
  41351=>"010011100",
  41352=>"000100001",
  41353=>"111100000",
  41354=>"011110100",
  41355=>"100101110",
  41356=>"001011110",
  41357=>"111010011",
  41358=>"000010110",
  41359=>"110111100",
  41360=>"001000110",
  41361=>"100011101",
  41362=>"001110110",
  41363=>"100001111",
  41364=>"100101001",
  41365=>"010111101",
  41366=>"111111010",
  41367=>"111100101",
  41368=>"111011110",
  41369=>"000000111",
  41370=>"111011100",
  41371=>"010101001",
  41372=>"010110010",
  41373=>"001000100",
  41374=>"111111000",
  41375=>"111001010",
  41376=>"010001100",
  41377=>"111111000",
  41378=>"101000110",
  41379=>"001100101",
  41380=>"001011001",
  41381=>"110100001",
  41382=>"100101011",
  41383=>"000111000",
  41384=>"110101010",
  41385=>"000011000",
  41386=>"111110000",
  41387=>"110000000",
  41388=>"010010111",
  41389=>"101100110",
  41390=>"001001001",
  41391=>"001000001",
  41392=>"101001001",
  41393=>"111101011",
  41394=>"001110010",
  41395=>"000011110",
  41396=>"100111100",
  41397=>"010000011",
  41398=>"100001111",
  41399=>"100101100",
  41400=>"111101001",
  41401=>"000000111",
  41402=>"100010100",
  41403=>"010000001",
  41404=>"011110111",
  41405=>"010101011",
  41406=>"000011001",
  41407=>"101110011",
  41408=>"001000001",
  41409=>"001100111",
  41410=>"111000001",
  41411=>"110111111",
  41412=>"101100101",
  41413=>"100000011",
  41414=>"011001110",
  41415=>"111111011",
  41416=>"110000110",
  41417=>"001010101",
  41418=>"110110110",
  41419=>"100111111",
  41420=>"000011110",
  41421=>"010100011",
  41422=>"101100111",
  41423=>"011010001",
  41424=>"100000100",
  41425=>"110100010",
  41426=>"100111001",
  41427=>"001010111",
  41428=>"101100110",
  41429=>"000011000",
  41430=>"010011001",
  41431=>"010101101",
  41432=>"111001001",
  41433=>"111000110",
  41434=>"101000000",
  41435=>"011011001",
  41436=>"010111110",
  41437=>"000100101",
  41438=>"111010100",
  41439=>"010011011",
  41440=>"010101100",
  41441=>"110011011",
  41442=>"010101001",
  41443=>"001100010",
  41444=>"100101000",
  41445=>"000100010",
  41446=>"110101010",
  41447=>"011110110",
  41448=>"100111010",
  41449=>"001001000",
  41450=>"101111111",
  41451=>"100110011",
  41452=>"000001010",
  41453=>"010000010",
  41454=>"101011111",
  41455=>"011101011",
  41456=>"111010000",
  41457=>"101111101",
  41458=>"110111010",
  41459=>"111110110",
  41460=>"001011111",
  41461=>"000100111",
  41462=>"111011111",
  41463=>"000011110",
  41464=>"000100000",
  41465=>"110111001",
  41466=>"010101110",
  41467=>"111101101",
  41468=>"011101101",
  41469=>"101011101",
  41470=>"000110010",
  41471=>"110111000",
  41472=>"011100110",
  41473=>"000000010",
  41474=>"000011100",
  41475=>"110010111",
  41476=>"000001000",
  41477=>"111101011",
  41478=>"010110110",
  41479=>"001101010",
  41480=>"010010001",
  41481=>"111011100",
  41482=>"111010111",
  41483=>"100110011",
  41484=>"100110101",
  41485=>"110111111",
  41486=>"011101000",
  41487=>"000000100",
  41488=>"100110101",
  41489=>"101000001",
  41490=>"000010000",
  41491=>"101000011",
  41492=>"010000011",
  41493=>"110011111",
  41494=>"101011011",
  41495=>"001110101",
  41496=>"000011011",
  41497=>"100010100",
  41498=>"000000110",
  41499=>"010010101",
  41500=>"100001000",
  41501=>"101001011",
  41502=>"101100110",
  41503=>"011010100",
  41504=>"000100000",
  41505=>"011000101",
  41506=>"011100100",
  41507=>"110011100",
  41508=>"010010001",
  41509=>"111001001",
  41510=>"011010111",
  41511=>"010010100",
  41512=>"110100011",
  41513=>"101001010",
  41514=>"000001100",
  41515=>"001001111",
  41516=>"100011000",
  41517=>"010111111",
  41518=>"110001010",
  41519=>"001101011",
  41520=>"110000010",
  41521=>"001010101",
  41522=>"111111011",
  41523=>"010010010",
  41524=>"100010000",
  41525=>"100011100",
  41526=>"010001001",
  41527=>"111001011",
  41528=>"110100011",
  41529=>"000100110",
  41530=>"111000100",
  41531=>"011011000",
  41532=>"011000110",
  41533=>"101001110",
  41534=>"011000010",
  41535=>"101010100",
  41536=>"010111011",
  41537=>"000001001",
  41538=>"100100000",
  41539=>"000000111",
  41540=>"000101111",
  41541=>"110001101",
  41542=>"011100000",
  41543=>"010010011",
  41544=>"110110000",
  41545=>"011001001",
  41546=>"001110100",
  41547=>"001101000",
  41548=>"001111001",
  41549=>"001110101",
  41550=>"101100100",
  41551=>"100100000",
  41552=>"110110010",
  41553=>"100001000",
  41554=>"001111100",
  41555=>"010011011",
  41556=>"101111000",
  41557=>"011110101",
  41558=>"100101101",
  41559=>"110110101",
  41560=>"101100110",
  41561=>"011101110",
  41562=>"110000000",
  41563=>"101010011",
  41564=>"101110001",
  41565=>"001000110",
  41566=>"000111110",
  41567=>"001000000",
  41568=>"011111001",
  41569=>"100000000",
  41570=>"110100111",
  41571=>"001000100",
  41572=>"011011110",
  41573=>"110100100",
  41574=>"101001001",
  41575=>"010101010",
  41576=>"010001011",
  41577=>"011101010",
  41578=>"111110101",
  41579=>"010101110",
  41580=>"110001011",
  41581=>"010000011",
  41582=>"110110111",
  41583=>"000100010",
  41584=>"011111100",
  41585=>"110011010",
  41586=>"111100011",
  41587=>"100100010",
  41588=>"010011000",
  41589=>"111000100",
  41590=>"000010101",
  41591=>"110010000",
  41592=>"010001001",
  41593=>"100001100",
  41594=>"011111110",
  41595=>"001000011",
  41596=>"101110000",
  41597=>"010110110",
  41598=>"010111001",
  41599=>"111111011",
  41600=>"110101011",
  41601=>"110101010",
  41602=>"001011110",
  41603=>"101111111",
  41604=>"001011111",
  41605=>"011001101",
  41606=>"001101111",
  41607=>"011100100",
  41608=>"111101100",
  41609=>"011101111",
  41610=>"101100000",
  41611=>"101111101",
  41612=>"000000100",
  41613=>"100111001",
  41614=>"110100011",
  41615=>"100010001",
  41616=>"100110011",
  41617=>"000011110",
  41618=>"111110100",
  41619=>"001111111",
  41620=>"000101100",
  41621=>"110111111",
  41622=>"001101001",
  41623=>"010101100",
  41624=>"000111111",
  41625=>"101001110",
  41626=>"110010110",
  41627=>"100100001",
  41628=>"110100000",
  41629=>"111110100",
  41630=>"101110001",
  41631=>"011001100",
  41632=>"000011001",
  41633=>"110110101",
  41634=>"010111100",
  41635=>"101001100",
  41636=>"111111100",
  41637=>"101100111",
  41638=>"110000111",
  41639=>"111001100",
  41640=>"111111111",
  41641=>"001010000",
  41642=>"110001010",
  41643=>"100010101",
  41644=>"000111111",
  41645=>"101011011",
  41646=>"011011010",
  41647=>"000100001",
  41648=>"001111000",
  41649=>"010000110",
  41650=>"001000101",
  41651=>"010110000",
  41652=>"000100100",
  41653=>"011001000",
  41654=>"000100000",
  41655=>"011111100",
  41656=>"000000010",
  41657=>"111011110",
  41658=>"010001111",
  41659=>"011101110",
  41660=>"100001110",
  41661=>"100111010",
  41662=>"100011011",
  41663=>"010111110",
  41664=>"010111100",
  41665=>"101100111",
  41666=>"101100001",
  41667=>"010001101",
  41668=>"111100100",
  41669=>"001000101",
  41670=>"101000000",
  41671=>"000111110",
  41672=>"100001000",
  41673=>"000000011",
  41674=>"101110111",
  41675=>"100001111",
  41676=>"111101100",
  41677=>"011011001",
  41678=>"000111010",
  41679=>"001010111",
  41680=>"101110010",
  41681=>"010000011",
  41682=>"011000011",
  41683=>"010101101",
  41684=>"000010110",
  41685=>"000000111",
  41686=>"111101001",
  41687=>"110001011",
  41688=>"100001000",
  41689=>"001101011",
  41690=>"110111010",
  41691=>"101000111",
  41692=>"001101011",
  41693=>"111110111",
  41694=>"111100111",
  41695=>"101100011",
  41696=>"110110000",
  41697=>"101111011",
  41698=>"100001101",
  41699=>"001100010",
  41700=>"101111001",
  41701=>"100101011",
  41702=>"001000100",
  41703=>"011000111",
  41704=>"000000001",
  41705=>"110111100",
  41706=>"110100100",
  41707=>"010101100",
  41708=>"111011100",
  41709=>"000110010",
  41710=>"100010011",
  41711=>"100000111",
  41712=>"000010110",
  41713=>"101011100",
  41714=>"011010010",
  41715=>"111011101",
  41716=>"111011001",
  41717=>"010100000",
  41718=>"000011010",
  41719=>"001101011",
  41720=>"111001011",
  41721=>"001010101",
  41722=>"001101000",
  41723=>"111111111",
  41724=>"101011011",
  41725=>"001001011",
  41726=>"001100001",
  41727=>"100111000",
  41728=>"001100111",
  41729=>"011101111",
  41730=>"000100110",
  41731=>"100000010",
  41732=>"000111011",
  41733=>"101100100",
  41734=>"100010001",
  41735=>"010101000",
  41736=>"101000010",
  41737=>"111111111",
  41738=>"001000001",
  41739=>"001010001",
  41740=>"100111010",
  41741=>"111010110",
  41742=>"000000011",
  41743=>"011110000",
  41744=>"101100100",
  41745=>"000110111",
  41746=>"110110111",
  41747=>"010001101",
  41748=>"011000001",
  41749=>"100000111",
  41750=>"111110001",
  41751=>"010110111",
  41752=>"101101101",
  41753=>"101100111",
  41754=>"000001111",
  41755=>"101101110",
  41756=>"011010110",
  41757=>"001110001",
  41758=>"010100000",
  41759=>"110010001",
  41760=>"010000010",
  41761=>"100011000",
  41762=>"001011001",
  41763=>"111111101",
  41764=>"001010110",
  41765=>"101000010",
  41766=>"101110000",
  41767=>"000110100",
  41768=>"100000001",
  41769=>"100110000",
  41770=>"111010110",
  41771=>"100000011",
  41772=>"011001011",
  41773=>"100100110",
  41774=>"001000001",
  41775=>"000110010",
  41776=>"010011110",
  41777=>"101110100",
  41778=>"010001111",
  41779=>"000000111",
  41780=>"001100000",
  41781=>"010110110",
  41782=>"101001000",
  41783=>"110110001",
  41784=>"111111110",
  41785=>"101101100",
  41786=>"000111001",
  41787=>"110011110",
  41788=>"111100101",
  41789=>"011001101",
  41790=>"110001001",
  41791=>"111110011",
  41792=>"101101110",
  41793=>"001110110",
  41794=>"101100010",
  41795=>"001111000",
  41796=>"010000100",
  41797=>"000000001",
  41798=>"001011000",
  41799=>"000011011",
  41800=>"010011101",
  41801=>"000111100",
  41802=>"011000110",
  41803=>"101001111",
  41804=>"000101101",
  41805=>"100001100",
  41806=>"001010000",
  41807=>"110011110",
  41808=>"011001001",
  41809=>"000001011",
  41810=>"101010000",
  41811=>"000011011",
  41812=>"000010101",
  41813=>"110110100",
  41814=>"010101111",
  41815=>"010101000",
  41816=>"001101000",
  41817=>"001000110",
  41818=>"001101000",
  41819=>"000100000",
  41820=>"111011100",
  41821=>"010001000",
  41822=>"000010100",
  41823=>"001000100",
  41824=>"100100111",
  41825=>"001010111",
  41826=>"011100111",
  41827=>"100010111",
  41828=>"001100111",
  41829=>"101010000",
  41830=>"000101101",
  41831=>"010001111",
  41832=>"101010101",
  41833=>"001010010",
  41834=>"100110010",
  41835=>"110111100",
  41836=>"000101110",
  41837=>"110111110",
  41838=>"110001100",
  41839=>"101011110",
  41840=>"000010011",
  41841=>"101000001",
  41842=>"011110001",
  41843=>"010100100",
  41844=>"110111011",
  41845=>"000001111",
  41846=>"001111001",
  41847=>"100001010",
  41848=>"000001000",
  41849=>"001100101",
  41850=>"000110100",
  41851=>"110011011",
  41852=>"001100010",
  41853=>"000010000",
  41854=>"001100110",
  41855=>"010110000",
  41856=>"010111000",
  41857=>"001100010",
  41858=>"000110110",
  41859=>"000101001",
  41860=>"111110101",
  41861=>"110001110",
  41862=>"100000001",
  41863=>"000001100",
  41864=>"111000111",
  41865=>"000001100",
  41866=>"111111101",
  41867=>"111011000",
  41868=>"101011100",
  41869=>"101110111",
  41870=>"000001011",
  41871=>"110010101",
  41872=>"110010010",
  41873=>"000001000",
  41874=>"111001100",
  41875=>"100100001",
  41876=>"111101110",
  41877=>"101110000",
  41878=>"110010011",
  41879=>"000000001",
  41880=>"100011111",
  41881=>"000001010",
  41882=>"000001000",
  41883=>"100001100",
  41884=>"011111110",
  41885=>"101001001",
  41886=>"010001011",
  41887=>"000000011",
  41888=>"111101101",
  41889=>"110010111",
  41890=>"011011010",
  41891=>"001010101",
  41892=>"000111010",
  41893=>"001110011",
  41894=>"101001110",
  41895=>"001000001",
  41896=>"001100001",
  41897=>"101001101",
  41898=>"100111111",
  41899=>"101101000",
  41900=>"000000100",
  41901=>"101111011",
  41902=>"111001000",
  41903=>"100011001",
  41904=>"100111000",
  41905=>"110011000",
  41906=>"100001101",
  41907=>"001001001",
  41908=>"110111001",
  41909=>"101001110",
  41910=>"000000111",
  41911=>"110111011",
  41912=>"011110010",
  41913=>"001011110",
  41914=>"011101010",
  41915=>"100001000",
  41916=>"101110011",
  41917=>"001000000",
  41918=>"110001010",
  41919=>"010011000",
  41920=>"011011111",
  41921=>"000101000",
  41922=>"011001101",
  41923=>"000011100",
  41924=>"001011101",
  41925=>"110110010",
  41926=>"110011111",
  41927=>"011111011",
  41928=>"100011111",
  41929=>"110111100",
  41930=>"111000010",
  41931=>"110111110",
  41932=>"101011000",
  41933=>"101100100",
  41934=>"000000111",
  41935=>"001000011",
  41936=>"110000101",
  41937=>"111011101",
  41938=>"011010100",
  41939=>"111101110",
  41940=>"101100110",
  41941=>"010111011",
  41942=>"010111100",
  41943=>"111110010",
  41944=>"011010111",
  41945=>"000000001",
  41946=>"010001000",
  41947=>"010101111",
  41948=>"001011100",
  41949=>"011111010",
  41950=>"111111101",
  41951=>"010010000",
  41952=>"110011011",
  41953=>"110010111",
  41954=>"001111101",
  41955=>"001100110",
  41956=>"001001001",
  41957=>"000000100",
  41958=>"100000011",
  41959=>"001110101",
  41960=>"101010100",
  41961=>"001011101",
  41962=>"000000001",
  41963=>"101010000",
  41964=>"111011110",
  41965=>"110110110",
  41966=>"101011011",
  41967=>"101011010",
  41968=>"001001100",
  41969=>"010000000",
  41970=>"111001001",
  41971=>"111111000",
  41972=>"010111010",
  41973=>"000010100",
  41974=>"101111011",
  41975=>"001000110",
  41976=>"110110000",
  41977=>"000101011",
  41978=>"010111100",
  41979=>"011000000",
  41980=>"001100110",
  41981=>"001100000",
  41982=>"110111100",
  41983=>"011011001",
  41984=>"010000111",
  41985=>"111111111",
  41986=>"111000100",
  41987=>"000110111",
  41988=>"111001011",
  41989=>"001011001",
  41990=>"101110010",
  41991=>"000001000",
  41992=>"111010000",
  41993=>"100001001",
  41994=>"101100110",
  41995=>"101101101",
  41996=>"110100100",
  41997=>"110101100",
  41998=>"001111011",
  41999=>"000010011",
  42000=>"110101011",
  42001=>"100110111",
  42002=>"101101111",
  42003=>"110001001",
  42004=>"000101010",
  42005=>"010100000",
  42006=>"010100011",
  42007=>"001100100",
  42008=>"000111000",
  42009=>"010100011",
  42010=>"001100000",
  42011=>"111010111",
  42012=>"000010100",
  42013=>"111110010",
  42014=>"110111111",
  42015=>"011011000",
  42016=>"011010101",
  42017=>"010100101",
  42018=>"101001001",
  42019=>"001011000",
  42020=>"111001111",
  42021=>"110100100",
  42022=>"011110110",
  42023=>"110101111",
  42024=>"000000001",
  42025=>"101010100",
  42026=>"001000101",
  42027=>"101011100",
  42028=>"011101110",
  42029=>"100010101",
  42030=>"010011100",
  42031=>"000101000",
  42032=>"011011110",
  42033=>"100111011",
  42034=>"101111110",
  42035=>"111110101",
  42036=>"100001000",
  42037=>"000111000",
  42038=>"001111000",
  42039=>"011010101",
  42040=>"100001101",
  42041=>"110011010",
  42042=>"111001111",
  42043=>"000000101",
  42044=>"001010010",
  42045=>"011101010",
  42046=>"011100100",
  42047=>"110000011",
  42048=>"001111110",
  42049=>"001111011",
  42050=>"001001010",
  42051=>"111110010",
  42052=>"100111101",
  42053=>"110010001",
  42054=>"000010001",
  42055=>"001101001",
  42056=>"101110100",
  42057=>"110111101",
  42058=>"100111000",
  42059=>"111011110",
  42060=>"011001110",
  42061=>"010011011",
  42062=>"100111010",
  42063=>"110111001",
  42064=>"010100101",
  42065=>"110111000",
  42066=>"001100110",
  42067=>"110000011",
  42068=>"011010111",
  42069=>"110101010",
  42070=>"101101001",
  42071=>"011100111",
  42072=>"010110100",
  42073=>"111100100",
  42074=>"101111011",
  42075=>"100101001",
  42076=>"000111111",
  42077=>"000100100",
  42078=>"001001010",
  42079=>"000010010",
  42080=>"100110110",
  42081=>"001010000",
  42082=>"001011111",
  42083=>"000001100",
  42084=>"111000010",
  42085=>"010001000",
  42086=>"000101101",
  42087=>"101110101",
  42088=>"000010100",
  42089=>"001110000",
  42090=>"101011011",
  42091=>"110101111",
  42092=>"000111000",
  42093=>"001100001",
  42094=>"001101011",
  42095=>"110010101",
  42096=>"000111011",
  42097=>"000011010",
  42098=>"111010010",
  42099=>"110100110",
  42100=>"101100111",
  42101=>"011110010",
  42102=>"100111111",
  42103=>"101101010",
  42104=>"100111000",
  42105=>"100101100",
  42106=>"111100000",
  42107=>"110000000",
  42108=>"010111001",
  42109=>"000111101",
  42110=>"101001000",
  42111=>"111110101",
  42112=>"000010010",
  42113=>"000000000",
  42114=>"111000101",
  42115=>"100111011",
  42116=>"010000100",
  42117=>"010111010",
  42118=>"110010000",
  42119=>"001011101",
  42120=>"100110100",
  42121=>"010100011",
  42122=>"000100010",
  42123=>"100101010",
  42124=>"100111100",
  42125=>"001011110",
  42126=>"011011110",
  42127=>"011011111",
  42128=>"101110101",
  42129=>"110110011",
  42130=>"000010010",
  42131=>"011101111",
  42132=>"101010111",
  42133=>"011000101",
  42134=>"001100100",
  42135=>"111000110",
  42136=>"111111101",
  42137=>"011000101",
  42138=>"111100111",
  42139=>"010010010",
  42140=>"110101101",
  42141=>"101111010",
  42142=>"111011110",
  42143=>"111101100",
  42144=>"110101001",
  42145=>"010100100",
  42146=>"110010110",
  42147=>"110101001",
  42148=>"111010101",
  42149=>"010010011",
  42150=>"000101110",
  42151=>"110010001",
  42152=>"010010001",
  42153=>"100010100",
  42154=>"000110111",
  42155=>"111101011",
  42156=>"011100010",
  42157=>"001011100",
  42158=>"110010011",
  42159=>"000100101",
  42160=>"000001000",
  42161=>"001000110",
  42162=>"101100011",
  42163=>"001000110",
  42164=>"101011000",
  42165=>"110011101",
  42166=>"000111100",
  42167=>"110111100",
  42168=>"101001000",
  42169=>"101001110",
  42170=>"000100000",
  42171=>"010110000",
  42172=>"010100111",
  42173=>"001010110",
  42174=>"010010001",
  42175=>"100110011",
  42176=>"110111000",
  42177=>"101011101",
  42178=>"001100000",
  42179=>"010001001",
  42180=>"000000111",
  42181=>"100001011",
  42182=>"001100101",
  42183=>"111010101",
  42184=>"000100010",
  42185=>"101111000",
  42186=>"111100110",
  42187=>"100110111",
  42188=>"111101110",
  42189=>"100100111",
  42190=>"000011011",
  42191=>"111000111",
  42192=>"010001000",
  42193=>"101001111",
  42194=>"110101101",
  42195=>"001111011",
  42196=>"000010101",
  42197=>"110010100",
  42198=>"001101111",
  42199=>"001001110",
  42200=>"010100001",
  42201=>"010000010",
  42202=>"010110101",
  42203=>"010111010",
  42204=>"110110000",
  42205=>"110111111",
  42206=>"001110010",
  42207=>"010010101",
  42208=>"110010110",
  42209=>"000011101",
  42210=>"110010011",
  42211=>"000000011",
  42212=>"100111110",
  42213=>"111001010",
  42214=>"110101111",
  42215=>"100011110",
  42216=>"010100101",
  42217=>"010001110",
  42218=>"111000001",
  42219=>"001000101",
  42220=>"101001100",
  42221=>"011111001",
  42222=>"010011000",
  42223=>"001100000",
  42224=>"010000010",
  42225=>"111010100",
  42226=>"101110110",
  42227=>"101010111",
  42228=>"101011111",
  42229=>"011000011",
  42230=>"010011110",
  42231=>"000100001",
  42232=>"001101111",
  42233=>"000010101",
  42234=>"010101111",
  42235=>"000100110",
  42236=>"001110011",
  42237=>"000011100",
  42238=>"000000000",
  42239=>"110101111",
  42240=>"110100000",
  42241=>"111100101",
  42242=>"000110000",
  42243=>"001111101",
  42244=>"010110100",
  42245=>"101100101",
  42246=>"100001100",
  42247=>"100000110",
  42248=>"000100101",
  42249=>"011100011",
  42250=>"101001110",
  42251=>"000001010",
  42252=>"110011111",
  42253=>"100001000",
  42254=>"111000001",
  42255=>"111101111",
  42256=>"101000010",
  42257=>"011011111",
  42258=>"010010111",
  42259=>"111100100",
  42260=>"011111010",
  42261=>"011011000",
  42262=>"001011010",
  42263=>"110000110",
  42264=>"100111101",
  42265=>"001000001",
  42266=>"000010011",
  42267=>"111101101",
  42268=>"111101100",
  42269=>"111101011",
  42270=>"001010101",
  42271=>"101001010",
  42272=>"100010101",
  42273=>"001110011",
  42274=>"110011101",
  42275=>"000001001",
  42276=>"111000011",
  42277=>"001001111",
  42278=>"001010100",
  42279=>"101000011",
  42280=>"001001011",
  42281=>"111101111",
  42282=>"110010111",
  42283=>"010100001",
  42284=>"011001111",
  42285=>"101010001",
  42286=>"110000011",
  42287=>"100101001",
  42288=>"001110100",
  42289=>"110010100",
  42290=>"010010001",
  42291=>"110100101",
  42292=>"110101111",
  42293=>"111000001",
  42294=>"100000011",
  42295=>"001000001",
  42296=>"010110000",
  42297=>"100111111",
  42298=>"000010110",
  42299=>"001111110",
  42300=>"000011101",
  42301=>"001101010",
  42302=>"001100101",
  42303=>"000101110",
  42304=>"001001001",
  42305=>"101010111",
  42306=>"010110111",
  42307=>"000010111",
  42308=>"100101001",
  42309=>"100101101",
  42310=>"010111000",
  42311=>"100011011",
  42312=>"110000100",
  42313=>"111000110",
  42314=>"010100110",
  42315=>"010111100",
  42316=>"000110100",
  42317=>"010001010",
  42318=>"111101001",
  42319=>"110010111",
  42320=>"100001010",
  42321=>"100110101",
  42322=>"111011101",
  42323=>"110000011",
  42324=>"110010110",
  42325=>"011101100",
  42326=>"011100011",
  42327=>"111010111",
  42328=>"101010110",
  42329=>"001111010",
  42330=>"010101100",
  42331=>"110011010",
  42332=>"011010000",
  42333=>"111001001",
  42334=>"100000110",
  42335=>"010001001",
  42336=>"110100100",
  42337=>"110111100",
  42338=>"001011101",
  42339=>"100001001",
  42340=>"100101101",
  42341=>"010000011",
  42342=>"100101100",
  42343=>"000010001",
  42344=>"011101101",
  42345=>"100100110",
  42346=>"101101001",
  42347=>"111000100",
  42348=>"010001100",
  42349=>"011111010",
  42350=>"001001010",
  42351=>"111010011",
  42352=>"011111000",
  42353=>"111011011",
  42354=>"011010111",
  42355=>"001101001",
  42356=>"100001111",
  42357=>"001000010",
  42358=>"011010011",
  42359=>"111011010",
  42360=>"011001110",
  42361=>"110001111",
  42362=>"100000010",
  42363=>"111011011",
  42364=>"011100101",
  42365=>"100101000",
  42366=>"000001011",
  42367=>"000000110",
  42368=>"011100110",
  42369=>"111000111",
  42370=>"100011111",
  42371=>"101001110",
  42372=>"011011111",
  42373=>"011100001",
  42374=>"100111001",
  42375=>"101001110",
  42376=>"000011000",
  42377=>"011111001",
  42378=>"101000000",
  42379=>"101001010",
  42380=>"011001110",
  42381=>"110011000",
  42382=>"001001110",
  42383=>"110000110",
  42384=>"000111001",
  42385=>"100001110",
  42386=>"011111011",
  42387=>"010101111",
  42388=>"110011110",
  42389=>"110001101",
  42390=>"110110110",
  42391=>"101110010",
  42392=>"011110110",
  42393=>"111001011",
  42394=>"011101001",
  42395=>"011000010",
  42396=>"110101000",
  42397=>"010100100",
  42398=>"111000011",
  42399=>"010100101",
  42400=>"111101000",
  42401=>"010010000",
  42402=>"101010111",
  42403=>"110000110",
  42404=>"010100110",
  42405=>"011001111",
  42406=>"100000100",
  42407=>"101111101",
  42408=>"011010111",
  42409=>"110100001",
  42410=>"010010001",
  42411=>"010010101",
  42412=>"101001010",
  42413=>"000100101",
  42414=>"010101001",
  42415=>"110110110",
  42416=>"000000110",
  42417=>"110111110",
  42418=>"100111100",
  42419=>"100100010",
  42420=>"000000010",
  42421=>"011011001",
  42422=>"000110110",
  42423=>"110000001",
  42424=>"011010010",
  42425=>"101011101",
  42426=>"110010011",
  42427=>"101101011",
  42428=>"110000000",
  42429=>"010000011",
  42430=>"101001010",
  42431=>"111010111",
  42432=>"001000000",
  42433=>"011011101",
  42434=>"101101010",
  42435=>"101100001",
  42436=>"101111011",
  42437=>"011001110",
  42438=>"111111011",
  42439=>"100000010",
  42440=>"001111101",
  42441=>"010100011",
  42442=>"011011001",
  42443=>"111110111",
  42444=>"001000101",
  42445=>"010100100",
  42446=>"010000000",
  42447=>"110011010",
  42448=>"101100000",
  42449=>"111100111",
  42450=>"001011111",
  42451=>"010010111",
  42452=>"011001000",
  42453=>"011010001",
  42454=>"011101100",
  42455=>"011100101",
  42456=>"110101111",
  42457=>"111100010",
  42458=>"001011111",
  42459=>"010000011",
  42460=>"011001001",
  42461=>"100011111",
  42462=>"010101101",
  42463=>"111100011",
  42464=>"111010011",
  42465=>"001111001",
  42466=>"101111101",
  42467=>"101111111",
  42468=>"101111111",
  42469=>"011101011",
  42470=>"001100100",
  42471=>"100010010",
  42472=>"101110101",
  42473=>"011101110",
  42474=>"001001001",
  42475=>"111101101",
  42476=>"001010100",
  42477=>"100000110",
  42478=>"110110010",
  42479=>"000101111",
  42480=>"000001110",
  42481=>"100101010",
  42482=>"001100010",
  42483=>"001010110",
  42484=>"001101101",
  42485=>"101011010",
  42486=>"001000010",
  42487=>"001001001",
  42488=>"111111110",
  42489=>"100100111",
  42490=>"000000011",
  42491=>"011111000",
  42492=>"000110010",
  42493=>"110110010",
  42494=>"011000100",
  42495=>"111001101",
  42496=>"100100101",
  42497=>"101011110",
  42498=>"000100000",
  42499=>"011110101",
  42500=>"011000000",
  42501=>"101110001",
  42502=>"111011010",
  42503=>"010111100",
  42504=>"000011011",
  42505=>"111011011",
  42506=>"100101101",
  42507=>"101101000",
  42508=>"010100101",
  42509=>"111101010",
  42510=>"100101001",
  42511=>"111000111",
  42512=>"111110010",
  42513=>"100101010",
  42514=>"110110100",
  42515=>"101010010",
  42516=>"110011111",
  42517=>"000000100",
  42518=>"110110100",
  42519=>"000101011",
  42520=>"001111000",
  42521=>"110111110",
  42522=>"000111110",
  42523=>"100101001",
  42524=>"001011000",
  42525=>"110001010",
  42526=>"010001000",
  42527=>"000101010",
  42528=>"111010011",
  42529=>"101100111",
  42530=>"101000111",
  42531=>"010111110",
  42532=>"000100011",
  42533=>"000100100",
  42534=>"111010000",
  42535=>"010000100",
  42536=>"110011111",
  42537=>"110000110",
  42538=>"111111100",
  42539=>"011110100",
  42540=>"110111111",
  42541=>"101011010",
  42542=>"111001011",
  42543=>"011100110",
  42544=>"001010010",
  42545=>"001011111",
  42546=>"111011101",
  42547=>"011001010",
  42548=>"011100011",
  42549=>"001010100",
  42550=>"010000011",
  42551=>"100110100",
  42552=>"110110000",
  42553=>"010000010",
  42554=>"111000000",
  42555=>"101100110",
  42556=>"100001100",
  42557=>"110000111",
  42558=>"100001011",
  42559=>"000111100",
  42560=>"001110001",
  42561=>"111011010",
  42562=>"000111001",
  42563=>"000010110",
  42564=>"010010111",
  42565=>"101100101",
  42566=>"000011001",
  42567=>"011101111",
  42568=>"000001001",
  42569=>"111101110",
  42570=>"110000010",
  42571=>"001110010",
  42572=>"111100011",
  42573=>"101111001",
  42574=>"000101111",
  42575=>"010010000",
  42576=>"010110111",
  42577=>"000000101",
  42578=>"011101001",
  42579=>"011111110",
  42580=>"111110100",
  42581=>"010111011",
  42582=>"110011011",
  42583=>"111111101",
  42584=>"101001100",
  42585=>"011101011",
  42586=>"100111010",
  42587=>"101110110",
  42588=>"011011010",
  42589=>"000101010",
  42590=>"011101001",
  42591=>"101100101",
  42592=>"011111010",
  42593=>"000100011",
  42594=>"000010110",
  42595=>"000001011",
  42596=>"010001110",
  42597=>"000010110",
  42598=>"000011001",
  42599=>"011100100",
  42600=>"000001010",
  42601=>"101001001",
  42602=>"110111011",
  42603=>"000111001",
  42604=>"100000101",
  42605=>"110110101",
  42606=>"101111000",
  42607=>"100001110",
  42608=>"101100010",
  42609=>"000001010",
  42610=>"010101110",
  42611=>"101100000",
  42612=>"001110010",
  42613=>"000011000",
  42614=>"000010011",
  42615=>"001001111",
  42616=>"110010010",
  42617=>"110011000",
  42618=>"100000101",
  42619=>"100000000",
  42620=>"100101000",
  42621=>"111010111",
  42622=>"011000000",
  42623=>"110110111",
  42624=>"011111001",
  42625=>"000000101",
  42626=>"011011101",
  42627=>"100000000",
  42628=>"000110011",
  42629=>"010110101",
  42630=>"110010111",
  42631=>"101100101",
  42632=>"101111111",
  42633=>"000001100",
  42634=>"000111110",
  42635=>"100101110",
  42636=>"101000011",
  42637=>"011011101",
  42638=>"001101010",
  42639=>"111000100",
  42640=>"111110100",
  42641=>"001011101",
  42642=>"111100110",
  42643=>"101010000",
  42644=>"110000010",
  42645=>"011011110",
  42646=>"001100001",
  42647=>"000110100",
  42648=>"110101101",
  42649=>"110111001",
  42650=>"001110100",
  42651=>"001110100",
  42652=>"100010111",
  42653=>"101110001",
  42654=>"101100101",
  42655=>"110001001",
  42656=>"011011010",
  42657=>"001101110",
  42658=>"100001110",
  42659=>"001101101",
  42660=>"000100100",
  42661=>"010011001",
  42662=>"010010011",
  42663=>"100000011",
  42664=>"111001011",
  42665=>"010010001",
  42666=>"110101111",
  42667=>"101100101",
  42668=>"010100000",
  42669=>"100001010",
  42670=>"110011001",
  42671=>"000000010",
  42672=>"010101111",
  42673=>"111101000",
  42674=>"110001101",
  42675=>"101011001",
  42676=>"001001111",
  42677=>"001010101",
  42678=>"010011001",
  42679=>"110010010",
  42680=>"110110000",
  42681=>"110010100",
  42682=>"110001011",
  42683=>"101011111",
  42684=>"000110000",
  42685=>"010100110",
  42686=>"100001001",
  42687=>"100010100",
  42688=>"100010000",
  42689=>"010110011",
  42690=>"111010001",
  42691=>"100111010",
  42692=>"000010010",
  42693=>"011100110",
  42694=>"100100010",
  42695=>"100111011",
  42696=>"100110111",
  42697=>"101000100",
  42698=>"100110010",
  42699=>"010000000",
  42700=>"100111101",
  42701=>"101111111",
  42702=>"010110100",
  42703=>"100010101",
  42704=>"111100001",
  42705=>"000000000",
  42706=>"011010111",
  42707=>"000101000",
  42708=>"110100001",
  42709=>"001101110",
  42710=>"100111100",
  42711=>"110101100",
  42712=>"101110000",
  42713=>"011001000",
  42714=>"100110001",
  42715=>"011010001",
  42716=>"001100101",
  42717=>"100100000",
  42718=>"000100100",
  42719=>"110010001",
  42720=>"010000001",
  42721=>"001111110",
  42722=>"001011110",
  42723=>"111101000",
  42724=>"110101000",
  42725=>"011111111",
  42726=>"100010101",
  42727=>"010011100",
  42728=>"010001011",
  42729=>"000001101",
  42730=>"101000110",
  42731=>"110110010",
  42732=>"100011000",
  42733=>"001101111",
  42734=>"010101010",
  42735=>"011001110",
  42736=>"111001011",
  42737=>"111010111",
  42738=>"010101000",
  42739=>"101110000",
  42740=>"000101111",
  42741=>"100100001",
  42742=>"101110100",
  42743=>"010111111",
  42744=>"011101001",
  42745=>"001111101",
  42746=>"100101011",
  42747=>"001000111",
  42748=>"101001001",
  42749=>"010111101",
  42750=>"101101001",
  42751=>"011111000",
  42752=>"000010001",
  42753=>"100101101",
  42754=>"110111011",
  42755=>"101000101",
  42756=>"010011111",
  42757=>"000101101",
  42758=>"101011010",
  42759=>"111000100",
  42760=>"111111110",
  42761=>"001000000",
  42762=>"100000100",
  42763=>"011010010",
  42764=>"001000000",
  42765=>"111110010",
  42766=>"111010100",
  42767=>"111111101",
  42768=>"001111111",
  42769=>"101010000",
  42770=>"111101100",
  42771=>"110001011",
  42772=>"101101001",
  42773=>"101111010",
  42774=>"110100001",
  42775=>"100001001",
  42776=>"100101111",
  42777=>"000110010",
  42778=>"001000011",
  42779=>"111010011",
  42780=>"000110000",
  42781=>"011000000",
  42782=>"110000110",
  42783=>"011111011",
  42784=>"110101110",
  42785=>"100010001",
  42786=>"000000000",
  42787=>"001111110",
  42788=>"100110011",
  42789=>"000111000",
  42790=>"010110111",
  42791=>"010100100",
  42792=>"000100010",
  42793=>"111100010",
  42794=>"101011111",
  42795=>"101101100",
  42796=>"001101001",
  42797=>"101001101",
  42798=>"010000000",
  42799=>"100100111",
  42800=>"001010110",
  42801=>"111000110",
  42802=>"111010100",
  42803=>"100111001",
  42804=>"010111001",
  42805=>"001010100",
  42806=>"101010101",
  42807=>"110101111",
  42808=>"001010100",
  42809=>"011000011",
  42810=>"010000011",
  42811=>"001111110",
  42812=>"110001000",
  42813=>"010011000",
  42814=>"001010101",
  42815=>"111001111",
  42816=>"011000010",
  42817=>"000011010",
  42818=>"111111110",
  42819=>"100110011",
  42820=>"000111110",
  42821=>"101000110",
  42822=>"010111100",
  42823=>"000110100",
  42824=>"111001001",
  42825=>"101111100",
  42826=>"000011100",
  42827=>"101010111",
  42828=>"100101100",
  42829=>"100101110",
  42830=>"000000100",
  42831=>"010001001",
  42832=>"001110101",
  42833=>"011000110",
  42834=>"011100101",
  42835=>"000110101",
  42836=>"100100010",
  42837=>"000110110",
  42838=>"110110011",
  42839=>"000001011",
  42840=>"011111000",
  42841=>"010011110",
  42842=>"011101001",
  42843=>"111010101",
  42844=>"010010101",
  42845=>"110101100",
  42846=>"111111111",
  42847=>"000100010",
  42848=>"100011001",
  42849=>"000010101",
  42850=>"111110010",
  42851=>"000001101",
  42852=>"000011000",
  42853=>"111110000",
  42854=>"101000010",
  42855=>"110101001",
  42856=>"110000000",
  42857=>"101110101",
  42858=>"011010010",
  42859=>"011111001",
  42860=>"110110010",
  42861=>"101011011",
  42862=>"000110111",
  42863=>"011001000",
  42864=>"110001010",
  42865=>"010101000",
  42866=>"001101000",
  42867=>"110110100",
  42868=>"001101100",
  42869=>"000110101",
  42870=>"101011100",
  42871=>"100110111",
  42872=>"110001110",
  42873=>"010100101",
  42874=>"010001000",
  42875=>"100111101",
  42876=>"111111011",
  42877=>"101111111",
  42878=>"011110100",
  42879=>"110111111",
  42880=>"010000001",
  42881=>"000001000",
  42882=>"000001111",
  42883=>"000001001",
  42884=>"100100011",
  42885=>"010010100",
  42886=>"010110011",
  42887=>"100111111",
  42888=>"001111000",
  42889=>"000110111",
  42890=>"000000010",
  42891=>"000111000",
  42892=>"100111011",
  42893=>"000100001",
  42894=>"100001110",
  42895=>"001010110",
  42896=>"000001000",
  42897=>"101000000",
  42898=>"010100001",
  42899=>"111101111",
  42900=>"010101010",
  42901=>"010000110",
  42902=>"101111001",
  42903=>"100000010",
  42904=>"001001010",
  42905=>"010110000",
  42906=>"101101000",
  42907=>"000100101",
  42908=>"111100110",
  42909=>"001000011",
  42910=>"101001110",
  42911=>"110111111",
  42912=>"001001110",
  42913=>"100110000",
  42914=>"010011101",
  42915=>"000001100",
  42916=>"100000010",
  42917=>"011111011",
  42918=>"001000111",
  42919=>"011010010",
  42920=>"110101010",
  42921=>"111110011",
  42922=>"111010001",
  42923=>"111100000",
  42924=>"100101110",
  42925=>"000011101",
  42926=>"001011110",
  42927=>"110011011",
  42928=>"000100000",
  42929=>"000111111",
  42930=>"000000100",
  42931=>"011110111",
  42932=>"111010001",
  42933=>"010101100",
  42934=>"000001001",
  42935=>"010101001",
  42936=>"111111101",
  42937=>"100110011",
  42938=>"011100011",
  42939=>"111011100",
  42940=>"101011010",
  42941=>"000100101",
  42942=>"101011001",
  42943=>"001111011",
  42944=>"011101110",
  42945=>"010100100",
  42946=>"001100100",
  42947=>"101101011",
  42948=>"011001010",
  42949=>"100111010",
  42950=>"100101110",
  42951=>"110011000",
  42952=>"101110001",
  42953=>"100111011",
  42954=>"100110100",
  42955=>"110010110",
  42956=>"010001100",
  42957=>"000000000",
  42958=>"001100101",
  42959=>"010000100",
  42960=>"010111111",
  42961=>"010000110",
  42962=>"111010100",
  42963=>"100000100",
  42964=>"010010000",
  42965=>"101100010",
  42966=>"101111001",
  42967=>"111011100",
  42968=>"001101000",
  42969=>"000011111",
  42970=>"001001000",
  42971=>"010101000",
  42972=>"001010100",
  42973=>"101111101",
  42974=>"101101011",
  42975=>"001000001",
  42976=>"011100001",
  42977=>"111000000",
  42978=>"110011101",
  42979=>"101101110",
  42980=>"010110001",
  42981=>"100101111",
  42982=>"110110101",
  42983=>"000011101",
  42984=>"111101010",
  42985=>"110010101",
  42986=>"010100011",
  42987=>"000101101",
  42988=>"001110101",
  42989=>"111100111",
  42990=>"100101101",
  42991=>"010100110",
  42992=>"110010100",
  42993=>"000111111",
  42994=>"001000000",
  42995=>"000111001",
  42996=>"110110110",
  42997=>"000001010",
  42998=>"111100011",
  42999=>"111101111",
  43000=>"111111110",
  43001=>"001101001",
  43002=>"001000010",
  43003=>"000101101",
  43004=>"101011100",
  43005=>"000110000",
  43006=>"100001000",
  43007=>"000111010",
  43008=>"111010011",
  43009=>"101000101",
  43010=>"010011100",
  43011=>"000000100",
  43012=>"110100100",
  43013=>"000100110",
  43014=>"000011010",
  43015=>"101100000",
  43016=>"011110000",
  43017=>"100100001",
  43018=>"000001111",
  43019=>"010111101",
  43020=>"010011011",
  43021=>"101000110",
  43022=>"011011000",
  43023=>"111110111",
  43024=>"111110111",
  43025=>"100111111",
  43026=>"100100011",
  43027=>"001100101",
  43028=>"111000111",
  43029=>"001011011",
  43030=>"010100010",
  43031=>"000011010",
  43032=>"101010011",
  43033=>"111110110",
  43034=>"110100110",
  43035=>"111100111",
  43036=>"110100001",
  43037=>"010100110",
  43038=>"011010010",
  43039=>"001000011",
  43040=>"110100011",
  43041=>"011101000",
  43042=>"111100100",
  43043=>"111000111",
  43044=>"011100010",
  43045=>"111101001",
  43046=>"011000001",
  43047=>"101101011",
  43048=>"101110101",
  43049=>"011100011",
  43050=>"110010000",
  43051=>"001011110",
  43052=>"011110100",
  43053=>"010000111",
  43054=>"110100100",
  43055=>"111000100",
  43056=>"111100100",
  43057=>"111111110",
  43058=>"000000000",
  43059=>"110101010",
  43060=>"110101100",
  43061=>"100101100",
  43062=>"110000011",
  43063=>"000010101",
  43064=>"010010101",
  43065=>"101000001",
  43066=>"100011100",
  43067=>"100000110",
  43068=>"100001011",
  43069=>"111000100",
  43070=>"010101000",
  43071=>"110111001",
  43072=>"110011000",
  43073=>"101011100",
  43074=>"000100010",
  43075=>"111101000",
  43076=>"011111111",
  43077=>"001010010",
  43078=>"100101101",
  43079=>"001110001",
  43080=>"111000100",
  43081=>"010000000",
  43082=>"010111000",
  43083=>"111101000",
  43084=>"000110111",
  43085=>"000100010",
  43086=>"111000100",
  43087=>"001010101",
  43088=>"101010101",
  43089=>"001000010",
  43090=>"001001001",
  43091=>"110111001",
  43092=>"100001011",
  43093=>"011010001",
  43094=>"011111100",
  43095=>"001001111",
  43096=>"110100010",
  43097=>"011110111",
  43098=>"000100000",
  43099=>"000100000",
  43100=>"000010110",
  43101=>"001010101",
  43102=>"111001100",
  43103=>"100011010",
  43104=>"110100001",
  43105=>"110000000",
  43106=>"010001110",
  43107=>"000111111",
  43108=>"010001111",
  43109=>"110111100",
  43110=>"011001101",
  43111=>"001011000",
  43112=>"111001100",
  43113=>"010000010",
  43114=>"001111111",
  43115=>"000100111",
  43116=>"101101001",
  43117=>"000110000",
  43118=>"110110011",
  43119=>"000010111",
  43120=>"011010010",
  43121=>"001100111",
  43122=>"001101010",
  43123=>"011011010",
  43124=>"011011010",
  43125=>"000010100",
  43126=>"111111101",
  43127=>"000010011",
  43128=>"001001000",
  43129=>"111001010",
  43130=>"100011110",
  43131=>"100100000",
  43132=>"011000000",
  43133=>"111000011",
  43134=>"001001110",
  43135=>"100100011",
  43136=>"100010111",
  43137=>"000110101",
  43138=>"000101001",
  43139=>"100111001",
  43140=>"001101000",
  43141=>"011110001",
  43142=>"110111111",
  43143=>"100001101",
  43144=>"101011110",
  43145=>"111110110",
  43146=>"000000101",
  43147=>"111000001",
  43148=>"110110100",
  43149=>"001000010",
  43150=>"110001000",
  43151=>"100100001",
  43152=>"011001110",
  43153=>"111111010",
  43154=>"000011000",
  43155=>"110111100",
  43156=>"001111111",
  43157=>"010100101",
  43158=>"100111011",
  43159=>"101111101",
  43160=>"100111101",
  43161=>"000010011",
  43162=>"110011100",
  43163=>"111111101",
  43164=>"001111011",
  43165=>"000000000",
  43166=>"101000011",
  43167=>"110110011",
  43168=>"111000000",
  43169=>"111111011",
  43170=>"111010101",
  43171=>"101101011",
  43172=>"111001110",
  43173=>"101101011",
  43174=>"001000110",
  43175=>"011000000",
  43176=>"101111111",
  43177=>"111111011",
  43178=>"011101000",
  43179=>"101100010",
  43180=>"111100010",
  43181=>"110100110",
  43182=>"000101101",
  43183=>"111010111",
  43184=>"011111111",
  43185=>"100001000",
  43186=>"000000101",
  43187=>"000000111",
  43188=>"110011110",
  43189=>"000010000",
  43190=>"100010111",
  43191=>"111000100",
  43192=>"101110011",
  43193=>"000110000",
  43194=>"011101111",
  43195=>"010100000",
  43196=>"111000101",
  43197=>"011011010",
  43198=>"100110001",
  43199=>"110111100",
  43200=>"111100110",
  43201=>"011010010",
  43202=>"011000011",
  43203=>"011111001",
  43204=>"110110100",
  43205=>"111010010",
  43206=>"100111110",
  43207=>"011000000",
  43208=>"110010110",
  43209=>"001100110",
  43210=>"101011101",
  43211=>"110011011",
  43212=>"100000111",
  43213=>"010011010",
  43214=>"000010011",
  43215=>"100001000",
  43216=>"100011101",
  43217=>"001110010",
  43218=>"001101010",
  43219=>"000100100",
  43220=>"110000010",
  43221=>"111100010",
  43222=>"111110110",
  43223=>"011001101",
  43224=>"101010001",
  43225=>"010000010",
  43226=>"111100111",
  43227=>"001011101",
  43228=>"000110000",
  43229=>"000000000",
  43230=>"010100100",
  43231=>"110001010",
  43232=>"000100101",
  43233=>"011011011",
  43234=>"111101101",
  43235=>"111110010",
  43236=>"000111110",
  43237=>"011111111",
  43238=>"001110000",
  43239=>"011001110",
  43240=>"101110101",
  43241=>"010010010",
  43242=>"111100000",
  43243=>"011001101",
  43244=>"001010001",
  43245=>"110101000",
  43246=>"000111011",
  43247=>"000000010",
  43248=>"111111101",
  43249=>"100110001",
  43250=>"111110111",
  43251=>"010100000",
  43252=>"000010000",
  43253=>"111000000",
  43254=>"100010111",
  43255=>"001001011",
  43256=>"101011000",
  43257=>"111001000",
  43258=>"111011100",
  43259=>"101001011",
  43260=>"110000110",
  43261=>"000110000",
  43262=>"000011100",
  43263=>"101100111",
  43264=>"110000110",
  43265=>"000000110",
  43266=>"100100110",
  43267=>"110011001",
  43268=>"111111101",
  43269=>"011011010",
  43270=>"000100100",
  43271=>"000110001",
  43272=>"101101001",
  43273=>"000111110",
  43274=>"001011111",
  43275=>"100000001",
  43276=>"001110100",
  43277=>"011010000",
  43278=>"011001010",
  43279=>"000001000",
  43280=>"110110110",
  43281=>"010001000",
  43282=>"100101110",
  43283=>"110111111",
  43284=>"000010010",
  43285=>"010000110",
  43286=>"001101010",
  43287=>"011110000",
  43288=>"000110010",
  43289=>"010101001",
  43290=>"001000000",
  43291=>"010101010",
  43292=>"001000011",
  43293=>"000100001",
  43294=>"000011111",
  43295=>"001001011",
  43296=>"001100010",
  43297=>"001000000",
  43298=>"101110001",
  43299=>"110111010",
  43300=>"111101001",
  43301=>"100100001",
  43302=>"110011101",
  43303=>"110000011",
  43304=>"011011111",
  43305=>"100110011",
  43306=>"010110000",
  43307=>"100000110",
  43308=>"101101001",
  43309=>"101000101",
  43310=>"101000101",
  43311=>"000100100",
  43312=>"010011101",
  43313=>"101100100",
  43314=>"000110101",
  43315=>"101011011",
  43316=>"100000100",
  43317=>"001000110",
  43318=>"001101101",
  43319=>"010001000",
  43320=>"001100101",
  43321=>"010000101",
  43322=>"111001101",
  43323=>"111111100",
  43324=>"101000000",
  43325=>"100000011",
  43326=>"110001100",
  43327=>"110001001",
  43328=>"100000000",
  43329=>"111001001",
  43330=>"001001100",
  43331=>"010011010",
  43332=>"100111100",
  43333=>"000111111",
  43334=>"010000111",
  43335=>"011111001",
  43336=>"111110011",
  43337=>"001010001",
  43338=>"101011000",
  43339=>"011010110",
  43340=>"011010100",
  43341=>"000101111",
  43342=>"100001101",
  43343=>"101111111",
  43344=>"011000010",
  43345=>"011101010",
  43346=>"001101111",
  43347=>"001100001",
  43348=>"011110111",
  43349=>"110011100",
  43350=>"111001101",
  43351=>"010111001",
  43352=>"000010000",
  43353=>"011000111",
  43354=>"100000101",
  43355=>"000111011",
  43356=>"000100000",
  43357=>"111010000",
  43358=>"011100111",
  43359=>"001011110",
  43360=>"111001001",
  43361=>"011111110",
  43362=>"100111111",
  43363=>"000100001",
  43364=>"001100000",
  43365=>"110001100",
  43366=>"010111011",
  43367=>"001000011",
  43368=>"101101001",
  43369=>"110001100",
  43370=>"000100110",
  43371=>"000110110",
  43372=>"101001011",
  43373=>"010110101",
  43374=>"110110010",
  43375=>"001101100",
  43376=>"000011100",
  43377=>"110010011",
  43378=>"111100100",
  43379=>"000110001",
  43380=>"000010110",
  43381=>"001000101",
  43382=>"110000111",
  43383=>"101101110",
  43384=>"010001111",
  43385=>"000001000",
  43386=>"010010100",
  43387=>"111101101",
  43388=>"000011110",
  43389=>"110000000",
  43390=>"100010100",
  43391=>"101001010",
  43392=>"100111000",
  43393=>"010000001",
  43394=>"000110010",
  43395=>"110010001",
  43396=>"001000101",
  43397=>"001110000",
  43398=>"001000110",
  43399=>"101011001",
  43400=>"010001000",
  43401=>"101101111",
  43402=>"000010100",
  43403=>"100100110",
  43404=>"000111001",
  43405=>"110010101",
  43406=>"101000001",
  43407=>"110010111",
  43408=>"000100010",
  43409=>"101001001",
  43410=>"111000101",
  43411=>"011011110",
  43412=>"110110011",
  43413=>"001011000",
  43414=>"001001101",
  43415=>"110101100",
  43416=>"000111100",
  43417=>"011111000",
  43418=>"111010000",
  43419=>"000011011",
  43420=>"110000101",
  43421=>"101101000",
  43422=>"101100001",
  43423=>"101110101",
  43424=>"001101001",
  43425=>"111100101",
  43426=>"101100000",
  43427=>"010100111",
  43428=>"010110011",
  43429=>"101100001",
  43430=>"111111111",
  43431=>"110100010",
  43432=>"001100111",
  43433=>"101010101",
  43434=>"011100001",
  43435=>"000010001",
  43436=>"111001111",
  43437=>"111110010",
  43438=>"001100101",
  43439=>"000000101",
  43440=>"111010001",
  43441=>"011001000",
  43442=>"001111001",
  43443=>"010011101",
  43444=>"101111101",
  43445=>"100101001",
  43446=>"001011001",
  43447=>"011110101",
  43448=>"111000101",
  43449=>"011010100",
  43450=>"001000101",
  43451=>"110111100",
  43452=>"110100000",
  43453=>"110011111",
  43454=>"101110100",
  43455=>"010111101",
  43456=>"100000001",
  43457=>"110001000",
  43458=>"110110000",
  43459=>"101101101",
  43460=>"110001110",
  43461=>"011000101",
  43462=>"011011000",
  43463=>"100101000",
  43464=>"101011100",
  43465=>"101100011",
  43466=>"101010010",
  43467=>"001101000",
  43468=>"001101110",
  43469=>"110010010",
  43470=>"011000011",
  43471=>"000011000",
  43472=>"100011101",
  43473=>"000010000",
  43474=>"010111111",
  43475=>"100100000",
  43476=>"110111101",
  43477=>"110100011",
  43478=>"111000011",
  43479=>"010010101",
  43480=>"110110110",
  43481=>"111100000",
  43482=>"110110100",
  43483=>"011100101",
  43484=>"010010100",
  43485=>"011111011",
  43486=>"101111001",
  43487=>"111010111",
  43488=>"100010001",
  43489=>"110101010",
  43490=>"001111010",
  43491=>"111010011",
  43492=>"100001111",
  43493=>"001010001",
  43494=>"000000001",
  43495=>"001001010",
  43496=>"111110101",
  43497=>"101111111",
  43498=>"000100000",
  43499=>"010111110",
  43500=>"111011010",
  43501=>"110010001",
  43502=>"000110001",
  43503=>"110010111",
  43504=>"101100101",
  43505=>"000111011",
  43506=>"011001010",
  43507=>"000110010",
  43508=>"111110111",
  43509=>"010100101",
  43510=>"001111111",
  43511=>"011110000",
  43512=>"001011111",
  43513=>"011010101",
  43514=>"111001111",
  43515=>"001110101",
  43516=>"110101100",
  43517=>"100110001",
  43518=>"000010011",
  43519=>"001101010",
  43520=>"110011100",
  43521=>"100110110",
  43522=>"011101111",
  43523=>"001011100",
  43524=>"011000001",
  43525=>"111010111",
  43526=>"111001011",
  43527=>"111000111",
  43528=>"110000111",
  43529=>"111100001",
  43530=>"001100101",
  43531=>"000010000",
  43532=>"000000001",
  43533=>"110011110",
  43534=>"011011111",
  43535=>"101001000",
  43536=>"000110101",
  43537=>"101110110",
  43538=>"000100000",
  43539=>"001110010",
  43540=>"000011010",
  43541=>"000110110",
  43542=>"101011000",
  43543=>"001110001",
  43544=>"101010000",
  43545=>"001000011",
  43546=>"011011111",
  43547=>"100101100",
  43548=>"001001000",
  43549=>"011011111",
  43550=>"101001100",
  43551=>"010110000",
  43552=>"001011010",
  43553=>"111010010",
  43554=>"001001111",
  43555=>"001000011",
  43556=>"011010100",
  43557=>"100011001",
  43558=>"100001011",
  43559=>"000001101",
  43560=>"011000101",
  43561=>"001001010",
  43562=>"111101011",
  43563=>"010100011",
  43564=>"111010110",
  43565=>"100101110",
  43566=>"101000100",
  43567=>"100011010",
  43568=>"110110010",
  43569=>"110101010",
  43570=>"001100010",
  43571=>"101011101",
  43572=>"111001100",
  43573=>"011010001",
  43574=>"011011001",
  43575=>"010110000",
  43576=>"110010101",
  43577=>"001000110",
  43578=>"000101110",
  43579=>"100100000",
  43580=>"011000101",
  43581=>"010001101",
  43582=>"011101101",
  43583=>"110101000",
  43584=>"111011111",
  43585=>"110011010",
  43586=>"001010010",
  43587=>"001000111",
  43588=>"001110101",
  43589=>"101011111",
  43590=>"000101000",
  43591=>"100101001",
  43592=>"001000100",
  43593=>"101101101",
  43594=>"010110001",
  43595=>"101010000",
  43596=>"100110101",
  43597=>"010101000",
  43598=>"000101100",
  43599=>"111101011",
  43600=>"101111110",
  43601=>"110111011",
  43602=>"000101001",
  43603=>"001000001",
  43604=>"010001100",
  43605=>"000011001",
  43606=>"100111100",
  43607=>"000111100",
  43608=>"010100010",
  43609=>"100101100",
  43610=>"001001001",
  43611=>"001101110",
  43612=>"011000101",
  43613=>"100000000",
  43614=>"111111001",
  43615=>"110001110",
  43616=>"100110001",
  43617=>"011000011",
  43618=>"100110110",
  43619=>"011001111",
  43620=>"111101010",
  43621=>"100110010",
  43622=>"100101100",
  43623=>"011011001",
  43624=>"000010010",
  43625=>"101111100",
  43626=>"001110000",
  43627=>"000101011",
  43628=>"101101010",
  43629=>"011000111",
  43630=>"001000101",
  43631=>"110101011",
  43632=>"011011001",
  43633=>"001110100",
  43634=>"100101111",
  43635=>"110010010",
  43636=>"111100111",
  43637=>"110010000",
  43638=>"000011111",
  43639=>"010010110",
  43640=>"110101100",
  43641=>"011001001",
  43642=>"000100001",
  43643=>"001100101",
  43644=>"110011101",
  43645=>"110100000",
  43646=>"001000011",
  43647=>"111001000",
  43648=>"101101000",
  43649=>"110011100",
  43650=>"001010010",
  43651=>"010000110",
  43652=>"010101111",
  43653=>"101110100",
  43654=>"110101111",
  43655=>"100000110",
  43656=>"011000111",
  43657=>"010000010",
  43658=>"011010001",
  43659=>"110101100",
  43660=>"100101011",
  43661=>"001010010",
  43662=>"100010000",
  43663=>"000010001",
  43664=>"111010010",
  43665=>"111100001",
  43666=>"010000110",
  43667=>"011000110",
  43668=>"000000001",
  43669=>"000000000",
  43670=>"110100010",
  43671=>"101001111",
  43672=>"011011100",
  43673=>"100000110",
  43674=>"100001100",
  43675=>"101001010",
  43676=>"001000110",
  43677=>"100100111",
  43678=>"010100111",
  43679=>"010000100",
  43680=>"000011011",
  43681=>"111010010",
  43682=>"001111111",
  43683=>"011110110",
  43684=>"000011101",
  43685=>"100001111",
  43686=>"011001010",
  43687=>"011111001",
  43688=>"011110010",
  43689=>"100110100",
  43690=>"000011101",
  43691=>"101011110",
  43692=>"010000000",
  43693=>"111011001",
  43694=>"010101000",
  43695=>"011010100",
  43696=>"010110110",
  43697=>"011010010",
  43698=>"000000001",
  43699=>"011001110",
  43700=>"000010000",
  43701=>"011111110",
  43702=>"110000000",
  43703=>"010100100",
  43704=>"110110101",
  43705=>"011111000",
  43706=>"000110100",
  43707=>"011000100",
  43708=>"011100000",
  43709=>"010011001",
  43710=>"001001000",
  43711=>"100100011",
  43712=>"101001010",
  43713=>"000111001",
  43714=>"101101111",
  43715=>"000001100",
  43716=>"111110101",
  43717=>"100001111",
  43718=>"111010000",
  43719=>"001010110",
  43720=>"100111111",
  43721=>"111010010",
  43722=>"001001001",
  43723=>"000001111",
  43724=>"011011110",
  43725=>"011100100",
  43726=>"010001011",
  43727=>"001010000",
  43728=>"111101100",
  43729=>"110101000",
  43730=>"111010101",
  43731=>"001011010",
  43732=>"000110010",
  43733=>"111000111",
  43734=>"111101111",
  43735=>"011111011",
  43736=>"011110011",
  43737=>"111110101",
  43738=>"011100000",
  43739=>"100001001",
  43740=>"101011011",
  43741=>"100101010",
  43742=>"010110101",
  43743=>"110100010",
  43744=>"101110101",
  43745=>"111111110",
  43746=>"000000011",
  43747=>"100111100",
  43748=>"100111100",
  43749=>"000011111",
  43750=>"000110001",
  43751=>"101111111",
  43752=>"001100101",
  43753=>"001101111",
  43754=>"101110001",
  43755=>"100000111",
  43756=>"111111011",
  43757=>"101001001",
  43758=>"110100101",
  43759=>"101000100",
  43760=>"101100011",
  43761=>"011100001",
  43762=>"100000101",
  43763=>"101010000",
  43764=>"010001000",
  43765=>"000010011",
  43766=>"110000000",
  43767=>"011101111",
  43768=>"111111011",
  43769=>"100011000",
  43770=>"001101011",
  43771=>"010001001",
  43772=>"001011111",
  43773=>"000000011",
  43774=>"111001001",
  43775=>"010100000",
  43776=>"100000111",
  43777=>"011010011",
  43778=>"101101111",
  43779=>"010111000",
  43780=>"111011000",
  43781=>"000000100",
  43782=>"000010110",
  43783=>"110111101",
  43784=>"001111110",
  43785=>"110001110",
  43786=>"111101010",
  43787=>"101010011",
  43788=>"001101111",
  43789=>"101011111",
  43790=>"111011100",
  43791=>"100101001",
  43792=>"111111111",
  43793=>"001100000",
  43794=>"010001010",
  43795=>"001100000",
  43796=>"011110111",
  43797=>"101001110",
  43798=>"110011111",
  43799=>"001011011",
  43800=>"011011011",
  43801=>"110010111",
  43802=>"111110101",
  43803=>"000110011",
  43804=>"100011001",
  43805=>"010001001",
  43806=>"011000001",
  43807=>"011001011",
  43808=>"001100100",
  43809=>"100110011",
  43810=>"011000000",
  43811=>"011111101",
  43812=>"101101110",
  43813=>"001111101",
  43814=>"000001000",
  43815=>"010101011",
  43816=>"010111110",
  43817=>"001010101",
  43818=>"000011101",
  43819=>"111110001",
  43820=>"110101101",
  43821=>"011010111",
  43822=>"000001110",
  43823=>"111111011",
  43824=>"001111110",
  43825=>"101111111",
  43826=>"001101000",
  43827=>"001110101",
  43828=>"101010011",
  43829=>"101111000",
  43830=>"010000010",
  43831=>"111000001",
  43832=>"010001100",
  43833=>"000011001",
  43834=>"011000110",
  43835=>"011000000",
  43836=>"100011111",
  43837=>"001011111",
  43838=>"110010100",
  43839=>"001001111",
  43840=>"000010111",
  43841=>"000111111",
  43842=>"011110000",
  43843=>"010100010",
  43844=>"001000100",
  43845=>"100101011",
  43846=>"011011010",
  43847=>"111111111",
  43848=>"110000010",
  43849=>"100111101",
  43850=>"111100001",
  43851=>"000011010",
  43852=>"011010000",
  43853=>"000111000",
  43854=>"000011011",
  43855=>"001110110",
  43856=>"111011011",
  43857=>"011000001",
  43858=>"001010101",
  43859=>"011011011",
  43860=>"011101000",
  43861=>"111100111",
  43862=>"101100111",
  43863=>"110011001",
  43864=>"110010011",
  43865=>"000000111",
  43866=>"000110001",
  43867=>"000000000",
  43868=>"111001000",
  43869=>"001000100",
  43870=>"100100001",
  43871=>"001000010",
  43872=>"001001011",
  43873=>"010010101",
  43874=>"111011011",
  43875=>"111011100",
  43876=>"101000110",
  43877=>"111110000",
  43878=>"001010100",
  43879=>"000110001",
  43880=>"111110001",
  43881=>"111110010",
  43882=>"100110101",
  43883=>"010100000",
  43884=>"110101101",
  43885=>"011101001",
  43886=>"110111111",
  43887=>"100111111",
  43888=>"100011110",
  43889=>"110010000",
  43890=>"111110110",
  43891=>"001011001",
  43892=>"000000010",
  43893=>"111110000",
  43894=>"100111001",
  43895=>"100000011",
  43896=>"101011100",
  43897=>"010001111",
  43898=>"100000001",
  43899=>"001001100",
  43900=>"001000111",
  43901=>"001111001",
  43902=>"000111001",
  43903=>"010111000",
  43904=>"101010000",
  43905=>"110111110",
  43906=>"001011101",
  43907=>"000000000",
  43908=>"011000000",
  43909=>"101010011",
  43910=>"101010100",
  43911=>"001011110",
  43912=>"000000011",
  43913=>"001010011",
  43914=>"001100001",
  43915=>"101101000",
  43916=>"011011001",
  43917=>"100000001",
  43918=>"000101000",
  43919=>"001100010",
  43920=>"001101101",
  43921=>"011100011",
  43922=>"001111011",
  43923=>"110111010",
  43924=>"101100101",
  43925=>"000101001",
  43926=>"000101011",
  43927=>"110010101",
  43928=>"001010100",
  43929=>"011000010",
  43930=>"000101100",
  43931=>"010001110",
  43932=>"000110000",
  43933=>"100101101",
  43934=>"100000001",
  43935=>"110110010",
  43936=>"110011110",
  43937=>"010000001",
  43938=>"100001000",
  43939=>"101101000",
  43940=>"001100001",
  43941=>"000001000",
  43942=>"011110111",
  43943=>"000001100",
  43944=>"000111010",
  43945=>"101001101",
  43946=>"010111100",
  43947=>"000100101",
  43948=>"001100010",
  43949=>"111110101",
  43950=>"011111100",
  43951=>"101100000",
  43952=>"110010101",
  43953=>"110101101",
  43954=>"110110111",
  43955=>"110001100",
  43956=>"100000111",
  43957=>"010101011",
  43958=>"010000001",
  43959=>"010000110",
  43960=>"001010010",
  43961=>"010101101",
  43962=>"010110101",
  43963=>"110000001",
  43964=>"011111011",
  43965=>"001010000",
  43966=>"100010010",
  43967=>"101001101",
  43968=>"000101010",
  43969=>"000100100",
  43970=>"000110011",
  43971=>"010101001",
  43972=>"000100001",
  43973=>"101001110",
  43974=>"111101001",
  43975=>"001111111",
  43976=>"001010010",
  43977=>"000011001",
  43978=>"101100110",
  43979=>"011000001",
  43980=>"011110101",
  43981=>"101000011",
  43982=>"001111101",
  43983=>"101001000",
  43984=>"101011000",
  43985=>"101010000",
  43986=>"010000011",
  43987=>"001100010",
  43988=>"010101010",
  43989=>"111110111",
  43990=>"101101110",
  43991=>"100110000",
  43992=>"110011100",
  43993=>"011011010",
  43994=>"101010111",
  43995=>"111000000",
  43996=>"100010010",
  43997=>"111010100",
  43998=>"111000001",
  43999=>"100101010",
  44000=>"110111111",
  44001=>"111111101",
  44002=>"010010100",
  44003=>"111001001",
  44004=>"011010011",
  44005=>"110101001",
  44006=>"100110101",
  44007=>"001001011",
  44008=>"001000000",
  44009=>"011000000",
  44010=>"010000001",
  44011=>"010001101",
  44012=>"010110011",
  44013=>"001011101",
  44014=>"101000111",
  44015=>"001100110",
  44016=>"000101110",
  44017=>"000000011",
  44018=>"110101111",
  44019=>"101011000",
  44020=>"101110001",
  44021=>"110100010",
  44022=>"101101000",
  44023=>"011000010",
  44024=>"110001110",
  44025=>"010100000",
  44026=>"000000111",
  44027=>"110001011",
  44028=>"001010111",
  44029=>"111000011",
  44030=>"000000101",
  44031=>"111000110",
  44032=>"011001111",
  44033=>"011000010",
  44034=>"101001011",
  44035=>"011111011",
  44036=>"111101011",
  44037=>"010101010",
  44038=>"011100100",
  44039=>"001001101",
  44040=>"001010110",
  44041=>"001001001",
  44042=>"110001000",
  44043=>"110101111",
  44044=>"100110100",
  44045=>"110110110",
  44046=>"001110011",
  44047=>"010111011",
  44048=>"010101010",
  44049=>"110100100",
  44050=>"111110000",
  44051=>"111001001",
  44052=>"011000101",
  44053=>"011110100",
  44054=>"111001010",
  44055=>"101100011",
  44056=>"101111110",
  44057=>"101000000",
  44058=>"000010101",
  44059=>"010111101",
  44060=>"010110001",
  44061=>"101001011",
  44062=>"100010001",
  44063=>"000111101",
  44064=>"001101100",
  44065=>"011000011",
  44066=>"100001000",
  44067=>"000011111",
  44068=>"000101000",
  44069=>"010001110",
  44070=>"001110110",
  44071=>"001001010",
  44072=>"001010011",
  44073=>"011111101",
  44074=>"001010100",
  44075=>"110100011",
  44076=>"001010100",
  44077=>"101111011",
  44078=>"011100111",
  44079=>"111101000",
  44080=>"101101010",
  44081=>"110001001",
  44082=>"010001101",
  44083=>"110110000",
  44084=>"011101110",
  44085=>"010000010",
  44086=>"011101000",
  44087=>"011000110",
  44088=>"000110011",
  44089=>"000000101",
  44090=>"001100011",
  44091=>"011100010",
  44092=>"011000111",
  44093=>"001111110",
  44094=>"010001010",
  44095=>"110100100",
  44096=>"111000111",
  44097=>"000010011",
  44098=>"100000110",
  44099=>"101011101",
  44100=>"011100000",
  44101=>"110111001",
  44102=>"010010100",
  44103=>"110010010",
  44104=>"000110111",
  44105=>"001111011",
  44106=>"001101001",
  44107=>"010001111",
  44108=>"000110101",
  44109=>"111001110",
  44110=>"111001101",
  44111=>"001001100",
  44112=>"110101011",
  44113=>"000000000",
  44114=>"111101010",
  44115=>"010111111",
  44116=>"110011101",
  44117=>"001101010",
  44118=>"001001011",
  44119=>"010101110",
  44120=>"111011011",
  44121=>"001001011",
  44122=>"101110000",
  44123=>"000111101",
  44124=>"000000111",
  44125=>"010010101",
  44126=>"000001101",
  44127=>"001000001",
  44128=>"100010101",
  44129=>"101100011",
  44130=>"100010111",
  44131=>"000111000",
  44132=>"010000000",
  44133=>"010001101",
  44134=>"010011011",
  44135=>"101011000",
  44136=>"101010101",
  44137=>"001100000",
  44138=>"111011011",
  44139=>"101011101",
  44140=>"101011000",
  44141=>"111010000",
  44142=>"110001000",
  44143=>"100000010",
  44144=>"001001101",
  44145=>"011111111",
  44146=>"000110010",
  44147=>"111110100",
  44148=>"101000011",
  44149=>"111011111",
  44150=>"100010010",
  44151=>"010100011",
  44152=>"111100011",
  44153=>"001001101",
  44154=>"000110000",
  44155=>"000001000",
  44156=>"111101011",
  44157=>"110111001",
  44158=>"010101101",
  44159=>"100001110",
  44160=>"001100010",
  44161=>"111000111",
  44162=>"011101101",
  44163=>"111010110",
  44164=>"011001001",
  44165=>"001010111",
  44166=>"010111011",
  44167=>"100110101",
  44168=>"011111101",
  44169=>"010100111",
  44170=>"001010010",
  44171=>"010001011",
  44172=>"011111000",
  44173=>"001010111",
  44174=>"010010100",
  44175=>"011110110",
  44176=>"010000001",
  44177=>"011011000",
  44178=>"000110110",
  44179=>"111011001",
  44180=>"101011010",
  44181=>"001100000",
  44182=>"011010010",
  44183=>"101110110",
  44184=>"011000011",
  44185=>"110101101",
  44186=>"011100100",
  44187=>"111100100",
  44188=>"010110110",
  44189=>"111101111",
  44190=>"100100000",
  44191=>"101001100",
  44192=>"001111111",
  44193=>"000001000",
  44194=>"010100001",
  44195=>"001101111",
  44196=>"001100100",
  44197=>"010111101",
  44198=>"010110000",
  44199=>"010000101",
  44200=>"110111000",
  44201=>"111110010",
  44202=>"001001111",
  44203=>"001100100",
  44204=>"001100100",
  44205=>"001001000",
  44206=>"111110110",
  44207=>"100011110",
  44208=>"000010001",
  44209=>"101010111",
  44210=>"011010101",
  44211=>"110101100",
  44212=>"001101101",
  44213=>"010000100",
  44214=>"100010110",
  44215=>"111011111",
  44216=>"100110100",
  44217=>"010111101",
  44218=>"100101000",
  44219=>"000011000",
  44220=>"001000100",
  44221=>"000001001",
  44222=>"000100111",
  44223=>"000100111",
  44224=>"010101111",
  44225=>"100011110",
  44226=>"111100101",
  44227=>"010100010",
  44228=>"000011000",
  44229=>"111101101",
  44230=>"001001001",
  44231=>"000110111",
  44232=>"001011101",
  44233=>"100110111",
  44234=>"001000101",
  44235=>"111100111",
  44236=>"010011000",
  44237=>"011101100",
  44238=>"100100101",
  44239=>"110111010",
  44240=>"101111110",
  44241=>"101101110",
  44242=>"110001101",
  44243=>"001111001",
  44244=>"000011101",
  44245=>"101100001",
  44246=>"001000100",
  44247=>"111011110",
  44248=>"001011111",
  44249=>"010100101",
  44250=>"001011000",
  44251=>"111001001",
  44252=>"101001101",
  44253=>"100100111",
  44254=>"011011000",
  44255=>"001101010",
  44256=>"100111111",
  44257=>"111100100",
  44258=>"010111111",
  44259=>"110110111",
  44260=>"110011100",
  44261=>"010010011",
  44262=>"110100010",
  44263=>"011100111",
  44264=>"110111001",
  44265=>"111100010",
  44266=>"001101100",
  44267=>"011000000",
  44268=>"010101010",
  44269=>"111101101",
  44270=>"010010011",
  44271=>"101001001",
  44272=>"111101110",
  44273=>"100001101",
  44274=>"101111101",
  44275=>"001000101",
  44276=>"110111001",
  44277=>"010110100",
  44278=>"010011010",
  44279=>"111111111",
  44280=>"011011010",
  44281=>"111110000",
  44282=>"100001000",
  44283=>"001010011",
  44284=>"011100001",
  44285=>"000110100",
  44286=>"101000000",
  44287=>"101011101",
  44288=>"101110101",
  44289=>"000110101",
  44290=>"101100101",
  44291=>"101110001",
  44292=>"001000000",
  44293=>"010010010",
  44294=>"111001101",
  44295=>"110001000",
  44296=>"111100110",
  44297=>"000111001",
  44298=>"010100010",
  44299=>"111100001",
  44300=>"101001010",
  44301=>"000000100",
  44302=>"110101011",
  44303=>"000011110",
  44304=>"001110011",
  44305=>"000100111",
  44306=>"101110011",
  44307=>"111010101",
  44308=>"001110000",
  44309=>"100010011",
  44310=>"011010010",
  44311=>"111000001",
  44312=>"000010100",
  44313=>"100110101",
  44314=>"011101001",
  44315=>"001011000",
  44316=>"100001101",
  44317=>"011100111",
  44318=>"111100000",
  44319=>"010111000",
  44320=>"011000110",
  44321=>"000111110",
  44322=>"101001011",
  44323=>"001100001",
  44324=>"101011001",
  44325=>"010010110",
  44326=>"000101110",
  44327=>"000111111",
  44328=>"011001000",
  44329=>"100011111",
  44330=>"001001101",
  44331=>"111000101",
  44332=>"111100011",
  44333=>"100111001",
  44334=>"000110110",
  44335=>"001101100",
  44336=>"100111000",
  44337=>"101101101",
  44338=>"001110100",
  44339=>"010111100",
  44340=>"101010111",
  44341=>"001010100",
  44342=>"011001010",
  44343=>"110000100",
  44344=>"001011001",
  44345=>"001101001",
  44346=>"000010000",
  44347=>"101001001",
  44348=>"100001001",
  44349=>"110101000",
  44350=>"010111101",
  44351=>"110011111",
  44352=>"101111001",
  44353=>"100000100",
  44354=>"010001110",
  44355=>"000110110",
  44356=>"011010010",
  44357=>"010110100",
  44358=>"111001101",
  44359=>"001010110",
  44360=>"001000000",
  44361=>"101100111",
  44362=>"100111000",
  44363=>"110100100",
  44364=>"000111011",
  44365=>"110111000",
  44366=>"110111101",
  44367=>"011010111",
  44368=>"011010001",
  44369=>"000101010",
  44370=>"010000000",
  44371=>"001000100",
  44372=>"000101001",
  44373=>"101011010",
  44374=>"001001100",
  44375=>"010100110",
  44376=>"000101000",
  44377=>"010010001",
  44378=>"001111101",
  44379=>"101011100",
  44380=>"010101011",
  44381=>"000100111",
  44382=>"110000010",
  44383=>"001011000",
  44384=>"000110001",
  44385=>"100010101",
  44386=>"000000001",
  44387=>"110111111",
  44388=>"000111010",
  44389=>"111101011",
  44390=>"000010010",
  44391=>"000010001",
  44392=>"001011111",
  44393=>"010000010",
  44394=>"101100101",
  44395=>"110111000",
  44396=>"011100001",
  44397=>"110100111",
  44398=>"111100100",
  44399=>"001010000",
  44400=>"111000101",
  44401=>"111010001",
  44402=>"101010100",
  44403=>"011110110",
  44404=>"100110011",
  44405=>"100001000",
  44406=>"001100000",
  44407=>"010111000",
  44408=>"000000000",
  44409=>"011001000",
  44410=>"111111110",
  44411=>"100101101",
  44412=>"110011110",
  44413=>"110010100",
  44414=>"010010111",
  44415=>"000001011",
  44416=>"000000101",
  44417=>"000001001",
  44418=>"110000000",
  44419=>"011110000",
  44420=>"001101000",
  44421=>"111010110",
  44422=>"101000001",
  44423=>"000000000",
  44424=>"000010100",
  44425=>"010010001",
  44426=>"000000011",
  44427=>"000101000",
  44428=>"101100010",
  44429=>"100000111",
  44430=>"111101010",
  44431=>"111011110",
  44432=>"010000111",
  44433=>"100100010",
  44434=>"110100001",
  44435=>"000100100",
  44436=>"110010000",
  44437=>"011100111",
  44438=>"101110000",
  44439=>"011101110",
  44440=>"001111111",
  44441=>"101000011",
  44442=>"000101000",
  44443=>"111000101",
  44444=>"011011000",
  44445=>"000010011",
  44446=>"111010011",
  44447=>"111001100",
  44448=>"110011010",
  44449=>"101001101",
  44450=>"010110100",
  44451=>"001010011",
  44452=>"101111011",
  44453=>"101100101",
  44454=>"111011100",
  44455=>"111111001",
  44456=>"000101111",
  44457=>"011101001",
  44458=>"101000010",
  44459=>"100000111",
  44460=>"000101100",
  44461=>"001001011",
  44462=>"111111101",
  44463=>"011011111",
  44464=>"111101101",
  44465=>"000010011",
  44466=>"101110010",
  44467=>"001110010",
  44468=>"111001101",
  44469=>"010001010",
  44470=>"101100110",
  44471=>"110000111",
  44472=>"110001100",
  44473=>"100010110",
  44474=>"001111111",
  44475=>"101011111",
  44476=>"000001110",
  44477=>"100101011",
  44478=>"110111100",
  44479=>"010001011",
  44480=>"100011111",
  44481=>"000010110",
  44482=>"000010111",
  44483=>"101111001",
  44484=>"100100010",
  44485=>"111100011",
  44486=>"000100000",
  44487=>"001001111",
  44488=>"100111100",
  44489=>"100110011",
  44490=>"100010111",
  44491=>"110110000",
  44492=>"000101110",
  44493=>"010100111",
  44494=>"000100000",
  44495=>"101111000",
  44496=>"100001000",
  44497=>"000110111",
  44498=>"111011101",
  44499=>"100100010",
  44500=>"001001100",
  44501=>"110111011",
  44502=>"000100001",
  44503=>"001000010",
  44504=>"001001000",
  44505=>"010001001",
  44506=>"000000001",
  44507=>"000100111",
  44508=>"100010010",
  44509=>"011101010",
  44510=>"101011001",
  44511=>"111011010",
  44512=>"100001100",
  44513=>"100011110",
  44514=>"000010101",
  44515=>"111001110",
  44516=>"000111001",
  44517=>"111111101",
  44518=>"111111010",
  44519=>"101011110",
  44520=>"011100010",
  44521=>"010110011",
  44522=>"011010110",
  44523=>"101001000",
  44524=>"110100000",
  44525=>"111111000",
  44526=>"111110101",
  44527=>"000111110",
  44528=>"100111001",
  44529=>"101011110",
  44530=>"101111100",
  44531=>"010100001",
  44532=>"110100110",
  44533=>"001100011",
  44534=>"011101111",
  44535=>"110110011",
  44536=>"100111111",
  44537=>"110011101",
  44538=>"000000111",
  44539=>"110000100",
  44540=>"000110000",
  44541=>"101001010",
  44542=>"100001110",
  44543=>"001001101",
  44544=>"001011100",
  44545=>"100001000",
  44546=>"000101001",
  44547=>"101001011",
  44548=>"111000110",
  44549=>"101001010",
  44550=>"111111100",
  44551=>"101000011",
  44552=>"001101001",
  44553=>"101101110",
  44554=>"111101110",
  44555=>"010011101",
  44556=>"011101011",
  44557=>"111000101",
  44558=>"100000000",
  44559=>"101001101",
  44560=>"110101010",
  44561=>"111011010",
  44562=>"001111101",
  44563=>"011001000",
  44564=>"000101001",
  44565=>"111101011",
  44566=>"100111111",
  44567=>"001010001",
  44568=>"100011101",
  44569=>"101000010",
  44570=>"001010101",
  44571=>"010100001",
  44572=>"001010100",
  44573=>"110001000",
  44574=>"000110010",
  44575=>"011011101",
  44576=>"011001000",
  44577=>"011100000",
  44578=>"101111011",
  44579=>"011111101",
  44580=>"110101111",
  44581=>"101110101",
  44582=>"011110010",
  44583=>"001100010",
  44584=>"100000100",
  44585=>"111100010",
  44586=>"101010111",
  44587=>"000101000",
  44588=>"000100110",
  44589=>"100011000",
  44590=>"010101000",
  44591=>"001011101",
  44592=>"111101111",
  44593=>"011101101",
  44594=>"100000001",
  44595=>"010001100",
  44596=>"110001111",
  44597=>"011110110",
  44598=>"101000001",
  44599=>"001101111",
  44600=>"111000000",
  44601=>"011101010",
  44602=>"011101111",
  44603=>"110000011",
  44604=>"101110001",
  44605=>"000000000",
  44606=>"010001110",
  44607=>"101111000",
  44608=>"110000111",
  44609=>"010110101",
  44610=>"001001011",
  44611=>"010101011",
  44612=>"111110100",
  44613=>"010100111",
  44614=>"100000001",
  44615=>"000001101",
  44616=>"101101000",
  44617=>"111000001",
  44618=>"111010011",
  44619=>"001001000",
  44620=>"000000000",
  44621=>"011100111",
  44622=>"101110010",
  44623=>"001100111",
  44624=>"000010001",
  44625=>"100011000",
  44626=>"011101010",
  44627=>"110101111",
  44628=>"110000111",
  44629=>"010001110",
  44630=>"001011101",
  44631=>"100000000",
  44632=>"000011100",
  44633=>"011001000",
  44634=>"000110000",
  44635=>"001101010",
  44636=>"001011101",
  44637=>"110011010",
  44638=>"111100100",
  44639=>"000000011",
  44640=>"010011111",
  44641=>"000101010",
  44642=>"111000010",
  44643=>"000011001",
  44644=>"011101111",
  44645=>"001100100",
  44646=>"011100110",
  44647=>"010010110",
  44648=>"101001001",
  44649=>"100000111",
  44650=>"101011011",
  44651=>"100100011",
  44652=>"110011001",
  44653=>"010110110",
  44654=>"101111010",
  44655=>"010000101",
  44656=>"011101001",
  44657=>"001001111",
  44658=>"110100011",
  44659=>"000101100",
  44660=>"111010100",
  44661=>"110100100",
  44662=>"010110111",
  44663=>"110000100",
  44664=>"110100011",
  44665=>"010011111",
  44666=>"110101100",
  44667=>"100011010",
  44668=>"001001011",
  44669=>"000110010",
  44670=>"001001001",
  44671=>"011001001",
  44672=>"010110011",
  44673=>"011110011",
  44674=>"110011101",
  44675=>"100101101",
  44676=>"011110110",
  44677=>"010100000",
  44678=>"000111000",
  44679=>"001001101",
  44680=>"000000000",
  44681=>"001000111",
  44682=>"010000101",
  44683=>"010010111",
  44684=>"100001011",
  44685=>"000010110",
  44686=>"100011011",
  44687=>"111101110",
  44688=>"100011110",
  44689=>"111100111",
  44690=>"111010101",
  44691=>"001101000",
  44692=>"100111111",
  44693=>"110110110",
  44694=>"000001100",
  44695=>"101001011",
  44696=>"011010101",
  44697=>"111110010",
  44698=>"011000100",
  44699=>"111100000",
  44700=>"111001001",
  44701=>"110010001",
  44702=>"000000010",
  44703=>"110110001",
  44704=>"010001111",
  44705=>"110000100",
  44706=>"001101010",
  44707=>"101110110",
  44708=>"101001011",
  44709=>"100111110",
  44710=>"100001011",
  44711=>"000000110",
  44712=>"110000101",
  44713=>"111011101",
  44714=>"001000010",
  44715=>"000110100",
  44716=>"111111001",
  44717=>"011000110",
  44718=>"011110010",
  44719=>"000100000",
  44720=>"010110010",
  44721=>"011000010",
  44722=>"100100011",
  44723=>"100101011",
  44724=>"001000010",
  44725=>"000110101",
  44726=>"010001001",
  44727=>"001111010",
  44728=>"100000011",
  44729=>"010011000",
  44730=>"000000100",
  44731=>"111000000",
  44732=>"010000101",
  44733=>"011000101",
  44734=>"000101000",
  44735=>"111000101",
  44736=>"101111111",
  44737=>"010101011",
  44738=>"100011101",
  44739=>"110010011",
  44740=>"011010011",
  44741=>"010110100",
  44742=>"100000111",
  44743=>"010011110",
  44744=>"001000100",
  44745=>"000001111",
  44746=>"100100101",
  44747=>"001100111",
  44748=>"011001110",
  44749=>"100111101",
  44750=>"000010110",
  44751=>"000110010",
  44752=>"011010101",
  44753=>"010100000",
  44754=>"000101010",
  44755=>"000100110",
  44756=>"100100011",
  44757=>"111111111",
  44758=>"011110100",
  44759=>"100011100",
  44760=>"001001100",
  44761=>"100111100",
  44762=>"011111001",
  44763=>"100111110",
  44764=>"111101100",
  44765=>"111010010",
  44766=>"111110010",
  44767=>"101011110",
  44768=>"010101111",
  44769=>"010110000",
  44770=>"101100110",
  44771=>"101111011",
  44772=>"100110001",
  44773=>"110101100",
  44774=>"111010011",
  44775=>"000000100",
  44776=>"100001111",
  44777=>"011001010",
  44778=>"011011111",
  44779=>"000000010",
  44780=>"110111100",
  44781=>"101001100",
  44782=>"011010011",
  44783=>"100101010",
  44784=>"101001100",
  44785=>"110100100",
  44786=>"011100000",
  44787=>"101100001",
  44788=>"101011011",
  44789=>"100100100",
  44790=>"101101101",
  44791=>"010110110",
  44792=>"001100010",
  44793=>"111101001",
  44794=>"001010000",
  44795=>"011110110",
  44796=>"101011101",
  44797=>"110010111",
  44798=>"000011101",
  44799=>"001010011",
  44800=>"110101111",
  44801=>"000110001",
  44802=>"010110110",
  44803=>"110001010",
  44804=>"010011110",
  44805=>"111110010",
  44806=>"101001001",
  44807=>"011011100",
  44808=>"000101001",
  44809=>"111101101",
  44810=>"010000000",
  44811=>"100011001",
  44812=>"011010111",
  44813=>"000011101",
  44814=>"100101010",
  44815=>"101110111",
  44816=>"100011001",
  44817=>"010011100",
  44818=>"011001100",
  44819=>"011100000",
  44820=>"010100001",
  44821=>"010001000",
  44822=>"100001001",
  44823=>"011101011",
  44824=>"010111111",
  44825=>"110001110",
  44826=>"100110000",
  44827=>"100000011",
  44828=>"001001010",
  44829=>"010001110",
  44830=>"110001010",
  44831=>"111010010",
  44832=>"101001111",
  44833=>"011010111",
  44834=>"000011101",
  44835=>"111000011",
  44836=>"100100011",
  44837=>"101001111",
  44838=>"011110110",
  44839=>"010000101",
  44840=>"101110000",
  44841=>"001100001",
  44842=>"101010001",
  44843=>"100100010",
  44844=>"001100011",
  44845=>"000000111",
  44846=>"110100001",
  44847=>"100100001",
  44848=>"000001100",
  44849=>"011011010",
  44850=>"110000101",
  44851=>"111001110",
  44852=>"100010110",
  44853=>"100111100",
  44854=>"010001111",
  44855=>"010111010",
  44856=>"110000010",
  44857=>"110101000",
  44858=>"010001101",
  44859=>"010000000",
  44860=>"000101100",
  44861=>"000100101",
  44862=>"100111111",
  44863=>"110001011",
  44864=>"001000001",
  44865=>"100000101",
  44866=>"001000100",
  44867=>"000110111",
  44868=>"010000000",
  44869=>"111100011",
  44870=>"101000001",
  44871=>"011100101",
  44872=>"011101110",
  44873=>"101011011",
  44874=>"101101111",
  44875=>"111010011",
  44876=>"001011101",
  44877=>"101111101",
  44878=>"111000010",
  44879=>"101110001",
  44880=>"100111110",
  44881=>"100111000",
  44882=>"110000000",
  44883=>"011000010",
  44884=>"111100000",
  44885=>"000000001",
  44886=>"000000011",
  44887=>"111110101",
  44888=>"111010000",
  44889=>"011010111",
  44890=>"100100011",
  44891=>"110110110",
  44892=>"100110000",
  44893=>"011000000",
  44894=>"100001100",
  44895=>"010010100",
  44896=>"100010101",
  44897=>"011001000",
  44898=>"000101001",
  44899=>"101100001",
  44900=>"010010000",
  44901=>"011011010",
  44902=>"011000000",
  44903=>"000100100",
  44904=>"110010010",
  44905=>"001011010",
  44906=>"111100000",
  44907=>"011100011",
  44908=>"001000111",
  44909=>"000010110",
  44910=>"110000110",
  44911=>"100100010",
  44912=>"100000010",
  44913=>"011110011",
  44914=>"001001010",
  44915=>"000111111",
  44916=>"111011111",
  44917=>"000011101",
  44918=>"101010001",
  44919=>"111010000",
  44920=>"111101000",
  44921=>"010011110",
  44922=>"000000110",
  44923=>"000110010",
  44924=>"100100000",
  44925=>"100100000",
  44926=>"000110000",
  44927=>"111101000",
  44928=>"101010000",
  44929=>"001100110",
  44930=>"001000001",
  44931=>"011100001",
  44932=>"010100110",
  44933=>"010010001",
  44934=>"000110001",
  44935=>"100011000",
  44936=>"001000010",
  44937=>"110101110",
  44938=>"001110011",
  44939=>"010011100",
  44940=>"010000010",
  44941=>"110011110",
  44942=>"101110010",
  44943=>"110111011",
  44944=>"001101101",
  44945=>"010111001",
  44946=>"110101101",
  44947=>"001001101",
  44948=>"011111001",
  44949=>"111110110",
  44950=>"100010001",
  44951=>"101101100",
  44952=>"010100111",
  44953=>"110001101",
  44954=>"001011110",
  44955=>"101010111",
  44956=>"101001100",
  44957=>"110011010",
  44958=>"111010001",
  44959=>"010001011",
  44960=>"110010100",
  44961=>"000000001",
  44962=>"001011111",
  44963=>"001111111",
  44964=>"000001010",
  44965=>"000011101",
  44966=>"010010110",
  44967=>"110011110",
  44968=>"111100000",
  44969=>"000000001",
  44970=>"101110001",
  44971=>"111000101",
  44972=>"010010101",
  44973=>"110100010",
  44974=>"101110111",
  44975=>"010010011",
  44976=>"110011001",
  44977=>"001111001",
  44978=>"101010111",
  44979=>"101110010",
  44980=>"111101100",
  44981=>"100011100",
  44982=>"110010110",
  44983=>"011011111",
  44984=>"101100001",
  44985=>"000011011",
  44986=>"111111101",
  44987=>"000010011",
  44988=>"001001010",
  44989=>"000111000",
  44990=>"011100101",
  44991=>"101100000",
  44992=>"110010011",
  44993=>"100100110",
  44994=>"100000011",
  44995=>"001100100",
  44996=>"001100011",
  44997=>"100110101",
  44998=>"001011101",
  44999=>"001000000",
  45000=>"000110000",
  45001=>"000001101",
  45002=>"000000001",
  45003=>"011110110",
  45004=>"011100000",
  45005=>"101100110",
  45006=>"011100110",
  45007=>"110001111",
  45008=>"010110100",
  45009=>"101001011",
  45010=>"101000000",
  45011=>"100100001",
  45012=>"100010101",
  45013=>"100011011",
  45014=>"000101010",
  45015=>"001000101",
  45016=>"001010101",
  45017=>"100001101",
  45018=>"111011000",
  45019=>"000000100",
  45020=>"100111000",
  45021=>"001101101",
  45022=>"100101001",
  45023=>"101100001",
  45024=>"000001011",
  45025=>"101010110",
  45026=>"111011110",
  45027=>"000101011",
  45028=>"110110110",
  45029=>"110110101",
  45030=>"000101101",
  45031=>"101001010",
  45032=>"100000111",
  45033=>"111101011",
  45034=>"011100100",
  45035=>"011011101",
  45036=>"011000100",
  45037=>"110011110",
  45038=>"101001110",
  45039=>"001010011",
  45040=>"110101101",
  45041=>"111100110",
  45042=>"000001001",
  45043=>"011000001",
  45044=>"101110011",
  45045=>"001000000",
  45046=>"111111000",
  45047=>"100100111",
  45048=>"110101011",
  45049=>"010111011",
  45050=>"111111000",
  45051=>"111000111",
  45052=>"001001010",
  45053=>"010110111",
  45054=>"101101100",
  45055=>"000110101",
  45056=>"110110111",
  45057=>"100101110",
  45058=>"001011011",
  45059=>"001010111",
  45060=>"100101111",
  45061=>"101000100",
  45062=>"101010001",
  45063=>"010000111",
  45064=>"000001001",
  45065=>"111110010",
  45066=>"100001111",
  45067=>"100100011",
  45068=>"011111000",
  45069=>"110100101",
  45070=>"111011000",
  45071=>"110110111",
  45072=>"001010110",
  45073=>"011000100",
  45074=>"110010011",
  45075=>"100001111",
  45076=>"010000000",
  45077=>"111101011",
  45078=>"010000111",
  45079=>"000110100",
  45080=>"110011001",
  45081=>"011101001",
  45082=>"101100011",
  45083=>"110010001",
  45084=>"000100000",
  45085=>"111101001",
  45086=>"001001110",
  45087=>"110011110",
  45088=>"100101100",
  45089=>"000011011",
  45090=>"000110100",
  45091=>"110101101",
  45092=>"100010101",
  45093=>"011011101",
  45094=>"101111000",
  45095=>"100111100",
  45096=>"010010101",
  45097=>"110010001",
  45098=>"111100011",
  45099=>"110011111",
  45100=>"101100101",
  45101=>"110001000",
  45102=>"000001000",
  45103=>"011100111",
  45104=>"010001110",
  45105=>"010010001",
  45106=>"001000001",
  45107=>"111010010",
  45108=>"000011001",
  45109=>"111100001",
  45110=>"100011000",
  45111=>"010001001",
  45112=>"111011000",
  45113=>"001001011",
  45114=>"001111011",
  45115=>"010101100",
  45116=>"101110000",
  45117=>"010110101",
  45118=>"110010011",
  45119=>"001110001",
  45120=>"010111011",
  45121=>"000100010",
  45122=>"111010001",
  45123=>"010000101",
  45124=>"000101000",
  45125=>"010001010",
  45126=>"011001101",
  45127=>"100000001",
  45128=>"100111000",
  45129=>"101001011",
  45130=>"100110100",
  45131=>"001100000",
  45132=>"000000011",
  45133=>"011111101",
  45134=>"110111111",
  45135=>"111010001",
  45136=>"010010100",
  45137=>"001000010",
  45138=>"000001101",
  45139=>"011001110",
  45140=>"110000000",
  45141=>"101010001",
  45142=>"000100111",
  45143=>"000001000",
  45144=>"110101101",
  45145=>"001001100",
  45146=>"111011101",
  45147=>"111101000",
  45148=>"010100000",
  45149=>"000000001",
  45150=>"010101010",
  45151=>"010010010",
  45152=>"100010001",
  45153=>"011011011",
  45154=>"010010111",
  45155=>"000001001",
  45156=>"100101010",
  45157=>"100011110",
  45158=>"000010010",
  45159=>"000101010",
  45160=>"100010001",
  45161=>"000110000",
  45162=>"000001001",
  45163=>"000101001",
  45164=>"000001111",
  45165=>"001100010",
  45166=>"101011101",
  45167=>"111110010",
  45168=>"000110011",
  45169=>"110011010",
  45170=>"001010010",
  45171=>"111111001",
  45172=>"001001110",
  45173=>"110111110",
  45174=>"101111010",
  45175=>"001100110",
  45176=>"001000000",
  45177=>"111001101",
  45178=>"001100000",
  45179=>"111100001",
  45180=>"111100101",
  45181=>"101010111",
  45182=>"000000001",
  45183=>"010111110",
  45184=>"111111010",
  45185=>"010010000",
  45186=>"011101000",
  45187=>"111001110",
  45188=>"111010000",
  45189=>"111011011",
  45190=>"011111010",
  45191=>"001000100",
  45192=>"011110011",
  45193=>"010010001",
  45194=>"110110110",
  45195=>"011000000",
  45196=>"011000010",
  45197=>"100001101",
  45198=>"111001010",
  45199=>"111001100",
  45200=>"011011110",
  45201=>"010101011",
  45202=>"100000000",
  45203=>"101111111",
  45204=>"001101111",
  45205=>"001011000",
  45206=>"000000111",
  45207=>"001000111",
  45208=>"110000010",
  45209=>"011011001",
  45210=>"101100100",
  45211=>"100111101",
  45212=>"000000111",
  45213=>"100100011",
  45214=>"101000111",
  45215=>"001100010",
  45216=>"010001011",
  45217=>"001100110",
  45218=>"001000001",
  45219=>"110111010",
  45220=>"100010100",
  45221=>"110000011",
  45222=>"010101011",
  45223=>"011011010",
  45224=>"111011111",
  45225=>"011000000",
  45226=>"000100011",
  45227=>"101110111",
  45228=>"011011110",
  45229=>"010101110",
  45230=>"101111111",
  45231=>"001010001",
  45232=>"101101011",
  45233=>"111001110",
  45234=>"110011000",
  45235=>"000000101",
  45236=>"001000101",
  45237=>"000001001",
  45238=>"111011110",
  45239=>"010110011",
  45240=>"010110101",
  45241=>"110001110",
  45242=>"110111011",
  45243=>"001000100",
  45244=>"101111111",
  45245=>"000000100",
  45246=>"100110101",
  45247=>"010110101",
  45248=>"011010001",
  45249=>"100100100",
  45250=>"011101110",
  45251=>"001001100",
  45252=>"001010011",
  45253=>"110110011",
  45254=>"110011100",
  45255=>"001100101",
  45256=>"001110000",
  45257=>"111101000",
  45258=>"111011110",
  45259=>"010101100",
  45260=>"101000011",
  45261=>"010011111",
  45262=>"111111011",
  45263=>"101000101",
  45264=>"001001100",
  45265=>"000010111",
  45266=>"011011110",
  45267=>"000111000",
  45268=>"111011111",
  45269=>"010001000",
  45270=>"001011101",
  45271=>"100101001",
  45272=>"100000111",
  45273=>"111010101",
  45274=>"010111011",
  45275=>"011110100",
  45276=>"000111111",
  45277=>"111101110",
  45278=>"100001001",
  45279=>"110010000",
  45280=>"110010010",
  45281=>"100000001",
  45282=>"111101100",
  45283=>"000101010",
  45284=>"011100000",
  45285=>"110100101",
  45286=>"001000101",
  45287=>"000101101",
  45288=>"100001010",
  45289=>"010110111",
  45290=>"011101010",
  45291=>"100111000",
  45292=>"100111010",
  45293=>"000010110",
  45294=>"100110010",
  45295=>"010111010",
  45296=>"110001111",
  45297=>"000100110",
  45298=>"100110001",
  45299=>"111101110",
  45300=>"101010110",
  45301=>"100001000",
  45302=>"111111000",
  45303=>"111000101",
  45304=>"011010101",
  45305=>"011001010",
  45306=>"101000101",
  45307=>"000100001",
  45308=>"101010011",
  45309=>"110110000",
  45310=>"111001011",
  45311=>"000011110",
  45312=>"010110000",
  45313=>"000100000",
  45314=>"101111011",
  45315=>"100000011",
  45316=>"001011111",
  45317=>"011110011",
  45318=>"110100010",
  45319=>"000100111",
  45320=>"010100011",
  45321=>"000010001",
  45322=>"111111111",
  45323=>"000101000",
  45324=>"001110011",
  45325=>"110001010",
  45326=>"110010101",
  45327=>"111111111",
  45328=>"101000010",
  45329=>"000111101",
  45330=>"010111101",
  45331=>"001011100",
  45332=>"001001100",
  45333=>"000100000",
  45334=>"000110001",
  45335=>"010111000",
  45336=>"110101000",
  45337=>"100001101",
  45338=>"011011001",
  45339=>"110101101",
  45340=>"011111010",
  45341=>"100101101",
  45342=>"110001100",
  45343=>"010100100",
  45344=>"111111010",
  45345=>"011100011",
  45346=>"101101001",
  45347=>"101111110",
  45348=>"111111011",
  45349=>"110011010",
  45350=>"111001001",
  45351=>"111100100",
  45352=>"001001000",
  45353=>"100101111",
  45354=>"110011110",
  45355=>"100101101",
  45356=>"001110100",
  45357=>"111111110",
  45358=>"011111110",
  45359=>"001100101",
  45360=>"000001010",
  45361=>"000000100",
  45362=>"111001001",
  45363=>"011000001",
  45364=>"100101110",
  45365=>"010000000",
  45366=>"011111111",
  45367=>"110111010",
  45368=>"100001110",
  45369=>"010100010",
  45370=>"001101111",
  45371=>"110111110",
  45372=>"011101011",
  45373=>"101110100",
  45374=>"100111110",
  45375=>"100011101",
  45376=>"111110001",
  45377=>"100011000",
  45378=>"111101011",
  45379=>"110100101",
  45380=>"110000001",
  45381=>"100101111",
  45382=>"000010010",
  45383=>"001000111",
  45384=>"100101101",
  45385=>"111001110",
  45386=>"110001000",
  45387=>"110110101",
  45388=>"001111001",
  45389=>"110100111",
  45390=>"110111101",
  45391=>"100000000",
  45392=>"100101011",
  45393=>"011001010",
  45394=>"111111101",
  45395=>"101100100",
  45396=>"001011010",
  45397=>"101001111",
  45398=>"011100101",
  45399=>"110000111",
  45400=>"001011011",
  45401=>"101100101",
  45402=>"000001000",
  45403=>"001001100",
  45404=>"111001100",
  45405=>"001001101",
  45406=>"001011000",
  45407=>"110001010",
  45408=>"110010101",
  45409=>"110111101",
  45410=>"111011101",
  45411=>"001110010",
  45412=>"111111111",
  45413=>"010101000",
  45414=>"100100011",
  45415=>"110111011",
  45416=>"011011001",
  45417=>"010011111",
  45418=>"100000001",
  45419=>"000010011",
  45420=>"000000000",
  45421=>"110110011",
  45422=>"010101000",
  45423=>"101111011",
  45424=>"000100110",
  45425=>"010000101",
  45426=>"110011110",
  45427=>"010010111",
  45428=>"000010111",
  45429=>"001100000",
  45430=>"011000110",
  45431=>"000100000",
  45432=>"100001001",
  45433=>"111101010",
  45434=>"011100101",
  45435=>"110010011",
  45436=>"111000001",
  45437=>"001000011",
  45438=>"000001000",
  45439=>"110001010",
  45440=>"101101101",
  45441=>"000110011",
  45442=>"101011001",
  45443=>"011011011",
  45444=>"001000100",
  45445=>"000001100",
  45446=>"001001110",
  45447=>"101110110",
  45448=>"000001110",
  45449=>"010101001",
  45450=>"101110001",
  45451=>"000101001",
  45452=>"010000110",
  45453=>"101101100",
  45454=>"100000111",
  45455=>"000100000",
  45456=>"000100000",
  45457=>"100111000",
  45458=>"110100110",
  45459=>"100001011",
  45460=>"001000101",
  45461=>"000100110",
  45462=>"110010111",
  45463=>"010101111",
  45464=>"110100101",
  45465=>"111010110",
  45466=>"101011111",
  45467=>"100101111",
  45468=>"011111011",
  45469=>"001010101",
  45470=>"100011011",
  45471=>"001000010",
  45472=>"101100000",
  45473=>"010011101",
  45474=>"010011010",
  45475=>"111110110",
  45476=>"001011101",
  45477=>"110101111",
  45478=>"010000001",
  45479=>"000111101",
  45480=>"111110000",
  45481=>"111011111",
  45482=>"100101001",
  45483=>"000101001",
  45484=>"111100011",
  45485=>"001001111",
  45486=>"010101010",
  45487=>"101110111",
  45488=>"100011011",
  45489=>"100000100",
  45490=>"100011101",
  45491=>"000101010",
  45492=>"111101001",
  45493=>"111010110",
  45494=>"010011001",
  45495=>"101110111",
  45496=>"011011010",
  45497=>"011000001",
  45498=>"001101001",
  45499=>"010010011",
  45500=>"101000000",
  45501=>"011010101",
  45502=>"111101100",
  45503=>"100100101",
  45504=>"101110011",
  45505=>"110001101",
  45506=>"000100010",
  45507=>"001101110",
  45508=>"001010010",
  45509=>"110100000",
  45510=>"000110010",
  45511=>"000010000",
  45512=>"010010010",
  45513=>"111000101",
  45514=>"011011101",
  45515=>"010010101",
  45516=>"100001100",
  45517=>"100101011",
  45518=>"000110000",
  45519=>"010001001",
  45520=>"000010100",
  45521=>"001010101",
  45522=>"111001001",
  45523=>"010010100",
  45524=>"110100011",
  45525=>"110011010",
  45526=>"100101011",
  45527=>"110001101",
  45528=>"100000001",
  45529=>"111111110",
  45530=>"010011010",
  45531=>"000100000",
  45532=>"101001110",
  45533=>"111001011",
  45534=>"000011010",
  45535=>"101011010",
  45536=>"111010100",
  45537=>"100001111",
  45538=>"110110000",
  45539=>"000100101",
  45540=>"001101000",
  45541=>"101010100",
  45542=>"000011011",
  45543=>"000000011",
  45544=>"100110101",
  45545=>"000110110",
  45546=>"000010000",
  45547=>"110110110",
  45548=>"000101110",
  45549=>"000001001",
  45550=>"010010101",
  45551=>"110011110",
  45552=>"111000000",
  45553=>"000001100",
  45554=>"111101010",
  45555=>"001000101",
  45556=>"111000010",
  45557=>"110101100",
  45558=>"011110011",
  45559=>"111011001",
  45560=>"111111110",
  45561=>"101100111",
  45562=>"000110110",
  45563=>"010001101",
  45564=>"010101000",
  45565=>"001000101",
  45566=>"001100101",
  45567=>"011101010",
  45568=>"000001000",
  45569=>"011111001",
  45570=>"110001100",
  45571=>"001010110",
  45572=>"000101000",
  45573=>"111101101",
  45574=>"111100110",
  45575=>"101010001",
  45576=>"001100000",
  45577=>"101011010",
  45578=>"011011001",
  45579=>"111011100",
  45580=>"000000010",
  45581=>"011101010",
  45582=>"011001000",
  45583=>"011011110",
  45584=>"101100110",
  45585=>"010111000",
  45586=>"011110001",
  45587=>"011010100",
  45588=>"011101100",
  45589=>"101000100",
  45590=>"010010101",
  45591=>"010001000",
  45592=>"110011010",
  45593=>"111100000",
  45594=>"000000011",
  45595=>"111110000",
  45596=>"110100110",
  45597=>"100010010",
  45598=>"101111011",
  45599=>"011010100",
  45600=>"010011110",
  45601=>"100001000",
  45602=>"010000000",
  45603=>"001110010",
  45604=>"001100011",
  45605=>"111011101",
  45606=>"110001000",
  45607=>"100110111",
  45608=>"111110000",
  45609=>"001011100",
  45610=>"001001001",
  45611=>"111111000",
  45612=>"101011111",
  45613=>"101000101",
  45614=>"110111000",
  45615=>"011110111",
  45616=>"011100100",
  45617=>"001111110",
  45618=>"001101000",
  45619=>"010101010",
  45620=>"110111000",
  45621=>"100001111",
  45622=>"100000000",
  45623=>"110101011",
  45624=>"000100001",
  45625=>"100110111",
  45626=>"101010010",
  45627=>"010111011",
  45628=>"010001010",
  45629=>"100010010",
  45630=>"101001111",
  45631=>"000011011",
  45632=>"100100010",
  45633=>"111101110",
  45634=>"100011011",
  45635=>"001111011",
  45636=>"011010000",
  45637=>"010011101",
  45638=>"110010000",
  45639=>"111111100",
  45640=>"101010000",
  45641=>"100111111",
  45642=>"001001100",
  45643=>"111111111",
  45644=>"001101111",
  45645=>"111010010",
  45646=>"111000110",
  45647=>"000010111",
  45648=>"100000010",
  45649=>"000110010",
  45650=>"101011001",
  45651=>"010110111",
  45652=>"001000100",
  45653=>"110001111",
  45654=>"011001001",
  45655=>"101111000",
  45656=>"110011110",
  45657=>"111101100",
  45658=>"101101011",
  45659=>"100000010",
  45660=>"110010010",
  45661=>"011100010",
  45662=>"111110010",
  45663=>"010010001",
  45664=>"000111001",
  45665=>"000100011",
  45666=>"001100000",
  45667=>"000011000",
  45668=>"110100010",
  45669=>"011100000",
  45670=>"101111011",
  45671=>"000101110",
  45672=>"011111010",
  45673=>"100001101",
  45674=>"100010110",
  45675=>"010111001",
  45676=>"011110110",
  45677=>"010111110",
  45678=>"010011001",
  45679=>"010000111",
  45680=>"101010000",
  45681=>"001000110",
  45682=>"101001101",
  45683=>"100000000",
  45684=>"001110101",
  45685=>"011000000",
  45686=>"111010010",
  45687=>"111000000",
  45688=>"110011001",
  45689=>"000010000",
  45690=>"110000100",
  45691=>"000010001",
  45692=>"111010100",
  45693=>"110011100",
  45694=>"101000100",
  45695=>"000001010",
  45696=>"001001110",
  45697=>"001110001",
  45698=>"001000100",
  45699=>"111010101",
  45700=>"110100110",
  45701=>"100011011",
  45702=>"010101101",
  45703=>"101010011",
  45704=>"000000101",
  45705=>"101111101",
  45706=>"110111011",
  45707=>"011000111",
  45708=>"011011111",
  45709=>"111110111",
  45710=>"010101010",
  45711=>"011001000",
  45712=>"000111001",
  45713=>"010001010",
  45714=>"000010000",
  45715=>"001001010",
  45716=>"000000110",
  45717=>"101010111",
  45718=>"101010110",
  45719=>"011011100",
  45720=>"111101100",
  45721=>"010110111",
  45722=>"100000010",
  45723=>"000110111",
  45724=>"010111111",
  45725=>"100000101",
  45726=>"111111001",
  45727=>"100010001",
  45728=>"010101000",
  45729=>"111010110",
  45730=>"010010111",
  45731=>"101001100",
  45732=>"101011101",
  45733=>"000000001",
  45734=>"100111100",
  45735=>"000000001",
  45736=>"110010001",
  45737=>"000000110",
  45738=>"100011100",
  45739=>"011010000",
  45740=>"000011010",
  45741=>"111100100",
  45742=>"101011000",
  45743=>"110101001",
  45744=>"110101100",
  45745=>"011101111",
  45746=>"011100001",
  45747=>"001111110",
  45748=>"111010000",
  45749=>"110001110",
  45750=>"011111101",
  45751=>"111000010",
  45752=>"001111111",
  45753=>"111011111",
  45754=>"010111110",
  45755=>"111101101",
  45756=>"000010110",
  45757=>"000010011",
  45758=>"011101111",
  45759=>"111111000",
  45760=>"000111111",
  45761=>"101101011",
  45762=>"000000110",
  45763=>"100011000",
  45764=>"010011001",
  45765=>"101100101",
  45766=>"100011010",
  45767=>"000010111",
  45768=>"000011101",
  45769=>"100000001",
  45770=>"011010011",
  45771=>"001111110",
  45772=>"001000010",
  45773=>"000001000",
  45774=>"000011101",
  45775=>"001110101",
  45776=>"101011000",
  45777=>"000111010",
  45778=>"000111011",
  45779=>"100100000",
  45780=>"001000001",
  45781=>"000000100",
  45782=>"111100101",
  45783=>"010111011",
  45784=>"010111000",
  45785=>"111010001",
  45786=>"000000001",
  45787=>"001000000",
  45788=>"111111110",
  45789=>"011000010",
  45790=>"100011010",
  45791=>"100010101",
  45792=>"101100100",
  45793=>"100001110",
  45794=>"100111101",
  45795=>"110001101",
  45796=>"000101100",
  45797=>"001100101",
  45798=>"111011000",
  45799=>"101001100",
  45800=>"100101100",
  45801=>"010111101",
  45802=>"111101001",
  45803=>"000011111",
  45804=>"110011011",
  45805=>"111100100",
  45806=>"000000000",
  45807=>"000000001",
  45808=>"111001100",
  45809=>"010111011",
  45810=>"000101000",
  45811=>"011101111",
  45812=>"010001011",
  45813=>"001100101",
  45814=>"101100000",
  45815=>"111111101",
  45816=>"000001100",
  45817=>"001111110",
  45818=>"110001111",
  45819=>"011010110",
  45820=>"110110110",
  45821=>"011011110",
  45822=>"110001001",
  45823=>"011100100",
  45824=>"011000000",
  45825=>"011111101",
  45826=>"001100000",
  45827=>"101101111",
  45828=>"000000010",
  45829=>"101010111",
  45830=>"011101000",
  45831=>"010110101",
  45832=>"101000100",
  45833=>"001111100",
  45834=>"110111101",
  45835=>"001010011",
  45836=>"110110111",
  45837=>"001010000",
  45838=>"000101110",
  45839=>"110101001",
  45840=>"010010100",
  45841=>"000000101",
  45842=>"111010111",
  45843=>"011001001",
  45844=>"101110001",
  45845=>"100111111",
  45846=>"100100000",
  45847=>"110111010",
  45848=>"011001111",
  45849=>"000010001",
  45850=>"111011101",
  45851=>"000101010",
  45852=>"000100100",
  45853=>"010100111",
  45854=>"101110001",
  45855=>"111110100",
  45856=>"001011100",
  45857=>"111010011",
  45858=>"000111101",
  45859=>"110000101",
  45860=>"011011000",
  45861=>"001101000",
  45862=>"110111110",
  45863=>"100010101",
  45864=>"101000101",
  45865=>"101101111",
  45866=>"111111100",
  45867=>"011011011",
  45868=>"000010001",
  45869=>"011100011",
  45870=>"111011100",
  45871=>"111010010",
  45872=>"111011110",
  45873=>"101001001",
  45874=>"001000011",
  45875=>"011100010",
  45876=>"000010100",
  45877=>"101101101",
  45878=>"110111110",
  45879=>"010100101",
  45880=>"100000100",
  45881=>"011010001",
  45882=>"000100010",
  45883=>"000001001",
  45884=>"100011111",
  45885=>"110011101",
  45886=>"101101001",
  45887=>"110100101",
  45888=>"110101001",
  45889=>"101010111",
  45890=>"111011011",
  45891=>"101001001",
  45892=>"000110101",
  45893=>"001111100",
  45894=>"010111100",
  45895=>"100001000",
  45896=>"111010000",
  45897=>"100011001",
  45898=>"101100000",
  45899=>"101000111",
  45900=>"011011010",
  45901=>"110110010",
  45902=>"010100100",
  45903=>"000000001",
  45904=>"111010010",
  45905=>"111000001",
  45906=>"111001100",
  45907=>"001010111",
  45908=>"000010000",
  45909=>"110100100",
  45910=>"100100000",
  45911=>"110000100",
  45912=>"100010010",
  45913=>"101111011",
  45914=>"010101010",
  45915=>"111110001",
  45916=>"001100011",
  45917=>"110111110",
  45918=>"111101101",
  45919=>"000010000",
  45920=>"010111001",
  45921=>"001011010",
  45922=>"001100010",
  45923=>"101000000",
  45924=>"000101110",
  45925=>"010101010",
  45926=>"010110010",
  45927=>"110110011",
  45928=>"110100111",
  45929=>"010000111",
  45930=>"111101000",
  45931=>"101101110",
  45932=>"011101110",
  45933=>"101000001",
  45934=>"101000010",
  45935=>"001001011",
  45936=>"000001111",
  45937=>"111000000",
  45938=>"011100110",
  45939=>"010111100",
  45940=>"001011000",
  45941=>"001111111",
  45942=>"100010100",
  45943=>"010001000",
  45944=>"000011001",
  45945=>"100101000",
  45946=>"010100000",
  45947=>"111010000",
  45948=>"000001110",
  45949=>"010000110",
  45950=>"111000011",
  45951=>"001010010",
  45952=>"011010000",
  45953=>"010011000",
  45954=>"001110101",
  45955=>"101100100",
  45956=>"010100111",
  45957=>"011100111",
  45958=>"101100000",
  45959=>"111111000",
  45960=>"010001101",
  45961=>"001110100",
  45962=>"111110110",
  45963=>"010100101",
  45964=>"100100000",
  45965=>"111001100",
  45966=>"000001100",
  45967=>"010001100",
  45968=>"100000001",
  45969=>"110010100",
  45970=>"010000000",
  45971=>"101010100",
  45972=>"001000011",
  45973=>"101101011",
  45974=>"000000010",
  45975=>"111011100",
  45976=>"010000110",
  45977=>"010000111",
  45978=>"001101001",
  45979=>"001000000",
  45980=>"100010000",
  45981=>"100001011",
  45982=>"111001000",
  45983=>"000010100",
  45984=>"110000000",
  45985=>"000100111",
  45986=>"110110100",
  45987=>"010010111",
  45988=>"000100010",
  45989=>"110010000",
  45990=>"000000111",
  45991=>"111010000",
  45992=>"000001100",
  45993=>"001000000",
  45994=>"110111001",
  45995=>"001000110",
  45996=>"110010000",
  45997=>"000110001",
  45998=>"111011100",
  45999=>"001011001",
  46000=>"101100100",
  46001=>"101101100",
  46002=>"001101111",
  46003=>"011001100",
  46004=>"001001011",
  46005=>"101111000",
  46006=>"000111010",
  46007=>"011001110",
  46008=>"110000000",
  46009=>"110111101",
  46010=>"011110111",
  46011=>"000001010",
  46012=>"110111011",
  46013=>"100101000",
  46014=>"101001010",
  46015=>"101101110",
  46016=>"100000111",
  46017=>"011110011",
  46018=>"111010000",
  46019=>"110110100",
  46020=>"010000101",
  46021=>"000110111",
  46022=>"110010000",
  46023=>"101001000",
  46024=>"100001100",
  46025=>"111011000",
  46026=>"001100101",
  46027=>"010000111",
  46028=>"101011001",
  46029=>"011110000",
  46030=>"110100110",
  46031=>"000101100",
  46032=>"100110010",
  46033=>"001011111",
  46034=>"110011111",
  46035=>"011110011",
  46036=>"001101010",
  46037=>"010001111",
  46038=>"000001010",
  46039=>"010000011",
  46040=>"000101101",
  46041=>"110000110",
  46042=>"010101001",
  46043=>"010110011",
  46044=>"001101101",
  46045=>"111010110",
  46046=>"010100000",
  46047=>"101001001",
  46048=>"111110001",
  46049=>"000100000",
  46050=>"111111011",
  46051=>"001011011",
  46052=>"110101000",
  46053=>"011100010",
  46054=>"000100000",
  46055=>"001000010",
  46056=>"011001011",
  46057=>"001011001",
  46058=>"011110000",
  46059=>"100100100",
  46060=>"010111110",
  46061=>"101010010",
  46062=>"110010001",
  46063=>"101011000",
  46064=>"010011001",
  46065=>"000110100",
  46066=>"101100101",
  46067=>"010011100",
  46068=>"010101111",
  46069=>"101110100",
  46070=>"111010000",
  46071=>"011010110",
  46072=>"100000100",
  46073=>"011011011",
  46074=>"000111110",
  46075=>"110001111",
  46076=>"101010000",
  46077=>"101110101",
  46078=>"000000001",
  46079=>"010011110",
  46080=>"111011000",
  46081=>"110101001",
  46082=>"101011100",
  46083=>"001111000",
  46084=>"110100010",
  46085=>"010011111",
  46086=>"001110101",
  46087=>"011111100",
  46088=>"111011101",
  46089=>"010101100",
  46090=>"111110100",
  46091=>"011011111",
  46092=>"101001000",
  46093=>"010101111",
  46094=>"100100011",
  46095=>"011001100",
  46096=>"100100010",
  46097=>"010000011",
  46098=>"000001010",
  46099=>"001001110",
  46100=>"100001101",
  46101=>"101110011",
  46102=>"000001001",
  46103=>"000010101",
  46104=>"111010000",
  46105=>"011010000",
  46106=>"110010100",
  46107=>"011100101",
  46108=>"110111111",
  46109=>"100011111",
  46110=>"100010000",
  46111=>"011110010",
  46112=>"110110111",
  46113=>"001000111",
  46114=>"011111011",
  46115=>"011111100",
  46116=>"000110000",
  46117=>"100000001",
  46118=>"001101010",
  46119=>"011010110",
  46120=>"111001110",
  46121=>"110100001",
  46122=>"010111001",
  46123=>"010110001",
  46124=>"111111101",
  46125=>"011101011",
  46126=>"001111011",
  46127=>"011011110",
  46128=>"001001011",
  46129=>"001101101",
  46130=>"000110011",
  46131=>"011001010",
  46132=>"111100010",
  46133=>"100011110",
  46134=>"111111111",
  46135=>"110101101",
  46136=>"000100001",
  46137=>"100110101",
  46138=>"010000001",
  46139=>"101010000",
  46140=>"011010010",
  46141=>"100110110",
  46142=>"100110110",
  46143=>"000010010",
  46144=>"111100111",
  46145=>"000001101",
  46146=>"011011000",
  46147=>"100011101",
  46148=>"000001010",
  46149=>"010000001",
  46150=>"010111110",
  46151=>"001111010",
  46152=>"000000000",
  46153=>"011010000",
  46154=>"001110011",
  46155=>"010111000",
  46156=>"000011001",
  46157=>"011110001",
  46158=>"010010111",
  46159=>"010111000",
  46160=>"101010000",
  46161=>"111000100",
  46162=>"001010110",
  46163=>"011111011",
  46164=>"001010110",
  46165=>"011010001",
  46166=>"111100111",
  46167=>"011101010",
  46168=>"110111011",
  46169=>"010010011",
  46170=>"100001001",
  46171=>"010100001",
  46172=>"001011000",
  46173=>"000110011",
  46174=>"111111010",
  46175=>"000001101",
  46176=>"010001101",
  46177=>"001001011",
  46178=>"101011011",
  46179=>"010010001",
  46180=>"111000000",
  46181=>"100001000",
  46182=>"100101010",
  46183=>"011111101",
  46184=>"100001110",
  46185=>"100010011",
  46186=>"000110001",
  46187=>"110110101",
  46188=>"101011010",
  46189=>"000101010",
  46190=>"011010000",
  46191=>"100010000",
  46192=>"101001101",
  46193=>"011001100",
  46194=>"011011101",
  46195=>"101001010",
  46196=>"001001111",
  46197=>"001111010",
  46198=>"000101000",
  46199=>"111111111",
  46200=>"000111100",
  46201=>"110110011",
  46202=>"000001000",
  46203=>"001000101",
  46204=>"100011111",
  46205=>"100100100",
  46206=>"011101110",
  46207=>"101101101",
  46208=>"100000011",
  46209=>"000100110",
  46210=>"110011111",
  46211=>"100101001",
  46212=>"010011111",
  46213=>"101010010",
  46214=>"111110000",
  46215=>"001010010",
  46216=>"001110101",
  46217=>"101111110",
  46218=>"111100101",
  46219=>"101000100",
  46220=>"100110110",
  46221=>"001110010",
  46222=>"001000101",
  46223=>"000001101",
  46224=>"110110100",
  46225=>"010101000",
  46226=>"111011010",
  46227=>"000111111",
  46228=>"000110100",
  46229=>"001010101",
  46230=>"110111101",
  46231=>"100000101",
  46232=>"111100101",
  46233=>"000111010",
  46234=>"001110101",
  46235=>"110001100",
  46236=>"000000010",
  46237=>"100001100",
  46238=>"011110011",
  46239=>"110110010",
  46240=>"110111011",
  46241=>"110010011",
  46242=>"010010010",
  46243=>"011101100",
  46244=>"110011111",
  46245=>"110111010",
  46246=>"001111000",
  46247=>"001000010",
  46248=>"010000001",
  46249=>"001011000",
  46250=>"011111011",
  46251=>"000100110",
  46252=>"001110101",
  46253=>"010001001",
  46254=>"011111011",
  46255=>"011110111",
  46256=>"110011101",
  46257=>"111100010",
  46258=>"111101011",
  46259=>"000011001",
  46260=>"001110001",
  46261=>"001101111",
  46262=>"001110000",
  46263=>"011111111",
  46264=>"010001100",
  46265=>"110101011",
  46266=>"000101000",
  46267=>"001101110",
  46268=>"000100110",
  46269=>"001010110",
  46270=>"011111000",
  46271=>"001010111",
  46272=>"110111100",
  46273=>"111100110",
  46274=>"001001101",
  46275=>"111101110",
  46276=>"000011110",
  46277=>"001100010",
  46278=>"101111111",
  46279=>"111000111",
  46280=>"001100111",
  46281=>"110101010",
  46282=>"111111110",
  46283=>"001000000",
  46284=>"000001000",
  46285=>"010111110",
  46286=>"101110000",
  46287=>"100110011",
  46288=>"101101110",
  46289=>"111010000",
  46290=>"100011111",
  46291=>"110011011",
  46292=>"011100011",
  46293=>"100000100",
  46294=>"100010101",
  46295=>"111010000",
  46296=>"001110110",
  46297=>"011101110",
  46298=>"011101111",
  46299=>"110010011",
  46300=>"011111010",
  46301=>"101001001",
  46302=>"001110001",
  46303=>"000010000",
  46304=>"111100111",
  46305=>"000000101",
  46306=>"000110111",
  46307=>"000010111",
  46308=>"110001000",
  46309=>"000001100",
  46310=>"110100100",
  46311=>"000101011",
  46312=>"110101011",
  46313=>"100011010",
  46314=>"100110000",
  46315=>"001001000",
  46316=>"001110011",
  46317=>"101010111",
  46318=>"110001010",
  46319=>"100100100",
  46320=>"100111111",
  46321=>"000001111",
  46322=>"010111100",
  46323=>"001100001",
  46324=>"111011110",
  46325=>"111111011",
  46326=>"001110010",
  46327=>"101111100",
  46328=>"101010010",
  46329=>"100101111",
  46330=>"100010000",
  46331=>"100111111",
  46332=>"110110010",
  46333=>"000101011",
  46334=>"111111011",
  46335=>"100000001",
  46336=>"010111101",
  46337=>"010111100",
  46338=>"000111101",
  46339=>"100011000",
  46340=>"000101000",
  46341=>"010000000",
  46342=>"000001000",
  46343=>"001101101",
  46344=>"111101101",
  46345=>"001000111",
  46346=>"000100110",
  46347=>"111000110",
  46348=>"010001000",
  46349=>"010000001",
  46350=>"111000100",
  46351=>"100000110",
  46352=>"111100011",
  46353=>"110000010",
  46354=>"001101000",
  46355=>"011111001",
  46356=>"100110001",
  46357=>"100011111",
  46358=>"110101010",
  46359=>"010101001",
  46360=>"011100011",
  46361=>"100010110",
  46362=>"000010110",
  46363=>"011110100",
  46364=>"111111001",
  46365=>"011110011",
  46366=>"001111011",
  46367=>"000101000",
  46368=>"001000000",
  46369=>"110111111",
  46370=>"000111110",
  46371=>"110000101",
  46372=>"000010100",
  46373=>"011100110",
  46374=>"010100100",
  46375=>"011000011",
  46376=>"100100100",
  46377=>"100011100",
  46378=>"001111111",
  46379=>"111101011",
  46380=>"001111000",
  46381=>"011000101",
  46382=>"010000101",
  46383=>"100010110",
  46384=>"110110111",
  46385=>"100010101",
  46386=>"101110111",
  46387=>"011000100",
  46388=>"111000100",
  46389=>"110110000",
  46390=>"101101010",
  46391=>"000001100",
  46392=>"110110000",
  46393=>"111001000",
  46394=>"010001101",
  46395=>"011110110",
  46396=>"000010000",
  46397=>"001100111",
  46398=>"001011100",
  46399=>"100111110",
  46400=>"100100011",
  46401=>"001110111",
  46402=>"010110001",
  46403=>"101111000",
  46404=>"101100000",
  46405=>"110001111",
  46406=>"101011001",
  46407=>"011011100",
  46408=>"010000110",
  46409=>"001101111",
  46410=>"000001010",
  46411=>"011001000",
  46412=>"110101101",
  46413=>"101001010",
  46414=>"000111110",
  46415=>"110100011",
  46416=>"100010101",
  46417=>"111010011",
  46418=>"011000100",
  46419=>"010110000",
  46420=>"000000010",
  46421=>"011111100",
  46422=>"010111111",
  46423=>"010100110",
  46424=>"011001111",
  46425=>"001100010",
  46426=>"110100101",
  46427=>"101010011",
  46428=>"011101011",
  46429=>"011010111",
  46430=>"000101000",
  46431=>"111010101",
  46432=>"100100110",
  46433=>"001110111",
  46434=>"110110001",
  46435=>"000010110",
  46436=>"000100101",
  46437=>"011101110",
  46438=>"110100010",
  46439=>"111001010",
  46440=>"110111000",
  46441=>"000100110",
  46442=>"000011111",
  46443=>"000110110",
  46444=>"111111111",
  46445=>"011111100",
  46446=>"111100000",
  46447=>"110101001",
  46448=>"110110101",
  46449=>"001001011",
  46450=>"101101001",
  46451=>"010111000",
  46452=>"111010000",
  46453=>"000001011",
  46454=>"100101001",
  46455=>"011101101",
  46456=>"100000110",
  46457=>"100110001",
  46458=>"011110010",
  46459=>"001000011",
  46460=>"001101101",
  46461=>"101000000",
  46462=>"111110001",
  46463=>"001001001",
  46464=>"011010001",
  46465=>"100110111",
  46466=>"001010101",
  46467=>"100100101",
  46468=>"110110110",
  46469=>"011100100",
  46470=>"000001011",
  46471=>"000001011",
  46472=>"010110110",
  46473=>"101101011",
  46474=>"110101100",
  46475=>"111101000",
  46476=>"011000111",
  46477=>"000000111",
  46478=>"111111101",
  46479=>"001101101",
  46480=>"001001011",
  46481=>"111110000",
  46482=>"011010010",
  46483=>"111011010",
  46484=>"001110011",
  46485=>"111000000",
  46486=>"011111101",
  46487=>"001101101",
  46488=>"111100010",
  46489=>"010000101",
  46490=>"011101010",
  46491=>"111001100",
  46492=>"111011101",
  46493=>"111101000",
  46494=>"010001100",
  46495=>"100101011",
  46496=>"100110101",
  46497=>"011111111",
  46498=>"101000011",
  46499=>"011011001",
  46500=>"111010101",
  46501=>"000011110",
  46502=>"101011010",
  46503=>"000000110",
  46504=>"001111001",
  46505=>"011010001",
  46506=>"100110010",
  46507=>"110010110",
  46508=>"111110001",
  46509=>"000111010",
  46510=>"100001001",
  46511=>"101010000",
  46512=>"100101101",
  46513=>"010000001",
  46514=>"111010011",
  46515=>"101000110",
  46516=>"010111001",
  46517=>"111000010",
  46518=>"011011000",
  46519=>"010011111",
  46520=>"111001110",
  46521=>"001000010",
  46522=>"110010100",
  46523=>"001100011",
  46524=>"001111001",
  46525=>"111000100",
  46526=>"110010111",
  46527=>"101010100",
  46528=>"000001010",
  46529=>"100010110",
  46530=>"011100111",
  46531=>"100101111",
  46532=>"010010110",
  46533=>"000000001",
  46534=>"011010010",
  46535=>"111000000",
  46536=>"111100011",
  46537=>"010111111",
  46538=>"110010101",
  46539=>"001011000",
  46540=>"000010000",
  46541=>"011001010",
  46542=>"110011101",
  46543=>"111100011",
  46544=>"100111111",
  46545=>"000111011",
  46546=>"011111000",
  46547=>"110000100",
  46548=>"111011111",
  46549=>"001100111",
  46550=>"100110001",
  46551=>"001000000",
  46552=>"010110010",
  46553=>"110100100",
  46554=>"001110000",
  46555=>"101100010",
  46556=>"000011000",
  46557=>"100001000",
  46558=>"111001100",
  46559=>"011010000",
  46560=>"110011001",
  46561=>"101010111",
  46562=>"010011111",
  46563=>"101111010",
  46564=>"000001010",
  46565=>"110111101",
  46566=>"110100000",
  46567=>"000000011",
  46568=>"111111111",
  46569=>"010011000",
  46570=>"111011101",
  46571=>"010110011",
  46572=>"111010010",
  46573=>"111001101",
  46574=>"111010010",
  46575=>"101010010",
  46576=>"110010001",
  46577=>"110110011",
  46578=>"011010101",
  46579=>"111101011",
  46580=>"101001110",
  46581=>"111111000",
  46582=>"111110111",
  46583=>"011000110",
  46584=>"001101011",
  46585=>"110000101",
  46586=>"010101100",
  46587=>"101110100",
  46588=>"111000000",
  46589=>"101001101",
  46590=>"110111100",
  46591=>"100001111",
  46592=>"101011001",
  46593=>"110110001",
  46594=>"111110100",
  46595=>"010011110",
  46596=>"001011100",
  46597=>"100100001",
  46598=>"011001110",
  46599=>"100000101",
  46600=>"101111101",
  46601=>"111110101",
  46602=>"001110110",
  46603=>"001001110",
  46604=>"111100101",
  46605=>"011101011",
  46606=>"001110000",
  46607=>"100110011",
  46608=>"101001011",
  46609=>"010101010",
  46610=>"110000111",
  46611=>"001111010",
  46612=>"000100110",
  46613=>"100011000",
  46614=>"110011100",
  46615=>"100100000",
  46616=>"011110010",
  46617=>"010000010",
  46618=>"111000010",
  46619=>"000000000",
  46620=>"001000011",
  46621=>"101100110",
  46622=>"000100111",
  46623=>"110111100",
  46624=>"010011101",
  46625=>"110001001",
  46626=>"010010000",
  46627=>"001000111",
  46628=>"000001110",
  46629=>"011101110",
  46630=>"111001010",
  46631=>"001010011",
  46632=>"000000000",
  46633=>"111111011",
  46634=>"010010011",
  46635=>"001011110",
  46636=>"100010101",
  46637=>"100000111",
  46638=>"100100111",
  46639=>"001111110",
  46640=>"100001000",
  46641=>"111000001",
  46642=>"000110111",
  46643=>"011010110",
  46644=>"000100011",
  46645=>"010010011",
  46646=>"011010101",
  46647=>"011001111",
  46648=>"000010011",
  46649=>"101110010",
  46650=>"010010101",
  46651=>"011001100",
  46652=>"100100110",
  46653=>"011001010",
  46654=>"010100010",
  46655=>"111011011",
  46656=>"001000111",
  46657=>"100101001",
  46658=>"010110010",
  46659=>"011110001",
  46660=>"100100101",
  46661=>"000010111",
  46662=>"101000101",
  46663=>"110101001",
  46664=>"011000100",
  46665=>"100100101",
  46666=>"110010011",
  46667=>"010000010",
  46668=>"110110110",
  46669=>"010100111",
  46670=>"000110001",
  46671=>"101100100",
  46672=>"101001010",
  46673=>"111110001",
  46674=>"011000100",
  46675=>"010011011",
  46676=>"101111110",
  46677=>"111000101",
  46678=>"011100010",
  46679=>"110110010",
  46680=>"101101111",
  46681=>"111101101",
  46682=>"011011111",
  46683=>"000001100",
  46684=>"010011110",
  46685=>"111110001",
  46686=>"011111111",
  46687=>"100010010",
  46688=>"011110000",
  46689=>"010110101",
  46690=>"000000000",
  46691=>"001111100",
  46692=>"000000101",
  46693=>"100000010",
  46694=>"101110101",
  46695=>"101100001",
  46696=>"111110111",
  46697=>"011111011",
  46698=>"110010010",
  46699=>"001111100",
  46700=>"110100010",
  46701=>"001010010",
  46702=>"110110111",
  46703=>"000101101",
  46704=>"001111110",
  46705=>"001001101",
  46706=>"110100111",
  46707=>"011100010",
  46708=>"000110011",
  46709=>"010101011",
  46710=>"101010000",
  46711=>"000101111",
  46712=>"100011000",
  46713=>"000011001",
  46714=>"001110000",
  46715=>"110011100",
  46716=>"000011101",
  46717=>"001110111",
  46718=>"011011100",
  46719=>"010001111",
  46720=>"001110111",
  46721=>"100000011",
  46722=>"110111010",
  46723=>"101011010",
  46724=>"101010001",
  46725=>"011000001",
  46726=>"001001110",
  46727=>"111110110",
  46728=>"110101000",
  46729=>"011011110",
  46730=>"000111010",
  46731=>"000101010",
  46732=>"010001100",
  46733=>"100100010",
  46734=>"100110011",
  46735=>"111010010",
  46736=>"111011000",
  46737=>"100000010",
  46738=>"110011100",
  46739=>"010100100",
  46740=>"100111001",
  46741=>"101001011",
  46742=>"101010010",
  46743=>"110001111",
  46744=>"001011110",
  46745=>"111000111",
  46746=>"000111111",
  46747=>"001101010",
  46748=>"110101000",
  46749=>"100110000",
  46750=>"100100000",
  46751=>"001110100",
  46752=>"101111010",
  46753=>"010010001",
  46754=>"110001010",
  46755=>"011000110",
  46756=>"111011010",
  46757=>"011001111",
  46758=>"001010010",
  46759=>"000000001",
  46760=>"011001101",
  46761=>"011011100",
  46762=>"011100000",
  46763=>"011011100",
  46764=>"001100110",
  46765=>"011001111",
  46766=>"100001111",
  46767=>"111010010",
  46768=>"000011111",
  46769=>"011001010",
  46770=>"010101100",
  46771=>"110000000",
  46772=>"111100111",
  46773=>"111011110",
  46774=>"000110010",
  46775=>"110010001",
  46776=>"100110010",
  46777=>"000000100",
  46778=>"101011000",
  46779=>"001000011",
  46780=>"101100111",
  46781=>"001000101",
  46782=>"111100100",
  46783=>"000010111",
  46784=>"101001011",
  46785=>"001100100",
  46786=>"010000100",
  46787=>"010010101",
  46788=>"000110010",
  46789=>"000010100",
  46790=>"000100110",
  46791=>"001010000",
  46792=>"111101100",
  46793=>"101001011",
  46794=>"010111010",
  46795=>"111100111",
  46796=>"011010011",
  46797=>"101110110",
  46798=>"100011101",
  46799=>"011100111",
  46800=>"111111010",
  46801=>"101101101",
  46802=>"101011110",
  46803=>"101101010",
  46804=>"100011011",
  46805=>"001110101",
  46806=>"110110010",
  46807=>"110010000",
  46808=>"000111101",
  46809=>"101011010",
  46810=>"011011101",
  46811=>"011010111",
  46812=>"000110000",
  46813=>"111001011",
  46814=>"000100101",
  46815=>"000001000",
  46816=>"110110011",
  46817=>"101000100",
  46818=>"101101010",
  46819=>"100010000",
  46820=>"110000011",
  46821=>"011110111",
  46822=>"011000100",
  46823=>"010011011",
  46824=>"011010101",
  46825=>"010111001",
  46826=>"000000111",
  46827=>"111000100",
  46828=>"000000100",
  46829=>"011011100",
  46830=>"011100101",
  46831=>"111100000",
  46832=>"100011001",
  46833=>"000001100",
  46834=>"010101111",
  46835=>"011111110",
  46836=>"101000111",
  46837=>"011000011",
  46838=>"011111000",
  46839=>"001010001",
  46840=>"111000010",
  46841=>"110000001",
  46842=>"100001011",
  46843=>"011001010",
  46844=>"101111010",
  46845=>"010111011",
  46846=>"101111110",
  46847=>"010010010",
  46848=>"011011011",
  46849=>"100100110",
  46850=>"111111010",
  46851=>"111111111",
  46852=>"001111000",
  46853=>"101100000",
  46854=>"001010010",
  46855=>"000110000",
  46856=>"001001000",
  46857=>"000110000",
  46858=>"111111010",
  46859=>"101000101",
  46860=>"101110000",
  46861=>"001100001",
  46862=>"000100101",
  46863=>"111000101",
  46864=>"001000001",
  46865=>"100111111",
  46866=>"101011010",
  46867=>"011100101",
  46868=>"010011001",
  46869=>"110110111",
  46870=>"011011011",
  46871=>"000100111",
  46872=>"010011011",
  46873=>"010000000",
  46874=>"000100001",
  46875=>"001011000",
  46876=>"001111000",
  46877=>"101010000",
  46878=>"111011001",
  46879=>"111000100",
  46880=>"000101100",
  46881=>"011000110",
  46882=>"000010010",
  46883=>"010111111",
  46884=>"000100000",
  46885=>"110110010",
  46886=>"010001111",
  46887=>"100110100",
  46888=>"100001111",
  46889=>"010010111",
  46890=>"100010001",
  46891=>"001010101",
  46892=>"110010101",
  46893=>"010100010",
  46894=>"110010010",
  46895=>"101010010",
  46896=>"101110000",
  46897=>"001111101",
  46898=>"101000000",
  46899=>"100001110",
  46900=>"011010010",
  46901=>"110101010",
  46902=>"100011011",
  46903=>"011010001",
  46904=>"001010111",
  46905=>"101010000",
  46906=>"100110010",
  46907=>"100101111",
  46908=>"000100000",
  46909=>"000001010",
  46910=>"100000100",
  46911=>"010011010",
  46912=>"110011010",
  46913=>"001000111",
  46914=>"010100101",
  46915=>"011110100",
  46916=>"110100111",
  46917=>"010011000",
  46918=>"001101010",
  46919=>"111111101",
  46920=>"010100011",
  46921=>"010010011",
  46922=>"000111010",
  46923=>"100111111",
  46924=>"110011111",
  46925=>"001101110",
  46926=>"101110011",
  46927=>"110001101",
  46928=>"000100011",
  46929=>"110000000",
  46930=>"111011010",
  46931=>"000010101",
  46932=>"111010100",
  46933=>"011111001",
  46934=>"001000101",
  46935=>"010110000",
  46936=>"000111001",
  46937=>"110111100",
  46938=>"110100011",
  46939=>"001100111",
  46940=>"100101111",
  46941=>"000100110",
  46942=>"110000010",
  46943=>"110110101",
  46944=>"101010111",
  46945=>"100100011",
  46946=>"000000111",
  46947=>"010101110",
  46948=>"101100010",
  46949=>"010001101",
  46950=>"111010101",
  46951=>"010001001",
  46952=>"011101101",
  46953=>"100101101",
  46954=>"110010110",
  46955=>"000001111",
  46956=>"010010010",
  46957=>"101100001",
  46958=>"001111010",
  46959=>"100101010",
  46960=>"010111011",
  46961=>"010010111",
  46962=>"111111100",
  46963=>"101010000",
  46964=>"000101101",
  46965=>"100011111",
  46966=>"011100110",
  46967=>"001100110",
  46968=>"111111100",
  46969=>"110000011",
  46970=>"000110001",
  46971=>"101110000",
  46972=>"110010000",
  46973=>"111010110",
  46974=>"011001001",
  46975=>"001101010",
  46976=>"000101111",
  46977=>"101010100",
  46978=>"100011011",
  46979=>"011011110",
  46980=>"011010111",
  46981=>"110000111",
  46982=>"100101001",
  46983=>"010000111",
  46984=>"111100100",
  46985=>"110110000",
  46986=>"100111100",
  46987=>"111110001",
  46988=>"001001110",
  46989=>"111010010",
  46990=>"110010101",
  46991=>"000000010",
  46992=>"000110100",
  46993=>"101001101",
  46994=>"101110111",
  46995=>"010100100",
  46996=>"110100110",
  46997=>"001111110",
  46998=>"001110100",
  46999=>"111000001",
  47000=>"000000100",
  47001=>"011110000",
  47002=>"110011111",
  47003=>"010111011",
  47004=>"000010101",
  47005=>"011001011",
  47006=>"110110011",
  47007=>"001010010",
  47008=>"101000000",
  47009=>"010101110",
  47010=>"111100100",
  47011=>"101110100",
  47012=>"111010001",
  47013=>"010110111",
  47014=>"101000000",
  47015=>"010101011",
  47016=>"111110000",
  47017=>"011010011",
  47018=>"011100010",
  47019=>"101010110",
  47020=>"001001111",
  47021=>"100000110",
  47022=>"111010100",
  47023=>"010100111",
  47024=>"000101011",
  47025=>"111000011",
  47026=>"001111010",
  47027=>"000011001",
  47028=>"011010111",
  47029=>"001110110",
  47030=>"001111100",
  47031=>"001111101",
  47032=>"010000011",
  47033=>"100110000",
  47034=>"010011011",
  47035=>"101001011",
  47036=>"101101111",
  47037=>"000001011",
  47038=>"111011110",
  47039=>"010100101",
  47040=>"001001000",
  47041=>"010101000",
  47042=>"100010011",
  47043=>"101010110",
  47044=>"000101110",
  47045=>"111010111",
  47046=>"111011011",
  47047=>"010010110",
  47048=>"111000110",
  47049=>"001111110",
  47050=>"100001011",
  47051=>"100001000",
  47052=>"101001101",
  47053=>"010111101",
  47054=>"011101010",
  47055=>"000011111",
  47056=>"110000110",
  47057=>"110011110",
  47058=>"101101001",
  47059=>"101110100",
  47060=>"010001111",
  47061=>"011001001",
  47062=>"001001101",
  47063=>"101101010",
  47064=>"001101000",
  47065=>"000111110",
  47066=>"110110010",
  47067=>"111011010",
  47068=>"100100000",
  47069=>"100100011",
  47070=>"010010111",
  47071=>"010110101",
  47072=>"010111011",
  47073=>"000010110",
  47074=>"011001010",
  47075=>"111000111",
  47076=>"111101000",
  47077=>"101100111",
  47078=>"000110110",
  47079=>"000100001",
  47080=>"100111000",
  47081=>"101110000",
  47082=>"101001010",
  47083=>"010111001",
  47084=>"011011010",
  47085=>"111101001",
  47086=>"011011110",
  47087=>"111110000",
  47088=>"001011010",
  47089=>"011100100",
  47090=>"000101010",
  47091=>"100001001",
  47092=>"111111000",
  47093=>"001010100",
  47094=>"110101000",
  47095=>"010001100",
  47096=>"010111001",
  47097=>"111110001",
  47098=>"110111111",
  47099=>"110110001",
  47100=>"110010000",
  47101=>"001001000",
  47102=>"000001010",
  47103=>"001010000",
  47104=>"001000000",
  47105=>"111011010",
  47106=>"010000000",
  47107=>"001110000",
  47108=>"000000111",
  47109=>"101101011",
  47110=>"010010001",
  47111=>"011001101",
  47112=>"110100001",
  47113=>"110000001",
  47114=>"100111110",
  47115=>"000101001",
  47116=>"110010101",
  47117=>"111111000",
  47118=>"101010001",
  47119=>"010111010",
  47120=>"010101110",
  47121=>"011010011",
  47122=>"001001000",
  47123=>"100100001",
  47124=>"111001111",
  47125=>"110001001",
  47126=>"111000001",
  47127=>"000000000",
  47128=>"100001110",
  47129=>"010010110",
  47130=>"111100111",
  47131=>"111010000",
  47132=>"011001100",
  47133=>"010110101",
  47134=>"111010000",
  47135=>"110110111",
  47136=>"010111010",
  47137=>"001101010",
  47138=>"110001000",
  47139=>"000111111",
  47140=>"110001001",
  47141=>"010110110",
  47142=>"111000100",
  47143=>"001010011",
  47144=>"101010111",
  47145=>"010010111",
  47146=>"111101111",
  47147=>"011111000",
  47148=>"110010101",
  47149=>"010110011",
  47150=>"000110011",
  47151=>"010101001",
  47152=>"001001101",
  47153=>"011100000",
  47154=>"001010000",
  47155=>"100110010",
  47156=>"001000101",
  47157=>"011010110",
  47158=>"010111100",
  47159=>"100010111",
  47160=>"011100100",
  47161=>"001010000",
  47162=>"010001000",
  47163=>"101001011",
  47164=>"101100101",
  47165=>"010011100",
  47166=>"001000111",
  47167=>"110001000",
  47168=>"110110101",
  47169=>"010001001",
  47170=>"010110001",
  47171=>"001001111",
  47172=>"101111100",
  47173=>"000011010",
  47174=>"000001001",
  47175=>"111000001",
  47176=>"010001100",
  47177=>"010000100",
  47178=>"000000111",
  47179=>"111101100",
  47180=>"010000000",
  47181=>"100110010",
  47182=>"110010000",
  47183=>"001010010",
  47184=>"000110101",
  47185=>"011000010",
  47186=>"110111010",
  47187=>"101111100",
  47188=>"001010110",
  47189=>"011001101",
  47190=>"111001010",
  47191=>"011011110",
  47192=>"100011000",
  47193=>"001111010",
  47194=>"100001100",
  47195=>"101010000",
  47196=>"010111000",
  47197=>"000001001",
  47198=>"000100100",
  47199=>"101010101",
  47200=>"001010110",
  47201=>"101011001",
  47202=>"110111011",
  47203=>"001100111",
  47204=>"110101110",
  47205=>"000011110",
  47206=>"010101100",
  47207=>"100111101",
  47208=>"011011100",
  47209=>"111001111",
  47210=>"011101110",
  47211=>"010000010",
  47212=>"110000010",
  47213=>"111110111",
  47214=>"001010100",
  47215=>"100011100",
  47216=>"001110111",
  47217=>"000111110",
  47218=>"011111111",
  47219=>"111000011",
  47220=>"011011110",
  47221=>"000100011",
  47222=>"010010001",
  47223=>"000010111",
  47224=>"110001010",
  47225=>"001011011",
  47226=>"001101000",
  47227=>"000011011",
  47228=>"100101100",
  47229=>"110001001",
  47230=>"000110101",
  47231=>"001101001",
  47232=>"000110010",
  47233=>"101100100",
  47234=>"110101000",
  47235=>"111011110",
  47236=>"100100000",
  47237=>"001101011",
  47238=>"001010110",
  47239=>"000110111",
  47240=>"010011110",
  47241=>"111000011",
  47242=>"100010000",
  47243=>"111110000",
  47244=>"111001111",
  47245=>"000111110",
  47246=>"101000101",
  47247=>"001001000",
  47248=>"100100000",
  47249=>"110010101",
  47250=>"100101111",
  47251=>"100011010",
  47252=>"111000110",
  47253=>"100100101",
  47254=>"011010110",
  47255=>"001010111",
  47256=>"100000011",
  47257=>"111001101",
  47258=>"000100000",
  47259=>"111010110",
  47260=>"001110101",
  47261=>"111000101",
  47262=>"011001010",
  47263=>"000110010",
  47264=>"111101001",
  47265=>"001001000",
  47266=>"110011000",
  47267=>"001000110",
  47268=>"110100111",
  47269=>"011010110",
  47270=>"000000010",
  47271=>"001001100",
  47272=>"111010001",
  47273=>"111010011",
  47274=>"000000011",
  47275=>"111100000",
  47276=>"100001001",
  47277=>"000100101",
  47278=>"010111001",
  47279=>"100110000",
  47280=>"100111100",
  47281=>"000001001",
  47282=>"001101101",
  47283=>"001100111",
  47284=>"010100101",
  47285=>"110100010",
  47286=>"111101101",
  47287=>"111110100",
  47288=>"001101011",
  47289=>"101111011",
  47290=>"110111111",
  47291=>"101010010",
  47292=>"110000011",
  47293=>"101101101",
  47294=>"110010000",
  47295=>"001101010",
  47296=>"011100100",
  47297=>"100101000",
  47298=>"011101110",
  47299=>"011001000",
  47300=>"001000010",
  47301=>"110010110",
  47302=>"100110111",
  47303=>"011101011",
  47304=>"111100101",
  47305=>"101010001",
  47306=>"011101011",
  47307=>"011010110",
  47308=>"011101110",
  47309=>"111101010",
  47310=>"110101000",
  47311=>"011011011",
  47312=>"111000010",
  47313=>"111111101",
  47314=>"000111100",
  47315=>"010011111",
  47316=>"010010111",
  47317=>"010000100",
  47318=>"010001010",
  47319=>"010110001",
  47320=>"101111101",
  47321=>"011001100",
  47322=>"111110010",
  47323=>"001011100",
  47324=>"011110100",
  47325=>"010000001",
  47326=>"000110110",
  47327=>"111100000",
  47328=>"010011101",
  47329=>"101110011",
  47330=>"010000100",
  47331=>"000010000",
  47332=>"110111110",
  47333=>"000000111",
  47334=>"101010101",
  47335=>"101001110",
  47336=>"010100010",
  47337=>"001110011",
  47338=>"010111111",
  47339=>"000100101",
  47340=>"110010000",
  47341=>"001001000",
  47342=>"001001110",
  47343=>"011010001",
  47344=>"101100100",
  47345=>"010001010",
  47346=>"011001000",
  47347=>"111101110",
  47348=>"101010000",
  47349=>"000010000",
  47350=>"011110001",
  47351=>"000101000",
  47352=>"010100000",
  47353=>"110101110",
  47354=>"000111010",
  47355=>"110000100",
  47356=>"011111111",
  47357=>"001000100",
  47358=>"001100011",
  47359=>"000110101",
  47360=>"011110101",
  47361=>"111100000",
  47362=>"101010100",
  47363=>"110110110",
  47364=>"100111000",
  47365=>"110100111",
  47366=>"011011110",
  47367=>"101101010",
  47368=>"101001110",
  47369=>"011100111",
  47370=>"100100101",
  47371=>"101001011",
  47372=>"111101001",
  47373=>"100011111",
  47374=>"101110010",
  47375=>"010110100",
  47376=>"111101010",
  47377=>"111101110",
  47378=>"101101100",
  47379=>"110110001",
  47380=>"100011100",
  47381=>"010110110",
  47382=>"000111110",
  47383=>"101110101",
  47384=>"111011101",
  47385=>"101001111",
  47386=>"011101011",
  47387=>"011111111",
  47388=>"101011100",
  47389=>"010101110",
  47390=>"111111110",
  47391=>"001100001",
  47392=>"100101101",
  47393=>"110111001",
  47394=>"010001010",
  47395=>"010000011",
  47396=>"111101011",
  47397=>"101100011",
  47398=>"010101011",
  47399=>"111110101",
  47400=>"001010101",
  47401=>"010011110",
  47402=>"111001010",
  47403=>"001010110",
  47404=>"100001010",
  47405=>"111100111",
  47406=>"111000100",
  47407=>"100000101",
  47408=>"111010100",
  47409=>"011010010",
  47410=>"111000010",
  47411=>"100001100",
  47412=>"100000011",
  47413=>"001010010",
  47414=>"011110011",
  47415=>"111110110",
  47416=>"100110111",
  47417=>"111101110",
  47418=>"000101010",
  47419=>"110110101",
  47420=>"001111111",
  47421=>"011110110",
  47422=>"000111001",
  47423=>"100101000",
  47424=>"100100110",
  47425=>"101111110",
  47426=>"101101100",
  47427=>"011101000",
  47428=>"011010110",
  47429=>"101100110",
  47430=>"010100011",
  47431=>"001001010",
  47432=>"111100010",
  47433=>"010000100",
  47434=>"110010000",
  47435=>"100011101",
  47436=>"101000000",
  47437=>"000111111",
  47438=>"011011010",
  47439=>"000101001",
  47440=>"111101011",
  47441=>"100100001",
  47442=>"010101000",
  47443=>"011000000",
  47444=>"101100011",
  47445=>"001001010",
  47446=>"010110010",
  47447=>"000111101",
  47448=>"011101100",
  47449=>"110100101",
  47450=>"100011111",
  47451=>"110011001",
  47452=>"000011100",
  47453=>"000101011",
  47454=>"000011110",
  47455=>"001001111",
  47456=>"101100000",
  47457=>"001100011",
  47458=>"101001111",
  47459=>"100011110",
  47460=>"011111010",
  47461=>"010011111",
  47462=>"010001110",
  47463=>"111011101",
  47464=>"110000001",
  47465=>"011011110",
  47466=>"011010000",
  47467=>"100011110",
  47468=>"000101100",
  47469=>"110110100",
  47470=>"010000010",
  47471=>"010011011",
  47472=>"010100000",
  47473=>"011100101",
  47474=>"000010110",
  47475=>"000001010",
  47476=>"111101011",
  47477=>"011010101",
  47478=>"011001100",
  47479=>"001100011",
  47480=>"100011010",
  47481=>"001001011",
  47482=>"101100100",
  47483=>"010111000",
  47484=>"100001000",
  47485=>"111010001",
  47486=>"000100001",
  47487=>"111000010",
  47488=>"100110000",
  47489=>"100111110",
  47490=>"111110011",
  47491=>"011010010",
  47492=>"010001011",
  47493=>"110000111",
  47494=>"100010110",
  47495=>"011000011",
  47496=>"111010110",
  47497=>"100001100",
  47498=>"101001010",
  47499=>"111011001",
  47500=>"000101010",
  47501=>"100000101",
  47502=>"101111000",
  47503=>"000100001",
  47504=>"010011110",
  47505=>"000101100",
  47506=>"111101010",
  47507=>"111011100",
  47508=>"001110101",
  47509=>"000011110",
  47510=>"001011101",
  47511=>"101110001",
  47512=>"101111111",
  47513=>"110100100",
  47514=>"000100110",
  47515=>"000001011",
  47516=>"111010110",
  47517=>"101001000",
  47518=>"011000110",
  47519=>"110111001",
  47520=>"111010110",
  47521=>"001000011",
  47522=>"110100100",
  47523=>"111000001",
  47524=>"001111000",
  47525=>"111001101",
  47526=>"110011001",
  47527=>"000000101",
  47528=>"110001101",
  47529=>"011011011",
  47530=>"111111111",
  47531=>"111100101",
  47532=>"000010010",
  47533=>"001101010",
  47534=>"001100110",
  47535=>"011100011",
  47536=>"111101000",
  47537=>"011000100",
  47538=>"010000010",
  47539=>"001011111",
  47540=>"101100010",
  47541=>"001111001",
  47542=>"000011011",
  47543=>"110001010",
  47544=>"111110010",
  47545=>"100111010",
  47546=>"100010101",
  47547=>"001010110",
  47548=>"001000111",
  47549=>"001111001",
  47550=>"011100001",
  47551=>"001111101",
  47552=>"111011001",
  47553=>"111111110",
  47554=>"100101110",
  47555=>"000010000",
  47556=>"100000011",
  47557=>"000000111",
  47558=>"100011100",
  47559=>"100000110",
  47560=>"000111001",
  47561=>"001110011",
  47562=>"111001110",
  47563=>"101001101",
  47564=>"111001000",
  47565=>"000001111",
  47566=>"100100011",
  47567=>"011110001",
  47568=>"000101101",
  47569=>"001000000",
  47570=>"110000000",
  47571=>"010011001",
  47572=>"110101001",
  47573=>"110001111",
  47574=>"101110010",
  47575=>"000010110",
  47576=>"101011111",
  47577=>"001001010",
  47578=>"110100010",
  47579=>"111001011",
  47580=>"000011001",
  47581=>"101011000",
  47582=>"110101010",
  47583=>"000100000",
  47584=>"010110110",
  47585=>"101110101",
  47586=>"100111111",
  47587=>"010110011",
  47588=>"010101000",
  47589=>"100011110",
  47590=>"011001110",
  47591=>"110001100",
  47592=>"000000110",
  47593=>"111111101",
  47594=>"011110111",
  47595=>"101110001",
  47596=>"000010101",
  47597=>"000111000",
  47598=>"100101011",
  47599=>"000110001",
  47600=>"010010001",
  47601=>"010100110",
  47602=>"110000001",
  47603=>"101110100",
  47604=>"011010001",
  47605=>"001100111",
  47606=>"001011000",
  47607=>"100101000",
  47608=>"101000010",
  47609=>"011100100",
  47610=>"001101001",
  47611=>"010001011",
  47612=>"011111111",
  47613=>"110100101",
  47614=>"001000011",
  47615=>"100110110",
  47616=>"000001000",
  47617=>"111001000",
  47618=>"110011100",
  47619=>"100001011",
  47620=>"010110011",
  47621=>"000111100",
  47622=>"111111010",
  47623=>"101111100",
  47624=>"101000111",
  47625=>"011101011",
  47626=>"000011010",
  47627=>"000111100",
  47628=>"110110000",
  47629=>"001110110",
  47630=>"010110000",
  47631=>"001100010",
  47632=>"000101010",
  47633=>"010000001",
  47634=>"110001010",
  47635=>"111110011",
  47636=>"011001100",
  47637=>"110100010",
  47638=>"110101011",
  47639=>"010000000",
  47640=>"101100011",
  47641=>"100110010",
  47642=>"000010010",
  47643=>"001111011",
  47644=>"111001101",
  47645=>"110010011",
  47646=>"001111000",
  47647=>"110111001",
  47648=>"010111110",
  47649=>"000000100",
  47650=>"100000000",
  47651=>"011101101",
  47652=>"111001000",
  47653=>"100100100",
  47654=>"111001101",
  47655=>"101011110",
  47656=>"001101001",
  47657=>"000110010",
  47658=>"111101111",
  47659=>"000010100",
  47660=>"100111100",
  47661=>"011010011",
  47662=>"101010001",
  47663=>"000011101",
  47664=>"000100110",
  47665=>"011111000",
  47666=>"001001100",
  47667=>"101011100",
  47668=>"011011000",
  47669=>"000110000",
  47670=>"111000111",
  47671=>"110101111",
  47672=>"111110010",
  47673=>"110001110",
  47674=>"100100100",
  47675=>"101111010",
  47676=>"110111110",
  47677=>"111111000",
  47678=>"010000001",
  47679=>"100011000",
  47680=>"011000101",
  47681=>"101101010",
  47682=>"010000111",
  47683=>"101100010",
  47684=>"110101101",
  47685=>"011110101",
  47686=>"000111100",
  47687=>"111110101",
  47688=>"010001111",
  47689=>"001010111",
  47690=>"100111100",
  47691=>"000110110",
  47692=>"011110101",
  47693=>"111001111",
  47694=>"000101010",
  47695=>"100111111",
  47696=>"001011100",
  47697=>"111001101",
  47698=>"010001000",
  47699=>"011101101",
  47700=>"010101110",
  47701=>"001010011",
  47702=>"101001011",
  47703=>"001111101",
  47704=>"111011110",
  47705=>"000101000",
  47706=>"111111011",
  47707=>"011000111",
  47708=>"111111011",
  47709=>"110111000",
  47710=>"010111100",
  47711=>"010100100",
  47712=>"001001011",
  47713=>"101001101",
  47714=>"001111001",
  47715=>"101111111",
  47716=>"010111100",
  47717=>"010100100",
  47718=>"011101100",
  47719=>"011101010",
  47720=>"101011000",
  47721=>"100100101",
  47722=>"011101111",
  47723=>"011010101",
  47724=>"100100011",
  47725=>"111111111",
  47726=>"101011110",
  47727=>"100101111",
  47728=>"001100110",
  47729=>"000110110",
  47730=>"111011101",
  47731=>"001010010",
  47732=>"010011110",
  47733=>"010010101",
  47734=>"110101000",
  47735=>"100111000",
  47736=>"111101011",
  47737=>"011010111",
  47738=>"011110001",
  47739=>"100001100",
  47740=>"100011000",
  47741=>"111001000",
  47742=>"000000000",
  47743=>"000110100",
  47744=>"111010000",
  47745=>"100011101",
  47746=>"110100110",
  47747=>"000001101",
  47748=>"101000000",
  47749=>"010111100",
  47750=>"001010101",
  47751=>"111000110",
  47752=>"100100101",
  47753=>"110011111",
  47754=>"110111101",
  47755=>"010001100",
  47756=>"011100000",
  47757=>"000100101",
  47758=>"000101011",
  47759=>"011010011",
  47760=>"010101000",
  47761=>"010011110",
  47762=>"101000110",
  47763=>"001111000",
  47764=>"110000110",
  47765=>"111100001",
  47766=>"101101110",
  47767=>"111110001",
  47768=>"010101111",
  47769=>"100010101",
  47770=>"100010110",
  47771=>"000010101",
  47772=>"010001110",
  47773=>"100100000",
  47774=>"000110010",
  47775=>"100010100",
  47776=>"111110101",
  47777=>"010111111",
  47778=>"000011101",
  47779=>"110101101",
  47780=>"000101110",
  47781=>"111111111",
  47782=>"010000001",
  47783=>"011100011",
  47784=>"111001100",
  47785=>"000011011",
  47786=>"110011111",
  47787=>"101110000",
  47788=>"110001001",
  47789=>"110110110",
  47790=>"110000111",
  47791=>"000011111",
  47792=>"001100011",
  47793=>"010000010",
  47794=>"010010000",
  47795=>"010100110",
  47796=>"110101000",
  47797=>"011111110",
  47798=>"111010010",
  47799=>"000101111",
  47800=>"110101110",
  47801=>"000101000",
  47802=>"011110100",
  47803=>"110111110",
  47804=>"101110001",
  47805=>"010100110",
  47806=>"010100110",
  47807=>"111100101",
  47808=>"000001110",
  47809=>"101011111",
  47810=>"101100000",
  47811=>"101110101",
  47812=>"010111010",
  47813=>"110100001",
  47814=>"011000111",
  47815=>"111011101",
  47816=>"110001011",
  47817=>"100001000",
  47818=>"101110001",
  47819=>"001100011",
  47820=>"101111101",
  47821=>"111101101",
  47822=>"011100111",
  47823=>"000100010",
  47824=>"110100001",
  47825=>"101011011",
  47826=>"001111001",
  47827=>"011101110",
  47828=>"001110111",
  47829=>"010001110",
  47830=>"001110000",
  47831=>"000110101",
  47832=>"000110000",
  47833=>"000110001",
  47834=>"010010011",
  47835=>"000010111",
  47836=>"110111100",
  47837=>"001110000",
  47838=>"111011001",
  47839=>"110010100",
  47840=>"101111111",
  47841=>"000100000",
  47842=>"011000110",
  47843=>"011100001",
  47844=>"110011010",
  47845=>"000010110",
  47846=>"010111011",
  47847=>"010001111",
  47848=>"000101000",
  47849=>"000111101",
  47850=>"000011110",
  47851=>"101011101",
  47852=>"000010110",
  47853=>"000011100",
  47854=>"110101101",
  47855=>"000001010",
  47856=>"101010001",
  47857=>"110011111",
  47858=>"100100100",
  47859=>"110010010",
  47860=>"010010001",
  47861=>"110110111",
  47862=>"100001011",
  47863=>"110110101",
  47864=>"000101011",
  47865=>"100000110",
  47866=>"011100000",
  47867=>"000000000",
  47868=>"000101001",
  47869=>"000110001",
  47870=>"100111010",
  47871=>"100001111",
  47872=>"000010101",
  47873=>"010001100",
  47874=>"000010100",
  47875=>"010100010",
  47876=>"000101111",
  47877=>"001000111",
  47878=>"110011011",
  47879=>"110111010",
  47880=>"110101110",
  47881=>"010011011",
  47882=>"001000100",
  47883=>"110001101",
  47884=>"001000010",
  47885=>"110100001",
  47886=>"100011100",
  47887=>"010001111",
  47888=>"110110100",
  47889=>"011010001",
  47890=>"110111001",
  47891=>"111100110",
  47892=>"010110010",
  47893=>"100101101",
  47894=>"001001111",
  47895=>"011010110",
  47896=>"001011101",
  47897=>"111010110",
  47898=>"101111111",
  47899=>"000110001",
  47900=>"100110010",
  47901=>"110111101",
  47902=>"010111010",
  47903=>"011001011",
  47904=>"111001101",
  47905=>"010011010",
  47906=>"010111011",
  47907=>"001010100",
  47908=>"010010001",
  47909=>"110001010",
  47910=>"000101110",
  47911=>"010001101",
  47912=>"101101111",
  47913=>"000110111",
  47914=>"001101101",
  47915=>"100001011",
  47916=>"111010101",
  47917=>"100011111",
  47918=>"010010100",
  47919=>"011000110",
  47920=>"011110101",
  47921=>"000110100",
  47922=>"010101000",
  47923=>"101000110",
  47924=>"010110000",
  47925=>"000100010",
  47926=>"111001101",
  47927=>"001100010",
  47928=>"101101001",
  47929=>"001110000",
  47930=>"101110011",
  47931=>"010000100",
  47932=>"010000100",
  47933=>"010101011",
  47934=>"110011110",
  47935=>"011010000",
  47936=>"100101011",
  47937=>"101010011",
  47938=>"101110011",
  47939=>"000010110",
  47940=>"001001000",
  47941=>"010000101",
  47942=>"101111101",
  47943=>"110101110",
  47944=>"110010001",
  47945=>"011000001",
  47946=>"111111010",
  47947=>"111101000",
  47948=>"010000111",
  47949=>"011101101",
  47950=>"100011010",
  47951=>"101000100",
  47952=>"100101000",
  47953=>"000100000",
  47954=>"000000001",
  47955=>"110011000",
  47956=>"111011010",
  47957=>"111101110",
  47958=>"110101110",
  47959=>"010000001",
  47960=>"110011001",
  47961=>"010001100",
  47962=>"101010101",
  47963=>"101101001",
  47964=>"111001001",
  47965=>"000111010",
  47966=>"011101110",
  47967=>"000110000",
  47968=>"101010001",
  47969=>"101110001",
  47970=>"100001110",
  47971=>"111000100",
  47972=>"100111110",
  47973=>"001111101",
  47974=>"001100001",
  47975=>"011111011",
  47976=>"000100000",
  47977=>"011100010",
  47978=>"101110100",
  47979=>"111011001",
  47980=>"100111111",
  47981=>"001011010",
  47982=>"001010111",
  47983=>"001010110",
  47984=>"100110000",
  47985=>"011110001",
  47986=>"000001111",
  47987=>"011101110",
  47988=>"101100110",
  47989=>"111101011",
  47990=>"100001001",
  47991=>"110000000",
  47992=>"100010101",
  47993=>"101000011",
  47994=>"101101010",
  47995=>"111001110",
  47996=>"011100111",
  47997=>"011001001",
  47998=>"111010111",
  47999=>"001000000",
  48000=>"111000110",
  48001=>"111100010",
  48002=>"100111000",
  48003=>"000010001",
  48004=>"100100011",
  48005=>"100111011",
  48006=>"101010110",
  48007=>"100111111",
  48008=>"000100010",
  48009=>"100010001",
  48010=>"011001101",
  48011=>"100001101",
  48012=>"001101001",
  48013=>"001000010",
  48014=>"000110111",
  48015=>"000000100",
  48016=>"110011000",
  48017=>"101101001",
  48018=>"010100000",
  48019=>"101010100",
  48020=>"011011100",
  48021=>"000010000",
  48022=>"110110101",
  48023=>"110011110",
  48024=>"010001101",
  48025=>"001000000",
  48026=>"011110100",
  48027=>"010111111",
  48028=>"100001000",
  48029=>"100010101",
  48030=>"111001010",
  48031=>"101101010",
  48032=>"010011000",
  48033=>"110011011",
  48034=>"100111110",
  48035=>"111111101",
  48036=>"011011101",
  48037=>"100111011",
  48038=>"001001001",
  48039=>"000111101",
  48040=>"101010001",
  48041=>"101010001",
  48042=>"101110111",
  48043=>"111001111",
  48044=>"000101111",
  48045=>"011100101",
  48046=>"111001000",
  48047=>"000011011",
  48048=>"000111000",
  48049=>"100100111",
  48050=>"100000001",
  48051=>"110001110",
  48052=>"111100010",
  48053=>"110110010",
  48054=>"001100000",
  48055=>"101010100",
  48056=>"000000111",
  48057=>"011011111",
  48058=>"010111010",
  48059=>"011110001",
  48060=>"000100110",
  48061=>"000001101",
  48062=>"111111001",
  48063=>"001111000",
  48064=>"110101010",
  48065=>"010100010",
  48066=>"000001001",
  48067=>"111001001",
  48068=>"000101001",
  48069=>"011010101",
  48070=>"100001001",
  48071=>"111100000",
  48072=>"000010001",
  48073=>"010010001",
  48074=>"010100100",
  48075=>"011111000",
  48076=>"000010000",
  48077=>"110011110",
  48078=>"100000100",
  48079=>"000111110",
  48080=>"110100000",
  48081=>"001000101",
  48082=>"100100011",
  48083=>"111000101",
  48084=>"010011001",
  48085=>"111111010",
  48086=>"110011111",
  48087=>"110000000",
  48088=>"110100110",
  48089=>"011000100",
  48090=>"000010000",
  48091=>"000000100",
  48092=>"100110101",
  48093=>"011000000",
  48094=>"110111000",
  48095=>"010011110",
  48096=>"111111011",
  48097=>"100101011",
  48098=>"100000111",
  48099=>"011111100",
  48100=>"010111001",
  48101=>"000101110",
  48102=>"101111010",
  48103=>"000000001",
  48104=>"101000111",
  48105=>"110110110",
  48106=>"011001100",
  48107=>"000000110",
  48108=>"110110100",
  48109=>"011001011",
  48110=>"010011101",
  48111=>"111000101",
  48112=>"010010001",
  48113=>"000010011",
  48114=>"100100111",
  48115=>"101101001",
  48116=>"001010110",
  48117=>"111110111",
  48118=>"100100110",
  48119=>"111100111",
  48120=>"001000010",
  48121=>"011011000",
  48122=>"100100100",
  48123=>"011100001",
  48124=>"000110011",
  48125=>"000010111",
  48126=>"100100100",
  48127=>"100010100",
  48128=>"011100100",
  48129=>"111101100",
  48130=>"110010010",
  48131=>"010010011",
  48132=>"110111110",
  48133=>"010111110",
  48134=>"010001110",
  48135=>"001001001",
  48136=>"110100001",
  48137=>"011111101",
  48138=>"011110110",
  48139=>"101111010",
  48140=>"101101010",
  48141=>"000011011",
  48142=>"011111101",
  48143=>"001001010",
  48144=>"011100110",
  48145=>"111001000",
  48146=>"110101011",
  48147=>"101100101",
  48148=>"100100111",
  48149=>"101111001",
  48150=>"111100001",
  48151=>"010000011",
  48152=>"111101010",
  48153=>"010111110",
  48154=>"100000101",
  48155=>"010100000",
  48156=>"110010010",
  48157=>"111110000",
  48158=>"010010000",
  48159=>"111100000",
  48160=>"000000011",
  48161=>"010101101",
  48162=>"010111110",
  48163=>"011100001",
  48164=>"010100110",
  48165=>"110110111",
  48166=>"100000100",
  48167=>"001100011",
  48168=>"011011100",
  48169=>"100010110",
  48170=>"100001101",
  48171=>"111011000",
  48172=>"111011000",
  48173=>"100001100",
  48174=>"111000111",
  48175=>"000110001",
  48176=>"100010010",
  48177=>"110101110",
  48178=>"100110101",
  48179=>"110000000",
  48180=>"110101100",
  48181=>"111010001",
  48182=>"011000000",
  48183=>"111000001",
  48184=>"000010101",
  48185=>"101001010",
  48186=>"110010111",
  48187=>"101001101",
  48188=>"011000110",
  48189=>"111101001",
  48190=>"000110011",
  48191=>"011010111",
  48192=>"110101010",
  48193=>"010010111",
  48194=>"111110110",
  48195=>"010111100",
  48196=>"100100111",
  48197=>"011000100",
  48198=>"111111100",
  48199=>"100101010",
  48200=>"010000101",
  48201=>"101111100",
  48202=>"101000100",
  48203=>"000100101",
  48204=>"010110100",
  48205=>"001101001",
  48206=>"111001110",
  48207=>"000100101",
  48208=>"010101011",
  48209=>"101111010",
  48210=>"000000100",
  48211=>"101001011",
  48212=>"010110100",
  48213=>"101010010",
  48214=>"001100000",
  48215=>"100110100",
  48216=>"011010001",
  48217=>"101010010",
  48218=>"001100110",
  48219=>"111001000",
  48220=>"110001010",
  48221=>"010101110",
  48222=>"110101111",
  48223=>"110101011",
  48224=>"110010110",
  48225=>"001100101",
  48226=>"110000111",
  48227=>"111010000",
  48228=>"011000010",
  48229=>"011000110",
  48230=>"011111000",
  48231=>"100110011",
  48232=>"011000001",
  48233=>"010011010",
  48234=>"101011000",
  48235=>"110011101",
  48236=>"011111100",
  48237=>"110000001",
  48238=>"010111011",
  48239=>"010111111",
  48240=>"000101111",
  48241=>"111111000",
  48242=>"111111111",
  48243=>"110101110",
  48244=>"001001001",
  48245=>"110111101",
  48246=>"111011101",
  48247=>"000001010",
  48248=>"010011000",
  48249=>"100110110",
  48250=>"000100001",
  48251=>"011000101",
  48252=>"100000101",
  48253=>"011001010",
  48254=>"101101011",
  48255=>"000111101",
  48256=>"110111001",
  48257=>"111101111",
  48258=>"011111011",
  48259=>"101101100",
  48260=>"111101010",
  48261=>"111111000",
  48262=>"010101101",
  48263=>"010110000",
  48264=>"011001001",
  48265=>"111010010",
  48266=>"000000101",
  48267=>"001100011",
  48268=>"011110110",
  48269=>"111001110",
  48270=>"000011000",
  48271=>"011111000",
  48272=>"101111000",
  48273=>"000001000",
  48274=>"101000000",
  48275=>"110100110",
  48276=>"101101000",
  48277=>"000101100",
  48278=>"001001001",
  48279=>"101011100",
  48280=>"010010000",
  48281=>"001100110",
  48282=>"000101100",
  48283=>"011000101",
  48284=>"000111000",
  48285=>"000101101",
  48286=>"000010000",
  48287=>"001000111",
  48288=>"110100010",
  48289=>"010011001",
  48290=>"010100100",
  48291=>"100010001",
  48292=>"000110000",
  48293=>"010001001",
  48294=>"010110001",
  48295=>"110001001",
  48296=>"001110110",
  48297=>"100110101",
  48298=>"111100101",
  48299=>"110001010",
  48300=>"110010101",
  48301=>"111111001",
  48302=>"100100110",
  48303=>"011001100",
  48304=>"110010001",
  48305=>"000100010",
  48306=>"001000011",
  48307=>"101001110",
  48308=>"100101011",
  48309=>"010000000",
  48310=>"001100110",
  48311=>"101011010",
  48312=>"000100010",
  48313=>"000101000",
  48314=>"101110100",
  48315=>"111111110",
  48316=>"011100001",
  48317=>"011000011",
  48318=>"001011010",
  48319=>"100110111",
  48320=>"011010000",
  48321=>"010000001",
  48322=>"111000000",
  48323=>"101001000",
  48324=>"111011001",
  48325=>"101110101",
  48326=>"110100111",
  48327=>"000110011",
  48328=>"011110100",
  48329=>"010101000",
  48330=>"011000111",
  48331=>"100110101",
  48332=>"110111010",
  48333=>"111101111",
  48334=>"101000111",
  48335=>"001100000",
  48336=>"101011110",
  48337=>"011000110",
  48338=>"011111101",
  48339=>"011000010",
  48340=>"100011110",
  48341=>"111110100",
  48342=>"001000011",
  48343=>"010010110",
  48344=>"000000001",
  48345=>"100110111",
  48346=>"000000000",
  48347=>"100001110",
  48348=>"111110011",
  48349=>"111111000",
  48350=>"110111111",
  48351=>"110100110",
  48352=>"001010010",
  48353=>"000001111",
  48354=>"011000100",
  48355=>"011010101",
  48356=>"110111110",
  48357=>"111110001",
  48358=>"011011001",
  48359=>"011010110",
  48360=>"100000000",
  48361=>"111001001",
  48362=>"011101110",
  48363=>"011000100",
  48364=>"010101010",
  48365=>"100110010",
  48366=>"101011111",
  48367=>"010111111",
  48368=>"100101010",
  48369=>"011110011",
  48370=>"111000110",
  48371=>"000100000",
  48372=>"000010001",
  48373=>"001001111",
  48374=>"001101000",
  48375=>"110010101",
  48376=>"100111111",
  48377=>"000011000",
  48378=>"011001110",
  48379=>"001101000",
  48380=>"101110110",
  48381=>"110111000",
  48382=>"001101100",
  48383=>"000001010",
  48384=>"110100000",
  48385=>"010100111",
  48386=>"111110001",
  48387=>"110010000",
  48388=>"100010000",
  48389=>"010001110",
  48390=>"010110001",
  48391=>"001000101",
  48392=>"001101001",
  48393=>"001100000",
  48394=>"101101011",
  48395=>"000000000",
  48396=>"000010101",
  48397=>"001010001",
  48398=>"100111101",
  48399=>"001000100",
  48400=>"001001101",
  48401=>"011000110",
  48402=>"000011011",
  48403=>"111111111",
  48404=>"110111101",
  48405=>"111100000",
  48406=>"010001011",
  48407=>"100110111",
  48408=>"100111001",
  48409=>"100001001",
  48410=>"001100001",
  48411=>"000010000",
  48412=>"001101001",
  48413=>"100111110",
  48414=>"111111100",
  48415=>"101000100",
  48416=>"000101111",
  48417=>"101111000",
  48418=>"111111111",
  48419=>"111011000",
  48420=>"100011010",
  48421=>"100000101",
  48422=>"111001001",
  48423=>"100111001",
  48424=>"101001101",
  48425=>"101010101",
  48426=>"001001010",
  48427=>"001111001",
  48428=>"010000010",
  48429=>"000000001",
  48430=>"011101000",
  48431=>"101110111",
  48432=>"111100001",
  48433=>"100010100",
  48434=>"000101010",
  48435=>"101001001",
  48436=>"001010001",
  48437=>"010100100",
  48438=>"111110100",
  48439=>"011011101",
  48440=>"001001100",
  48441=>"000110110",
  48442=>"100011011",
  48443=>"011110111",
  48444=>"010111001",
  48445=>"010001111",
  48446=>"111111110",
  48447=>"101110000",
  48448=>"100011100",
  48449=>"001001110",
  48450=>"000001000",
  48451=>"101100011",
  48452=>"001011011",
  48453=>"010101111",
  48454=>"000011110",
  48455=>"111111001",
  48456=>"111010101",
  48457=>"010110001",
  48458=>"111111010",
  48459=>"001110001",
  48460=>"110111111",
  48461=>"111111111",
  48462=>"001101001",
  48463=>"111001111",
  48464=>"010011011",
  48465=>"100100011",
  48466=>"011100111",
  48467=>"111100101",
  48468=>"100101110",
  48469=>"100010010",
  48470=>"100011010",
  48471=>"010000111",
  48472=>"110101110",
  48473=>"101000110",
  48474=>"001010011",
  48475=>"111101101",
  48476=>"101101101",
  48477=>"011100001",
  48478=>"001011100",
  48479=>"100010011",
  48480=>"110101110",
  48481=>"101111011",
  48482=>"000000010",
  48483=>"111010010",
  48484=>"001000111",
  48485=>"010100101",
  48486=>"111011101",
  48487=>"111111101",
  48488=>"100010010",
  48489=>"111100111",
  48490=>"001111010",
  48491=>"111011101",
  48492=>"010101010",
  48493=>"101101100",
  48494=>"011100000",
  48495=>"000001000",
  48496=>"010000000",
  48497=>"101000100",
  48498=>"000011010",
  48499=>"001100101",
  48500=>"100100011",
  48501=>"011110011",
  48502=>"000111000",
  48503=>"100110101",
  48504=>"001010100",
  48505=>"111110001",
  48506=>"010101110",
  48507=>"010001100",
  48508=>"001010010",
  48509=>"101001111",
  48510=>"011011110",
  48511=>"000111100",
  48512=>"010001011",
  48513=>"001100111",
  48514=>"111000000",
  48515=>"010101111",
  48516=>"001101100",
  48517=>"100111011",
  48518=>"100101110",
  48519=>"001001101",
  48520=>"010000100",
  48521=>"111110101",
  48522=>"000110101",
  48523=>"011001101",
  48524=>"111100101",
  48525=>"110000010",
  48526=>"011111110",
  48527=>"100010101",
  48528=>"101011111",
  48529=>"111000011",
  48530=>"111100110",
  48531=>"010000100",
  48532=>"101111011",
  48533=>"011010001",
  48534=>"000110110",
  48535=>"001111100",
  48536=>"100000011",
  48537=>"100000010",
  48538=>"011000001",
  48539=>"110000010",
  48540=>"111000111",
  48541=>"010010101",
  48542=>"101101100",
  48543=>"010011100",
  48544=>"011111001",
  48545=>"011110000",
  48546=>"001001001",
  48547=>"000000101",
  48548=>"110001001",
  48549=>"010110110",
  48550=>"110010111",
  48551=>"010100010",
  48552=>"000100100",
  48553=>"000000101",
  48554=>"001100011",
  48555=>"011101010",
  48556=>"011010100",
  48557=>"111101010",
  48558=>"111001001",
  48559=>"001101011",
  48560=>"101100010",
  48561=>"010100010",
  48562=>"001011101",
  48563=>"010001001",
  48564=>"110001010",
  48565=>"100011110",
  48566=>"111011110",
  48567=>"011100110",
  48568=>"111110011",
  48569=>"111000100",
  48570=>"000110111",
  48571=>"100100101",
  48572=>"000000101",
  48573=>"001010110",
  48574=>"111000000",
  48575=>"101000000",
  48576=>"110111011",
  48577=>"101100111",
  48578=>"111001010",
  48579=>"001000111",
  48580=>"001011111",
  48581=>"100100011",
  48582=>"111010000",
  48583=>"000010001",
  48584=>"111001111",
  48585=>"010010110",
  48586=>"110000000",
  48587=>"001010100",
  48588=>"000011110",
  48589=>"110101011",
  48590=>"100010111",
  48591=>"000110111",
  48592=>"000101100",
  48593=>"110110111",
  48594=>"111111101",
  48595=>"011100010",
  48596=>"111011101",
  48597=>"111111010",
  48598=>"000110111",
  48599=>"111111111",
  48600=>"110011011",
  48601=>"110000101",
  48602=>"011100001",
  48603=>"100100101",
  48604=>"110010111",
  48605=>"010010110",
  48606=>"100000001",
  48607=>"000010101",
  48608=>"101000111",
  48609=>"000110011",
  48610=>"011101011",
  48611=>"100101010",
  48612=>"111111000",
  48613=>"000000001",
  48614=>"100101001",
  48615=>"110101000",
  48616=>"101011010",
  48617=>"010011110",
  48618=>"011000101",
  48619=>"001110111",
  48620=>"001011101",
  48621=>"010101001",
  48622=>"111001101",
  48623=>"110110010",
  48624=>"110100110",
  48625=>"011000010",
  48626=>"101100111",
  48627=>"101010000",
  48628=>"110100111",
  48629=>"100010101",
  48630=>"110010010",
  48631=>"111001101",
  48632=>"010000000",
  48633=>"001101011",
  48634=>"101010110",
  48635=>"001000111",
  48636=>"000111110",
  48637=>"100011000",
  48638=>"001100011",
  48639=>"111111011",
  48640=>"110010000",
  48641=>"100110001",
  48642=>"100100101",
  48643=>"101001011",
  48644=>"010000111",
  48645=>"101111110",
  48646=>"011010111",
  48647=>"010000000",
  48648=>"110011000",
  48649=>"100001110",
  48650=>"000011101",
  48651=>"010000111",
  48652=>"101110101",
  48653=>"110010000",
  48654=>"011111000",
  48655=>"000110110",
  48656=>"110110000",
  48657=>"101000000",
  48658=>"110111011",
  48659=>"110110100",
  48660=>"000110001",
  48661=>"100111011",
  48662=>"000110001",
  48663=>"101111111",
  48664=>"100000110",
  48665=>"100110011",
  48666=>"101010000",
  48667=>"010011000",
  48668=>"111111111",
  48669=>"011110111",
  48670=>"110010110",
  48671=>"101111011",
  48672=>"000011110",
  48673=>"101101000",
  48674=>"010001100",
  48675=>"101110010",
  48676=>"111000100",
  48677=>"001110011",
  48678=>"010100100",
  48679=>"001000001",
  48680=>"000011110",
  48681=>"010001010",
  48682=>"111011100",
  48683=>"011010001",
  48684=>"100001001",
  48685=>"011111111",
  48686=>"011111001",
  48687=>"000000001",
  48688=>"110101010",
  48689=>"011110100",
  48690=>"000111111",
  48691=>"011110110",
  48692=>"101001011",
  48693=>"101000001",
  48694=>"011010010",
  48695=>"111101101",
  48696=>"011101110",
  48697=>"000100000",
  48698=>"111001100",
  48699=>"010001100",
  48700=>"101001101",
  48701=>"000011110",
  48702=>"000110101",
  48703=>"101111110",
  48704=>"000000001",
  48705=>"000111111",
  48706=>"011101111",
  48707=>"101010011",
  48708=>"001110000",
  48709=>"100111010",
  48710=>"011101100",
  48711=>"010101100",
  48712=>"001001010",
  48713=>"001000101",
  48714=>"000101011",
  48715=>"001100010",
  48716=>"000100111",
  48717=>"110000000",
  48718=>"010101110",
  48719=>"101010001",
  48720=>"100000010",
  48721=>"100111010",
  48722=>"100110110",
  48723=>"100111001",
  48724=>"111101000",
  48725=>"011000111",
  48726=>"100101101",
  48727=>"100001111",
  48728=>"100101011",
  48729=>"111010111",
  48730=>"110101111",
  48731=>"111001011",
  48732=>"110110010",
  48733=>"111101100",
  48734=>"000110100",
  48735=>"101010110",
  48736=>"011010011",
  48737=>"000011011",
  48738=>"101110101",
  48739=>"101110110",
  48740=>"011000110",
  48741=>"101111011",
  48742=>"100001100",
  48743=>"011001000",
  48744=>"101101100",
  48745=>"101100100",
  48746=>"010100111",
  48747=>"000010111",
  48748=>"100000011",
  48749=>"011011101",
  48750=>"001111111",
  48751=>"010111010",
  48752=>"010000000",
  48753=>"001000101",
  48754=>"011001000",
  48755=>"001001111",
  48756=>"110001001",
  48757=>"011001001",
  48758=>"110110100",
  48759=>"110110110",
  48760=>"000001010",
  48761=>"101100110",
  48762=>"100000101",
  48763=>"101110111",
  48764=>"111011011",
  48765=>"111101010",
  48766=>"111101010",
  48767=>"010110011",
  48768=>"000100111",
  48769=>"001110110",
  48770=>"010011111",
  48771=>"000001111",
  48772=>"011001110",
  48773=>"000000000",
  48774=>"011100001",
  48775=>"111111011",
  48776=>"111111111",
  48777=>"011011011",
  48778=>"000001110",
  48779=>"111010101",
  48780=>"000111111",
  48781=>"101011110",
  48782=>"011000000",
  48783=>"001111110",
  48784=>"100110010",
  48785=>"011011101",
  48786=>"000011110",
  48787=>"101111110",
  48788=>"010011000",
  48789=>"010001010",
  48790=>"101000111",
  48791=>"110010000",
  48792=>"100110010",
  48793=>"011101001",
  48794=>"101010010",
  48795=>"111011111",
  48796=>"010101010",
  48797=>"001010111",
  48798=>"001100000",
  48799=>"011101101",
  48800=>"000100100",
  48801=>"110100001",
  48802=>"100011110",
  48803=>"010010111",
  48804=>"011010010",
  48805=>"000100100",
  48806=>"101110110",
  48807=>"000001000",
  48808=>"100001011",
  48809=>"011001010",
  48810=>"111111010",
  48811=>"101101101",
  48812=>"111001101",
  48813=>"101010111",
  48814=>"111110001",
  48815=>"000010011",
  48816=>"111001111",
  48817=>"100101000",
  48818=>"101010001",
  48819=>"001010101",
  48820=>"010011111",
  48821=>"011110010",
  48822=>"001010010",
  48823=>"100010100",
  48824=>"001010000",
  48825=>"100010100",
  48826=>"010001111",
  48827=>"100111011",
  48828=>"110100111",
  48829=>"010011011",
  48830=>"000101010",
  48831=>"001101110",
  48832=>"010100011",
  48833=>"101101111",
  48834=>"011011011",
  48835=>"001111011",
  48836=>"011111001",
  48837=>"000100011",
  48838=>"000000001",
  48839=>"101101100",
  48840=>"001111000",
  48841=>"010001101",
  48842=>"001010111",
  48843=>"111110111",
  48844=>"001101011",
  48845=>"110000000",
  48846=>"001110000",
  48847=>"001000001",
  48848=>"110100110",
  48849=>"111011011",
  48850=>"100111110",
  48851=>"111010110",
  48852=>"111000110",
  48853=>"111101011",
  48854=>"001010101",
  48855=>"011010101",
  48856=>"001101111",
  48857=>"110101110",
  48858=>"111110000",
  48859=>"100100010",
  48860=>"010011011",
  48861=>"011110000",
  48862=>"100110110",
  48863=>"011110111",
  48864=>"010000000",
  48865=>"011101001",
  48866=>"000000111",
  48867=>"100111000",
  48868=>"101111111",
  48869=>"011001000",
  48870=>"111010110",
  48871=>"110000110",
  48872=>"001010010",
  48873=>"001001010",
  48874=>"011101111",
  48875=>"001100101",
  48876=>"001010110",
  48877=>"001000001",
  48878=>"100111000",
  48879=>"100111000",
  48880=>"010110101",
  48881=>"001000111",
  48882=>"000011001",
  48883=>"010001010",
  48884=>"011100101",
  48885=>"110001010",
  48886=>"001000000",
  48887=>"100010010",
  48888=>"000100010",
  48889=>"110110010",
  48890=>"110011010",
  48891=>"000101101",
  48892=>"000110101",
  48893=>"111001110",
  48894=>"010100010",
  48895=>"111011111",
  48896=>"101100001",
  48897=>"000110010",
  48898=>"010001011",
  48899=>"110100011",
  48900=>"001010010",
  48901=>"110110110",
  48902=>"110011101",
  48903=>"001011001",
  48904=>"011010010",
  48905=>"010100010",
  48906=>"000001110",
  48907=>"110010101",
  48908=>"111101100",
  48909=>"101011111",
  48910=>"010101011",
  48911=>"010000100",
  48912=>"110101001",
  48913=>"001110111",
  48914=>"101100010",
  48915=>"010000100",
  48916=>"110010111",
  48917=>"001001100",
  48918=>"000100011",
  48919=>"011101111",
  48920=>"010111100",
  48921=>"001100011",
  48922=>"010101101",
  48923=>"011000001",
  48924=>"010000110",
  48925=>"010100010",
  48926=>"100110000",
  48927=>"111000010",
  48928=>"000100100",
  48929=>"101000000",
  48930=>"110100110",
  48931=>"001100110",
  48932=>"101000110",
  48933=>"010011110",
  48934=>"011011110",
  48935=>"100000001",
  48936=>"001011111",
  48937=>"100111010",
  48938=>"011010010",
  48939=>"011101000",
  48940=>"101111111",
  48941=>"000000000",
  48942=>"010110111",
  48943=>"111100101",
  48944=>"000110001",
  48945=>"010111011",
  48946=>"000010000",
  48947=>"011101111",
  48948=>"101011011",
  48949=>"010100100",
  48950=>"000000000",
  48951=>"110111000",
  48952=>"000111111",
  48953=>"010111100",
  48954=>"011011010",
  48955=>"100011001",
  48956=>"010101110",
  48957=>"000101010",
  48958=>"011010010",
  48959=>"001010000",
  48960=>"111000111",
  48961=>"000000011",
  48962=>"011110011",
  48963=>"101011010",
  48964=>"000010111",
  48965=>"101101101",
  48966=>"101100001",
  48967=>"111111111",
  48968=>"001011110",
  48969=>"100101111",
  48970=>"110100111",
  48971=>"110000001",
  48972=>"011001100",
  48973=>"010001111",
  48974=>"101011001",
  48975=>"111101010",
  48976=>"100111000",
  48977=>"111110011",
  48978=>"100011000",
  48979=>"111100001",
  48980=>"000101111",
  48981=>"000001011",
  48982=>"010011101",
  48983=>"001110000",
  48984=>"100000110",
  48985=>"110000001",
  48986=>"100001001",
  48987=>"000011100",
  48988=>"000011001",
  48989=>"110000010",
  48990=>"000110010",
  48991=>"100001010",
  48992=>"010001010",
  48993=>"000000000",
  48994=>"100101110",
  48995=>"110011100",
  48996=>"001110101",
  48997=>"011001000",
  48998=>"111110010",
  48999=>"100000000",
  49000=>"010101001",
  49001=>"011101000",
  49002=>"010011010",
  49003=>"110110110",
  49004=>"111000011",
  49005=>"100011010",
  49006=>"100011000",
  49007=>"110000110",
  49008=>"010010001",
  49009=>"111011011",
  49010=>"000111100",
  49011=>"110010100",
  49012=>"010101000",
  49013=>"101001001",
  49014=>"101101111",
  49015=>"001110000",
  49016=>"001100101",
  49017=>"110010010",
  49018=>"001111010",
  49019=>"100010000",
  49020=>"110111101",
  49021=>"000011001",
  49022=>"110001000",
  49023=>"111001010",
  49024=>"110001010",
  49025=>"011010111",
  49026=>"111100010",
  49027=>"100000011",
  49028=>"000000110",
  49029=>"110100001",
  49030=>"000000001",
  49031=>"111111000",
  49032=>"110111010",
  49033=>"000110101",
  49034=>"110010000",
  49035=>"010000001",
  49036=>"101100000",
  49037=>"001110100",
  49038=>"011010000",
  49039=>"011001010",
  49040=>"111011110",
  49041=>"111111011",
  49042=>"011101001",
  49043=>"111011111",
  49044=>"010001000",
  49045=>"001111111",
  49046=>"010010111",
  49047=>"001101001",
  49048=>"000001011",
  49049=>"111111110",
  49050=>"110010001",
  49051=>"100000100",
  49052=>"000111101",
  49053=>"100111101",
  49054=>"100000011",
  49055=>"000110000",
  49056=>"101001000",
  49057=>"011111011",
  49058=>"001000011",
  49059=>"100011100",
  49060=>"110000001",
  49061=>"111110000",
  49062=>"011001001",
  49063=>"010000101",
  49064=>"111001111",
  49065=>"000001010",
  49066=>"011010000",
  49067=>"101110000",
  49068=>"001100000",
  49069=>"000011011",
  49070=>"110100011",
  49071=>"100100111",
  49072=>"000001110",
  49073=>"111011011",
  49074=>"000010001",
  49075=>"111111100",
  49076=>"011101111",
  49077=>"111011000",
  49078=>"010110000",
  49079=>"001011101",
  49080=>"110000011",
  49081=>"100101000",
  49082=>"110010100",
  49083=>"010001111",
  49084=>"101111110",
  49085=>"000001100",
  49086=>"000011110",
  49087=>"010000100",
  49088=>"111100110",
  49089=>"000010111",
  49090=>"011010001",
  49091=>"001110101",
  49092=>"000110110",
  49093=>"000000110",
  49094=>"101101010",
  49095=>"100010000",
  49096=>"001010011",
  49097=>"111000100",
  49098=>"010101000",
  49099=>"001100001",
  49100=>"111000001",
  49101=>"001000110",
  49102=>"101011100",
  49103=>"110111100",
  49104=>"101111000",
  49105=>"011101010",
  49106=>"001001010",
  49107=>"000111000",
  49108=>"111110101",
  49109=>"000011100",
  49110=>"011000010",
  49111=>"001111111",
  49112=>"111001110",
  49113=>"110101110",
  49114=>"110100101",
  49115=>"010100110",
  49116=>"001001111",
  49117=>"111100101",
  49118=>"011110111",
  49119=>"110111001",
  49120=>"011010010",
  49121=>"101101101",
  49122=>"001110000",
  49123=>"100110001",
  49124=>"000111111",
  49125=>"001001100",
  49126=>"100000011",
  49127=>"100110101",
  49128=>"100010110",
  49129=>"000000011",
  49130=>"101011100",
  49131=>"101111001",
  49132=>"010110011",
  49133=>"101011000",
  49134=>"111111101",
  49135=>"111011101",
  49136=>"011000110",
  49137=>"110001100",
  49138=>"101110100",
  49139=>"110001100",
  49140=>"111011011",
  49141=>"000100110",
  49142=>"000000100",
  49143=>"110111011",
  49144=>"111101110",
  49145=>"010011011",
  49146=>"100101010",
  49147=>"101101010",
  49148=>"111011011",
  49149=>"100101101",
  49150=>"100111100",
  49151=>"101101100",
  49152=>"010111001",
  49153=>"010100001",
  49154=>"000010000",
  49155=>"101010101",
  49156=>"011110011",
  49157=>"010000111",
  49158=>"111011110",
  49159=>"110011111",
  49160=>"010010000",
  49161=>"011011110",
  49162=>"010011100",
  49163=>"111000000",
  49164=>"100110100",
  49165=>"010100111",
  49166=>"001011001",
  49167=>"000001101",
  49168=>"111001100",
  49169=>"111101011",
  49170=>"011000000",
  49171=>"100110000",
  49172=>"010010111",
  49173=>"101001001",
  49174=>"000000101",
  49175=>"001111011",
  49176=>"110110111",
  49177=>"011100111",
  49178=>"011011101",
  49179=>"111111110",
  49180=>"001001010",
  49181=>"011100001",
  49182=>"000111000",
  49183=>"000000010",
  49184=>"110100110",
  49185=>"110011011",
  49186=>"001101000",
  49187=>"001101001",
  49188=>"110000110",
  49189=>"001101001",
  49190=>"001010010",
  49191=>"011010111",
  49192=>"100100011",
  49193=>"101101000",
  49194=>"010100001",
  49195=>"111001100",
  49196=>"000000100",
  49197=>"111001010",
  49198=>"000011100",
  49199=>"101010010",
  49200=>"111110100",
  49201=>"110101111",
  49202=>"110010011",
  49203=>"001111000",
  49204=>"001000111",
  49205=>"010010010",
  49206=>"011010001",
  49207=>"011110110",
  49208=>"110001100",
  49209=>"010000010",
  49210=>"111011111",
  49211=>"100010001",
  49212=>"010101010",
  49213=>"110101010",
  49214=>"010100000",
  49215=>"100010001",
  49216=>"000100110",
  49217=>"010100101",
  49218=>"010001110",
  49219=>"101010100",
  49220=>"100010000",
  49221=>"100011000",
  49222=>"000000111",
  49223=>"000010111",
  49224=>"010111111",
  49225=>"100100110",
  49226=>"011011000",
  49227=>"101000101",
  49228=>"101111001",
  49229=>"101100111",
  49230=>"010010001",
  49231=>"100100000",
  49232=>"000111110",
  49233=>"000000000",
  49234=>"011001111",
  49235=>"010000110",
  49236=>"000000010",
  49237=>"000101000",
  49238=>"100110110",
  49239=>"010100111",
  49240=>"000111111",
  49241=>"011011000",
  49242=>"110100101",
  49243=>"010010001",
  49244=>"111100001",
  49245=>"111101000",
  49246=>"010000100",
  49247=>"010110001",
  49248=>"010000001",
  49249=>"001111100",
  49250=>"111111111",
  49251=>"111101010",
  49252=>"000001010",
  49253=>"101001100",
  49254=>"010001100",
  49255=>"100000100",
  49256=>"101010001",
  49257=>"001010011",
  49258=>"010011011",
  49259=>"100101100",
  49260=>"011101001",
  49261=>"000000111",
  49262=>"011000000",
  49263=>"111111111",
  49264=>"010100011",
  49265=>"110110001",
  49266=>"011111101",
  49267=>"110010110",
  49268=>"000011001",
  49269=>"101110100",
  49270=>"101000100",
  49271=>"101000111",
  49272=>"101000010",
  49273=>"001111001",
  49274=>"100110100",
  49275=>"111100110",
  49276=>"110101011",
  49277=>"001111011",
  49278=>"011011000",
  49279=>"101101101",
  49280=>"111111011",
  49281=>"111011001",
  49282=>"110111101",
  49283=>"101000100",
  49284=>"111010000",
  49285=>"101011111",
  49286=>"010000101",
  49287=>"011100110",
  49288=>"110000110",
  49289=>"000011011",
  49290=>"001010101",
  49291=>"010001110",
  49292=>"000010000",
  49293=>"101110010",
  49294=>"010111000",
  49295=>"010111101",
  49296=>"101001111",
  49297=>"001001000",
  49298=>"001110100",
  49299=>"011011110",
  49300=>"100000000",
  49301=>"010101001",
  49302=>"111011110",
  49303=>"111100111",
  49304=>"111101110",
  49305=>"000100101",
  49306=>"000011110",
  49307=>"101010000",
  49308=>"000001101",
  49309=>"110100000",
  49310=>"101100111",
  49311=>"111111001",
  49312=>"110001101",
  49313=>"000000001",
  49314=>"110110010",
  49315=>"000000101",
  49316=>"111100110",
  49317=>"010100010",
  49318=>"011011100",
  49319=>"110000010",
  49320=>"001011100",
  49321=>"000001100",
  49322=>"101111111",
  49323=>"111111101",
  49324=>"011000001",
  49325=>"000010100",
  49326=>"011011011",
  49327=>"001101100",
  49328=>"001010110",
  49329=>"000010011",
  49330=>"100111010",
  49331=>"010011011",
  49332=>"111011100",
  49333=>"111111001",
  49334=>"110101011",
  49335=>"110001000",
  49336=>"001101110",
  49337=>"110010011",
  49338=>"110000110",
  49339=>"111000010",
  49340=>"110100001",
  49341=>"100010010",
  49342=>"000101100",
  49343=>"101000101",
  49344=>"100010001",
  49345=>"000011110",
  49346=>"001100000",
  49347=>"101011001",
  49348=>"001000110",
  49349=>"101100111",
  49350=>"000110000",
  49351=>"000101100",
  49352=>"011000001",
  49353=>"110010101",
  49354=>"010010110",
  49355=>"111111001",
  49356=>"111001010",
  49357=>"011010000",
  49358=>"111000010",
  49359=>"100111100",
  49360=>"101111000",
  49361=>"100111000",
  49362=>"101001111",
  49363=>"001010111",
  49364=>"001000010",
  49365=>"110001010",
  49366=>"101001101",
  49367=>"100111101",
  49368=>"111100011",
  49369=>"000010101",
  49370=>"101000110",
  49371=>"000000011",
  49372=>"001001001",
  49373=>"101011001",
  49374=>"001100000",
  49375=>"010000101",
  49376=>"111011101",
  49377=>"101101001",
  49378=>"100010100",
  49379=>"010001001",
  49380=>"001001101",
  49381=>"111111001",
  49382=>"111110001",
  49383=>"010111111",
  49384=>"100011011",
  49385=>"101000100",
  49386=>"000101001",
  49387=>"101010101",
  49388=>"100000000",
  49389=>"100101001",
  49390=>"100010001",
  49391=>"010001111",
  49392=>"010011001",
  49393=>"001101011",
  49394=>"011011001",
  49395=>"011011000",
  49396=>"111010010",
  49397=>"110011001",
  49398=>"101111110",
  49399=>"010111010",
  49400=>"000111101",
  49401=>"100101001",
  49402=>"110011000",
  49403=>"000110010",
  49404=>"001000111",
  49405=>"111000011",
  49406=>"101000100",
  49407=>"000101100",
  49408=>"111111000",
  49409=>"001101110",
  49410=>"001110101",
  49411=>"111110101",
  49412=>"000001001",
  49413=>"011100001",
  49414=>"110011111",
  49415=>"001101000",
  49416=>"100100110",
  49417=>"101010010",
  49418=>"001111011",
  49419=>"010010010",
  49420=>"000110001",
  49421=>"111110000",
  49422=>"010001101",
  49423=>"010001001",
  49424=>"001001100",
  49425=>"011101111",
  49426=>"111011101",
  49427=>"111010000",
  49428=>"100000110",
  49429=>"110000000",
  49430=>"000011011",
  49431=>"000110111",
  49432=>"110000000",
  49433=>"101111001",
  49434=>"010001010",
  49435=>"111111010",
  49436=>"000001010",
  49437=>"001111011",
  49438=>"000111001",
  49439=>"100010100",
  49440=>"111001100",
  49441=>"011011001",
  49442=>"010111001",
  49443=>"111010111",
  49444=>"001111110",
  49445=>"101010101",
  49446=>"001111100",
  49447=>"110101011",
  49448=>"101011101",
  49449=>"011010010",
  49450=>"000101101",
  49451=>"011011101",
  49452=>"100011010",
  49453=>"011001010",
  49454=>"011001000",
  49455=>"001001010",
  49456=>"010000011",
  49457=>"011000001",
  49458=>"110111110",
  49459=>"101011101",
  49460=>"110100011",
  49461=>"111000110",
  49462=>"111110110",
  49463=>"011011111",
  49464=>"101001100",
  49465=>"010110011",
  49466=>"101100111",
  49467=>"001000111",
  49468=>"111011100",
  49469=>"111100100",
  49470=>"000010111",
  49471=>"110111010",
  49472=>"011100101",
  49473=>"101011010",
  49474=>"001011000",
  49475=>"101010001",
  49476=>"100010100",
  49477=>"001011011",
  49478=>"111110101",
  49479=>"100110100",
  49480=>"010000000",
  49481=>"010101101",
  49482=>"111110000",
  49483=>"110110000",
  49484=>"101010001",
  49485=>"001011010",
  49486=>"001010110",
  49487=>"000101000",
  49488=>"011111101",
  49489=>"000101110",
  49490=>"100110011",
  49491=>"111010110",
  49492=>"110100001",
  49493=>"110011001",
  49494=>"111010111",
  49495=>"011000111",
  49496=>"000110001",
  49497=>"100001001",
  49498=>"001011110",
  49499=>"000000001",
  49500=>"011000001",
  49501=>"000100111",
  49502=>"000010011",
  49503=>"101011010",
  49504=>"110011011",
  49505=>"100010110",
  49506=>"101110001",
  49507=>"000000000",
  49508=>"110101111",
  49509=>"101000101",
  49510=>"001100001",
  49511=>"101111100",
  49512=>"011010011",
  49513=>"010111000",
  49514=>"101111111",
  49515=>"101111001",
  49516=>"000000110",
  49517=>"001111010",
  49518=>"111001011",
  49519=>"001100001",
  49520=>"011000011",
  49521=>"000111110",
  49522=>"111101111",
  49523=>"100000011",
  49524=>"000000110",
  49525=>"111111101",
  49526=>"011001010",
  49527=>"111000010",
  49528=>"110110111",
  49529=>"000101100",
  49530=>"011001011",
  49531=>"011000101",
  49532=>"110010010",
  49533=>"011011111",
  49534=>"101000011",
  49535=>"001010000",
  49536=>"111111001",
  49537=>"001011100",
  49538=>"101111011",
  49539=>"110011111",
  49540=>"111001011",
  49541=>"111110100",
  49542=>"100100100",
  49543=>"100110001",
  49544=>"001100101",
  49545=>"011000100",
  49546=>"111111111",
  49547=>"111111011",
  49548=>"001101110",
  49549=>"110100000",
  49550=>"000101010",
  49551=>"110101101",
  49552=>"011111111",
  49553=>"100001110",
  49554=>"000110110",
  49555=>"000010011",
  49556=>"100000110",
  49557=>"110000000",
  49558=>"010001011",
  49559=>"100010001",
  49560=>"011101001",
  49561=>"001001110",
  49562=>"000100101",
  49563=>"001110000",
  49564=>"001010111",
  49565=>"100011001",
  49566=>"100100100",
  49567=>"100011010",
  49568=>"010100000",
  49569=>"010011000",
  49570=>"111110000",
  49571=>"110010010",
  49572=>"100000101",
  49573=>"111011011",
  49574=>"000100100",
  49575=>"000000101",
  49576=>"010100111",
  49577=>"110100111",
  49578=>"010010100",
  49579=>"001110001",
  49580=>"000011000",
  49581=>"111111111",
  49582=>"100101101",
  49583=>"100110101",
  49584=>"010011001",
  49585=>"101001101",
  49586=>"111111000",
  49587=>"100010010",
  49588=>"010011110",
  49589=>"100000010",
  49590=>"001001010",
  49591=>"100011111",
  49592=>"000101111",
  49593=>"001000010",
  49594=>"101010010",
  49595=>"000111010",
  49596=>"111111100",
  49597=>"101000001",
  49598=>"011110001",
  49599=>"110101101",
  49600=>"101111100",
  49601=>"101010001",
  49602=>"011010111",
  49603=>"001101011",
  49604=>"100111100",
  49605=>"110110001",
  49606=>"111001011",
  49607=>"000000010",
  49608=>"010110010",
  49609=>"011010110",
  49610=>"000000101",
  49611=>"101000110",
  49612=>"010100010",
  49613=>"000000011",
  49614=>"010000110",
  49615=>"001001110",
  49616=>"101011110",
  49617=>"100011001",
  49618=>"000001001",
  49619=>"011001000",
  49620=>"010101010",
  49621=>"111001101",
  49622=>"110101110",
  49623=>"110001000",
  49624=>"001100001",
  49625=>"010010100",
  49626=>"001110111",
  49627=>"111010100",
  49628=>"111001100",
  49629=>"101010000",
  49630=>"100111100",
  49631=>"101110000",
  49632=>"011011000",
  49633=>"010110100",
  49634=>"011111100",
  49635=>"101101111",
  49636=>"001111000",
  49637=>"100010110",
  49638=>"011001100",
  49639=>"011100111",
  49640=>"110100011",
  49641=>"111100101",
  49642=>"010100101",
  49643=>"101110111",
  49644=>"100011110",
  49645=>"110000111",
  49646=>"011000011",
  49647=>"110000100",
  49648=>"100111010",
  49649=>"000010111",
  49650=>"101100011",
  49651=>"111011111",
  49652=>"011100100",
  49653=>"001000111",
  49654=>"001110001",
  49655=>"001010001",
  49656=>"110100100",
  49657=>"110010111",
  49658=>"001000010",
  49659=>"001111101",
  49660=>"011110110",
  49661=>"111101100",
  49662=>"011010011",
  49663=>"110011000",
  49664=>"110100100",
  49665=>"010110100",
  49666=>"100101111",
  49667=>"001110111",
  49668=>"101011110",
  49669=>"010101000",
  49670=>"110000111",
  49671=>"010110111",
  49672=>"000111010",
  49673=>"010000110",
  49674=>"110010011",
  49675=>"001110100",
  49676=>"100101000",
  49677=>"010111100",
  49678=>"101110001",
  49679=>"101011010",
  49680=>"111000001",
  49681=>"100101110",
  49682=>"100010100",
  49683=>"100010100",
  49684=>"101101111",
  49685=>"001000000",
  49686=>"100010010",
  49687=>"010001101",
  49688=>"101100111",
  49689=>"101100101",
  49690=>"011000111",
  49691=>"000000111",
  49692=>"000011111",
  49693=>"100101010",
  49694=>"111111111",
  49695=>"110001100",
  49696=>"000011000",
  49697=>"001010110",
  49698=>"100001010",
  49699=>"101111111",
  49700=>"000110100",
  49701=>"001000011",
  49702=>"010011100",
  49703=>"101011111",
  49704=>"100011111",
  49705=>"000100001",
  49706=>"110000100",
  49707=>"100011100",
  49708=>"000100001",
  49709=>"000010111",
  49710=>"010100111",
  49711=>"110000011",
  49712=>"101011111",
  49713=>"010100010",
  49714=>"111101101",
  49715=>"001001010",
  49716=>"100000000",
  49717=>"110100011",
  49718=>"010011110",
  49719=>"110010001",
  49720=>"110110110",
  49721=>"110110010",
  49722=>"101101101",
  49723=>"010001111",
  49724=>"100001111",
  49725=>"011010111",
  49726=>"100011111",
  49727=>"000101010",
  49728=>"101101000",
  49729=>"101010001",
  49730=>"001100010",
  49731=>"011000110",
  49732=>"000110100",
  49733=>"101101101",
  49734=>"100011011",
  49735=>"001001111",
  49736=>"111011110",
  49737=>"111111110",
  49738=>"011000111",
  49739=>"111110111",
  49740=>"100101011",
  49741=>"001000110",
  49742=>"111101100",
  49743=>"000110111",
  49744=>"000000111",
  49745=>"000000010",
  49746=>"101111111",
  49747=>"000000010",
  49748=>"000100010",
  49749=>"010100100",
  49750=>"001010110",
  49751=>"000101100",
  49752=>"011101110",
  49753=>"001100101",
  49754=>"010110000",
  49755=>"000111111",
  49756=>"001100000",
  49757=>"110000100",
  49758=>"111000111",
  49759=>"000000000",
  49760=>"111010101",
  49761=>"010111011",
  49762=>"101010100",
  49763=>"000000001",
  49764=>"101101000",
  49765=>"100100010",
  49766=>"110011101",
  49767=>"101101100",
  49768=>"001100110",
  49769=>"010011011",
  49770=>"110011010",
  49771=>"000011101",
  49772=>"111010101",
  49773=>"001010100",
  49774=>"001101011",
  49775=>"111111011",
  49776=>"101100011",
  49777=>"001010000",
  49778=>"101110101",
  49779=>"010000000",
  49780=>"110110101",
  49781=>"101000010",
  49782=>"000000001",
  49783=>"100000011",
  49784=>"100100000",
  49785=>"010110110",
  49786=>"101001111",
  49787=>"111110101",
  49788=>"000011000",
  49789=>"100001001",
  49790=>"101101110",
  49791=>"110011100",
  49792=>"111010110",
  49793=>"011011111",
  49794=>"001000010",
  49795=>"110110011",
  49796=>"011101101",
  49797=>"100010111",
  49798=>"000011101",
  49799=>"000101000",
  49800=>"010010101",
  49801=>"001100001",
  49802=>"100100101",
  49803=>"111101110",
  49804=>"001100001",
  49805=>"111111100",
  49806=>"001111101",
  49807=>"000100001",
  49808=>"110000101",
  49809=>"110000111",
  49810=>"010111101",
  49811=>"010001000",
  49812=>"001001011",
  49813=>"001010100",
  49814=>"011110010",
  49815=>"100111011",
  49816=>"110001000",
  49817=>"001001001",
  49818=>"000101111",
  49819=>"010110000",
  49820=>"101010110",
  49821=>"100101111",
  49822=>"010011010",
  49823=>"010111101",
  49824=>"110010101",
  49825=>"010101000",
  49826=>"011101001",
  49827=>"001101100",
  49828=>"011111011",
  49829=>"110011000",
  49830=>"011110100",
  49831=>"000100000",
  49832=>"000001011",
  49833=>"001110001",
  49834=>"100100010",
  49835=>"110001001",
  49836=>"010101100",
  49837=>"110100100",
  49838=>"111010011",
  49839=>"000101110",
  49840=>"100000010",
  49841=>"011000001",
  49842=>"111011011",
  49843=>"011101101",
  49844=>"111010101",
  49845=>"110100010",
  49846=>"001010111",
  49847=>"010010111",
  49848=>"000100011",
  49849=>"011011110",
  49850=>"100011100",
  49851=>"100101000",
  49852=>"000000000",
  49853=>"001001111",
  49854=>"111000000",
  49855=>"011010110",
  49856=>"000010011",
  49857=>"000001000",
  49858=>"011111101",
  49859=>"111110101",
  49860=>"001010100",
  49861=>"100101001",
  49862=>"011000100",
  49863=>"100111001",
  49864=>"111110101",
  49865=>"110001000",
  49866=>"011010101",
  49867=>"101010000",
  49868=>"100010000",
  49869=>"001111100",
  49870=>"010011000",
  49871=>"101101000",
  49872=>"110111010",
  49873=>"101111100",
  49874=>"000110011",
  49875=>"100011001",
  49876=>"010101010",
  49877=>"000010000",
  49878=>"000100101",
  49879=>"111000100",
  49880=>"010011101",
  49881=>"000001001",
  49882=>"010001110",
  49883=>"101000010",
  49884=>"111001101",
  49885=>"010000000",
  49886=>"000000011",
  49887=>"111100000",
  49888=>"011010000",
  49889=>"001100100",
  49890=>"001011110",
  49891=>"011000000",
  49892=>"011101101",
  49893=>"111001000",
  49894=>"000101010",
  49895=>"011110011",
  49896=>"001100011",
  49897=>"100010011",
  49898=>"010111001",
  49899=>"001010101",
  49900=>"010001010",
  49901=>"101011110",
  49902=>"000010011",
  49903=>"111101000",
  49904=>"000100101",
  49905=>"000111000",
  49906=>"000010100",
  49907=>"000010000",
  49908=>"110101011",
  49909=>"101010011",
  49910=>"001101011",
  49911=>"001111011",
  49912=>"111110011",
  49913=>"001010101",
  49914=>"111001100",
  49915=>"010101111",
  49916=>"101110101",
  49917=>"100100011",
  49918=>"100001000",
  49919=>"010010110",
  49920=>"100101011",
  49921=>"110110111",
  49922=>"101001001",
  49923=>"100011101",
  49924=>"110111001",
  49925=>"010000010",
  49926=>"111011001",
  49927=>"100010101",
  49928=>"001101010",
  49929=>"010100011",
  49930=>"001101101",
  49931=>"000101010",
  49932=>"010010101",
  49933=>"110010000",
  49934=>"001000001",
  49935=>"110011101",
  49936=>"011100111",
  49937=>"010100111",
  49938=>"111110111",
  49939=>"001100011",
  49940=>"010000000",
  49941=>"111111101",
  49942=>"011001110",
  49943=>"011101001",
  49944=>"000011011",
  49945=>"000010010",
  49946=>"001000011",
  49947=>"110100110",
  49948=>"101101111",
  49949=>"110100100",
  49950=>"100111010",
  49951=>"101100010",
  49952=>"111011100",
  49953=>"100110010",
  49954=>"100011011",
  49955=>"001100001",
  49956=>"111100001",
  49957=>"100011011",
  49958=>"111110010",
  49959=>"110000011",
  49960=>"110011111",
  49961=>"101101001",
  49962=>"111100010",
  49963=>"010100101",
  49964=>"001011100",
  49965=>"110101010",
  49966=>"011111010",
  49967=>"001101010",
  49968=>"000101101",
  49969=>"101001001",
  49970=>"000101000",
  49971=>"100010110",
  49972=>"011000010",
  49973=>"111111111",
  49974=>"110111111",
  49975=>"010111000",
  49976=>"000101011",
  49977=>"010001000",
  49978=>"100000110",
  49979=>"101011000",
  49980=>"000101110",
  49981=>"110111100",
  49982=>"000110011",
  49983=>"010000111",
  49984=>"010000101",
  49985=>"010110011",
  49986=>"011001111",
  49987=>"000000011",
  49988=>"101010110",
  49989=>"110100010",
  49990=>"101010110",
  49991=>"100011000",
  49992=>"001101111",
  49993=>"110001111",
  49994=>"101001100",
  49995=>"000010010",
  49996=>"101001000",
  49997=>"101101001",
  49998=>"110001111",
  49999=>"110011001",
  50000=>"101100110",
  50001=>"001000100",
  50002=>"100000111",
  50003=>"000101101",
  50004=>"111000110",
  50005=>"001000000",
  50006=>"010010010",
  50007=>"011010010",
  50008=>"000011011",
  50009=>"000111011",
  50010=>"000111110",
  50011=>"010110000",
  50012=>"011101110",
  50013=>"100011100",
  50014=>"100100110",
  50015=>"001001101",
  50016=>"000111100",
  50017=>"111111011",
  50018=>"001011000",
  50019=>"111001101",
  50020=>"010100001",
  50021=>"000111110",
  50022=>"010100011",
  50023=>"111111100",
  50024=>"100010111",
  50025=>"100011000",
  50026=>"100011010",
  50027=>"111100111",
  50028=>"110111010",
  50029=>"101011100",
  50030=>"000101100",
  50031=>"111101000",
  50032=>"100000100",
  50033=>"111001101",
  50034=>"111111101",
  50035=>"011101100",
  50036=>"100010101",
  50037=>"010010001",
  50038=>"100101111",
  50039=>"100000100",
  50040=>"011100011",
  50041=>"011001001",
  50042=>"111101110",
  50043=>"111000101",
  50044=>"100101000",
  50045=>"110111000",
  50046=>"110011010",
  50047=>"110000101",
  50048=>"000101110",
  50049=>"101010000",
  50050=>"110101001",
  50051=>"010001000",
  50052=>"100100000",
  50053=>"100101000",
  50054=>"101110111",
  50055=>"111100100",
  50056=>"110100000",
  50057=>"101011010",
  50058=>"111101010",
  50059=>"111010111",
  50060=>"111010110",
  50061=>"101000011",
  50062=>"110100011",
  50063=>"111100111",
  50064=>"100001111",
  50065=>"010000100",
  50066=>"000011001",
  50067=>"100100000",
  50068=>"101101111",
  50069=>"010101100",
  50070=>"111110000",
  50071=>"011110110",
  50072=>"110011101",
  50073=>"010100011",
  50074=>"011000001",
  50075=>"000111001",
  50076=>"110111001",
  50077=>"011000001",
  50078=>"010100001",
  50079=>"101000100",
  50080=>"000000000",
  50081=>"101101101",
  50082=>"001001111",
  50083=>"001110010",
  50084=>"101001110",
  50085=>"010010010",
  50086=>"010010011",
  50087=>"111111101",
  50088=>"001000100",
  50089=>"111100101",
  50090=>"000010111",
  50091=>"100011101",
  50092=>"000010110",
  50093=>"000011101",
  50094=>"110000111",
  50095=>"000011110",
  50096=>"011101110",
  50097=>"100000000",
  50098=>"000001111",
  50099=>"100010100",
  50100=>"001110100",
  50101=>"111000000",
  50102=>"101010110",
  50103=>"100110101",
  50104=>"010001001",
  50105=>"110100011",
  50106=>"111100101",
  50107=>"000001010",
  50108=>"010100010",
  50109=>"010010000",
  50110=>"100111110",
  50111=>"101100000",
  50112=>"101100111",
  50113=>"110111000",
  50114=>"010000001",
  50115=>"101001110",
  50116=>"011110011",
  50117=>"011000000",
  50118=>"111000110",
  50119=>"111111111",
  50120=>"011111001",
  50121=>"110001101",
  50122=>"101010000",
  50123=>"100101011",
  50124=>"101110110",
  50125=>"001000110",
  50126=>"110000010",
  50127=>"000110101",
  50128=>"111000001",
  50129=>"000010001",
  50130=>"011011011",
  50131=>"001001101",
  50132=>"010110000",
  50133=>"100001011",
  50134=>"000011001",
  50135=>"010101011",
  50136=>"001010000",
  50137=>"110010100",
  50138=>"010001010",
  50139=>"000000000",
  50140=>"010101100",
  50141=>"010000000",
  50142=>"011011011",
  50143=>"100101011",
  50144=>"010011011",
  50145=>"110001100",
  50146=>"010110101",
  50147=>"100111111",
  50148=>"000010000",
  50149=>"101001001",
  50150=>"110011010",
  50151=>"000100011",
  50152=>"111010010",
  50153=>"101111010",
  50154=>"000010111",
  50155=>"101110001",
  50156=>"111011011",
  50157=>"101101111",
  50158=>"010000000",
  50159=>"011000110",
  50160=>"011110000",
  50161=>"111111011",
  50162=>"100010111",
  50163=>"010100001",
  50164=>"110111111",
  50165=>"100110011",
  50166=>"001111000",
  50167=>"000110011",
  50168=>"111001101",
  50169=>"100101101",
  50170=>"000100000",
  50171=>"001100111",
  50172=>"111011100",
  50173=>"100011101",
  50174=>"000001001",
  50175=>"100110100",
  50176=>"111101010",
  50177=>"111110011",
  50178=>"110100010",
  50179=>"000000110",
  50180=>"100001011",
  50181=>"000011010",
  50182=>"001111001",
  50183=>"001011100",
  50184=>"100110101",
  50185=>"011001001",
  50186=>"001100110",
  50187=>"010111111",
  50188=>"111101011",
  50189=>"000111101",
  50190=>"111100011",
  50191=>"101010011",
  50192=>"010110001",
  50193=>"101000100",
  50194=>"100100011",
  50195=>"101000001",
  50196=>"101101000",
  50197=>"101010111",
  50198=>"110111110",
  50199=>"010011011",
  50200=>"100100000",
  50201=>"110101011",
  50202=>"010010111",
  50203=>"111001111",
  50204=>"110001010",
  50205=>"001100100",
  50206=>"111000100",
  50207=>"110011011",
  50208=>"000001100",
  50209=>"101101111",
  50210=>"111000010",
  50211=>"000100101",
  50212=>"000100000",
  50213=>"011010001",
  50214=>"010110111",
  50215=>"110101111",
  50216=>"110110100",
  50217=>"000110101",
  50218=>"001000010",
  50219=>"110101100",
  50220=>"110001011",
  50221=>"111110001",
  50222=>"001100100",
  50223=>"111110011",
  50224=>"100011001",
  50225=>"010010101",
  50226=>"101001110",
  50227=>"011011100",
  50228=>"100011011",
  50229=>"010101011",
  50230=>"000000010",
  50231=>"110001110",
  50232=>"110010001",
  50233=>"000101011",
  50234=>"111010000",
  50235=>"010100110",
  50236=>"000000100",
  50237=>"011010110",
  50238=>"110010100",
  50239=>"100111101",
  50240=>"010101000",
  50241=>"110011001",
  50242=>"110101111",
  50243=>"011001011",
  50244=>"100011011",
  50245=>"100001111",
  50246=>"111111001",
  50247=>"000011011",
  50248=>"101001110",
  50249=>"011101111",
  50250=>"001111001",
  50251=>"011111000",
  50252=>"001000101",
  50253=>"001100000",
  50254=>"011010111",
  50255=>"111101111",
  50256=>"100100001",
  50257=>"111111001",
  50258=>"010011000",
  50259=>"110110101",
  50260=>"011101101",
  50261=>"001111100",
  50262=>"000100010",
  50263=>"001010000",
  50264=>"000001100",
  50265=>"011000101",
  50266=>"100010110",
  50267=>"110000101",
  50268=>"001001100",
  50269=>"000101000",
  50270=>"100000011",
  50271=>"000011010",
  50272=>"111111011",
  50273=>"110011110",
  50274=>"111101101",
  50275=>"010110011",
  50276=>"011011000",
  50277=>"111111100",
  50278=>"101011110",
  50279=>"111101101",
  50280=>"001001001",
  50281=>"111100111",
  50282=>"100001101",
  50283=>"111010010",
  50284=>"001110011",
  50285=>"000010110",
  50286=>"011100011",
  50287=>"001001101",
  50288=>"000110101",
  50289=>"010010011",
  50290=>"110111000",
  50291=>"110111010",
  50292=>"000010110",
  50293=>"001100010",
  50294=>"110111001",
  50295=>"000101111",
  50296=>"101110100",
  50297=>"110111111",
  50298=>"111001010",
  50299=>"110010111",
  50300=>"000001001",
  50301=>"000010010",
  50302=>"101001010",
  50303=>"000101100",
  50304=>"100110010",
  50305=>"000100000",
  50306=>"010011110",
  50307=>"010111001",
  50308=>"000000011",
  50309=>"000001111",
  50310=>"001000110",
  50311=>"101001111",
  50312=>"001001010",
  50313=>"010011101",
  50314=>"001000011",
  50315=>"110111101",
  50316=>"001110000",
  50317=>"110100111",
  50318=>"111010010",
  50319=>"010101101",
  50320=>"001011011",
  50321=>"001001111",
  50322=>"000100101",
  50323=>"111101001",
  50324=>"110111110",
  50325=>"011111100",
  50326=>"001100011",
  50327=>"111011100",
  50328=>"101100111",
  50329=>"100111001",
  50330=>"100110001",
  50331=>"010101100",
  50332=>"011000001",
  50333=>"101011100",
  50334=>"101001110",
  50335=>"011010010",
  50336=>"001011101",
  50337=>"110011001",
  50338=>"101100100",
  50339=>"000010010",
  50340=>"010001110",
  50341=>"000100001",
  50342=>"011110111",
  50343=>"101010010",
  50344=>"101100001",
  50345=>"111001100",
  50346=>"010010110",
  50347=>"000101101",
  50348=>"101010011",
  50349=>"111011011",
  50350=>"110111100",
  50351=>"010001110",
  50352=>"000011101",
  50353=>"100000110",
  50354=>"110100001",
  50355=>"100011010",
  50356=>"110001011",
  50357=>"011001000",
  50358=>"000011100",
  50359=>"000001110",
  50360=>"010111111",
  50361=>"011010110",
  50362=>"010000100",
  50363=>"001110100",
  50364=>"111111100",
  50365=>"110101110",
  50366=>"001010000",
  50367=>"111001011",
  50368=>"101011010",
  50369=>"011011101",
  50370=>"111110100",
  50371=>"111000000",
  50372=>"011010000",
  50373=>"001001110",
  50374=>"110001010",
  50375=>"001000110",
  50376=>"010010100",
  50377=>"010001010",
  50378=>"011001100",
  50379=>"110111010",
  50380=>"111111110",
  50381=>"001001001",
  50382=>"000101111",
  50383=>"111110101",
  50384=>"111001010",
  50385=>"011010010",
  50386=>"001111011",
  50387=>"001011000",
  50388=>"010011010",
  50389=>"001010011",
  50390=>"011100111",
  50391=>"010110100",
  50392=>"100000110",
  50393=>"001001111",
  50394=>"100100010",
  50395=>"010001000",
  50396=>"001111010",
  50397=>"000111101",
  50398=>"110010111",
  50399=>"101110000",
  50400=>"000000001",
  50401=>"011111010",
  50402=>"000110000",
  50403=>"001011000",
  50404=>"010000111",
  50405=>"001101000",
  50406=>"001000000",
  50407=>"101110011",
  50408=>"000010011",
  50409=>"111000111",
  50410=>"011011110",
  50411=>"010101100",
  50412=>"110101100",
  50413=>"101001110",
  50414=>"000110110",
  50415=>"001111111",
  50416=>"000101111",
  50417=>"111010010",
  50418=>"001011011",
  50419=>"101011110",
  50420=>"001010100",
  50421=>"000011010",
  50422=>"101110111",
  50423=>"000111001",
  50424=>"111000000",
  50425=>"100000000",
  50426=>"010001111",
  50427=>"101001011",
  50428=>"010010001",
  50429=>"000101100",
  50430=>"000011101",
  50431=>"001001010",
  50432=>"111100010",
  50433=>"111001000",
  50434=>"100111001",
  50435=>"101000001",
  50436=>"011100011",
  50437=>"010000111",
  50438=>"110011100",
  50439=>"001010110",
  50440=>"011110100",
  50441=>"000001011",
  50442=>"100010100",
  50443=>"111001100",
  50444=>"001111110",
  50445=>"111111111",
  50446=>"000110110",
  50447=>"011000101",
  50448=>"010111000",
  50449=>"000110000",
  50450=>"100010010",
  50451=>"001111110",
  50452=>"100010001",
  50453=>"000010100",
  50454=>"000101001",
  50455=>"010011111",
  50456=>"011000000",
  50457=>"110100001",
  50458=>"001011000",
  50459=>"111001000",
  50460=>"100100110",
  50461=>"001100100",
  50462=>"010100110",
  50463=>"011000000",
  50464=>"111100010",
  50465=>"011110111",
  50466=>"001100011",
  50467=>"000010000",
  50468=>"111100110",
  50469=>"101111000",
  50470=>"000011100",
  50471=>"000110010",
  50472=>"000000011",
  50473=>"101110011",
  50474=>"100001100",
  50475=>"100100010",
  50476=>"110000001",
  50477=>"000011010",
  50478=>"000010011",
  50479=>"101110111",
  50480=>"001001110",
  50481=>"111110110",
  50482=>"001101011",
  50483=>"010001101",
  50484=>"000000001",
  50485=>"001001000",
  50486=>"000111011",
  50487=>"110100011",
  50488=>"000100011",
  50489=>"011001111",
  50490=>"011010111",
  50491=>"011011000",
  50492=>"000000100",
  50493=>"101111000",
  50494=>"010011000",
  50495=>"001111101",
  50496=>"110110100",
  50497=>"000110110",
  50498=>"100111111",
  50499=>"100010100",
  50500=>"010101111",
  50501=>"000001011",
  50502=>"010010001",
  50503=>"101001011",
  50504=>"011110000",
  50505=>"101011101",
  50506=>"100100000",
  50507=>"010001110",
  50508=>"110010001",
  50509=>"110000101",
  50510=>"100001001",
  50511=>"011111010",
  50512=>"011110001",
  50513=>"100011101",
  50514=>"000010100",
  50515=>"010111010",
  50516=>"111011101",
  50517=>"011000110",
  50518=>"101010000",
  50519=>"110100101",
  50520=>"010001011",
  50521=>"010100110",
  50522=>"001101001",
  50523=>"100011000",
  50524=>"001111100",
  50525=>"101101010",
  50526=>"111001010",
  50527=>"010010010",
  50528=>"000011111",
  50529=>"101010100",
  50530=>"010010010",
  50531=>"001000101",
  50532=>"001101111",
  50533=>"010010000",
  50534=>"000001111",
  50535=>"101100000",
  50536=>"010111001",
  50537=>"001001000",
  50538=>"101001100",
  50539=>"000001011",
  50540=>"011011100",
  50541=>"000001000",
  50542=>"000011010",
  50543=>"001110010",
  50544=>"000010100",
  50545=>"111010100",
  50546=>"010010010",
  50547=>"111110000",
  50548=>"001011101",
  50549=>"110111111",
  50550=>"011010000",
  50551=>"110101101",
  50552=>"101010100",
  50553=>"001001110",
  50554=>"111001100",
  50555=>"001111000",
  50556=>"010101110",
  50557=>"001100001",
  50558=>"111011110",
  50559=>"111001101",
  50560=>"000100010",
  50561=>"001101100",
  50562=>"110011110",
  50563=>"001011010",
  50564=>"101010000",
  50565=>"101010011",
  50566=>"010101001",
  50567=>"100000001",
  50568=>"000000000",
  50569=>"110101011",
  50570=>"100101101",
  50571=>"001000100",
  50572=>"011111101",
  50573=>"000000010",
  50574=>"110001101",
  50575=>"110111010",
  50576=>"000000111",
  50577=>"010100100",
  50578=>"000100101",
  50579=>"001110101",
  50580=>"011110010",
  50581=>"001010011",
  50582=>"111001001",
  50583=>"111000000",
  50584=>"001111110",
  50585=>"000001010",
  50586=>"000110100",
  50587=>"001101101",
  50588=>"001111100",
  50589=>"001101001",
  50590=>"101100011",
  50591=>"010110100",
  50592=>"010100011",
  50593=>"011111000",
  50594=>"110011010",
  50595=>"000000101",
  50596=>"011100110",
  50597=>"111100111",
  50598=>"101111001",
  50599=>"101101101",
  50600=>"111000001",
  50601=>"000010111",
  50602=>"000110110",
  50603=>"000010111",
  50604=>"010101000",
  50605=>"011001001",
  50606=>"011101000",
  50607=>"001100101",
  50608=>"000010000",
  50609=>"010010110",
  50610=>"011101100",
  50611=>"011001011",
  50612=>"001000100",
  50613=>"101011110",
  50614=>"100010000",
  50615=>"100000101",
  50616=>"010011000",
  50617=>"010011101",
  50618=>"101000000",
  50619=>"101110110",
  50620=>"010110110",
  50621=>"100100011",
  50622=>"011101010",
  50623=>"110110001",
  50624=>"101010100",
  50625=>"001101100",
  50626=>"001000111",
  50627=>"100110000",
  50628=>"010110000",
  50629=>"001010010",
  50630=>"110100111",
  50631=>"011001000",
  50632=>"100100011",
  50633=>"101110101",
  50634=>"000010110",
  50635=>"101000111",
  50636=>"000010011",
  50637=>"110010111",
  50638=>"110000011",
  50639=>"010111001",
  50640=>"100110111",
  50641=>"000000011",
  50642=>"110100000",
  50643=>"110100111",
  50644=>"101110011",
  50645=>"000000010",
  50646=>"001111100",
  50647=>"101110110",
  50648=>"110100111",
  50649=>"111101011",
  50650=>"010110001",
  50651=>"100000000",
  50652=>"100110111",
  50653=>"100111100",
  50654=>"101101001",
  50655=>"001001101",
  50656=>"101110111",
  50657=>"001010111",
  50658=>"111000001",
  50659=>"110110000",
  50660=>"011111111",
  50661=>"001110111",
  50662=>"000100110",
  50663=>"000000001",
  50664=>"000100000",
  50665=>"001100011",
  50666=>"110100111",
  50667=>"110101110",
  50668=>"000111001",
  50669=>"101011111",
  50670=>"000000110",
  50671=>"010011100",
  50672=>"010100001",
  50673=>"100111010",
  50674=>"000111000",
  50675=>"111110100",
  50676=>"010011110",
  50677=>"000101100",
  50678=>"100000101",
  50679=>"000000100",
  50680=>"101110110",
  50681=>"000101000",
  50682=>"101000011",
  50683=>"110100000",
  50684=>"111000100",
  50685=>"001000101",
  50686=>"001010111",
  50687=>"011001101",
  50688=>"011000010",
  50689=>"110000101",
  50690=>"110000000",
  50691=>"001001110",
  50692=>"001110111",
  50693=>"011101001",
  50694=>"111111110",
  50695=>"000010000",
  50696=>"100001000",
  50697=>"000011110",
  50698=>"001000000",
  50699=>"010101111",
  50700=>"000101100",
  50701=>"110011011",
  50702=>"100000101",
  50703=>"100000101",
  50704=>"001100100",
  50705=>"100010001",
  50706=>"100010001",
  50707=>"011100110",
  50708=>"100000000",
  50709=>"010001010",
  50710=>"001111100",
  50711=>"110011011",
  50712=>"010000101",
  50713=>"000111001",
  50714=>"100001100",
  50715=>"010010111",
  50716=>"111010001",
  50717=>"101100100",
  50718=>"100001011",
  50719=>"000111101",
  50720=>"111010001",
  50721=>"000010011",
  50722=>"000110010",
  50723=>"000110101",
  50724=>"001101010",
  50725=>"000000101",
  50726=>"101001111",
  50727=>"000010100",
  50728=>"100010000",
  50729=>"111111011",
  50730=>"111001010",
  50731=>"011100100",
  50732=>"110001110",
  50733=>"010011100",
  50734=>"101010100",
  50735=>"001001011",
  50736=>"010101101",
  50737=>"111000111",
  50738=>"010010111",
  50739=>"100111001",
  50740=>"000101100",
  50741=>"101101111",
  50742=>"000111010",
  50743=>"111101011",
  50744=>"100000011",
  50745=>"100001100",
  50746=>"101000110",
  50747=>"110111101",
  50748=>"100101110",
  50749=>"100010100",
  50750=>"010110101",
  50751=>"100000100",
  50752=>"011000110",
  50753=>"110010001",
  50754=>"000010000",
  50755=>"111001011",
  50756=>"010011000",
  50757=>"011001011",
  50758=>"000000000",
  50759=>"101101111",
  50760=>"111100001",
  50761=>"100010000",
  50762=>"111110110",
  50763=>"001111111",
  50764=>"101011101",
  50765=>"110000001",
  50766=>"010101111",
  50767=>"000101010",
  50768=>"000000010",
  50769=>"010010000",
  50770=>"010111001",
  50771=>"111001000",
  50772=>"001100001",
  50773=>"000000000",
  50774=>"000000100",
  50775=>"110101011",
  50776=>"000000010",
  50777=>"110101001",
  50778=>"101011001",
  50779=>"011010000",
  50780=>"000110110",
  50781=>"101001000",
  50782=>"000000001",
  50783=>"011010100",
  50784=>"001000110",
  50785=>"001111001",
  50786=>"000010011",
  50787=>"011001000",
  50788=>"101011001",
  50789=>"111110000",
  50790=>"000101111",
  50791=>"111011110",
  50792=>"010110110",
  50793=>"000000000",
  50794=>"100110001",
  50795=>"010000000",
  50796=>"100100111",
  50797=>"001101111",
  50798=>"011101010",
  50799=>"111011000",
  50800=>"000011100",
  50801=>"101111101",
  50802=>"101110010",
  50803=>"001011111",
  50804=>"011010011",
  50805=>"001100001",
  50806=>"011100011",
  50807=>"001100110",
  50808=>"100000011",
  50809=>"000010010",
  50810=>"010101110",
  50811=>"001000110",
  50812=>"010100000",
  50813=>"001111001",
  50814=>"111100100",
  50815=>"100000000",
  50816=>"101010001",
  50817=>"111111101",
  50818=>"000111001",
  50819=>"001000000",
  50820=>"000101000",
  50821=>"010001100",
  50822=>"100111100",
  50823=>"100100010",
  50824=>"000011110",
  50825=>"001101011",
  50826=>"111101101",
  50827=>"101000001",
  50828=>"111111000",
  50829=>"000001000",
  50830=>"110001000",
  50831=>"000110101",
  50832=>"101100110",
  50833=>"101110000",
  50834=>"101110010",
  50835=>"010011100",
  50836=>"101110010",
  50837=>"011110101",
  50838=>"111100101",
  50839=>"010011101",
  50840=>"100111010",
  50841=>"001010000",
  50842=>"000110111",
  50843=>"000110111",
  50844=>"111000101",
  50845=>"011101111",
  50846=>"111111111",
  50847=>"000010110",
  50848=>"111010100",
  50849=>"001100101",
  50850=>"110000000",
  50851=>"000111001",
  50852=>"100010100",
  50853=>"110100111",
  50854=>"111001011",
  50855=>"101100101",
  50856=>"111001010",
  50857=>"000000101",
  50858=>"100000000",
  50859=>"011110110",
  50860=>"001010000",
  50861=>"111000001",
  50862=>"110011010",
  50863=>"100000001",
  50864=>"101010010",
  50865=>"001000011",
  50866=>"010000110",
  50867=>"110110000",
  50868=>"001010001",
  50869=>"000010101",
  50870=>"000001011",
  50871=>"011001001",
  50872=>"101010111",
  50873=>"111111011",
  50874=>"011101101",
  50875=>"110001111",
  50876=>"001000101",
  50877=>"011110111",
  50878=>"000011100",
  50879=>"000001100",
  50880=>"011010111",
  50881=>"000111110",
  50882=>"100001011",
  50883=>"110111111",
  50884=>"011011101",
  50885=>"000000000",
  50886=>"111101100",
  50887=>"100111000",
  50888=>"011110000",
  50889=>"111101101",
  50890=>"001110010",
  50891=>"000000000",
  50892=>"111000101",
  50893=>"001011011",
  50894=>"000000111",
  50895=>"001010011",
  50896=>"010110100",
  50897=>"001010001",
  50898=>"101101110",
  50899=>"010111011",
  50900=>"111101101",
  50901=>"101001000",
  50902=>"111010010",
  50903=>"000111011",
  50904=>"001001010",
  50905=>"000000010",
  50906=>"000100101",
  50907=>"111001001",
  50908=>"101001111",
  50909=>"110110101",
  50910=>"001010110",
  50911=>"001000001",
  50912=>"010111001",
  50913=>"111011110",
  50914=>"000111101",
  50915=>"010110111",
  50916=>"110101100",
  50917=>"001001000",
  50918=>"010111101",
  50919=>"100101100",
  50920=>"000001010",
  50921=>"100000101",
  50922=>"100001111",
  50923=>"010000000",
  50924=>"100001010",
  50925=>"000000111",
  50926=>"110100100",
  50927=>"001100101",
  50928=>"111111101",
  50929=>"010011101",
  50930=>"011010000",
  50931=>"001100010",
  50932=>"010110001",
  50933=>"101110110",
  50934=>"111110110",
  50935=>"100101001",
  50936=>"011010100",
  50937=>"111100000",
  50938=>"110010001",
  50939=>"001000010",
  50940=>"110110110",
  50941=>"100000001",
  50942=>"110011000",
  50943=>"010011101",
  50944=>"101101001",
  50945=>"110001111",
  50946=>"000000011",
  50947=>"000010111",
  50948=>"000110101",
  50949=>"000011010",
  50950=>"101010010",
  50951=>"110100000",
  50952=>"101010011",
  50953=>"001011010",
  50954=>"101110010",
  50955=>"100110111",
  50956=>"001001101",
  50957=>"110100110",
  50958=>"011101101",
  50959=>"000001000",
  50960=>"000001100",
  50961=>"001000011",
  50962=>"010100001",
  50963=>"100100000",
  50964=>"111001100",
  50965=>"010011000",
  50966=>"111000000",
  50967=>"000100110",
  50968=>"111101101",
  50969=>"100011101",
  50970=>"000101011",
  50971=>"011110100",
  50972=>"101101001",
  50973=>"110101111",
  50974=>"111100001",
  50975=>"110010110",
  50976=>"010010001",
  50977=>"000100111",
  50978=>"011111011",
  50979=>"000100011",
  50980=>"010001011",
  50981=>"111010001",
  50982=>"011101010",
  50983=>"001011011",
  50984=>"101000100",
  50985=>"111110000",
  50986=>"010011001",
  50987=>"100100010",
  50988=>"101101110",
  50989=>"001101011",
  50990=>"101000100",
  50991=>"011000000",
  50992=>"110000010",
  50993=>"111010101",
  50994=>"110001101",
  50995=>"111011001",
  50996=>"001110100",
  50997=>"001011001",
  50998=>"010010101",
  50999=>"101100001",
  51000=>"100000100",
  51001=>"000100010",
  51002=>"010100101",
  51003=>"101111110",
  51004=>"111110011",
  51005=>"001000101",
  51006=>"111010010",
  51007=>"000001001",
  51008=>"101101011",
  51009=>"010000011",
  51010=>"000001111",
  51011=>"101101111",
  51012=>"011111000",
  51013=>"000100011",
  51014=>"110101111",
  51015=>"101101101",
  51016=>"001001100",
  51017=>"110101101",
  51018=>"111011011",
  51019=>"000010001",
  51020=>"010011100",
  51021=>"100011011",
  51022=>"000101010",
  51023=>"010010000",
  51024=>"101110011",
  51025=>"001101000",
  51026=>"101011101",
  51027=>"111011111",
  51028=>"011111011",
  51029=>"110010000",
  51030=>"100000010",
  51031=>"010110011",
  51032=>"110010010",
  51033=>"100111100",
  51034=>"100000010",
  51035=>"011001101",
  51036=>"011011011",
  51037=>"000111010",
  51038=>"100110101",
  51039=>"101001100",
  51040=>"110101001",
  51041=>"011001011",
  51042=>"011010111",
  51043=>"011001110",
  51044=>"000111011",
  51045=>"001000101",
  51046=>"000110010",
  51047=>"011000101",
  51048=>"011111010",
  51049=>"010111110",
  51050=>"000001001",
  51051=>"101111111",
  51052=>"000100000",
  51053=>"111000001",
  51054=>"011010000",
  51055=>"110001000",
  51056=>"100110100",
  51057=>"111101100",
  51058=>"011000100",
  51059=>"010010100",
  51060=>"100010100",
  51061=>"101011111",
  51062=>"100010001",
  51063=>"101110000",
  51064=>"101110010",
  51065=>"100001111",
  51066=>"111011011",
  51067=>"111000011",
  51068=>"001111100",
  51069=>"011101111",
  51070=>"000010101",
  51071=>"100110000",
  51072=>"001110001",
  51073=>"111001101",
  51074=>"000101110",
  51075=>"000001111",
  51076=>"000110100",
  51077=>"000001011",
  51078=>"000011100",
  51079=>"001010100",
  51080=>"110000110",
  51081=>"001100010",
  51082=>"100001011",
  51083=>"000010010",
  51084=>"101010000",
  51085=>"111111111",
  51086=>"011010011",
  51087=>"011100111",
  51088=>"111000001",
  51089=>"010110101",
  51090=>"001100100",
  51091=>"000100101",
  51092=>"001011111",
  51093=>"110111111",
  51094=>"010111010",
  51095=>"000011010",
  51096=>"100001111",
  51097=>"000001100",
  51098=>"001000111",
  51099=>"011111110",
  51100=>"011101101",
  51101=>"010101110",
  51102=>"110110010",
  51103=>"001100010",
  51104=>"111111101",
  51105=>"101101010",
  51106=>"101011100",
  51107=>"010111111",
  51108=>"010001001",
  51109=>"101101000",
  51110=>"110111011",
  51111=>"100111000",
  51112=>"100010000",
  51113=>"001110100",
  51114=>"110111101",
  51115=>"101111110",
  51116=>"001010001",
  51117=>"000001010",
  51118=>"011110101",
  51119=>"101011010",
  51120=>"001110010",
  51121=>"101010001",
  51122=>"010010011",
  51123=>"111110111",
  51124=>"111111010",
  51125=>"010000001",
  51126=>"101110011",
  51127=>"101100011",
  51128=>"101111001",
  51129=>"111100010",
  51130=>"000001111",
  51131=>"010101101",
  51132=>"010011011",
  51133=>"001000100",
  51134=>"110111110",
  51135=>"101000010",
  51136=>"000010001",
  51137=>"000110001",
  51138=>"110000010",
  51139=>"110011111",
  51140=>"110110100",
  51141=>"010010111",
  51142=>"101010111",
  51143=>"001001110",
  51144=>"001010111",
  51145=>"100010100",
  51146=>"000001100",
  51147=>"101000100",
  51148=>"101011101",
  51149=>"000000110",
  51150=>"001100000",
  51151=>"111111101",
  51152=>"000010001",
  51153=>"010000010",
  51154=>"001110011",
  51155=>"111101110",
  51156=>"011010001",
  51157=>"110110100",
  51158=>"101010001",
  51159=>"100011101",
  51160=>"100011010",
  51161=>"001011000",
  51162=>"101101100",
  51163=>"010111111",
  51164=>"111001010",
  51165=>"011110000",
  51166=>"111001101",
  51167=>"100010100",
  51168=>"111011111",
  51169=>"000010001",
  51170=>"000111001",
  51171=>"000111011",
  51172=>"011101011",
  51173=>"111010111",
  51174=>"110001111",
  51175=>"000111100",
  51176=>"111000000",
  51177=>"110001110",
  51178=>"001100100",
  51179=>"111001010",
  51180=>"111001001",
  51181=>"011011101",
  51182=>"010111001",
  51183=>"100011001",
  51184=>"100101010",
  51185=>"010100110",
  51186=>"010011000",
  51187=>"001010111",
  51188=>"010011111",
  51189=>"010100100",
  51190=>"110111000",
  51191=>"101011001",
  51192=>"000000101",
  51193=>"000010110",
  51194=>"000011000",
  51195=>"001010001",
  51196=>"111010001",
  51197=>"100101110",
  51198=>"111100001",
  51199=>"011011000",
  51200=>"110100111",
  51201=>"110000100",
  51202=>"110110111",
  51203=>"000001010",
  51204=>"011110111",
  51205=>"111110011",
  51206=>"001010110",
  51207=>"111100000",
  51208=>"101001110",
  51209=>"001010111",
  51210=>"000000010",
  51211=>"001010100",
  51212=>"010100001",
  51213=>"011000110",
  51214=>"000100000",
  51215=>"000000100",
  51216=>"110000001",
  51217=>"000010000",
  51218=>"110100110",
  51219=>"001000110",
  51220=>"110011001",
  51221=>"000111011",
  51222=>"111010010",
  51223=>"111100001",
  51224=>"111000010",
  51225=>"001000000",
  51226=>"011010101",
  51227=>"000111100",
  51228=>"011000100",
  51229=>"010010011",
  51230=>"111010001",
  51231=>"000000110",
  51232=>"011010100",
  51233=>"001110100",
  51234=>"111100001",
  51235=>"001000011",
  51236=>"111100010",
  51237=>"010011000",
  51238=>"101100011",
  51239=>"011111100",
  51240=>"010010100",
  51241=>"101100110",
  51242=>"110110011",
  51243=>"111011101",
  51244=>"100011010",
  51245=>"011101101",
  51246=>"000110100",
  51247=>"010111001",
  51248=>"001010101",
  51249=>"001100000",
  51250=>"110000111",
  51251=>"111000100",
  51252=>"111011000",
  51253=>"010000010",
  51254=>"110100000",
  51255=>"010110101",
  51256=>"000000111",
  51257=>"011000111",
  51258=>"100111011",
  51259=>"111011111",
  51260=>"101110101",
  51261=>"010001001",
  51262=>"010110000",
  51263=>"010111010",
  51264=>"010100000",
  51265=>"101000010",
  51266=>"110011000",
  51267=>"110011101",
  51268=>"111100100",
  51269=>"111101100",
  51270=>"101001010",
  51271=>"000111110",
  51272=>"100010001",
  51273=>"100010010",
  51274=>"101001100",
  51275=>"110110110",
  51276=>"000111101",
  51277=>"010110111",
  51278=>"001010000",
  51279=>"000100010",
  51280=>"110110111",
  51281=>"000110010",
  51282=>"101111100",
  51283=>"011001011",
  51284=>"110011101",
  51285=>"010100000",
  51286=>"101100101",
  51287=>"000100001",
  51288=>"110110100",
  51289=>"000111110",
  51290=>"100011111",
  51291=>"100111101",
  51292=>"110111010",
  51293=>"011000010",
  51294=>"011011011",
  51295=>"000101110",
  51296=>"011110110",
  51297=>"001011010",
  51298=>"000101010",
  51299=>"011101001",
  51300=>"011000001",
  51301=>"001101000",
  51302=>"000111110",
  51303=>"000110110",
  51304=>"111011000",
  51305=>"010011101",
  51306=>"000111011",
  51307=>"110010111",
  51308=>"111100000",
  51309=>"111000010",
  51310=>"000110011",
  51311=>"111101111",
  51312=>"010101010",
  51313=>"000010011",
  51314=>"011001001",
  51315=>"111101110",
  51316=>"001110101",
  51317=>"100111001",
  51318=>"011001100",
  51319=>"110100110",
  51320=>"110001100",
  51321=>"001000000",
  51322=>"100001010",
  51323=>"000001110",
  51324=>"000111111",
  51325=>"010011001",
  51326=>"111100111",
  51327=>"101111000",
  51328=>"100100111",
  51329=>"100110011",
  51330=>"111000111",
  51331=>"011000010",
  51332=>"010000100",
  51333=>"101010010",
  51334=>"000101100",
  51335=>"110110011",
  51336=>"111101111",
  51337=>"111000000",
  51338=>"100011001",
  51339=>"011010101",
  51340=>"010010010",
  51341=>"110111011",
  51342=>"001111011",
  51343=>"000110011",
  51344=>"000101111",
  51345=>"100101010",
  51346=>"101010000",
  51347=>"110000011",
  51348=>"101001000",
  51349=>"010001011",
  51350=>"001110100",
  51351=>"011100110",
  51352=>"000000100",
  51353=>"010000110",
  51354=>"111010111",
  51355=>"000010010",
  51356=>"111011011",
  51357=>"111010100",
  51358=>"001100000",
  51359=>"001110101",
  51360=>"101100001",
  51361=>"110111010",
  51362=>"111101111",
  51363=>"101100110",
  51364=>"100111001",
  51365=>"111100100",
  51366=>"000000101",
  51367=>"110010001",
  51368=>"000001111",
  51369=>"010101100",
  51370=>"000101100",
  51371=>"000011011",
  51372=>"011010010",
  51373=>"101111000",
  51374=>"100011100",
  51375=>"110010000",
  51376=>"101100101",
  51377=>"000101110",
  51378=>"000011101",
  51379=>"111100100",
  51380=>"110000110",
  51381=>"011000101",
  51382=>"010011111",
  51383=>"100011000",
  51384=>"011010000",
  51385=>"000010011",
  51386=>"010110000",
  51387=>"101011110",
  51388=>"010001001",
  51389=>"001000000",
  51390=>"010100111",
  51391=>"100010000",
  51392=>"001011110",
  51393=>"000001100",
  51394=>"111100100",
  51395=>"010000101",
  51396=>"110000111",
  51397=>"011010001",
  51398=>"000010000",
  51399=>"100010100",
  51400=>"111101001",
  51401=>"110111001",
  51402=>"011010101",
  51403=>"010010000",
  51404=>"111110101",
  51405=>"111110100",
  51406=>"111110111",
  51407=>"100010111",
  51408=>"111100110",
  51409=>"101001110",
  51410=>"100100100",
  51411=>"001110101",
  51412=>"110010111",
  51413=>"001100011",
  51414=>"010110110",
  51415=>"101001100",
  51416=>"010100000",
  51417=>"111110110",
  51418=>"001000110",
  51419=>"011101111",
  51420=>"010111001",
  51421=>"110111101",
  51422=>"101000101",
  51423=>"000000001",
  51424=>"011101011",
  51425=>"101100101",
  51426=>"100010011",
  51427=>"100001100",
  51428=>"110001101",
  51429=>"010101110",
  51430=>"011100010",
  51431=>"011000101",
  51432=>"001010100",
  51433=>"001000000",
  51434=>"001111100",
  51435=>"111100000",
  51436=>"001111011",
  51437=>"100101100",
  51438=>"000001011",
  51439=>"000100000",
  51440=>"000000101",
  51441=>"000010001",
  51442=>"001101011",
  51443=>"101110100",
  51444=>"111011010",
  51445=>"000000100",
  51446=>"100001101",
  51447=>"011011000",
  51448=>"100010000",
  51449=>"111000110",
  51450=>"110010001",
  51451=>"100111011",
  51452=>"001011001",
  51453=>"101110101",
  51454=>"010001000",
  51455=>"001010101",
  51456=>"010010110",
  51457=>"100101100",
  51458=>"010001000",
  51459=>"001010010",
  51460=>"111010101",
  51461=>"000000110",
  51462=>"110101000",
  51463=>"010001111",
  51464=>"000111101",
  51465=>"101001001",
  51466=>"000011111",
  51467=>"011011001",
  51468=>"001000101",
  51469=>"111010001",
  51470=>"000110011",
  51471=>"000111101",
  51472=>"100010000",
  51473=>"010111010",
  51474=>"010001110",
  51475=>"111111101",
  51476=>"101110010",
  51477=>"111011011",
  51478=>"011000110",
  51479=>"100100100",
  51480=>"100010101",
  51481=>"001000011",
  51482=>"111110111",
  51483=>"001010110",
  51484=>"010000000",
  51485=>"111001001",
  51486=>"000100100",
  51487=>"100111110",
  51488=>"111100000",
  51489=>"000110100",
  51490=>"100010011",
  51491=>"101010101",
  51492=>"011011101",
  51493=>"100100101",
  51494=>"100001001",
  51495=>"001011100",
  51496=>"111010100",
  51497=>"011010001",
  51498=>"000110100",
  51499=>"000100011",
  51500=>"000110101",
  51501=>"100011111",
  51502=>"001001111",
  51503=>"011101100",
  51504=>"111111100",
  51505=>"101110010",
  51506=>"001101100",
  51507=>"000110110",
  51508=>"011100011",
  51509=>"110111111",
  51510=>"000001010",
  51511=>"100001101",
  51512=>"101100011",
  51513=>"011011000",
  51514=>"100110101",
  51515=>"111010110",
  51516=>"110001011",
  51517=>"110110100",
  51518=>"010000111",
  51519=>"000110011",
  51520=>"010100111",
  51521=>"101101101",
  51522=>"000110010",
  51523=>"000100110",
  51524=>"010100101",
  51525=>"100101111",
  51526=>"001001101",
  51527=>"001100110",
  51528=>"100101111",
  51529=>"110011110",
  51530=>"110010101",
  51531=>"100001100",
  51532=>"001111000",
  51533=>"000111001",
  51534=>"110111001",
  51535=>"100110110",
  51536=>"000100100",
  51537=>"101000010",
  51538=>"011011000",
  51539=>"101001000",
  51540=>"000110100",
  51541=>"011001110",
  51542=>"111111110",
  51543=>"100000111",
  51544=>"110010110",
  51545=>"011101000",
  51546=>"100110001",
  51547=>"010010010",
  51548=>"010101110",
  51549=>"001011011",
  51550=>"011011000",
  51551=>"100001011",
  51552=>"011001001",
  51553=>"110001011",
  51554=>"011010100",
  51555=>"001000111",
  51556=>"110011000",
  51557=>"011011100",
  51558=>"010111000",
  51559=>"010100010",
  51560=>"100001100",
  51561=>"011110000",
  51562=>"110000101",
  51563=>"101111000",
  51564=>"011000111",
  51565=>"011011101",
  51566=>"111010110",
  51567=>"101100001",
  51568=>"100100010",
  51569=>"101110000",
  51570=>"100010010",
  51571=>"101010100",
  51572=>"100000010",
  51573=>"100101111",
  51574=>"000001100",
  51575=>"110011001",
  51576=>"100111001",
  51577=>"110011101",
  51578=>"111111001",
  51579=>"011110111",
  51580=>"011110011",
  51581=>"001101001",
  51582=>"010111111",
  51583=>"100100011",
  51584=>"111111110",
  51585=>"011010010",
  51586=>"010111100",
  51587=>"111011101",
  51588=>"110010110",
  51589=>"101101110",
  51590=>"111100110",
  51591=>"010111010",
  51592=>"110100111",
  51593=>"010001110",
  51594=>"000000111",
  51595=>"001111100",
  51596=>"011100111",
  51597=>"111110100",
  51598=>"010100101",
  51599=>"100110110",
  51600=>"111011010",
  51601=>"000000101",
  51602=>"100110011",
  51603=>"001110100",
  51604=>"001110111",
  51605=>"000110010",
  51606=>"111001101",
  51607=>"101010001",
  51608=>"111110110",
  51609=>"110000111",
  51610=>"101000111",
  51611=>"001110100",
  51612=>"010011110",
  51613=>"011100100",
  51614=>"100000100",
  51615=>"000110110",
  51616=>"100100100",
  51617=>"101111000",
  51618=>"000010101",
  51619=>"000000101",
  51620=>"110000100",
  51621=>"100000011",
  51622=>"000000011",
  51623=>"000001001",
  51624=>"001111110",
  51625=>"001000111",
  51626=>"101110000",
  51627=>"111001001",
  51628=>"100101110",
  51629=>"001101101",
  51630=>"000011100",
  51631=>"111001000",
  51632=>"111111110",
  51633=>"110110111",
  51634=>"110110110",
  51635=>"010000000",
  51636=>"001001011",
  51637=>"001010001",
  51638=>"000101010",
  51639=>"111111101",
  51640=>"001001100",
  51641=>"001111110",
  51642=>"101011110",
  51643=>"101000011",
  51644=>"011111110",
  51645=>"000100010",
  51646=>"011110111",
  51647=>"111101010",
  51648=>"101000001",
  51649=>"000010011",
  51650=>"010000010",
  51651=>"101110111",
  51652=>"111000011",
  51653=>"000000111",
  51654=>"111001001",
  51655=>"000100101",
  51656=>"101101010",
  51657=>"101000111",
  51658=>"101101000",
  51659=>"000001100",
  51660=>"000001000",
  51661=>"000110111",
  51662=>"110100100",
  51663=>"011101100",
  51664=>"100111111",
  51665=>"001111111",
  51666=>"000000100",
  51667=>"101111111",
  51668=>"001010101",
  51669=>"000000110",
  51670=>"110010011",
  51671=>"100100111",
  51672=>"000110001",
  51673=>"111111000",
  51674=>"000010111",
  51675=>"010111000",
  51676=>"100111111",
  51677=>"011100110",
  51678=>"111111111",
  51679=>"110010000",
  51680=>"000000101",
  51681=>"000011111",
  51682=>"000010101",
  51683=>"010100101",
  51684=>"000100100",
  51685=>"101001101",
  51686=>"100101111",
  51687=>"011011011",
  51688=>"110101010",
  51689=>"011001010",
  51690=>"010011111",
  51691=>"100111010",
  51692=>"001010111",
  51693=>"100100001",
  51694=>"111110010",
  51695=>"000001000",
  51696=>"010110011",
  51697=>"011011010",
  51698=>"011111001",
  51699=>"001111110",
  51700=>"110001000",
  51701=>"111001000",
  51702=>"110010001",
  51703=>"100100110",
  51704=>"011111011",
  51705=>"110011100",
  51706=>"001001111",
  51707=>"100000101",
  51708=>"110000011",
  51709=>"101010110",
  51710=>"100100101",
  51711=>"101010111",
  51712=>"011110111",
  51713=>"011101110",
  51714=>"011111110",
  51715=>"010011110",
  51716=>"110101000",
  51717=>"010011111",
  51718=>"010111111",
  51719=>"110001000",
  51720=>"000001101",
  51721=>"111000110",
  51722=>"100101101",
  51723=>"011011001",
  51724=>"101000111",
  51725=>"000011001",
  51726=>"111110100",
  51727=>"011000000",
  51728=>"101010100",
  51729=>"010000000",
  51730=>"111110100",
  51731=>"111100100",
  51732=>"110100000",
  51733=>"101110010",
  51734=>"111111010",
  51735=>"110100011",
  51736=>"010000000",
  51737=>"110000100",
  51738=>"110111001",
  51739=>"010111101",
  51740=>"110101110",
  51741=>"000001100",
  51742=>"111011010",
  51743=>"010100110",
  51744=>"100100111",
  51745=>"100010100",
  51746=>"101100001",
  51747=>"000110100",
  51748=>"000011101",
  51749=>"111100101",
  51750=>"011111011",
  51751=>"000010100",
  51752=>"010110001",
  51753=>"001100100",
  51754=>"101001010",
  51755=>"101100010",
  51756=>"111011011",
  51757=>"001100011",
  51758=>"010101101",
  51759=>"001010001",
  51760=>"010001101",
  51761=>"110111101",
  51762=>"011000000",
  51763=>"011100001",
  51764=>"101100111",
  51765=>"110000000",
  51766=>"000100101",
  51767=>"110000000",
  51768=>"100011111",
  51769=>"110001100",
  51770=>"011011000",
  51771=>"010101110",
  51772=>"001010110",
  51773=>"000010010",
  51774=>"111100010",
  51775=>"101111101",
  51776=>"101111001",
  51777=>"000110010",
  51778=>"011000001",
  51779=>"001111001",
  51780=>"101100000",
  51781=>"001001010",
  51782=>"000000011",
  51783=>"010110110",
  51784=>"010011010",
  51785=>"011100110",
  51786=>"010010010",
  51787=>"101111010",
  51788=>"101001011",
  51789=>"011111101",
  51790=>"100100101",
  51791=>"001001001",
  51792=>"001000010",
  51793=>"111111010",
  51794=>"100101011",
  51795=>"000001100",
  51796=>"110101000",
  51797=>"000001011",
  51798=>"101100101",
  51799=>"100110110",
  51800=>"001001110",
  51801=>"001001010",
  51802=>"111000100",
  51803=>"111101011",
  51804=>"011001011",
  51805=>"101010001",
  51806=>"011001111",
  51807=>"000100010",
  51808=>"110010000",
  51809=>"001000110",
  51810=>"100000111",
  51811=>"110000100",
  51812=>"000010111",
  51813=>"000100110",
  51814=>"010110001",
  51815=>"011010101",
  51816=>"110111011",
  51817=>"000000101",
  51818=>"101010000",
  51819=>"100000110",
  51820=>"101100011",
  51821=>"000100010",
  51822=>"001101011",
  51823=>"100000101",
  51824=>"000101000",
  51825=>"000101001",
  51826=>"010011110",
  51827=>"010100001",
  51828=>"001110100",
  51829=>"010000110",
  51830=>"001011101",
  51831=>"101111000",
  51832=>"101111010",
  51833=>"111100101",
  51834=>"001111110",
  51835=>"110100100",
  51836=>"011001011",
  51837=>"000100100",
  51838=>"101111010",
  51839=>"100111111",
  51840=>"001000101",
  51841=>"100110111",
  51842=>"011011010",
  51843=>"011001111",
  51844=>"110000100",
  51845=>"011011100",
  51846=>"000101101",
  51847=>"001000011",
  51848=>"110010110",
  51849=>"000011001",
  51850=>"100111011",
  51851=>"101010101",
  51852=>"010011110",
  51853=>"111111010",
  51854=>"110111001",
  51855=>"000000001",
  51856=>"110010101",
  51857=>"111011100",
  51858=>"010110010",
  51859=>"100100001",
  51860=>"001010111",
  51861=>"110111111",
  51862=>"100011111",
  51863=>"100110000",
  51864=>"000011000",
  51865=>"111010111",
  51866=>"111111101",
  51867=>"001011011",
  51868=>"100000010",
  51869=>"011011110",
  51870=>"101000000",
  51871=>"000000000",
  51872=>"001000101",
  51873=>"001011000",
  51874=>"001001010",
  51875=>"110101111",
  51876=>"000101111",
  51877=>"001010101",
  51878=>"101100001",
  51879=>"101101110",
  51880=>"011111100",
  51881=>"001100001",
  51882=>"101101111",
  51883=>"001110111",
  51884=>"010111111",
  51885=>"111011101",
  51886=>"011000010",
  51887=>"101001100",
  51888=>"001100110",
  51889=>"000010000",
  51890=>"010001010",
  51891=>"110001110",
  51892=>"001010101",
  51893=>"000111110",
  51894=>"110111011",
  51895=>"001000011",
  51896=>"000111000",
  51897=>"101000000",
  51898=>"001111110",
  51899=>"110110010",
  51900=>"110110111",
  51901=>"010011110",
  51902=>"001100100",
  51903=>"000010111",
  51904=>"000000000",
  51905=>"100111100",
  51906=>"000001111",
  51907=>"110111011",
  51908=>"010010111",
  51909=>"101111100",
  51910=>"011000101",
  51911=>"001110101",
  51912=>"110101100",
  51913=>"000100110",
  51914=>"100111011",
  51915=>"101100011",
  51916=>"111000111",
  51917=>"100100010",
  51918=>"111111100",
  51919=>"101010001",
  51920=>"111000100",
  51921=>"111111100",
  51922=>"010000000",
  51923=>"101011011",
  51924=>"001000101",
  51925=>"110100010",
  51926=>"110011101",
  51927=>"000111010",
  51928=>"111111010",
  51929=>"111001011",
  51930=>"101110110",
  51931=>"000110011",
  51932=>"000010011",
  51933=>"011101000",
  51934=>"001001101",
  51935=>"101111111",
  51936=>"011111000",
  51937=>"101000010",
  51938=>"000101110",
  51939=>"011010110",
  51940=>"100001101",
  51941=>"011000000",
  51942=>"100010110",
  51943=>"011011011",
  51944=>"000011110",
  51945=>"001101000",
  51946=>"000001000",
  51947=>"000011000",
  51948=>"010001110",
  51949=>"010101011",
  51950=>"000111111",
  51951=>"101101011",
  51952=>"100000101",
  51953=>"000001000",
  51954=>"100010111",
  51955=>"010111001",
  51956=>"110110001",
  51957=>"000111100",
  51958=>"010101101",
  51959=>"101111101",
  51960=>"100011001",
  51961=>"111011001",
  51962=>"001010001",
  51963=>"011000000",
  51964=>"000001001",
  51965=>"000110110",
  51966=>"010110011",
  51967=>"011100100",
  51968=>"010010011",
  51969=>"110110101",
  51970=>"111110100",
  51971=>"101000100",
  51972=>"111001110",
  51973=>"111000000",
  51974=>"001110101",
  51975=>"011001011",
  51976=>"010100011",
  51977=>"011110001",
  51978=>"101011110",
  51979=>"111100000",
  51980=>"000111111",
  51981=>"111110111",
  51982=>"000000011",
  51983=>"101111111",
  51984=>"011111100",
  51985=>"111100100",
  51986=>"000101000",
  51987=>"011001000",
  51988=>"010110111",
  51989=>"101010100",
  51990=>"111101001",
  51991=>"001001101",
  51992=>"100101101",
  51993=>"110101111",
  51994=>"000101101",
  51995=>"101011000",
  51996=>"111100101",
  51997=>"111111000",
  51998=>"000010100",
  51999=>"011101001",
  52000=>"111111011",
  52001=>"011011110",
  52002=>"000000000",
  52003=>"110001111",
  52004=>"010001000",
  52005=>"000000011",
  52006=>"011100010",
  52007=>"111101101",
  52008=>"110010011",
  52009=>"000010001",
  52010=>"001000010",
  52011=>"100110001",
  52012=>"101010111",
  52013=>"010100001",
  52014=>"111111001",
  52015=>"111010011",
  52016=>"010000000",
  52017=>"111000100",
  52018=>"111111011",
  52019=>"011000001",
  52020=>"000110101",
  52021=>"010000110",
  52022=>"000011111",
  52023=>"010010100",
  52024=>"010010011",
  52025=>"111000101",
  52026=>"000000011",
  52027=>"111010110",
  52028=>"100101111",
  52029=>"110100011",
  52030=>"000111010",
  52031=>"000001011",
  52032=>"000010000",
  52033=>"111010011",
  52034=>"001100010",
  52035=>"110000100",
  52036=>"101110100",
  52037=>"111100000",
  52038=>"000100100",
  52039=>"010100000",
  52040=>"011010001",
  52041=>"010000000",
  52042=>"001011111",
  52043=>"000011011",
  52044=>"100011000",
  52045=>"110001001",
  52046=>"111110111",
  52047=>"101011100",
  52048=>"110111111",
  52049=>"000010011",
  52050=>"110001001",
  52051=>"111001110",
  52052=>"010000110",
  52053=>"100101001",
  52054=>"101001010",
  52055=>"101011011",
  52056=>"001110110",
  52057=>"010101110",
  52058=>"001000000",
  52059=>"110100000",
  52060=>"100101010",
  52061=>"000010000",
  52062=>"111101001",
  52063=>"110000100",
  52064=>"100001010",
  52065=>"000100111",
  52066=>"011100001",
  52067=>"010110111",
  52068=>"011101010",
  52069=>"011101000",
  52070=>"100100110",
  52071=>"011011001",
  52072=>"111010100",
  52073=>"010010101",
  52074=>"000010100",
  52075=>"101010110",
  52076=>"011010101",
  52077=>"110011101",
  52078=>"111111110",
  52079=>"110111001",
  52080=>"101101001",
  52081=>"101001000",
  52082=>"011011100",
  52083=>"111011100",
  52084=>"001001100",
  52085=>"010111100",
  52086=>"101010101",
  52087=>"110111111",
  52088=>"011011001",
  52089=>"000010110",
  52090=>"011000101",
  52091=>"101111011",
  52092=>"101100110",
  52093=>"001001111",
  52094=>"111100111",
  52095=>"001101110",
  52096=>"011001011",
  52097=>"101101000",
  52098=>"011000000",
  52099=>"101000101",
  52100=>"100011111",
  52101=>"110101110",
  52102=>"100001101",
  52103=>"011100000",
  52104=>"101111110",
  52105=>"111110000",
  52106=>"100001000",
  52107=>"101100111",
  52108=>"101100100",
  52109=>"101100011",
  52110=>"001010110",
  52111=>"010111111",
  52112=>"101000101",
  52113=>"001101111",
  52114=>"111011000",
  52115=>"001010100",
  52116=>"010011110",
  52117=>"101101010",
  52118=>"101101101",
  52119=>"101111011",
  52120=>"100000111",
  52121=>"000010011",
  52122=>"001000011",
  52123=>"101000100",
  52124=>"000111000",
  52125=>"001000010",
  52126=>"110110001",
  52127=>"001101101",
  52128=>"011001000",
  52129=>"010101111",
  52130=>"111001110",
  52131=>"100011000",
  52132=>"110010111",
  52133=>"011101101",
  52134=>"100100010",
  52135=>"110010110",
  52136=>"100111111",
  52137=>"001000110",
  52138=>"111111010",
  52139=>"100111111",
  52140=>"110001101",
  52141=>"101110110",
  52142=>"100110100",
  52143=>"110110011",
  52144=>"111100000",
  52145=>"001110001",
  52146=>"011101101",
  52147=>"000001011",
  52148=>"000010010",
  52149=>"011101100",
  52150=>"000111111",
  52151=>"010001000",
  52152=>"001100101",
  52153=>"010000111",
  52154=>"011011101",
  52155=>"000111110",
  52156=>"011010000",
  52157=>"011000100",
  52158=>"010101101",
  52159=>"100100101",
  52160=>"011110010",
  52161=>"001000101",
  52162=>"011101111",
  52163=>"001110010",
  52164=>"110110001",
  52165=>"010100111",
  52166=>"100011100",
  52167=>"011101101",
  52168=>"011111011",
  52169=>"100001000",
  52170=>"001000011",
  52171=>"101110100",
  52172=>"001110000",
  52173=>"111000101",
  52174=>"001100111",
  52175=>"101100100",
  52176=>"100101011",
  52177=>"111111010",
  52178=>"001001111",
  52179=>"000000011",
  52180=>"111010100",
  52181=>"100110111",
  52182=>"011010010",
  52183=>"111111111",
  52184=>"111010000",
  52185=>"100001111",
  52186=>"111000100",
  52187=>"110011010",
  52188=>"101001011",
  52189=>"000000101",
  52190=>"001001010",
  52191=>"010011011",
  52192=>"000100001",
  52193=>"001001000",
  52194=>"111010100",
  52195=>"011101110",
  52196=>"011010110",
  52197=>"101111010",
  52198=>"100000100",
  52199=>"100010011",
  52200=>"011101100",
  52201=>"010011110",
  52202=>"010010101",
  52203=>"101100011",
  52204=>"100000110",
  52205=>"010110101",
  52206=>"001011110",
  52207=>"010110001",
  52208=>"011100100",
  52209=>"111111001",
  52210=>"010000011",
  52211=>"101111000",
  52212=>"100010110",
  52213=>"000000110",
  52214=>"100000000",
  52215=>"011101100",
  52216=>"000000111",
  52217=>"001010111",
  52218=>"011001111",
  52219=>"111010000",
  52220=>"101101011",
  52221=>"000100010",
  52222=>"100111101",
  52223=>"010101011",
  52224=>"000001011",
  52225=>"111001001",
  52226=>"010011000",
  52227=>"100100010",
  52228=>"100101000",
  52229=>"011001000",
  52230=>"110111110",
  52231=>"010000001",
  52232=>"001000011",
  52233=>"111011010",
  52234=>"011001111",
  52235=>"001010001",
  52236=>"010111111",
  52237=>"110101111",
  52238=>"001100111",
  52239=>"100001110",
  52240=>"001111110",
  52241=>"000001011",
  52242=>"010000010",
  52243=>"100001001",
  52244=>"000011101",
  52245=>"001110011",
  52246=>"010110101",
  52247=>"001000110",
  52248=>"000110111",
  52249=>"111010000",
  52250=>"110001010",
  52251=>"101110100",
  52252=>"011000110",
  52253=>"100000010",
  52254=>"111000011",
  52255=>"101111010",
  52256=>"011011010",
  52257=>"000011000",
  52258=>"011000100",
  52259=>"100100111",
  52260=>"011111100",
  52261=>"101110111",
  52262=>"110011111",
  52263=>"111100010",
  52264=>"011100110",
  52265=>"000001011",
  52266=>"101011000",
  52267=>"010111010",
  52268=>"001000001",
  52269=>"010101111",
  52270=>"111101011",
  52271=>"100101110",
  52272=>"001000101",
  52273=>"011111111",
  52274=>"011101010",
  52275=>"111101000",
  52276=>"110101010",
  52277=>"101111100",
  52278=>"110101101",
  52279=>"111011001",
  52280=>"011110011",
  52281=>"100011001",
  52282=>"101011000",
  52283=>"111111010",
  52284=>"000111111",
  52285=>"000010100",
  52286=>"110011010",
  52287=>"000001110",
  52288=>"110000100",
  52289=>"000111010",
  52290=>"100010000",
  52291=>"110111000",
  52292=>"010000000",
  52293=>"000010000",
  52294=>"100000101",
  52295=>"100001101",
  52296=>"100000010",
  52297=>"110101111",
  52298=>"101111110",
  52299=>"001011010",
  52300=>"111111000",
  52301=>"101101110",
  52302=>"010101000",
  52303=>"011011000",
  52304=>"101101000",
  52305=>"010001101",
  52306=>"111111110",
  52307=>"111100111",
  52308=>"111101111",
  52309=>"111100101",
  52310=>"011010100",
  52311=>"101011000",
  52312=>"101110001",
  52313=>"011000101",
  52314=>"110110100",
  52315=>"100111101",
  52316=>"000110000",
  52317=>"110110110",
  52318=>"011001100",
  52319=>"100001111",
  52320=>"111011001",
  52321=>"010101100",
  52322=>"011011011",
  52323=>"000100111",
  52324=>"100001111",
  52325=>"010111011",
  52326=>"111111110",
  52327=>"001111100",
  52328=>"110101010",
  52329=>"110001110",
  52330=>"001101001",
  52331=>"000100100",
  52332=>"101111011",
  52333=>"000111010",
  52334=>"010001011",
  52335=>"011000001",
  52336=>"101110001",
  52337=>"110100000",
  52338=>"111110101",
  52339=>"111101001",
  52340=>"001011101",
  52341=>"110001100",
  52342=>"011100101",
  52343=>"001110100",
  52344=>"011010001",
  52345=>"111000111",
  52346=>"001100111",
  52347=>"100111011",
  52348=>"101011101",
  52349=>"010101011",
  52350=>"111100100",
  52351=>"010000110",
  52352=>"000010010",
  52353=>"000111110",
  52354=>"111100011",
  52355=>"111100001",
  52356=>"000100011",
  52357=>"100010101",
  52358=>"000001011",
  52359=>"100111110",
  52360=>"101011001",
  52361=>"110001101",
  52362=>"110101011",
  52363=>"111101011",
  52364=>"111011001",
  52365=>"001101000",
  52366=>"001111100",
  52367=>"001101100",
  52368=>"110010110",
  52369=>"010010011",
  52370=>"100000101",
  52371=>"000011101",
  52372=>"010010110",
  52373=>"011011010",
  52374=>"111001011",
  52375=>"001000110",
  52376=>"110100001",
  52377=>"111100100",
  52378=>"010001101",
  52379=>"101101101",
  52380=>"111111010",
  52381=>"100110111",
  52382=>"010001011",
  52383=>"110111101",
  52384=>"000000010",
  52385=>"010101000",
  52386=>"110011110",
  52387=>"101000000",
  52388=>"010011110",
  52389=>"010111010",
  52390=>"101011000",
  52391=>"000110101",
  52392=>"101111101",
  52393=>"011100001",
  52394=>"001000101",
  52395=>"101111010",
  52396=>"001010001",
  52397=>"111111001",
  52398=>"111001101",
  52399=>"010111000",
  52400=>"110000101",
  52401=>"101110000",
  52402=>"000000101",
  52403=>"101011111",
  52404=>"110110000",
  52405=>"010000000",
  52406=>"101100101",
  52407=>"001111011",
  52408=>"100101110",
  52409=>"011111111",
  52410=>"110110011",
  52411=>"011111100",
  52412=>"100101011",
  52413=>"101011100",
  52414=>"110111011",
  52415=>"101111001",
  52416=>"001101111",
  52417=>"001101110",
  52418=>"111011110",
  52419=>"101111000",
  52420=>"111100010",
  52421=>"011101101",
  52422=>"001110101",
  52423=>"000000010",
  52424=>"011010010",
  52425=>"111101001",
  52426=>"011000011",
  52427=>"000111000",
  52428=>"100001111",
  52429=>"001110111",
  52430=>"110001110",
  52431=>"000111101",
  52432=>"111100111",
  52433=>"000100000",
  52434=>"010010000",
  52435=>"000000000",
  52436=>"011110011",
  52437=>"101000010",
  52438=>"111010101",
  52439=>"111110110",
  52440=>"010100001",
  52441=>"101110000",
  52442=>"110011101",
  52443=>"000000101",
  52444=>"000100000",
  52445=>"111100001",
  52446=>"100000110",
  52447=>"111010110",
  52448=>"100011101",
  52449=>"010010011",
  52450=>"101000101",
  52451=>"100011111",
  52452=>"010011010",
  52453=>"101100110",
  52454=>"100100011",
  52455=>"100101101",
  52456=>"110000100",
  52457=>"011010101",
  52458=>"100100111",
  52459=>"101101110",
  52460=>"100001010",
  52461=>"000000011",
  52462=>"100001011",
  52463=>"111110010",
  52464=>"110000000",
  52465=>"111100100",
  52466=>"010001000",
  52467=>"000100100",
  52468=>"010010000",
  52469=>"001111011",
  52470=>"101001100",
  52471=>"100000111",
  52472=>"110000000",
  52473=>"100000011",
  52474=>"000010000",
  52475=>"110010001",
  52476=>"101010101",
  52477=>"100100000",
  52478=>"110000010",
  52479=>"111011010",
  52480=>"001111000",
  52481=>"010110011",
  52482=>"111001100",
  52483=>"000010111",
  52484=>"010000101",
  52485=>"011100111",
  52486=>"111110110",
  52487=>"011011010",
  52488=>"111011000",
  52489=>"101010110",
  52490=>"110111111",
  52491=>"000011100",
  52492=>"001101101",
  52493=>"110010010",
  52494=>"011001000",
  52495=>"000011001",
  52496=>"111101111",
  52497=>"100001110",
  52498=>"010111000",
  52499=>"000101110",
  52500=>"101001000",
  52501=>"011000100",
  52502=>"001001100",
  52503=>"101010110",
  52504=>"101011111",
  52505=>"011110000",
  52506=>"001001000",
  52507=>"000011111",
  52508=>"110000010",
  52509=>"000101001",
  52510=>"011111001",
  52511=>"001101011",
  52512=>"111100001",
  52513=>"111111100",
  52514=>"110110001",
  52515=>"010110111",
  52516=>"111011000",
  52517=>"100111010",
  52518=>"011000100",
  52519=>"111110111",
  52520=>"111110001",
  52521=>"010100000",
  52522=>"110110001",
  52523=>"111111110",
  52524=>"101100000",
  52525=>"111001100",
  52526=>"001001111",
  52527=>"011111110",
  52528=>"111010001",
  52529=>"110011001",
  52530=>"011100000",
  52531=>"001011000",
  52532=>"000000010",
  52533=>"100100011",
  52534=>"101100100",
  52535=>"001110001",
  52536=>"101101101",
  52537=>"101001101",
  52538=>"110000110",
  52539=>"011101010",
  52540=>"000100111",
  52541=>"001100100",
  52542=>"000100100",
  52543=>"110111010",
  52544=>"100011101",
  52545=>"000100111",
  52546=>"011010000",
  52547=>"011100100",
  52548=>"001001110",
  52549=>"110110101",
  52550=>"110001101",
  52551=>"100010000",
  52552=>"010010101",
  52553=>"110010011",
  52554=>"111010001",
  52555=>"000101110",
  52556=>"011000011",
  52557=>"101010000",
  52558=>"101110101",
  52559=>"000100100",
  52560=>"111110000",
  52561=>"010001110",
  52562=>"101000101",
  52563=>"110111100",
  52564=>"111110111",
  52565=>"100011101",
  52566=>"011111110",
  52567=>"101011100",
  52568=>"001001101",
  52569=>"101101110",
  52570=>"011110110",
  52571=>"111110010",
  52572=>"000110111",
  52573=>"111110101",
  52574=>"000001011",
  52575=>"001101101",
  52576=>"100011101",
  52577=>"000100011",
  52578=>"011101010",
  52579=>"011101011",
  52580=>"101100100",
  52581=>"011101001",
  52582=>"101111111",
  52583=>"001101010",
  52584=>"101100100",
  52585=>"010101001",
  52586=>"111011011",
  52587=>"100011110",
  52588=>"101000100",
  52589=>"111100010",
  52590=>"011011111",
  52591=>"110011110",
  52592=>"000001000",
  52593=>"111100001",
  52594=>"001100101",
  52595=>"101101111",
  52596=>"110101010",
  52597=>"001001100",
  52598=>"001111111",
  52599=>"010100010",
  52600=>"000011110",
  52601=>"110000111",
  52602=>"011110010",
  52603=>"010010101",
  52604=>"101001001",
  52605=>"011000011",
  52606=>"010000000",
  52607=>"100001011",
  52608=>"100110000",
  52609=>"110110000",
  52610=>"111101010",
  52611=>"011111011",
  52612=>"010011000",
  52613=>"000010000",
  52614=>"111111111",
  52615=>"010010101",
  52616=>"000111000",
  52617=>"101100111",
  52618=>"101110011",
  52619=>"011010110",
  52620=>"001100010",
  52621=>"010110101",
  52622=>"101110100",
  52623=>"011100010",
  52624=>"010100111",
  52625=>"100101011",
  52626=>"111111100",
  52627=>"011110110",
  52628=>"101100110",
  52629=>"100011011",
  52630=>"000001110",
  52631=>"000101111",
  52632=>"110101110",
  52633=>"110011100",
  52634=>"011110000",
  52635=>"001010001",
  52636=>"001110000",
  52637=>"110110000",
  52638=>"100001100",
  52639=>"011011101",
  52640=>"010101010",
  52641=>"010101011",
  52642=>"111011100",
  52643=>"110101111",
  52644=>"111000001",
  52645=>"000000010",
  52646=>"110011001",
  52647=>"101101110",
  52648=>"000110011",
  52649=>"010011000",
  52650=>"001001110",
  52651=>"110111100",
  52652=>"010010001",
  52653=>"011100001",
  52654=>"001010111",
  52655=>"000011111",
  52656=>"110111101",
  52657=>"100001001",
  52658=>"000001111",
  52659=>"000001000",
  52660=>"010000011",
  52661=>"101011111",
  52662=>"000011011",
  52663=>"001000011",
  52664=>"111011001",
  52665=>"100010111",
  52666=>"101100001",
  52667=>"101111010",
  52668=>"111001000",
  52669=>"111110100",
  52670=>"111001101",
  52671=>"000111100",
  52672=>"011100101",
  52673=>"000101110",
  52674=>"111101111",
  52675=>"101100000",
  52676=>"011000001",
  52677=>"011100011",
  52678=>"011101010",
  52679=>"100010100",
  52680=>"010100111",
  52681=>"001100111",
  52682=>"000111001",
  52683=>"001101101",
  52684=>"010101011",
  52685=>"111001111",
  52686=>"111101000",
  52687=>"100000000",
  52688=>"010101001",
  52689=>"001001111",
  52690=>"110110111",
  52691=>"000101101",
  52692=>"111000100",
  52693=>"100110000",
  52694=>"100100111",
  52695=>"000010100",
  52696=>"101010111",
  52697=>"100010101",
  52698=>"010111000",
  52699=>"100001000",
  52700=>"100010011",
  52701=>"110011111",
  52702=>"011010000",
  52703=>"111011110",
  52704=>"100111111",
  52705=>"100111101",
  52706=>"101100001",
  52707=>"111011011",
  52708=>"011101110",
  52709=>"101011011",
  52710=>"010010110",
  52711=>"111000111",
  52712=>"001001111",
  52713=>"010100011",
  52714=>"000000000",
  52715=>"100001100",
  52716=>"111101001",
  52717=>"000111010",
  52718=>"010100010",
  52719=>"110110110",
  52720=>"010010111",
  52721=>"101111010",
  52722=>"011011110",
  52723=>"100011001",
  52724=>"111001000",
  52725=>"111111100",
  52726=>"111010010",
  52727=>"110111001",
  52728=>"100001011",
  52729=>"011001110",
  52730=>"011011110",
  52731=>"011001001",
  52732=>"011101101",
  52733=>"000010011",
  52734=>"000111010",
  52735=>"111100011",
  52736=>"101110111",
  52737=>"000011000",
  52738=>"110100110",
  52739=>"110000010",
  52740=>"010100001",
  52741=>"000101101",
  52742=>"011000001",
  52743=>"111111110",
  52744=>"011010101",
  52745=>"000001111",
  52746=>"010011111",
  52747=>"000111010",
  52748=>"100110110",
  52749=>"000010111",
  52750=>"010000000",
  52751=>"010001000",
  52752=>"010101000",
  52753=>"010100011",
  52754=>"100111010",
  52755=>"110001000",
  52756=>"101000101",
  52757=>"100101110",
  52758=>"110111110",
  52759=>"110110001",
  52760=>"101001110",
  52761=>"110111001",
  52762=>"010010010",
  52763=>"111001111",
  52764=>"111011011",
  52765=>"011101100",
  52766=>"110101100",
  52767=>"100111011",
  52768=>"101101101",
  52769=>"001100110",
  52770=>"000001011",
  52771=>"011111100",
  52772=>"010100111",
  52773=>"000001010",
  52774=>"111101101",
  52775=>"011111110",
  52776=>"010111000",
  52777=>"101101111",
  52778=>"100011001",
  52779=>"100000101",
  52780=>"101101101",
  52781=>"011010111",
  52782=>"010110011",
  52783=>"010000001",
  52784=>"111111110",
  52785=>"100010001",
  52786=>"111100111",
  52787=>"010011000",
  52788=>"100010001",
  52789=>"111001011",
  52790=>"110010001",
  52791=>"110100110",
  52792=>"100111001",
  52793=>"101010100",
  52794=>"100111000",
  52795=>"100100111",
  52796=>"001111100",
  52797=>"010010001",
  52798=>"011101111",
  52799=>"100111011",
  52800=>"001101111",
  52801=>"111100011",
  52802=>"101010101",
  52803=>"010001100",
  52804=>"110100000",
  52805=>"101010010",
  52806=>"010000000",
  52807=>"001011111",
  52808=>"110000010",
  52809=>"010001101",
  52810=>"011101101",
  52811=>"000010000",
  52812=>"000110110",
  52813=>"010000000",
  52814=>"010010000",
  52815=>"100011000",
  52816=>"100010000",
  52817=>"111101101",
  52818=>"111011100",
  52819=>"111010010",
  52820=>"101010110",
  52821=>"011110010",
  52822=>"110110111",
  52823=>"001010111",
  52824=>"010100010",
  52825=>"110111000",
  52826=>"101101001",
  52827=>"111010111",
  52828=>"101111110",
  52829=>"010100111",
  52830=>"110110011",
  52831=>"011101011",
  52832=>"110001101",
  52833=>"000100101",
  52834=>"001010110",
  52835=>"010010011",
  52836=>"001100000",
  52837=>"101010010",
  52838=>"101011010",
  52839=>"101000000",
  52840=>"001000000",
  52841=>"001010011",
  52842=>"101110100",
  52843=>"101010001",
  52844=>"011110100",
  52845=>"111100100",
  52846=>"100101010",
  52847=>"011000011",
  52848=>"100100011",
  52849=>"110110101",
  52850=>"100011111",
  52851=>"101110001",
  52852=>"011110101",
  52853=>"001100101",
  52854=>"101111110",
  52855=>"100001000",
  52856=>"000011011",
  52857=>"011101101",
  52858=>"011101000",
  52859=>"011100011",
  52860=>"110111110",
  52861=>"000000000",
  52862=>"001001001",
  52863=>"000001101",
  52864=>"110000111",
  52865=>"111010101",
  52866=>"101010110",
  52867=>"111010110",
  52868=>"101101100",
  52869=>"110010111",
  52870=>"101011110",
  52871=>"010000010",
  52872=>"000000101",
  52873=>"100101100",
  52874=>"111111111",
  52875=>"001000110",
  52876=>"111000100",
  52877=>"010101000",
  52878=>"010010101",
  52879=>"101110111",
  52880=>"110000010",
  52881=>"101001100",
  52882=>"111010011",
  52883=>"010110110",
  52884=>"000100000",
  52885=>"010010001",
  52886=>"001110111",
  52887=>"111001001",
  52888=>"110110101",
  52889=>"011111000",
  52890=>"101101000",
  52891=>"010001001",
  52892=>"001110101",
  52893=>"011001011",
  52894=>"000010010",
  52895=>"001000101",
  52896=>"010001100",
  52897=>"010010100",
  52898=>"111101100",
  52899=>"101100101",
  52900=>"111001011",
  52901=>"101100100",
  52902=>"011111011",
  52903=>"100001111",
  52904=>"001000110",
  52905=>"100010100",
  52906=>"011100110",
  52907=>"110001100",
  52908=>"101001000",
  52909=>"101100001",
  52910=>"000100000",
  52911=>"001101000",
  52912=>"010110101",
  52913=>"011100000",
  52914=>"100000000",
  52915=>"001010101",
  52916=>"110110110",
  52917=>"100111100",
  52918=>"001001101",
  52919=>"011011011",
  52920=>"001111001",
  52921=>"000100011",
  52922=>"100110011",
  52923=>"000010110",
  52924=>"110100111",
  52925=>"011110101",
  52926=>"110100010",
  52927=>"111111011",
  52928=>"100000001",
  52929=>"000101110",
  52930=>"001110001",
  52931=>"110001110",
  52932=>"110100111",
  52933=>"100001010",
  52934=>"001101111",
  52935=>"111111101",
  52936=>"011000111",
  52937=>"011101011",
  52938=>"110101110",
  52939=>"110101101",
  52940=>"110000111",
  52941=>"110011100",
  52942=>"101101111",
  52943=>"110001111",
  52944=>"100100100",
  52945=>"101000100",
  52946=>"011001010",
  52947=>"001100010",
  52948=>"111110110",
  52949=>"000010001",
  52950=>"100001101",
  52951=>"110100001",
  52952=>"100000110",
  52953=>"010110000",
  52954=>"101100001",
  52955=>"010001011",
  52956=>"010010011",
  52957=>"000101110",
  52958=>"010000111",
  52959=>"010111011",
  52960=>"101000101",
  52961=>"100100100",
  52962=>"011011110",
  52963=>"100011011",
  52964=>"110000110",
  52965=>"111010010",
  52966=>"111001111",
  52967=>"000010000",
  52968=>"111110010",
  52969=>"111111011",
  52970=>"001101101",
  52971=>"110011010",
  52972=>"100111100",
  52973=>"001011110",
  52974=>"101110100",
  52975=>"000100101",
  52976=>"010000001",
  52977=>"001011101",
  52978=>"011000000",
  52979=>"011001111",
  52980=>"100100010",
  52981=>"111110110",
  52982=>"101010110",
  52983=>"111111101",
  52984=>"111101000",
  52985=>"111111111",
  52986=>"111000110",
  52987=>"101000110",
  52988=>"101001100",
  52989=>"110010101",
  52990=>"011101010",
  52991=>"001001000",
  52992=>"110000010",
  52993=>"000000000",
  52994=>"010001100",
  52995=>"100000101",
  52996=>"010010011",
  52997=>"111111111",
  52998=>"010000111",
  52999=>"111100000",
  53000=>"011001100",
  53001=>"010011011",
  53002=>"110010000",
  53003=>"111100101",
  53004=>"101011010",
  53005=>"010111010",
  53006=>"010000110",
  53007=>"000100101",
  53008=>"010101111",
  53009=>"011010011",
  53010=>"111111010",
  53011=>"000010100",
  53012=>"100101000",
  53013=>"110110001",
  53014=>"100010110",
  53015=>"100001001",
  53016=>"010000101",
  53017=>"100101111",
  53018=>"100101000",
  53019=>"111111111",
  53020=>"000101000",
  53021=>"101111111",
  53022=>"110001110",
  53023=>"011010110",
  53024=>"010001001",
  53025=>"001000001",
  53026=>"001100011",
  53027=>"101110101",
  53028=>"001111100",
  53029=>"001011100",
  53030=>"101110001",
  53031=>"001000001",
  53032=>"100000101",
  53033=>"101100111",
  53034=>"100110101",
  53035=>"110110111",
  53036=>"001010010",
  53037=>"000000000",
  53038=>"001100101",
  53039=>"011101111",
  53040=>"110111100",
  53041=>"001001011",
  53042=>"001011110",
  53043=>"001110010",
  53044=>"001001011",
  53045=>"111100100",
  53046=>"011101011",
  53047=>"100001111",
  53048=>"111010100",
  53049=>"001010011",
  53050=>"000101001",
  53051=>"100110001",
  53052=>"111010001",
  53053=>"101001100",
  53054=>"011100111",
  53055=>"001011011",
  53056=>"011111010",
  53057=>"100111111",
  53058=>"001011011",
  53059=>"100001010",
  53060=>"000000100",
  53061=>"010100000",
  53062=>"010100010",
  53063=>"010111111",
  53064=>"011010111",
  53065=>"100101100",
  53066=>"001001011",
  53067=>"101001110",
  53068=>"110000101",
  53069=>"001000000",
  53070=>"110101000",
  53071=>"000111101",
  53072=>"010100110",
  53073=>"111011001",
  53074=>"010011000",
  53075=>"100100100",
  53076=>"011011010",
  53077=>"111110000",
  53078=>"100111111",
  53079=>"000100110",
  53080=>"000101011",
  53081=>"000111110",
  53082=>"001010100",
  53083=>"110101011",
  53084=>"111101111",
  53085=>"110001111",
  53086=>"100000100",
  53087=>"000000001",
  53088=>"000110010",
  53089=>"110000111",
  53090=>"000011100",
  53091=>"001011101",
  53092=>"111000001",
  53093=>"011010000",
  53094=>"010001001",
  53095=>"100101110",
  53096=>"100000000",
  53097=>"101000111",
  53098=>"110010000",
  53099=>"011111001",
  53100=>"110000110",
  53101=>"110001000",
  53102=>"111001001",
  53103=>"101000000",
  53104=>"110011100",
  53105=>"010110100",
  53106=>"101101111",
  53107=>"010111110",
  53108=>"100110010",
  53109=>"000100000",
  53110=>"011011000",
  53111=>"111000110",
  53112=>"111100001",
  53113=>"001010110",
  53114=>"011010000",
  53115=>"111111011",
  53116=>"110010111",
  53117=>"001111101",
  53118=>"011001000",
  53119=>"010101011",
  53120=>"010010010",
  53121=>"100011010",
  53122=>"100001100",
  53123=>"001110011",
  53124=>"011110111",
  53125=>"101101001",
  53126=>"111111110",
  53127=>"110000001",
  53128=>"111011111",
  53129=>"110111011",
  53130=>"011111101",
  53131=>"101011001",
  53132=>"100111100",
  53133=>"110010101",
  53134=>"101000011",
  53135=>"110110100",
  53136=>"101011000",
  53137=>"001111110",
  53138=>"111110100",
  53139=>"000101110",
  53140=>"001111111",
  53141=>"000110011",
  53142=>"000110011",
  53143=>"101001000",
  53144=>"001011101",
  53145=>"100000100",
  53146=>"000111110",
  53147=>"110111101",
  53148=>"011101011",
  53149=>"111111011",
  53150=>"100111010",
  53151=>"100010000",
  53152=>"011100101",
  53153=>"001010110",
  53154=>"010010000",
  53155=>"101010111",
  53156=>"101111101",
  53157=>"111100111",
  53158=>"111010011",
  53159=>"000000100",
  53160=>"110111110",
  53161=>"001111100",
  53162=>"101110101",
  53163=>"011011000",
  53164=>"011000011",
  53165=>"110101011",
  53166=>"110110000",
  53167=>"000001010",
  53168=>"011000001",
  53169=>"111111001",
  53170=>"111111100",
  53171=>"100110111",
  53172=>"001000101",
  53173=>"011101010",
  53174=>"011000101",
  53175=>"111011011",
  53176=>"110000010",
  53177=>"100001110",
  53178=>"100101011",
  53179=>"101110000",
  53180=>"000000100",
  53181=>"110100111",
  53182=>"001000011",
  53183=>"110111101",
  53184=>"010110111",
  53185=>"111101111",
  53186=>"111001000",
  53187=>"101000001",
  53188=>"011011001",
  53189=>"111101000",
  53190=>"000110000",
  53191=>"111101010",
  53192=>"100100101",
  53193=>"000010010",
  53194=>"101010111",
  53195=>"110011111",
  53196=>"011010000",
  53197=>"011110110",
  53198=>"111101101",
  53199=>"100000111",
  53200=>"010000001",
  53201=>"111110001",
  53202=>"100010110",
  53203=>"111111100",
  53204=>"010100100",
  53205=>"111101110",
  53206=>"100000010",
  53207=>"000011011",
  53208=>"000001110",
  53209=>"111000010",
  53210=>"100101001",
  53211=>"101110000",
  53212=>"000111010",
  53213=>"100000000",
  53214=>"001010110",
  53215=>"111001111",
  53216=>"111110110",
  53217=>"000101011",
  53218=>"000000010",
  53219=>"101111111",
  53220=>"000010000",
  53221=>"010000011",
  53222=>"110011100",
  53223=>"110001000",
  53224=>"001111111",
  53225=>"000111010",
  53226=>"110011110",
  53227=>"011001011",
  53228=>"100000101",
  53229=>"001101111",
  53230=>"100010100",
  53231=>"110110001",
  53232=>"011010010",
  53233=>"000101000",
  53234=>"101011010",
  53235=>"011000101",
  53236=>"100001100",
  53237=>"001011011",
  53238=>"111001001",
  53239=>"101000100",
  53240=>"000001011",
  53241=>"100110011",
  53242=>"111110101",
  53243=>"111001010",
  53244=>"010000100",
  53245=>"010110100",
  53246=>"110000110",
  53247=>"111011010",
  53248=>"111101010",
  53249=>"101101000",
  53250=>"111110110",
  53251=>"000100101",
  53252=>"101011011",
  53253=>"110101001",
  53254=>"111000010",
  53255=>"110001100",
  53256=>"111101111",
  53257=>"100011000",
  53258=>"011100000",
  53259=>"101111111",
  53260=>"001011001",
  53261=>"011000110",
  53262=>"111111101",
  53263=>"010000000",
  53264=>"110010010",
  53265=>"110011000",
  53266=>"111101111",
  53267=>"010101011",
  53268=>"000000001",
  53269=>"001100100",
  53270=>"100001100",
  53271=>"001011001",
  53272=>"110100111",
  53273=>"101001010",
  53274=>"010101000",
  53275=>"110111110",
  53276=>"000101111",
  53277=>"101100001",
  53278=>"001101111",
  53279=>"110011011",
  53280=>"110101000",
  53281=>"100010001",
  53282=>"101100100",
  53283=>"111100111",
  53284=>"101101100",
  53285=>"001100011",
  53286=>"111100111",
  53287=>"011100110",
  53288=>"011111111",
  53289=>"001111001",
  53290=>"001100101",
  53291=>"101010100",
  53292=>"001000010",
  53293=>"101101000",
  53294=>"110011010",
  53295=>"011011101",
  53296=>"000011000",
  53297=>"100010001",
  53298=>"111010101",
  53299=>"110010000",
  53300=>"100001001",
  53301=>"111000100",
  53302=>"100101111",
  53303=>"010010111",
  53304=>"000101110",
  53305=>"000101101",
  53306=>"101000110",
  53307=>"001001000",
  53308=>"111110100",
  53309=>"101011000",
  53310=>"111000101",
  53311=>"000101010",
  53312=>"010111000",
  53313=>"000011011",
  53314=>"001101111",
  53315=>"001100000",
  53316=>"011111000",
  53317=>"100000000",
  53318=>"001111111",
  53319=>"101000000",
  53320=>"000101001",
  53321=>"000100011",
  53322=>"000000001",
  53323=>"000000111",
  53324=>"010010010",
  53325=>"110000101",
  53326=>"111111001",
  53327=>"110001000",
  53328=>"010110010",
  53329=>"101000101",
  53330=>"010111110",
  53331=>"011001000",
  53332=>"100111000",
  53333=>"111111001",
  53334=>"010001010",
  53335=>"010100101",
  53336=>"110001110",
  53337=>"001111000",
  53338=>"101000001",
  53339=>"010001110",
  53340=>"011101000",
  53341=>"000000101",
  53342=>"001011010",
  53343=>"111110111",
  53344=>"001101010",
  53345=>"010011110",
  53346=>"010111011",
  53347=>"000011010",
  53348=>"011001100",
  53349=>"001011101",
  53350=>"011111010",
  53351=>"000010010",
  53352=>"101111111",
  53353=>"101000000",
  53354=>"110110111",
  53355=>"100011110",
  53356=>"100011010",
  53357=>"101000001",
  53358=>"101011101",
  53359=>"010111011",
  53360=>"110010100",
  53361=>"000110100",
  53362=>"000100010",
  53363=>"101110000",
  53364=>"110011011",
  53365=>"111100101",
  53366=>"100101011",
  53367=>"111000000",
  53368=>"000100111",
  53369=>"001100010",
  53370=>"101011001",
  53371=>"110011110",
  53372=>"001111101",
  53373=>"111101101",
  53374=>"001000000",
  53375=>"110110111",
  53376=>"010001101",
  53377=>"110101110",
  53378=>"001010001",
  53379=>"101101110",
  53380=>"110100010",
  53381=>"000000111",
  53382=>"000001110",
  53383=>"111100100",
  53384=>"110011001",
  53385=>"101100110",
  53386=>"001010001",
  53387=>"000001111",
  53388=>"011010100",
  53389=>"101100111",
  53390=>"010001000",
  53391=>"111101000",
  53392=>"010110001",
  53393=>"101111111",
  53394=>"110110000",
  53395=>"111100001",
  53396=>"111110000",
  53397=>"000110110",
  53398=>"001011011",
  53399=>"100111011",
  53400=>"010111111",
  53401=>"110010101",
  53402=>"011001011",
  53403=>"101000100",
  53404=>"000001111",
  53405=>"101000101",
  53406=>"111001110",
  53407=>"110010011",
  53408=>"010100101",
  53409=>"011100111",
  53410=>"110111001",
  53411=>"000101111",
  53412=>"000011100",
  53413=>"101010111",
  53414=>"111101101",
  53415=>"101000011",
  53416=>"010000000",
  53417=>"111010100",
  53418=>"100000001",
  53419=>"011110111",
  53420=>"011101111",
  53421=>"011101010",
  53422=>"111111111",
  53423=>"111111100",
  53424=>"001000101",
  53425=>"101110000",
  53426=>"011110101",
  53427=>"000011010",
  53428=>"111001010",
  53429=>"111010100",
  53430=>"100101110",
  53431=>"111000101",
  53432=>"011001110",
  53433=>"001000010",
  53434=>"010001011",
  53435=>"111011000",
  53436=>"001100010",
  53437=>"100100110",
  53438=>"110010000",
  53439=>"001001111",
  53440=>"100000001",
  53441=>"100111000",
  53442=>"011011111",
  53443=>"000001010",
  53444=>"000100110",
  53445=>"000011101",
  53446=>"000011000",
  53447=>"110010011",
  53448=>"100111010",
  53449=>"011001111",
  53450=>"101101101",
  53451=>"001000001",
  53452=>"101001111",
  53453=>"001011101",
  53454=>"111110100",
  53455=>"110101000",
  53456=>"001111111",
  53457=>"110101100",
  53458=>"101011110",
  53459=>"101101001",
  53460=>"111010000",
  53461=>"011001011",
  53462=>"110101101",
  53463=>"011101010",
  53464=>"111010000",
  53465=>"000111010",
  53466=>"001000001",
  53467=>"010100010",
  53468=>"111111010",
  53469=>"010100011",
  53470=>"101101111",
  53471=>"100100001",
  53472=>"000001010",
  53473=>"011010110",
  53474=>"100100111",
  53475=>"000011011",
  53476=>"110100100",
  53477=>"000100000",
  53478=>"000000010",
  53479=>"010101010",
  53480=>"001000100",
  53481=>"011110110",
  53482=>"000100100",
  53483=>"001111101",
  53484=>"110011110",
  53485=>"110010111",
  53486=>"101110111",
  53487=>"001100000",
  53488=>"000111001",
  53489=>"110000000",
  53490=>"000010111",
  53491=>"010100100",
  53492=>"110001110",
  53493=>"110001001",
  53494=>"100010001",
  53495=>"100111110",
  53496=>"001111111",
  53497=>"010111011",
  53498=>"110100101",
  53499=>"100110110",
  53500=>"000010001",
  53501=>"111110101",
  53502=>"111110111",
  53503=>"000101100",
  53504=>"111111110",
  53505=>"100000111",
  53506=>"100110001",
  53507=>"000000011",
  53508=>"100111001",
  53509=>"000000111",
  53510=>"100000101",
  53511=>"111111001",
  53512=>"001111111",
  53513=>"001001110",
  53514=>"001100111",
  53515=>"100001001",
  53516=>"010001100",
  53517=>"101100101",
  53518=>"111101111",
  53519=>"000000110",
  53520=>"001100100",
  53521=>"011000001",
  53522=>"000011100",
  53523=>"010111011",
  53524=>"000011101",
  53525=>"000000111",
  53526=>"011010000",
  53527=>"011000001",
  53528=>"101111011",
  53529=>"100101010",
  53530=>"000000000",
  53531=>"111110111",
  53532=>"011101011",
  53533=>"111000101",
  53534=>"010111111",
  53535=>"000011011",
  53536=>"001100011",
  53537=>"110010001",
  53538=>"000111101",
  53539=>"101110010",
  53540=>"111101110",
  53541=>"000000000",
  53542=>"111110100",
  53543=>"000101101",
  53544=>"010101100",
  53545=>"010001101",
  53546=>"011100110",
  53547=>"000000011",
  53548=>"010011000",
  53549=>"011110111",
  53550=>"101011111",
  53551=>"000010001",
  53552=>"001111000",
  53553=>"100010110",
  53554=>"010001100",
  53555=>"010011000",
  53556=>"110100101",
  53557=>"000000011",
  53558=>"001111001",
  53559=>"100011111",
  53560=>"000010001",
  53561=>"011101111",
  53562=>"011110100",
  53563=>"100110110",
  53564=>"001000101",
  53565=>"010000000",
  53566=>"100011000",
  53567=>"010000000",
  53568=>"110101011",
  53569=>"011001000",
  53570=>"011111001",
  53571=>"001000111",
  53572=>"111000110",
  53573=>"101110100",
  53574=>"011111111",
  53575=>"010000101",
  53576=>"100011010",
  53577=>"101100101",
  53578=>"001111011",
  53579=>"101001011",
  53580=>"001010010",
  53581=>"001111100",
  53582=>"010000001",
  53583=>"111010000",
  53584=>"100111010",
  53585=>"001100001",
  53586=>"010111111",
  53587=>"000111000",
  53588=>"100000111",
  53589=>"010010000",
  53590=>"111001000",
  53591=>"010010011",
  53592=>"111000101",
  53593=>"001011001",
  53594=>"100100011",
  53595=>"111101001",
  53596=>"101011010",
  53597=>"011010010",
  53598=>"010001001",
  53599=>"000111101",
  53600=>"000111010",
  53601=>"101000101",
  53602=>"111000100",
  53603=>"000000011",
  53604=>"001001000",
  53605=>"100101010",
  53606=>"100100100",
  53607=>"110000110",
  53608=>"001001110",
  53609=>"001111110",
  53610=>"101011011",
  53611=>"000011001",
  53612=>"010001100",
  53613=>"101100001",
  53614=>"000101000",
  53615=>"011001101",
  53616=>"000011100",
  53617=>"011100110",
  53618=>"111011001",
  53619=>"100110011",
  53620=>"111011001",
  53621=>"000101101",
  53622=>"000000011",
  53623=>"010000111",
  53624=>"010000001",
  53625=>"011110011",
  53626=>"010001011",
  53627=>"000000001",
  53628=>"000100001",
  53629=>"111011001",
  53630=>"000110111",
  53631=>"101000111",
  53632=>"100100001",
  53633=>"010110001",
  53634=>"001011101",
  53635=>"110010100",
  53636=>"100100101",
  53637=>"000010110",
  53638=>"110110101",
  53639=>"111111011",
  53640=>"111000001",
  53641=>"001000110",
  53642=>"110100000",
  53643=>"110101010",
  53644=>"011000110",
  53645=>"010111111",
  53646=>"010001001",
  53647=>"001111010",
  53648=>"010001111",
  53649=>"111001001",
  53650=>"001111101",
  53651=>"100100011",
  53652=>"100010101",
  53653=>"101000101",
  53654=>"101010010",
  53655=>"111010001",
  53656=>"011000011",
  53657=>"000001000",
  53658=>"000110011",
  53659=>"000010001",
  53660=>"111010010",
  53661=>"001000010",
  53662=>"101100001",
  53663=>"010000100",
  53664=>"110010000",
  53665=>"000010011",
  53666=>"011000010",
  53667=>"000000000",
  53668=>"111000110",
  53669=>"000000100",
  53670=>"101010100",
  53671=>"101001100",
  53672=>"000000100",
  53673=>"101001000",
  53674=>"000111011",
  53675=>"110110100",
  53676=>"011010010",
  53677=>"000100110",
  53678=>"100001010",
  53679=>"111111110",
  53680=>"000110000",
  53681=>"000101011",
  53682=>"101001100",
  53683=>"000101100",
  53684=>"111010110",
  53685=>"011011110",
  53686=>"001101110",
  53687=>"010000001",
  53688=>"001100100",
  53689=>"000111100",
  53690=>"000101000",
  53691=>"100010011",
  53692=>"101111101",
  53693=>"111101100",
  53694=>"110000100",
  53695=>"111001010",
  53696=>"111001111",
  53697=>"110101001",
  53698=>"111110101",
  53699=>"111100011",
  53700=>"010100100",
  53701=>"001011011",
  53702=>"010001101",
  53703=>"001000000",
  53704=>"001011010",
  53705=>"100101101",
  53706=>"000011100",
  53707=>"100000011",
  53708=>"000011100",
  53709=>"111100001",
  53710=>"101011110",
  53711=>"111000111",
  53712=>"110000010",
  53713=>"001010000",
  53714=>"000010110",
  53715=>"111110011",
  53716=>"010100010",
  53717=>"011011000",
  53718=>"111011100",
  53719=>"111000111",
  53720=>"000110010",
  53721=>"111100101",
  53722=>"010011110",
  53723=>"001110001",
  53724=>"111110010",
  53725=>"001101010",
  53726=>"001000000",
  53727=>"000000000",
  53728=>"011110010",
  53729=>"110100101",
  53730=>"110001111",
  53731=>"110111110",
  53732=>"100001010",
  53733=>"101101001",
  53734=>"100101101",
  53735=>"010000010",
  53736=>"110101001",
  53737=>"010011100",
  53738=>"010000111",
  53739=>"111111000",
  53740=>"000000111",
  53741=>"110100110",
  53742=>"101100001",
  53743=>"000011010",
  53744=>"001011001",
  53745=>"001101111",
  53746=>"111110101",
  53747=>"100010010",
  53748=>"100011101",
  53749=>"110000100",
  53750=>"110001010",
  53751=>"010101010",
  53752=>"111100001",
  53753=>"011001000",
  53754=>"110000101",
  53755=>"101011110",
  53756=>"000111101",
  53757=>"010101000",
  53758=>"001101100",
  53759=>"111111101",
  53760=>"101010001",
  53761=>"001011111",
  53762=>"001111101",
  53763=>"011111000",
  53764=>"101110101",
  53765=>"111101000",
  53766=>"110110101",
  53767=>"001100110",
  53768=>"110110101",
  53769=>"111100000",
  53770=>"010001001",
  53771=>"110111000",
  53772=>"111100001",
  53773=>"110001000",
  53774=>"111111000",
  53775=>"001100001",
  53776=>"100110101",
  53777=>"010010110",
  53778=>"001111010",
  53779=>"111111101",
  53780=>"111000000",
  53781=>"100111111",
  53782=>"101110001",
  53783=>"010111101",
  53784=>"001000100",
  53785=>"011100001",
  53786=>"001011001",
  53787=>"000101100",
  53788=>"010001000",
  53789=>"000011000",
  53790=>"111101101",
  53791=>"110100011",
  53792=>"111000001",
  53793=>"000001000",
  53794=>"000000000",
  53795=>"101001101",
  53796=>"110111101",
  53797=>"111111110",
  53798=>"001011010",
  53799=>"111101001",
  53800=>"111010101",
  53801=>"001001111",
  53802=>"001000011",
  53803=>"110000101",
  53804=>"000101111",
  53805=>"001001001",
  53806=>"101101101",
  53807=>"100000101",
  53808=>"000000111",
  53809=>"100111011",
  53810=>"100101011",
  53811=>"000000000",
  53812=>"101100111",
  53813=>"000111111",
  53814=>"000011101",
  53815=>"010011001",
  53816=>"001011111",
  53817=>"101101000",
  53818=>"101110001",
  53819=>"000001100",
  53820=>"000001111",
  53821=>"000001000",
  53822=>"101100010",
  53823=>"111100100",
  53824=>"000001001",
  53825=>"001100001",
  53826=>"101100111",
  53827=>"001111010",
  53828=>"101000100",
  53829=>"000110011",
  53830=>"010000001",
  53831=>"001011110",
  53832=>"010011010",
  53833=>"111111110",
  53834=>"010010100",
  53835=>"010101001",
  53836=>"110100100",
  53837=>"110100000",
  53838=>"110001000",
  53839=>"001011110",
  53840=>"111010100",
  53841=>"000010101",
  53842=>"110101101",
  53843=>"010010100",
  53844=>"011100010",
  53845=>"000011001",
  53846=>"000000010",
  53847=>"110101011",
  53848=>"011001000",
  53849=>"101101110",
  53850=>"100110000",
  53851=>"101100001",
  53852=>"110011101",
  53853=>"101011010",
  53854=>"001111011",
  53855=>"001101101",
  53856=>"101111001",
  53857=>"111011001",
  53858=>"101101101",
  53859=>"010000110",
  53860=>"000001011",
  53861=>"100100100",
  53862=>"011000010",
  53863=>"101111001",
  53864=>"000001101",
  53865=>"010010101",
  53866=>"110000100",
  53867=>"001100011",
  53868=>"101000110",
  53869=>"111000011",
  53870=>"100010111",
  53871=>"010111010",
  53872=>"000100101",
  53873=>"011010000",
  53874=>"110000111",
  53875=>"101011110",
  53876=>"000000010",
  53877=>"111111010",
  53878=>"010011110",
  53879=>"111100011",
  53880=>"110000111",
  53881=>"011100101",
  53882=>"101110101",
  53883=>"101100010",
  53884=>"101101011",
  53885=>"111111011",
  53886=>"101000111",
  53887=>"010100111",
  53888=>"001111111",
  53889=>"110110010",
  53890=>"111011010",
  53891=>"000100010",
  53892=>"001101100",
  53893=>"110100001",
  53894=>"000111101",
  53895=>"110011001",
  53896=>"000011101",
  53897=>"101110001",
  53898=>"000101001",
  53899=>"101011001",
  53900=>"010111110",
  53901=>"111110000",
  53902=>"111100001",
  53903=>"001001011",
  53904=>"110001000",
  53905=>"011010110",
  53906=>"100110000",
  53907=>"000101010",
  53908=>"100011101",
  53909=>"001001111",
  53910=>"011110101",
  53911=>"100001111",
  53912=>"000010100",
  53913=>"111101111",
  53914=>"101101100",
  53915=>"111111101",
  53916=>"101110000",
  53917=>"000101111",
  53918=>"011100010",
  53919=>"101101101",
  53920=>"111101001",
  53921=>"111110001",
  53922=>"100001010",
  53923=>"000110011",
  53924=>"111111001",
  53925=>"000001010",
  53926=>"111111111",
  53927=>"010010010",
  53928=>"100111110",
  53929=>"100010100",
  53930=>"001101011",
  53931=>"100100100",
  53932=>"001111100",
  53933=>"011001100",
  53934=>"110000100",
  53935=>"001011111",
  53936=>"100110011",
  53937=>"001000011",
  53938=>"111011101",
  53939=>"100011000",
  53940=>"110001010",
  53941=>"011001010",
  53942=>"010100110",
  53943=>"110000000",
  53944=>"100111110",
  53945=>"001101010",
  53946=>"111010110",
  53947=>"101001000",
  53948=>"101000000",
  53949=>"011011010",
  53950=>"010101101",
  53951=>"111110000",
  53952=>"111011000",
  53953=>"000010101",
  53954=>"001011011",
  53955=>"001110110",
  53956=>"010001010",
  53957=>"100000001",
  53958=>"111011000",
  53959=>"001100110",
  53960=>"101011101",
  53961=>"110111000",
  53962=>"001110001",
  53963=>"100001000",
  53964=>"011011001",
  53965=>"111100101",
  53966=>"110011111",
  53967=>"001100100",
  53968=>"101000001",
  53969=>"010111000",
  53970=>"110000111",
  53971=>"011010111",
  53972=>"110000000",
  53973=>"000011111",
  53974=>"001110001",
  53975=>"101011011",
  53976=>"001000101",
  53977=>"111110110",
  53978=>"010100000",
  53979=>"100110110",
  53980=>"100100001",
  53981=>"111110011",
  53982=>"000010010",
  53983=>"101100010",
  53984=>"000001001",
  53985=>"110000011",
  53986=>"010001000",
  53987=>"101110011",
  53988=>"000111100",
  53989=>"111000111",
  53990=>"110111110",
  53991=>"110010010",
  53992=>"001100000",
  53993=>"110101111",
  53994=>"010100100",
  53995=>"010100001",
  53996=>"000000011",
  53997=>"000010111",
  53998=>"111010011",
  53999=>"011010101",
  54000=>"111011101",
  54001=>"111000100",
  54002=>"011101100",
  54003=>"111110001",
  54004=>"110000011",
  54005=>"100111110",
  54006=>"001111110",
  54007=>"111110101",
  54008=>"010011000",
  54009=>"010101101",
  54010=>"100111101",
  54011=>"111011111",
  54012=>"100010010",
  54013=>"111001001",
  54014=>"010001001",
  54015=>"000100101",
  54016=>"011100110",
  54017=>"101110010",
  54018=>"111010101",
  54019=>"011110001",
  54020=>"100011101",
  54021=>"110000001",
  54022=>"001101111",
  54023=>"100011111",
  54024=>"011111001",
  54025=>"100110111",
  54026=>"101101000",
  54027=>"111001000",
  54028=>"010010000",
  54029=>"101000110",
  54030=>"111011100",
  54031=>"010011010",
  54032=>"101110010",
  54033=>"000100101",
  54034=>"100111110",
  54035=>"100110110",
  54036=>"101011011",
  54037=>"110011000",
  54038=>"000110000",
  54039=>"101100100",
  54040=>"111100110",
  54041=>"001111110",
  54042=>"100001001",
  54043=>"000011100",
  54044=>"011000101",
  54045=>"111010111",
  54046=>"110100000",
  54047=>"001001010",
  54048=>"110111110",
  54049=>"010100100",
  54050=>"110000011",
  54051=>"110001000",
  54052=>"101011001",
  54053=>"110111001",
  54054=>"010010110",
  54055=>"111010101",
  54056=>"010011000",
  54057=>"111100000",
  54058=>"101011011",
  54059=>"010000111",
  54060=>"110111010",
  54061=>"000001101",
  54062=>"001011001",
  54063=>"011100000",
  54064=>"000011011",
  54065=>"100100000",
  54066=>"100111010",
  54067=>"110101110",
  54068=>"111011111",
  54069=>"111110001",
  54070=>"001011001",
  54071=>"000011111",
  54072=>"101001100",
  54073=>"000001000",
  54074=>"011101100",
  54075=>"110001001",
  54076=>"101100101",
  54077=>"000001100",
  54078=>"101110101",
  54079=>"100001010",
  54080=>"111000111",
  54081=>"111100111",
  54082=>"010100010",
  54083=>"100010110",
  54084=>"000101110",
  54085=>"110110110",
  54086=>"010100000",
  54087=>"000111111",
  54088=>"001100100",
  54089=>"111001100",
  54090=>"001010110",
  54091=>"001110101",
  54092=>"001011001",
  54093=>"110001010",
  54094=>"100100000",
  54095=>"010011101",
  54096=>"010100010",
  54097=>"111000010",
  54098=>"101010011",
  54099=>"011010000",
  54100=>"111000010",
  54101=>"000101000",
  54102=>"100000001",
  54103=>"010010100",
  54104=>"101111000",
  54105=>"111011010",
  54106=>"100000110",
  54107=>"100001111",
  54108=>"111100110",
  54109=>"001000100",
  54110=>"001001001",
  54111=>"000000001",
  54112=>"111100111",
  54113=>"111010000",
  54114=>"000011101",
  54115=>"100110000",
  54116=>"110111111",
  54117=>"000111110",
  54118=>"001001011",
  54119=>"001011011",
  54120=>"111111111",
  54121=>"001000100",
  54122=>"110101100",
  54123=>"110101110",
  54124=>"011000001",
  54125=>"011001101",
  54126=>"001100110",
  54127=>"010100110",
  54128=>"111111000",
  54129=>"110001000",
  54130=>"100101101",
  54131=>"111011001",
  54132=>"111101001",
  54133=>"010010001",
  54134=>"000001111",
  54135=>"111000001",
  54136=>"110111001",
  54137=>"000010001",
  54138=>"111010111",
  54139=>"001110010",
  54140=>"000000000",
  54141=>"100000001",
  54142=>"011111100",
  54143=>"010011011",
  54144=>"010011000",
  54145=>"001111010",
  54146=>"101010000",
  54147=>"001001100",
  54148=>"001110111",
  54149=>"011011110",
  54150=>"000010010",
  54151=>"001110011",
  54152=>"111110000",
  54153=>"100000111",
  54154=>"000000001",
  54155=>"011000110",
  54156=>"111011101",
  54157=>"111111110",
  54158=>"000001011",
  54159=>"000100110",
  54160=>"000011000",
  54161=>"001010011",
  54162=>"001000000",
  54163=>"011001111",
  54164=>"101001000",
  54165=>"000000101",
  54166=>"101001010",
  54167=>"100101001",
  54168=>"111100101",
  54169=>"111001000",
  54170=>"011010000",
  54171=>"100010010",
  54172=>"000000111",
  54173=>"101000101",
  54174=>"000010100",
  54175=>"011110000",
  54176=>"100000101",
  54177=>"001101011",
  54178=>"101100000",
  54179=>"110101001",
  54180=>"001000000",
  54181=>"000111010",
  54182=>"101010111",
  54183=>"011000100",
  54184=>"010111000",
  54185=>"111001111",
  54186=>"000111111",
  54187=>"110111001",
  54188=>"110010011",
  54189=>"100011000",
  54190=>"010011001",
  54191=>"110111111",
  54192=>"110011101",
  54193=>"011101100",
  54194=>"101101110",
  54195=>"110110001",
  54196=>"010101100",
  54197=>"010111101",
  54198=>"101010011",
  54199=>"111001011",
  54200=>"111111111",
  54201=>"011000100",
  54202=>"011001001",
  54203=>"111100100",
  54204=>"111111101",
  54205=>"100101111",
  54206=>"111001001",
  54207=>"111110000",
  54208=>"110100101",
  54209=>"111101110",
  54210=>"110110001",
  54211=>"110010100",
  54212=>"000011000",
  54213=>"001101111",
  54214=>"000000011",
  54215=>"001001101",
  54216=>"111000111",
  54217=>"011111011",
  54218=>"011101110",
  54219=>"100100000",
  54220=>"100011011",
  54221=>"110100001",
  54222=>"000001110",
  54223=>"110110010",
  54224=>"101011111",
  54225=>"000000000",
  54226=>"011001001",
  54227=>"101010101",
  54228=>"001011011",
  54229=>"011011011",
  54230=>"111111010",
  54231=>"001110011",
  54232=>"101100100",
  54233=>"010100111",
  54234=>"011111110",
  54235=>"110010011",
  54236=>"000101110",
  54237=>"000111100",
  54238=>"010001000",
  54239=>"101011100",
  54240=>"000101001",
  54241=>"100000001",
  54242=>"001101010",
  54243=>"111100000",
  54244=>"111101101",
  54245=>"100000001",
  54246=>"010000010",
  54247=>"011111000",
  54248=>"000101111",
  54249=>"100001111",
  54250=>"111000110",
  54251=>"011110000",
  54252=>"110101111",
  54253=>"111101001",
  54254=>"100110101",
  54255=>"101001010",
  54256=>"101111010",
  54257=>"011001000",
  54258=>"000001000",
  54259=>"110111001",
  54260=>"000011110",
  54261=>"000010100",
  54262=>"001111110",
  54263=>"000001010",
  54264=>"010001111",
  54265=>"111011111",
  54266=>"000100001",
  54267=>"011110011",
  54268=>"100001000",
  54269=>"000010101",
  54270=>"101000000",
  54271=>"100011001",
  54272=>"000110111",
  54273=>"000000001",
  54274=>"110101110",
  54275=>"111001011",
  54276=>"011000111",
  54277=>"110100100",
  54278=>"001111010",
  54279=>"001001100",
  54280=>"110010101",
  54281=>"101011000",
  54282=>"110101100",
  54283=>"110110000",
  54284=>"000100001",
  54285=>"110000000",
  54286=>"000010100",
  54287=>"000010000",
  54288=>"001100010",
  54289=>"001001110",
  54290=>"111101111",
  54291=>"001100001",
  54292=>"111110100",
  54293=>"010001110",
  54294=>"111111010",
  54295=>"110101101",
  54296=>"010110000",
  54297=>"000011001",
  54298=>"110100001",
  54299=>"110111101",
  54300=>"001001111",
  54301=>"100011100",
  54302=>"111100101",
  54303=>"010011000",
  54304=>"011000011",
  54305=>"110001111",
  54306=>"010100101",
  54307=>"101111110",
  54308=>"111010101",
  54309=>"110110010",
  54310=>"000111100",
  54311=>"100111101",
  54312=>"001101000",
  54313=>"001101100",
  54314=>"110010010",
  54315=>"000000010",
  54316=>"110000011",
  54317=>"001101100",
  54318=>"011000001",
  54319=>"100101000",
  54320=>"001111110",
  54321=>"001000001",
  54322=>"110011101",
  54323=>"110100000",
  54324=>"111111000",
  54325=>"111011110",
  54326=>"010111100",
  54327=>"010011111",
  54328=>"100100110",
  54329=>"001110111",
  54330=>"010011001",
  54331=>"100011011",
  54332=>"000111101",
  54333=>"011000000",
  54334=>"010101101",
  54335=>"110011011",
  54336=>"101000110",
  54337=>"000001010",
  54338=>"010110010",
  54339=>"001101101",
  54340=>"000101111",
  54341=>"101111000",
  54342=>"101100100",
  54343=>"010011010",
  54344=>"001000101",
  54345=>"011000111",
  54346=>"001010010",
  54347=>"110111010",
  54348=>"110010000",
  54349=>"010100110",
  54350=>"010001100",
  54351=>"010001101",
  54352=>"101011001",
  54353=>"100100001",
  54354=>"101110101",
  54355=>"111010000",
  54356=>"111001001",
  54357=>"001001110",
  54358=>"010100101",
  54359=>"101111001",
  54360=>"100111011",
  54361=>"111000100",
  54362=>"110000010",
  54363=>"111110010",
  54364=>"010010001",
  54365=>"101001101",
  54366=>"010110110",
  54367=>"011101000",
  54368=>"011110000",
  54369=>"011011100",
  54370=>"111111101",
  54371=>"000111001",
  54372=>"111101001",
  54373=>"010111110",
  54374=>"001010011",
  54375=>"110001000",
  54376=>"111011001",
  54377=>"000111010",
  54378=>"001001010",
  54379=>"110110001",
  54380=>"000101101",
  54381=>"000100110",
  54382=>"001100010",
  54383=>"010100010",
  54384=>"011001110",
  54385=>"111110001",
  54386=>"110010100",
  54387=>"001011001",
  54388=>"001110100",
  54389=>"110101110",
  54390=>"011000011",
  54391=>"110110110",
  54392=>"101110011",
  54393=>"010110000",
  54394=>"000001101",
  54395=>"111010100",
  54396=>"001101111",
  54397=>"000010001",
  54398=>"111001100",
  54399=>"100010001",
  54400=>"100101101",
  54401=>"010100110",
  54402=>"111010011",
  54403=>"111011001",
  54404=>"110100101",
  54405=>"100011111",
  54406=>"000101000",
  54407=>"011010101",
  54408=>"011111011",
  54409=>"011110110",
  54410=>"110100001",
  54411=>"001001001",
  54412=>"111100100",
  54413=>"110100100",
  54414=>"011111100",
  54415=>"110010111",
  54416=>"001001010",
  54417=>"111011100",
  54418=>"100100100",
  54419=>"011111001",
  54420=>"100101000",
  54421=>"111110010",
  54422=>"001011001",
  54423=>"100011100",
  54424=>"010101000",
  54425=>"111100111",
  54426=>"000110101",
  54427=>"010101000",
  54428=>"111000100",
  54429=>"111001101",
  54430=>"100000100",
  54431=>"110000001",
  54432=>"000100100",
  54433=>"110011100",
  54434=>"101000100",
  54435=>"001110000",
  54436=>"001111011",
  54437=>"110111011",
  54438=>"010111110",
  54439=>"111011101",
  54440=>"110100101",
  54441=>"001011111",
  54442=>"000011010",
  54443=>"011100100",
  54444=>"011101111",
  54445=>"100100110",
  54446=>"110010010",
  54447=>"000100001",
  54448=>"000000001",
  54449=>"101011110",
  54450=>"110011110",
  54451=>"111001000",
  54452=>"101101101",
  54453=>"010000111",
  54454=>"001001111",
  54455=>"010111010",
  54456=>"000001011",
  54457=>"100100100",
  54458=>"001111010",
  54459=>"000000011",
  54460=>"000100100",
  54461=>"011000010",
  54462=>"110000001",
  54463=>"101111110",
  54464=>"011110101",
  54465=>"100000011",
  54466=>"000001111",
  54467=>"011101010",
  54468=>"111100101",
  54469=>"001110010",
  54470=>"111000110",
  54471=>"100011000",
  54472=>"101111101",
  54473=>"011110100",
  54474=>"110010101",
  54475=>"101001111",
  54476=>"001110010",
  54477=>"100000001",
  54478=>"011001101",
  54479=>"011101101",
  54480=>"010101011",
  54481=>"000010010",
  54482=>"101010110",
  54483=>"111010110",
  54484=>"011110111",
  54485=>"011111011",
  54486=>"101010100",
  54487=>"000110110",
  54488=>"111010111",
  54489=>"100101101",
  54490=>"011000101",
  54491=>"101010000",
  54492=>"101100110",
  54493=>"100010110",
  54494=>"001010111",
  54495=>"100101101",
  54496=>"100001001",
  54497=>"101000110",
  54498=>"001100000",
  54499=>"101100000",
  54500=>"111011110",
  54501=>"011000011",
  54502=>"001101111",
  54503=>"101011000",
  54504=>"100000010",
  54505=>"100011111",
  54506=>"101101111",
  54507=>"010010110",
  54508=>"100011111",
  54509=>"010010101",
  54510=>"101100001",
  54511=>"000000000",
  54512=>"101000001",
  54513=>"100110101",
  54514=>"111100010",
  54515=>"111011110",
  54516=>"100010100",
  54517=>"000101010",
  54518=>"111110110",
  54519=>"101100101",
  54520=>"011011011",
  54521=>"001111011",
  54522=>"101100110",
  54523=>"101110001",
  54524=>"111101001",
  54525=>"111010110",
  54526=>"101100111",
  54527=>"110001100",
  54528=>"110100000",
  54529=>"001111001",
  54530=>"101010001",
  54531=>"010011100",
  54532=>"011011010",
  54533=>"101111001",
  54534=>"101011100",
  54535=>"100101111",
  54536=>"011111000",
  54537=>"111111111",
  54538=>"001011100",
  54539=>"000011001",
  54540=>"110000101",
  54541=>"111101101",
  54542=>"001110101",
  54543=>"100010000",
  54544=>"011010111",
  54545=>"111000011",
  54546=>"001110010",
  54547=>"000011011",
  54548=>"000000010",
  54549=>"010000100",
  54550=>"000001000",
  54551=>"010101000",
  54552=>"111010011",
  54553=>"111011101",
  54554=>"111000001",
  54555=>"000001101",
  54556=>"010000110",
  54557=>"110111010",
  54558=>"111010000",
  54559=>"101000000",
  54560=>"100101011",
  54561=>"111000011",
  54562=>"111011101",
  54563=>"000101011",
  54564=>"000110001",
  54565=>"110000000",
  54566=>"001101101",
  54567=>"111101001",
  54568=>"001011110",
  54569=>"100001111",
  54570=>"110110101",
  54571=>"001010011",
  54572=>"000001001",
  54573=>"001111100",
  54574=>"000100110",
  54575=>"100100001",
  54576=>"100010000",
  54577=>"101110011",
  54578=>"110100110",
  54579=>"010000110",
  54580=>"101010101",
  54581=>"000101011",
  54582=>"111110011",
  54583=>"111101001",
  54584=>"000001001",
  54585=>"001010010",
  54586=>"001110111",
  54587=>"010000101",
  54588=>"111110010",
  54589=>"010010010",
  54590=>"101111011",
  54591=>"000011000",
  54592=>"110111100",
  54593=>"001001001",
  54594=>"110101101",
  54595=>"110101001",
  54596=>"101000111",
  54597=>"101011110",
  54598=>"001001011",
  54599=>"000111111",
  54600=>"011001011",
  54601=>"101011111",
  54602=>"101101101",
  54603=>"011011101",
  54604=>"111010111",
  54605=>"101111000",
  54606=>"110100101",
  54607=>"010111110",
  54608=>"000001001",
  54609=>"010001100",
  54610=>"110110111",
  54611=>"101111001",
  54612=>"100111101",
  54613=>"111111100",
  54614=>"101000101",
  54615=>"100101111",
  54616=>"101101100",
  54617=>"011010001",
  54618=>"011010000",
  54619=>"101110111",
  54620=>"001101110",
  54621=>"111001000",
  54622=>"011000000",
  54623=>"001010010",
  54624=>"101011011",
  54625=>"110011100",
  54626=>"000111101",
  54627=>"111001111",
  54628=>"010010010",
  54629=>"000001101",
  54630=>"011010111",
  54631=>"011101010",
  54632=>"000101011",
  54633=>"111011000",
  54634=>"110111101",
  54635=>"001111110",
  54636=>"110011000",
  54637=>"000001001",
  54638=>"110110000",
  54639=>"011000000",
  54640=>"110011010",
  54641=>"101110110",
  54642=>"001111001",
  54643=>"110101111",
  54644=>"100001111",
  54645=>"010001011",
  54646=>"101010111",
  54647=>"100001111",
  54648=>"101001101",
  54649=>"011001111",
  54650=>"100001100",
  54651=>"011110111",
  54652=>"010001100",
  54653=>"111111011",
  54654=>"010011110",
  54655=>"000001010",
  54656=>"000100111",
  54657=>"101101101",
  54658=>"001101101",
  54659=>"110011101",
  54660=>"101111101",
  54661=>"010000101",
  54662=>"111010000",
  54663=>"000000000",
  54664=>"111111111",
  54665=>"101011011",
  54666=>"101110101",
  54667=>"101011111",
  54668=>"100001110",
  54669=>"110110001",
  54670=>"001111110",
  54671=>"101010100",
  54672=>"010110101",
  54673=>"001111110",
  54674=>"011011000",
  54675=>"011101110",
  54676=>"111111010",
  54677=>"001001011",
  54678=>"100010000",
  54679=>"101000111",
  54680=>"101001000",
  54681=>"001001001",
  54682=>"010011000",
  54683=>"111110001",
  54684=>"101000010",
  54685=>"100010001",
  54686=>"011011011",
  54687=>"110011010",
  54688=>"000000101",
  54689=>"101110111",
  54690=>"100001110",
  54691=>"111000000",
  54692=>"000000101",
  54693=>"010011010",
  54694=>"010011110",
  54695=>"011101101",
  54696=>"101101000",
  54697=>"010110101",
  54698=>"100101011",
  54699=>"001001000",
  54700=>"101000000",
  54701=>"100010001",
  54702=>"111100101",
  54703=>"001101011",
  54704=>"001011101",
  54705=>"100000110",
  54706=>"001111110",
  54707=>"001001011",
  54708=>"011101101",
  54709=>"011111001",
  54710=>"101010111",
  54711=>"100100110",
  54712=>"110111010",
  54713=>"110100100",
  54714=>"100000110",
  54715=>"010110100",
  54716=>"100111010",
  54717=>"100101111",
  54718=>"101000100",
  54719=>"000110101",
  54720=>"101111001",
  54721=>"111101100",
  54722=>"111101010",
  54723=>"111011101",
  54724=>"100000111",
  54725=>"101101100",
  54726=>"011111001",
  54727=>"100111101",
  54728=>"001000111",
  54729=>"001100110",
  54730=>"010111001",
  54731=>"110110111",
  54732=>"011001011",
  54733=>"101110001",
  54734=>"101100101",
  54735=>"101100000",
  54736=>"110001110",
  54737=>"100111011",
  54738=>"001001100",
  54739=>"001101101",
  54740=>"001101101",
  54741=>"000001010",
  54742=>"000010011",
  54743=>"111111001",
  54744=>"001101010",
  54745=>"111110001",
  54746=>"111011000",
  54747=>"010111011",
  54748=>"111110000",
  54749=>"011000001",
  54750=>"110101011",
  54751=>"100100011",
  54752=>"100001110",
  54753=>"011010001",
  54754=>"110101111",
  54755=>"111110111",
  54756=>"111011110",
  54757=>"001110000",
  54758=>"101011010",
  54759=>"000101001",
  54760=>"010010000",
  54761=>"001101111",
  54762=>"010101010",
  54763=>"000101110",
  54764=>"001110101",
  54765=>"101010110",
  54766=>"100011100",
  54767=>"001111001",
  54768=>"001111000",
  54769=>"010011000",
  54770=>"000010100",
  54771=>"111111001",
  54772=>"001011110",
  54773=>"000000111",
  54774=>"001000110",
  54775=>"001101011",
  54776=>"111111100",
  54777=>"010010111",
  54778=>"101111000",
  54779=>"000111011",
  54780=>"111001010",
  54781=>"100110000",
  54782=>"000110000",
  54783=>"101101110",
  54784=>"011111101",
  54785=>"011000111",
  54786=>"111111101",
  54787=>"001000011",
  54788=>"111110110",
  54789=>"101101110",
  54790=>"000010001",
  54791=>"111110001",
  54792=>"011011101",
  54793=>"011000100",
  54794=>"101111010",
  54795=>"010011111",
  54796=>"111110100",
  54797=>"001111101",
  54798=>"000000010",
  54799=>"011110010",
  54800=>"000111100",
  54801=>"110011010",
  54802=>"000000001",
  54803=>"000101000",
  54804=>"110000001",
  54805=>"001111010",
  54806=>"000111000",
  54807=>"111011110",
  54808=>"110111010",
  54809=>"001011111",
  54810=>"111011110",
  54811=>"101111000",
  54812=>"111101110",
  54813=>"011011011",
  54814=>"111101001",
  54815=>"001111111",
  54816=>"000010011",
  54817=>"011110011",
  54818=>"011101111",
  54819=>"000100011",
  54820=>"101001100",
  54821=>"100010100",
  54822=>"110000111",
  54823=>"101111001",
  54824=>"010000100",
  54825=>"010110100",
  54826=>"000000110",
  54827=>"100100111",
  54828=>"001011101",
  54829=>"110010000",
  54830=>"110100100",
  54831=>"111110101",
  54832=>"111010110",
  54833=>"111111110",
  54834=>"010111011",
  54835=>"000010100",
  54836=>"011101000",
  54837=>"111001010",
  54838=>"000100110",
  54839=>"010110011",
  54840=>"000100101",
  54841=>"001011010",
  54842=>"000100001",
  54843=>"001011100",
  54844=>"010101000",
  54845=>"111100000",
  54846=>"000000001",
  54847=>"000000001",
  54848=>"000000001",
  54849=>"010101011",
  54850=>"110000101",
  54851=>"011110011",
  54852=>"001101001",
  54853=>"111101110",
  54854=>"001100101",
  54855=>"100001001",
  54856=>"100101010",
  54857=>"101000100",
  54858=>"010111100",
  54859=>"000101011",
  54860=>"110100100",
  54861=>"101000101",
  54862=>"111111101",
  54863=>"111010000",
  54864=>"001111010",
  54865=>"000010111",
  54866=>"000111010",
  54867=>"000100000",
  54868=>"001010010",
  54869=>"111000100",
  54870=>"000000111",
  54871=>"001000101",
  54872=>"101111101",
  54873=>"001011100",
  54874=>"110100000",
  54875=>"110111110",
  54876=>"000101011",
  54877=>"101101011",
  54878=>"001010110",
  54879=>"101100011",
  54880=>"011100100",
  54881=>"000000000",
  54882=>"101111111",
  54883=>"001000101",
  54884=>"111010011",
  54885=>"000000000",
  54886=>"000100100",
  54887=>"000010011",
  54888=>"111110110",
  54889=>"001001001",
  54890=>"010100000",
  54891=>"100010001",
  54892=>"100001111",
  54893=>"011001101",
  54894=>"110000010",
  54895=>"111111110",
  54896=>"111111001",
  54897=>"111110110",
  54898=>"001011110",
  54899=>"001011011",
  54900=>"011011111",
  54901=>"111111110",
  54902=>"000000110",
  54903=>"111000000",
  54904=>"001110001",
  54905=>"110010011",
  54906=>"011011101",
  54907=>"000110101",
  54908=>"001000000",
  54909=>"010010101",
  54910=>"101010001",
  54911=>"111000001",
  54912=>"101010000",
  54913=>"001001110",
  54914=>"000100100",
  54915=>"001110111",
  54916=>"000100111",
  54917=>"011111000",
  54918=>"001101000",
  54919=>"011010111",
  54920=>"110011011",
  54921=>"010001111",
  54922=>"101111100",
  54923=>"111111110",
  54924=>"101000101",
  54925=>"101111100",
  54926=>"001100101",
  54927=>"001001010",
  54928=>"100000110",
  54929=>"111100110",
  54930=>"011010101",
  54931=>"001111101",
  54932=>"101001111",
  54933=>"101100111",
  54934=>"111000110",
  54935=>"111111101",
  54936=>"001111010",
  54937=>"101101100",
  54938=>"101000011",
  54939=>"010011111",
  54940=>"000000111",
  54941=>"111100111",
  54942=>"100110011",
  54943=>"101010010",
  54944=>"010001000",
  54945=>"110011110",
  54946=>"110110100",
  54947=>"100000001",
  54948=>"101001111",
  54949=>"000100100",
  54950=>"011010111",
  54951=>"100011010",
  54952=>"101010110",
  54953=>"100100101",
  54954=>"001000111",
  54955=>"011110001",
  54956=>"110110000",
  54957=>"100110111",
  54958=>"000000100",
  54959=>"000100001",
  54960=>"000000000",
  54961=>"010001101",
  54962=>"011001001",
  54963=>"011000111",
  54964=>"010100100",
  54965=>"101100111",
  54966=>"011101101",
  54967=>"010110111",
  54968=>"110000110",
  54969=>"010110110",
  54970=>"000010110",
  54971=>"001100111",
  54972=>"111111101",
  54973=>"010001101",
  54974=>"100001101",
  54975=>"000100011",
  54976=>"110000100",
  54977=>"101011101",
  54978=>"110110000",
  54979=>"000000010",
  54980=>"011101011",
  54981=>"100100100",
  54982=>"011100101",
  54983=>"011010101",
  54984=>"000000101",
  54985=>"000100010",
  54986=>"111000110",
  54987=>"000000111",
  54988=>"001110000",
  54989=>"100111111",
  54990=>"011110011",
  54991=>"001000000",
  54992=>"011110100",
  54993=>"100010100",
  54994=>"101001010",
  54995=>"001111011",
  54996=>"110111110",
  54997=>"111011110",
  54998=>"100011101",
  54999=>"010001110",
  55000=>"010011010",
  55001=>"100001000",
  55002=>"100000110",
  55003=>"010000101",
  55004=>"111000000",
  55005=>"011111000",
  55006=>"010010110",
  55007=>"110111101",
  55008=>"100010001",
  55009=>"100001111",
  55010=>"100100101",
  55011=>"111011010",
  55012=>"011010101",
  55013=>"110001000",
  55014=>"001111000",
  55015=>"010011001",
  55016=>"110111100",
  55017=>"000101101",
  55018=>"011010001",
  55019=>"010001000",
  55020=>"111110010",
  55021=>"100000101",
  55022=>"111110110",
  55023=>"110011111",
  55024=>"010111110",
  55025=>"111110001",
  55026=>"001101110",
  55027=>"110000111",
  55028=>"111110100",
  55029=>"011001100",
  55030=>"010011011",
  55031=>"000010000",
  55032=>"000011010",
  55033=>"000010001",
  55034=>"011101111",
  55035=>"110010001",
  55036=>"000001111",
  55037=>"101110010",
  55038=>"011100101",
  55039=>"000100011",
  55040=>"111010101",
  55041=>"010011110",
  55042=>"110110111",
  55043=>"011000000",
  55044=>"011110110",
  55045=>"111010100",
  55046=>"101110001",
  55047=>"100100001",
  55048=>"101110001",
  55049=>"100111110",
  55050=>"010101111",
  55051=>"011000001",
  55052=>"010010010",
  55053=>"001100110",
  55054=>"011101110",
  55055=>"111101000",
  55056=>"010110000",
  55057=>"111100111",
  55058=>"111010010",
  55059=>"011101110",
  55060=>"100010110",
  55061=>"010110000",
  55062=>"000101110",
  55063=>"010110001",
  55064=>"011111001",
  55065=>"000111110",
  55066=>"100101110",
  55067=>"000000100",
  55068=>"011101010",
  55069=>"011100110",
  55070=>"110000101",
  55071=>"010011001",
  55072=>"111101110",
  55073=>"100101000",
  55074=>"100001010",
  55075=>"011101001",
  55076=>"110001000",
  55077=>"100101100",
  55078=>"001001000",
  55079=>"110100110",
  55080=>"101110000",
  55081=>"101111110",
  55082=>"111110000",
  55083=>"010110000",
  55084=>"000100100",
  55085=>"111111101",
  55086=>"000100101",
  55087=>"011000000",
  55088=>"011001001",
  55089=>"110000100",
  55090=>"011101110",
  55091=>"110011100",
  55092=>"101111001",
  55093=>"011011010",
  55094=>"111101100",
  55095=>"110100000",
  55096=>"100100110",
  55097=>"100101001",
  55098=>"110001100",
  55099=>"101001100",
  55100=>"011110111",
  55101=>"000101010",
  55102=>"111010110",
  55103=>"111100111",
  55104=>"000000001",
  55105=>"000100011",
  55106=>"001101110",
  55107=>"001110001",
  55108=>"000101000",
  55109=>"001010100",
  55110=>"000101001",
  55111=>"100100001",
  55112=>"101010111",
  55113=>"111000010",
  55114=>"110000001",
  55115=>"101000000",
  55116=>"000001101",
  55117=>"011000111",
  55118=>"011110100",
  55119=>"000011010",
  55120=>"001001101",
  55121=>"011111001",
  55122=>"001100001",
  55123=>"100010011",
  55124=>"101100001",
  55125=>"100011000",
  55126=>"001010101",
  55127=>"101000011",
  55128=>"111110111",
  55129=>"011101111",
  55130=>"101111101",
  55131=>"101111100",
  55132=>"101001010",
  55133=>"101011011",
  55134=>"001000111",
  55135=>"100101110",
  55136=>"000100010",
  55137=>"101101100",
  55138=>"100111011",
  55139=>"000011010",
  55140=>"110101001",
  55141=>"010000000",
  55142=>"101110111",
  55143=>"110101000",
  55144=>"000001000",
  55145=>"111110111",
  55146=>"100101101",
  55147=>"100110011",
  55148=>"100010010",
  55149=>"001000000",
  55150=>"100011010",
  55151=>"110011110",
  55152=>"100100101",
  55153=>"111110001",
  55154=>"111001010",
  55155=>"000000111",
  55156=>"001100100",
  55157=>"111100110",
  55158=>"000001111",
  55159=>"110011101",
  55160=>"101000111",
  55161=>"110011011",
  55162=>"101001110",
  55163=>"001000100",
  55164=>"010111100",
  55165=>"011011110",
  55166=>"000000010",
  55167=>"111110001",
  55168=>"101001010",
  55169=>"001010101",
  55170=>"111000101",
  55171=>"100010010",
  55172=>"001000000",
  55173=>"001000100",
  55174=>"100000100",
  55175=>"100010010",
  55176=>"001101001",
  55177=>"000011101",
  55178=>"001010001",
  55179=>"001101100",
  55180=>"011011001",
  55181=>"100110110",
  55182=>"100001010",
  55183=>"100111101",
  55184=>"111001101",
  55185=>"111001101",
  55186=>"101101001",
  55187=>"000101000",
  55188=>"100100001",
  55189=>"101011111",
  55190=>"011001001",
  55191=>"000000000",
  55192=>"111000100",
  55193=>"111101111",
  55194=>"111110111",
  55195=>"001100110",
  55196=>"100100110",
  55197=>"001011010",
  55198=>"010100011",
  55199=>"011111010",
  55200=>"101011011",
  55201=>"110100010",
  55202=>"000010110",
  55203=>"110101101",
  55204=>"001100010",
  55205=>"010101110",
  55206=>"111111010",
  55207=>"001111011",
  55208=>"001111110",
  55209=>"001100001",
  55210=>"000001100",
  55211=>"110100011",
  55212=>"111010110",
  55213=>"100001110",
  55214=>"000100101",
  55215=>"111010010",
  55216=>"111111000",
  55217=>"111100010",
  55218=>"111001100",
  55219=>"110001011",
  55220=>"000001000",
  55221=>"101010110",
  55222=>"101001011",
  55223=>"011010000",
  55224=>"000100001",
  55225=>"001010011",
  55226=>"100111000",
  55227=>"101110100",
  55228=>"011010111",
  55229=>"111010001",
  55230=>"110100110",
  55231=>"100001111",
  55232=>"010100110",
  55233=>"011011000",
  55234=>"111101000",
  55235=>"100001101",
  55236=>"000001100",
  55237=>"101110010",
  55238=>"111011110",
  55239=>"110111101",
  55240=>"101110000",
  55241=>"101100011",
  55242=>"101110101",
  55243=>"000101110",
  55244=>"111100001",
  55245=>"111000000",
  55246=>"010000000",
  55247=>"110001100",
  55248=>"011011101",
  55249=>"100000000",
  55250=>"000100001",
  55251=>"000111010",
  55252=>"001011011",
  55253=>"100111001",
  55254=>"110010001",
  55255=>"010111110",
  55256=>"000000001",
  55257=>"100101000",
  55258=>"010010111",
  55259=>"100110100",
  55260=>"110111111",
  55261=>"000100001",
  55262=>"000101001",
  55263=>"100101000",
  55264=>"101101111",
  55265=>"111100010",
  55266=>"011001011",
  55267=>"110010001",
  55268=>"000100001",
  55269=>"100011110",
  55270=>"111011111",
  55271=>"111100000",
  55272=>"010101010",
  55273=>"011000010",
  55274=>"001001010",
  55275=>"111100100",
  55276=>"111111101",
  55277=>"010010000",
  55278=>"010011000",
  55279=>"000110100",
  55280=>"011101000",
  55281=>"001110001",
  55282=>"001000101",
  55283=>"110111010",
  55284=>"010101000",
  55285=>"111000010",
  55286=>"000000011",
  55287=>"000000010",
  55288=>"010101010",
  55289=>"111100000",
  55290=>"000000000",
  55291=>"111101000",
  55292=>"001001001",
  55293=>"011111110",
  55294=>"101011011",
  55295=>"011010001",
  55296=>"101100001",
  55297=>"010011000",
  55298=>"001000011",
  55299=>"111010001",
  55300=>"011010100",
  55301=>"101111101",
  55302=>"001000000",
  55303=>"011000100",
  55304=>"000111011",
  55305=>"110100011",
  55306=>"100010110",
  55307=>"111010110",
  55308=>"111111110",
  55309=>"100011110",
  55310=>"010101001",
  55311=>"111111100",
  55312=>"010100100",
  55313=>"000110101",
  55314=>"110100011",
  55315=>"011111111",
  55316=>"110111001",
  55317=>"100101100",
  55318=>"110111111",
  55319=>"000001110",
  55320=>"010111101",
  55321=>"110111001",
  55322=>"100011110",
  55323=>"001011100",
  55324=>"001010010",
  55325=>"011111000",
  55326=>"110101101",
  55327=>"111101011",
  55328=>"101011100",
  55329=>"111011111",
  55330=>"100010100",
  55331=>"110111010",
  55332=>"111011010",
  55333=>"101101101",
  55334=>"100001110",
  55335=>"000001011",
  55336=>"110111100",
  55337=>"111011011",
  55338=>"011111101",
  55339=>"100010110",
  55340=>"011100011",
  55341=>"001101110",
  55342=>"010000110",
  55343=>"000101011",
  55344=>"100100101",
  55345=>"000110101",
  55346=>"001010000",
  55347=>"001111100",
  55348=>"010101011",
  55349=>"011010001",
  55350=>"001010100",
  55351=>"101100101",
  55352=>"000110100",
  55353=>"100100010",
  55354=>"001100000",
  55355=>"011111111",
  55356=>"100101110",
  55357=>"001110000",
  55358=>"100110011",
  55359=>"010100010",
  55360=>"110100111",
  55361=>"001110000",
  55362=>"110010000",
  55363=>"100001001",
  55364=>"111011110",
  55365=>"001110100",
  55366=>"111010000",
  55367=>"001010110",
  55368=>"111000101",
  55369=>"000010100",
  55370=>"010011001",
  55371=>"000010010",
  55372=>"011011011",
  55373=>"011110100",
  55374=>"001001011",
  55375=>"111101100",
  55376=>"000010101",
  55377=>"000010010",
  55378=>"001111111",
  55379=>"011000101",
  55380=>"100110100",
  55381=>"001001001",
  55382=>"111101011",
  55383=>"000101110",
  55384=>"000011010",
  55385=>"001110101",
  55386=>"010001011",
  55387=>"111011101",
  55388=>"001011111",
  55389=>"111001101",
  55390=>"001101001",
  55391=>"011100000",
  55392=>"111010111",
  55393=>"001010010",
  55394=>"001110100",
  55395=>"110001010",
  55396=>"110011001",
  55397=>"110111010",
  55398=>"000100001",
  55399=>"110011001",
  55400=>"000110000",
  55401=>"111100001",
  55402=>"101000101",
  55403=>"110110111",
  55404=>"010011001",
  55405=>"001100000",
  55406=>"101110100",
  55407=>"001001010",
  55408=>"111110110",
  55409=>"101101100",
  55410=>"111101000",
  55411=>"001111001",
  55412=>"010101001",
  55413=>"111001111",
  55414=>"101101101",
  55415=>"000001110",
  55416=>"011110110",
  55417=>"001000101",
  55418=>"111111100",
  55419=>"110011110",
  55420=>"110110110",
  55421=>"111100000",
  55422=>"010101100",
  55423=>"100011011",
  55424=>"100000111",
  55425=>"000011011",
  55426=>"111111011",
  55427=>"000101101",
  55428=>"101110111",
  55429=>"111010000",
  55430=>"111110000",
  55431=>"001110010",
  55432=>"110101011",
  55433=>"011110111",
  55434=>"100000110",
  55435=>"111111100",
  55436=>"000010000",
  55437=>"011011111",
  55438=>"011001011",
  55439=>"001001101",
  55440=>"100110101",
  55441=>"000010111",
  55442=>"000000110",
  55443=>"101001101",
  55444=>"110111010",
  55445=>"000110001",
  55446=>"010101000",
  55447=>"110111101",
  55448=>"000011001",
  55449=>"111001110",
  55450=>"111111000",
  55451=>"101001110",
  55452=>"101110001",
  55453=>"110001101",
  55454=>"000101010",
  55455=>"001100001",
  55456=>"110011000",
  55457=>"001001101",
  55458=>"000011001",
  55459=>"010010001",
  55460=>"010000101",
  55461=>"101000111",
  55462=>"110000000",
  55463=>"110110100",
  55464=>"110000001",
  55465=>"011000110",
  55466=>"101110001",
  55467=>"001011111",
  55468=>"011001111",
  55469=>"001101110",
  55470=>"101101111",
  55471=>"110001110",
  55472=>"001010110",
  55473=>"100110000",
  55474=>"000101001",
  55475=>"001011001",
  55476=>"011010001",
  55477=>"100001000",
  55478=>"001000111",
  55479=>"111101000",
  55480=>"101010100",
  55481=>"110001011",
  55482=>"101000010",
  55483=>"001111100",
  55484=>"111110000",
  55485=>"001111000",
  55486=>"011111111",
  55487=>"000111011",
  55488=>"001100100",
  55489=>"100110001",
  55490=>"000011000",
  55491=>"110010101",
  55492=>"000111000",
  55493=>"111100011",
  55494=>"110100001",
  55495=>"000010011",
  55496=>"110001001",
  55497=>"000010111",
  55498=>"110111100",
  55499=>"101011000",
  55500=>"001011100",
  55501=>"010011011",
  55502=>"101001001",
  55503=>"001100011",
  55504=>"000111111",
  55505=>"000001000",
  55506=>"110000001",
  55507=>"010011001",
  55508=>"001101000",
  55509=>"111001111",
  55510=>"111011100",
  55511=>"101000100",
  55512=>"101101000",
  55513=>"110101111",
  55514=>"011111010",
  55515=>"011011101",
  55516=>"110011000",
  55517=>"001100111",
  55518=>"111111000",
  55519=>"101101110",
  55520=>"111110110",
  55521=>"000011110",
  55522=>"111011000",
  55523=>"010000001",
  55524=>"000101101",
  55525=>"000110000",
  55526=>"100100001",
  55527=>"001011100",
  55528=>"110010010",
  55529=>"101110000",
  55530=>"010101100",
  55531=>"100111011",
  55532=>"101011101",
  55533=>"110011011",
  55534=>"100100001",
  55535=>"100101001",
  55536=>"000101101",
  55537=>"111000001",
  55538=>"111110000",
  55539=>"111011110",
  55540=>"010001100",
  55541=>"111000011",
  55542=>"010101011",
  55543=>"011000101",
  55544=>"101001111",
  55545=>"010010001",
  55546=>"011010110",
  55547=>"011100000",
  55548=>"000111111",
  55549=>"011000001",
  55550=>"011100111",
  55551=>"100001000",
  55552=>"110000010",
  55553=>"111101000",
  55554=>"110100010",
  55555=>"110010000",
  55556=>"110101010",
  55557=>"100001010",
  55558=>"011011101",
  55559=>"101111111",
  55560=>"110011011",
  55561=>"001011010",
  55562=>"001111111",
  55563=>"000100001",
  55564=>"011011101",
  55565=>"000011100",
  55566=>"110011100",
  55567=>"001000100",
  55568=>"101100111",
  55569=>"101001011",
  55570=>"100000111",
  55571=>"011001110",
  55572=>"111000000",
  55573=>"011110111",
  55574=>"000101110",
  55575=>"110101110",
  55576=>"101001010",
  55577=>"101010111",
  55578=>"100001011",
  55579=>"011111001",
  55580=>"001000001",
  55581=>"000100101",
  55582=>"111100001",
  55583=>"011110010",
  55584=>"101001010",
  55585=>"011001111",
  55586=>"001101100",
  55587=>"110100111",
  55588=>"000100011",
  55589=>"111011010",
  55590=>"100011010",
  55591=>"101010100",
  55592=>"100001011",
  55593=>"010010010",
  55594=>"101111110",
  55595=>"111010000",
  55596=>"001100110",
  55597=>"001011100",
  55598=>"101000000",
  55599=>"011101010",
  55600=>"111110111",
  55601=>"010101010",
  55602=>"011001111",
  55603=>"010101100",
  55604=>"000111110",
  55605=>"010000100",
  55606=>"010000000",
  55607=>"000001101",
  55608=>"110100000",
  55609=>"001011110",
  55610=>"101001110",
  55611=>"010000000",
  55612=>"001100001",
  55613=>"001010101",
  55614=>"111100000",
  55615=>"111001100",
  55616=>"101101111",
  55617=>"100010110",
  55618=>"001111111",
  55619=>"011010001",
  55620=>"100011101",
  55621=>"100010000",
  55622=>"110011000",
  55623=>"111101101",
  55624=>"011010101",
  55625=>"101001010",
  55626=>"111010000",
  55627=>"111111111",
  55628=>"111000110",
  55629=>"111111110",
  55630=>"010110001",
  55631=>"011110111",
  55632=>"110111011",
  55633=>"100010001",
  55634=>"010110100",
  55635=>"011111110",
  55636=>"110111100",
  55637=>"011010011",
  55638=>"000100101",
  55639=>"000100111",
  55640=>"111110010",
  55641=>"101100101",
  55642=>"001100010",
  55643=>"011000001",
  55644=>"111101110",
  55645=>"011111001",
  55646=>"111100000",
  55647=>"101110111",
  55648=>"101000101",
  55649=>"111010000",
  55650=>"000011001",
  55651=>"111111100",
  55652=>"010010101",
  55653=>"100000100",
  55654=>"101100001",
  55655=>"011010111",
  55656=>"001100001",
  55657=>"001100010",
  55658=>"001001010",
  55659=>"110010000",
  55660=>"011000110",
  55661=>"000111111",
  55662=>"000011100",
  55663=>"100111111",
  55664=>"111001011",
  55665=>"101110101",
  55666=>"111110001",
  55667=>"011001101",
  55668=>"111110001",
  55669=>"001001010",
  55670=>"000000110",
  55671=>"111001100",
  55672=>"101100010",
  55673=>"010010101",
  55674=>"100011110",
  55675=>"000100010",
  55676=>"001100110",
  55677=>"010000001",
  55678=>"001011101",
  55679=>"011000111",
  55680=>"010001000",
  55681=>"111101100",
  55682=>"101100001",
  55683=>"001000011",
  55684=>"010011101",
  55685=>"111011111",
  55686=>"000111110",
  55687=>"101101110",
  55688=>"101100011",
  55689=>"100110101",
  55690=>"011011010",
  55691=>"111100001",
  55692=>"110000010",
  55693=>"000111011",
  55694=>"000011000",
  55695=>"101010001",
  55696=>"101101110",
  55697=>"110010000",
  55698=>"001011001",
  55699=>"111100000",
  55700=>"011111111",
  55701=>"001001011",
  55702=>"001100100",
  55703=>"001001000",
  55704=>"000001010",
  55705=>"001001101",
  55706=>"000100110",
  55707=>"000100011",
  55708=>"101100110",
  55709=>"111111101",
  55710=>"010101111",
  55711=>"001111111",
  55712=>"101010111",
  55713=>"000000000",
  55714=>"110110110",
  55715=>"001000100",
  55716=>"000010001",
  55717=>"001110110",
  55718=>"010011111",
  55719=>"110100001",
  55720=>"001011111",
  55721=>"011111111",
  55722=>"000000001",
  55723=>"000001011",
  55724=>"011111111",
  55725=>"001000100",
  55726=>"110010000",
  55727=>"001001111",
  55728=>"111011101",
  55729=>"100010100",
  55730=>"010010000",
  55731=>"000111001",
  55732=>"110110001",
  55733=>"000001011",
  55734=>"001100100",
  55735=>"000010001",
  55736=>"001001101",
  55737=>"010000111",
  55738=>"101001011",
  55739=>"000010001",
  55740=>"000110010",
  55741=>"110011010",
  55742=>"010100110",
  55743=>"001001100",
  55744=>"100011000",
  55745=>"001000000",
  55746=>"101111010",
  55747=>"100000000",
  55748=>"000100011",
  55749=>"101100101",
  55750=>"101101000",
  55751=>"011011000",
  55752=>"110010011",
  55753=>"000011111",
  55754=>"110101000",
  55755=>"110010000",
  55756=>"100110100",
  55757=>"110111111",
  55758=>"110010110",
  55759=>"100011111",
  55760=>"011101110",
  55761=>"001000101",
  55762=>"111100010",
  55763=>"101110010",
  55764=>"101110110",
  55765=>"100101100",
  55766=>"100101111",
  55767=>"111011011",
  55768=>"001001100",
  55769=>"110011011",
  55770=>"101000101",
  55771=>"100010110",
  55772=>"100000111",
  55773=>"010001111",
  55774=>"100000010",
  55775=>"011110010",
  55776=>"000001011",
  55777=>"100111101",
  55778=>"011110011",
  55779=>"010100101",
  55780=>"110000100",
  55781=>"010010100",
  55782=>"000100001",
  55783=>"001010111",
  55784=>"101111000",
  55785=>"100001100",
  55786=>"100011101",
  55787=>"010001000",
  55788=>"101001111",
  55789=>"000101001",
  55790=>"101110111",
  55791=>"111110011",
  55792=>"010001011",
  55793=>"111010000",
  55794=>"000110110",
  55795=>"101101100",
  55796=>"110010101",
  55797=>"101010100",
  55798=>"011010001",
  55799=>"100011110",
  55800=>"111010010",
  55801=>"111100100",
  55802=>"000101110",
  55803=>"100001010",
  55804=>"000100000",
  55805=>"110101010",
  55806=>"111010001",
  55807=>"000111001",
  55808=>"000000110",
  55809=>"111101010",
  55810=>"100011100",
  55811=>"110011001",
  55812=>"000110111",
  55813=>"000010000",
  55814=>"110101010",
  55815=>"111110010",
  55816=>"001010000",
  55817=>"110000001",
  55818=>"001110100",
  55819=>"100111110",
  55820=>"111100000",
  55821=>"010110110",
  55822=>"111100001",
  55823=>"001010110",
  55824=>"111010110",
  55825=>"110001110",
  55826=>"101101111",
  55827=>"110011111",
  55828=>"001010110",
  55829=>"010001001",
  55830=>"101011010",
  55831=>"010110100",
  55832=>"110001110",
  55833=>"011001100",
  55834=>"110000000",
  55835=>"111111001",
  55836=>"111010110",
  55837=>"100001110",
  55838=>"110010111",
  55839=>"011111000",
  55840=>"000100111",
  55841=>"100111010",
  55842=>"001010010",
  55843=>"101001000",
  55844=>"101110010",
  55845=>"101101110",
  55846=>"000100011",
  55847=>"100011010",
  55848=>"001011011",
  55849=>"100010011",
  55850=>"110110000",
  55851=>"101110011",
  55852=>"101101001",
  55853=>"011111011",
  55854=>"000101010",
  55855=>"100000110",
  55856=>"101101101",
  55857=>"100011101",
  55858=>"101011001",
  55859=>"111001000",
  55860=>"101010001",
  55861=>"010110010",
  55862=>"000001101",
  55863=>"101100011",
  55864=>"010010101",
  55865=>"111101001",
  55866=>"100001010",
  55867=>"011000001",
  55868=>"010010110",
  55869=>"010011101",
  55870=>"001100111",
  55871=>"111101001",
  55872=>"010101000",
  55873=>"111101000",
  55874=>"111011010",
  55875=>"110000110",
  55876=>"000000111",
  55877=>"100101111",
  55878=>"110110000",
  55879=>"010101111",
  55880=>"101101001",
  55881=>"001100011",
  55882=>"001101001",
  55883=>"110010111",
  55884=>"111111011",
  55885=>"011111100",
  55886=>"000000000",
  55887=>"101101010",
  55888=>"001111100",
  55889=>"001100011",
  55890=>"000101101",
  55891=>"011011000",
  55892=>"000100000",
  55893=>"001010000",
  55894=>"111110001",
  55895=>"010010111",
  55896=>"001000010",
  55897=>"111111001",
  55898=>"111110100",
  55899=>"011111110",
  55900=>"010000001",
  55901=>"000010101",
  55902=>"000010011",
  55903=>"100010010",
  55904=>"110101110",
  55905=>"001010011",
  55906=>"010111010",
  55907=>"001001110",
  55908=>"111010111",
  55909=>"000010001",
  55910=>"001010100",
  55911=>"100111111",
  55912=>"011000001",
  55913=>"110011010",
  55914=>"010000000",
  55915=>"011011101",
  55916=>"101100100",
  55917=>"110100001",
  55918=>"111010110",
  55919=>"010111111",
  55920=>"000000111",
  55921=>"100001100",
  55922=>"100100010",
  55923=>"100100011",
  55924=>"001111101",
  55925=>"110010111",
  55926=>"010110000",
  55927=>"000110010",
  55928=>"011101010",
  55929=>"101000010",
  55930=>"110001000",
  55931=>"001111011",
  55932=>"010101011",
  55933=>"111110011",
  55934=>"111110100",
  55935=>"000011100",
  55936=>"001011110",
  55937=>"010101100",
  55938=>"000110110",
  55939=>"100110110",
  55940=>"001010100",
  55941=>"011111010",
  55942=>"111101100",
  55943=>"111110001",
  55944=>"010000110",
  55945=>"000011010",
  55946=>"110010011",
  55947=>"110010111",
  55948=>"001011000",
  55949=>"010011011",
  55950=>"010000011",
  55951=>"100001010",
  55952=>"101001100",
  55953=>"000001010",
  55954=>"100001110",
  55955=>"111000010",
  55956=>"100011010",
  55957=>"000010001",
  55958=>"000011110",
  55959=>"100011010",
  55960=>"011101100",
  55961=>"011111000",
  55962=>"110010100",
  55963=>"011011101",
  55964=>"010010110",
  55965=>"010110011",
  55966=>"111110110",
  55967=>"010101101",
  55968=>"000011011",
  55969=>"000010001",
  55970=>"010100110",
  55971=>"111111101",
  55972=>"100000101",
  55973=>"100000110",
  55974=>"010000010",
  55975=>"100000101",
  55976=>"001010001",
  55977=>"100001110",
  55978=>"110110101",
  55979=>"000000100",
  55980=>"010111011",
  55981=>"000010010",
  55982=>"010101011",
  55983=>"110111110",
  55984=>"110101011",
  55985=>"000001100",
  55986=>"111001010",
  55987=>"010110110",
  55988=>"001100100",
  55989=>"111000100",
  55990=>"010111101",
  55991=>"100101100",
  55992=>"100010100",
  55993=>"101000010",
  55994=>"000101011",
  55995=>"111001001",
  55996=>"000100000",
  55997=>"110111001",
  55998=>"101100101",
  55999=>"010000010",
  56000=>"111111011",
  56001=>"110111111",
  56002=>"000010000",
  56003=>"111001010",
  56004=>"100010010",
  56005=>"001111001",
  56006=>"111111111",
  56007=>"111011110",
  56008=>"100011111",
  56009=>"101111000",
  56010=>"100110001",
  56011=>"011010011",
  56012=>"111101010",
  56013=>"000100100",
  56014=>"011001000",
  56015=>"000001110",
  56016=>"001110000",
  56017=>"001010110",
  56018=>"011101000",
  56019=>"100110110",
  56020=>"011000001",
  56021=>"111010111",
  56022=>"110101101",
  56023=>"000001010",
  56024=>"001011111",
  56025=>"000011110",
  56026=>"000111100",
  56027=>"100100000",
  56028=>"001000010",
  56029=>"101100010",
  56030=>"011011010",
  56031=>"111101000",
  56032=>"101101000",
  56033=>"111010110",
  56034=>"101101010",
  56035=>"000101000",
  56036=>"010000011",
  56037=>"011001001",
  56038=>"000010000",
  56039=>"010000110",
  56040=>"110101010",
  56041=>"000001101",
  56042=>"010010100",
  56043=>"111111111",
  56044=>"010110010",
  56045=>"001010010",
  56046=>"111111111",
  56047=>"000100111",
  56048=>"000011010",
  56049=>"000110010",
  56050=>"000001100",
  56051=>"111100011",
  56052=>"111000100",
  56053=>"111010010",
  56054=>"011011101",
  56055=>"000001000",
  56056=>"000011001",
  56057=>"011110111",
  56058=>"010100000",
  56059=>"001011101",
  56060=>"001010100",
  56061=>"011101111",
  56062=>"000100000",
  56063=>"010111010",
  56064=>"110010110",
  56065=>"000000100",
  56066=>"100010100",
  56067=>"000011011",
  56068=>"010000011",
  56069=>"101010111",
  56070=>"100100010",
  56071=>"111110101",
  56072=>"011100101",
  56073=>"001011010",
  56074=>"111010000",
  56075=>"111110111",
  56076=>"110010011",
  56077=>"101010000",
  56078=>"110010000",
  56079=>"101111111",
  56080=>"000001111",
  56081=>"011011110",
  56082=>"101001011",
  56083=>"101011111",
  56084=>"000101010",
  56085=>"101001100",
  56086=>"101000101",
  56087=>"010101010",
  56088=>"101000110",
  56089=>"101100000",
  56090=>"111101101",
  56091=>"101000000",
  56092=>"001110110",
  56093=>"010110011",
  56094=>"111100100",
  56095=>"111001100",
  56096=>"011001110",
  56097=>"101100000",
  56098=>"101000100",
  56099=>"111111111",
  56100=>"100001010",
  56101=>"000110101",
  56102=>"000100000",
  56103=>"000101001",
  56104=>"110011001",
  56105=>"011001111",
  56106=>"100011111",
  56107=>"010000110",
  56108=>"101011011",
  56109=>"010011000",
  56110=>"110100111",
  56111=>"110001010",
  56112=>"100010111",
  56113=>"110011000",
  56114=>"101100001",
  56115=>"110001110",
  56116=>"000101111",
  56117=>"111010000",
  56118=>"101010110",
  56119=>"010111111",
  56120=>"110000011",
  56121=>"010101010",
  56122=>"110001010",
  56123=>"000110000",
  56124=>"101011000",
  56125=>"010011001",
  56126=>"011011111",
  56127=>"001000111",
  56128=>"100100111",
  56129=>"100001011",
  56130=>"001101110",
  56131=>"111100110",
  56132=>"100100110",
  56133=>"110010011",
  56134=>"111110100",
  56135=>"111010000",
  56136=>"110111111",
  56137=>"001010111",
  56138=>"110001000",
  56139=>"010100011",
  56140=>"011001101",
  56141=>"000111100",
  56142=>"101011111",
  56143=>"011011011",
  56144=>"111011111",
  56145=>"110001110",
  56146=>"001011000",
  56147=>"101100110",
  56148=>"001000000",
  56149=>"000011100",
  56150=>"100010100",
  56151=>"010011100",
  56152=>"011110010",
  56153=>"110100011",
  56154=>"101001010",
  56155=>"000010011",
  56156=>"011000101",
  56157=>"100000001",
  56158=>"011100000",
  56159=>"011101100",
  56160=>"100001010",
  56161=>"001100010",
  56162=>"101001101",
  56163=>"110101111",
  56164=>"110100001",
  56165=>"101011000",
  56166=>"100110101",
  56167=>"001010111",
  56168=>"001100000",
  56169=>"110100101",
  56170=>"010100010",
  56171=>"000100100",
  56172=>"110000001",
  56173=>"001001011",
  56174=>"000011110",
  56175=>"011001011",
  56176=>"010110010",
  56177=>"000011110",
  56178=>"001100011",
  56179=>"010110111",
  56180=>"101000001",
  56181=>"000111111",
  56182=>"111001111",
  56183=>"110111100",
  56184=>"111101101",
  56185=>"001000101",
  56186=>"001100011",
  56187=>"111110001",
  56188=>"001110000",
  56189=>"101100000",
  56190=>"000001000",
  56191=>"000010100",
  56192=>"010010000",
  56193=>"000111101",
  56194=>"100010010",
  56195=>"111110101",
  56196=>"000110100",
  56197=>"011000011",
  56198=>"111111000",
  56199=>"111010001",
  56200=>"101011110",
  56201=>"101110111",
  56202=>"100011101",
  56203=>"110111010",
  56204=>"111011100",
  56205=>"011001011",
  56206=>"111011100",
  56207=>"100001111",
  56208=>"011011000",
  56209=>"000111110",
  56210=>"001001100",
  56211=>"001000001",
  56212=>"110100110",
  56213=>"110011101",
  56214=>"110100100",
  56215=>"111101101",
  56216=>"001000000",
  56217=>"000010011",
  56218=>"101000011",
  56219=>"111010000",
  56220=>"010000000",
  56221=>"100100000",
  56222=>"000011001",
  56223=>"010110000",
  56224=>"110111001",
  56225=>"000110110",
  56226=>"111000111",
  56227=>"110101011",
  56228=>"111111010",
  56229=>"110010011",
  56230=>"010010001",
  56231=>"010100010",
  56232=>"101001111",
  56233=>"011101000",
  56234=>"011000110",
  56235=>"100111100",
  56236=>"001101111",
  56237=>"011001111",
  56238=>"111011011",
  56239=>"101100100",
  56240=>"010000101",
  56241=>"000011110",
  56242=>"011111111",
  56243=>"100010010",
  56244=>"111001100",
  56245=>"111101011",
  56246=>"110111110",
  56247=>"000010100",
  56248=>"010100101",
  56249=>"101000010",
  56250=>"010000100",
  56251=>"110000111",
  56252=>"001010110",
  56253=>"000100010",
  56254=>"001001101",
  56255=>"001101101",
  56256=>"000100011",
  56257=>"010001111",
  56258=>"010110000",
  56259=>"001110010",
  56260=>"110111100",
  56261=>"011001010",
  56262=>"101010010",
  56263=>"011011001",
  56264=>"000010010",
  56265=>"100011000",
  56266=>"011011010",
  56267=>"101101010",
  56268=>"110011010",
  56269=>"001111111",
  56270=>"110101101",
  56271=>"101000010",
  56272=>"000000011",
  56273=>"100000111",
  56274=>"011010000",
  56275=>"000001101",
  56276=>"000101001",
  56277=>"110010111",
  56278=>"110111101",
  56279=>"011110010",
  56280=>"000110110",
  56281=>"010111011",
  56282=>"111111111",
  56283=>"010100011",
  56284=>"101000001",
  56285=>"010010101",
  56286=>"100010110",
  56287=>"001010101",
  56288=>"000110011",
  56289=>"011000111",
  56290=>"101001101",
  56291=>"001000001",
  56292=>"001000101",
  56293=>"100101100",
  56294=>"001000100",
  56295=>"010001100",
  56296=>"001000100",
  56297=>"110001001",
  56298=>"000001000",
  56299=>"101101111",
  56300=>"111101111",
  56301=>"010110100",
  56302=>"111101100",
  56303=>"100011011",
  56304=>"010110101",
  56305=>"000111100",
  56306=>"101111000",
  56307=>"110111000",
  56308=>"011011101",
  56309=>"001000000",
  56310=>"000101010",
  56311=>"101000111",
  56312=>"100110000",
  56313=>"101111110",
  56314=>"110000101",
  56315=>"000001110",
  56316=>"000100010",
  56317=>"001011011",
  56318=>"010001101",
  56319=>"010001101",
  56320=>"111010101",
  56321=>"111001101",
  56322=>"000000010",
  56323=>"001001101",
  56324=>"101111101",
  56325=>"011011110",
  56326=>"111101000",
  56327=>"010010001",
  56328=>"111101010",
  56329=>"000011110",
  56330=>"100101000",
  56331=>"001000110",
  56332=>"101101101",
  56333=>"100001001",
  56334=>"111011110",
  56335=>"010000000",
  56336=>"001100010",
  56337=>"100110011",
  56338=>"011010001",
  56339=>"111111100",
  56340=>"101000101",
  56341=>"101000010",
  56342=>"110101100",
  56343=>"101010100",
  56344=>"010001100",
  56345=>"001111100",
  56346=>"001001101",
  56347=>"111011000",
  56348=>"000000010",
  56349=>"111010100",
  56350=>"111010011",
  56351=>"100110001",
  56352=>"011110011",
  56353=>"001001010",
  56354=>"011011011",
  56355=>"110000101",
  56356=>"100000000",
  56357=>"011111000",
  56358=>"010010011",
  56359=>"100101010",
  56360=>"010101001",
  56361=>"010100101",
  56362=>"111110110",
  56363=>"011101011",
  56364=>"000000110",
  56365=>"110111101",
  56366=>"100111111",
  56367=>"011001101",
  56368=>"011011111",
  56369=>"001001001",
  56370=>"110111010",
  56371=>"000110100",
  56372=>"001010011",
  56373=>"110010011",
  56374=>"001000100",
  56375=>"011001001",
  56376=>"100100011",
  56377=>"111101111",
  56378=>"100011100",
  56379=>"110011010",
  56380=>"100011001",
  56381=>"010000011",
  56382=>"110111011",
  56383=>"100110100",
  56384=>"111010001",
  56385=>"011101000",
  56386=>"010001011",
  56387=>"011101010",
  56388=>"001001101",
  56389=>"000010110",
  56390=>"100010010",
  56391=>"000100010",
  56392=>"111111100",
  56393=>"010001101",
  56394=>"111011100",
  56395=>"010111101",
  56396=>"000000110",
  56397=>"001001011",
  56398=>"001100100",
  56399=>"010001111",
  56400=>"011110100",
  56401=>"011011111",
  56402=>"101011111",
  56403=>"011000110",
  56404=>"100111101",
  56405=>"010010010",
  56406=>"100100100",
  56407=>"000111011",
  56408=>"001111100",
  56409=>"000000111",
  56410=>"000100111",
  56411=>"101001111",
  56412=>"111110000",
  56413=>"111000010",
  56414=>"010000101",
  56415=>"100111011",
  56416=>"000001011",
  56417=>"111000001",
  56418=>"100011000",
  56419=>"011001010",
  56420=>"100110111",
  56421=>"000110110",
  56422=>"000110011",
  56423=>"100100010",
  56424=>"100100101",
  56425=>"011101011",
  56426=>"101011100",
  56427=>"110011000",
  56428=>"010010001",
  56429=>"001111010",
  56430=>"101000111",
  56431=>"110111111",
  56432=>"000101100",
  56433=>"000001000",
  56434=>"111101110",
  56435=>"010000011",
  56436=>"001110110",
  56437=>"101110001",
  56438=>"101010000",
  56439=>"010110001",
  56440=>"111101011",
  56441=>"110011110",
  56442=>"000101101",
  56443=>"010010100",
  56444=>"100101001",
  56445=>"101111000",
  56446=>"000100011",
  56447=>"111000000",
  56448=>"001111010",
  56449=>"001011101",
  56450=>"111111010",
  56451=>"010011110",
  56452=>"011101101",
  56453=>"011111010",
  56454=>"011100000",
  56455=>"100010101",
  56456=>"111111010",
  56457=>"000011100",
  56458=>"000001100",
  56459=>"001100110",
  56460=>"000001100",
  56461=>"111110010",
  56462=>"111111010",
  56463=>"111011111",
  56464=>"011111000",
  56465=>"101100010",
  56466=>"100101010",
  56467=>"001101100",
  56468=>"011111001",
  56469=>"111111100",
  56470=>"011111110",
  56471=>"110110011",
  56472=>"000011010",
  56473=>"010010110",
  56474=>"100011001",
  56475=>"010001011",
  56476=>"110011011",
  56477=>"110001000",
  56478=>"010101000",
  56479=>"111100101",
  56480=>"111111010",
  56481=>"110111101",
  56482=>"100101010",
  56483=>"110100100",
  56484=>"001101110",
  56485=>"110111111",
  56486=>"110110001",
  56487=>"111100011",
  56488=>"100001011",
  56489=>"000010001",
  56490=>"100010110",
  56491=>"000000100",
  56492=>"101011111",
  56493=>"001010010",
  56494=>"001000110",
  56495=>"010011100",
  56496=>"110000001",
  56497=>"000000010",
  56498=>"111110000",
  56499=>"110010110",
  56500=>"100111100",
  56501=>"010000000",
  56502=>"111111011",
  56503=>"000000101",
  56504=>"010101000",
  56505=>"011110110",
  56506=>"010101110",
  56507=>"000010110",
  56508=>"011101000",
  56509=>"000111001",
  56510=>"011011011",
  56511=>"000111110",
  56512=>"000010010",
  56513=>"101001100",
  56514=>"111101001",
  56515=>"111111110",
  56516=>"100110010",
  56517=>"010100000",
  56518=>"111110100",
  56519=>"001111110",
  56520=>"110001110",
  56521=>"010111000",
  56522=>"111110101",
  56523=>"001000000",
  56524=>"110011001",
  56525=>"010101001",
  56526=>"111001011",
  56527=>"000111000",
  56528=>"010111110",
  56529=>"110100111",
  56530=>"110101100",
  56531=>"001100001",
  56532=>"000011110",
  56533=>"100011000",
  56534=>"110000111",
  56535=>"110010101",
  56536=>"011001011",
  56537=>"010110110",
  56538=>"100111001",
  56539=>"101111000",
  56540=>"011001010",
  56541=>"001100111",
  56542=>"101010100",
  56543=>"000001011",
  56544=>"111000110",
  56545=>"111111111",
  56546=>"001000010",
  56547=>"000110111",
  56548=>"011010011",
  56549=>"100000000",
  56550=>"111110000",
  56551=>"001101010",
  56552=>"111001011",
  56553=>"000111011",
  56554=>"000000101",
  56555=>"010101000",
  56556=>"000110000",
  56557=>"010010010",
  56558=>"011000010",
  56559=>"010010010",
  56560=>"100000000",
  56561=>"001010011",
  56562=>"100100001",
  56563=>"111101001",
  56564=>"110110010",
  56565=>"010100101",
  56566=>"001110111",
  56567=>"000011001",
  56568=>"101100101",
  56569=>"001000000",
  56570=>"111101111",
  56571=>"111100000",
  56572=>"101101000",
  56573=>"110101110",
  56574=>"110000101",
  56575=>"001100000",
  56576=>"011001000",
  56577=>"000011100",
  56578=>"001100111",
  56579=>"100010000",
  56580=>"111001001",
  56581=>"000000001",
  56582=>"010101011",
  56583=>"011110010",
  56584=>"011000000",
  56585=>"001010100",
  56586=>"011001110",
  56587=>"000110010",
  56588=>"111000100",
  56589=>"001010010",
  56590=>"010110100",
  56591=>"001111010",
  56592=>"110100001",
  56593=>"111010000",
  56594=>"101101111",
  56595=>"111010110",
  56596=>"011010110",
  56597=>"010010001",
  56598=>"101111100",
  56599=>"001001100",
  56600=>"000001100",
  56601=>"011110011",
  56602=>"110010000",
  56603=>"001001110",
  56604=>"001101110",
  56605=>"000100001",
  56606=>"010110000",
  56607=>"011001000",
  56608=>"011000010",
  56609=>"100001111",
  56610=>"011110101",
  56611=>"011111111",
  56612=>"101011101",
  56613=>"110000001",
  56614=>"110011101",
  56615=>"011100111",
  56616=>"010110000",
  56617=>"101111110",
  56618=>"000000001",
  56619=>"001001001",
  56620=>"111011100",
  56621=>"001110000",
  56622=>"100000010",
  56623=>"101010110",
  56624=>"011101110",
  56625=>"111111110",
  56626=>"100000000",
  56627=>"101011111",
  56628=>"100000111",
  56629=>"101001011",
  56630=>"100011011",
  56631=>"110001001",
  56632=>"001011100",
  56633=>"100110100",
  56634=>"010100011",
  56635=>"101000011",
  56636=>"110000010",
  56637=>"100011010",
  56638=>"110110101",
  56639=>"100101101",
  56640=>"010001111",
  56641=>"010100001",
  56642=>"000110111",
  56643=>"110110001",
  56644=>"110000110",
  56645=>"101111101",
  56646=>"101010110",
  56647=>"110000011",
  56648=>"010111100",
  56649=>"000011101",
  56650=>"010011110",
  56651=>"001111010",
  56652=>"101010111",
  56653=>"010110111",
  56654=>"011011011",
  56655=>"110010111",
  56656=>"100110001",
  56657=>"001100010",
  56658=>"101001001",
  56659=>"101011111",
  56660=>"110010001",
  56661=>"001101001",
  56662=>"000100001",
  56663=>"001001011",
  56664=>"000001000",
  56665=>"010111011",
  56666=>"000011110",
  56667=>"010100111",
  56668=>"101101001",
  56669=>"100100000",
  56670=>"001110101",
  56671=>"011110110",
  56672=>"001011010",
  56673=>"001011100",
  56674=>"001001101",
  56675=>"101011111",
  56676=>"100101000",
  56677=>"001001101",
  56678=>"100100100",
  56679=>"111010101",
  56680=>"011111000",
  56681=>"100100010",
  56682=>"111111100",
  56683=>"010100110",
  56684=>"000100100",
  56685=>"110101011",
  56686=>"011010101",
  56687=>"001010000",
  56688=>"000110110",
  56689=>"100001101",
  56690=>"100011010",
  56691=>"010001000",
  56692=>"001001010",
  56693=>"011101000",
  56694=>"110111110",
  56695=>"101101110",
  56696=>"111110000",
  56697=>"111111000",
  56698=>"000010011",
  56699=>"101101100",
  56700=>"110000001",
  56701=>"101001110",
  56702=>"000111011",
  56703=>"100001100",
  56704=>"100001110",
  56705=>"010010000",
  56706=>"101101111",
  56707=>"000100001",
  56708=>"000110101",
  56709=>"000000111",
  56710=>"110101001",
  56711=>"011110010",
  56712=>"110010100",
  56713=>"100111110",
  56714=>"010000010",
  56715=>"000010010",
  56716=>"110011000",
  56717=>"101101011",
  56718=>"001110001",
  56719=>"011100010",
  56720=>"110001001",
  56721=>"110100001",
  56722=>"010000101",
  56723=>"000110110",
  56724=>"000011111",
  56725=>"110100111",
  56726=>"101001111",
  56727=>"101011001",
  56728=>"111000111",
  56729=>"000001111",
  56730=>"111110111",
  56731=>"001111001",
  56732=>"111000111",
  56733=>"101100010",
  56734=>"001000100",
  56735=>"010000110",
  56736=>"011100010",
  56737=>"010010000",
  56738=>"111111010",
  56739=>"000001011",
  56740=>"011100010",
  56741=>"100101111",
  56742=>"101000110",
  56743=>"000010010",
  56744=>"110010000",
  56745=>"100100011",
  56746=>"001001110",
  56747=>"000001001",
  56748=>"011000110",
  56749=>"010100000",
  56750=>"000111101",
  56751=>"110111101",
  56752=>"100000100",
  56753=>"010001010",
  56754=>"111111011",
  56755=>"001111110",
  56756=>"111010101",
  56757=>"101000111",
  56758=>"001101000",
  56759=>"001000110",
  56760=>"010101000",
  56761=>"110110100",
  56762=>"011111101",
  56763=>"011000110",
  56764=>"100110100",
  56765=>"101000100",
  56766=>"110110000",
  56767=>"111111001",
  56768=>"001001000",
  56769=>"110111001",
  56770=>"001000000",
  56771=>"000111110",
  56772=>"111101101",
  56773=>"101000101",
  56774=>"001110010",
  56775=>"001011101",
  56776=>"110111110",
  56777=>"010101110",
  56778=>"011110001",
  56779=>"010001010",
  56780=>"110110100",
  56781=>"010101001",
  56782=>"101100101",
  56783=>"100011110",
  56784=>"001111101",
  56785=>"110110111",
  56786=>"001110000",
  56787=>"011100011",
  56788=>"110000100",
  56789=>"010110110",
  56790=>"010110000",
  56791=>"111101111",
  56792=>"100011111",
  56793=>"010000111",
  56794=>"100011001",
  56795=>"110100111",
  56796=>"000001011",
  56797=>"011010111",
  56798=>"010011100",
  56799=>"010100101",
  56800=>"111100011",
  56801=>"101011010",
  56802=>"010011000",
  56803=>"111111011",
  56804=>"010000110",
  56805=>"000101111",
  56806=>"101000110",
  56807=>"010100001",
  56808=>"100111101",
  56809=>"100111011",
  56810=>"010110010",
  56811=>"111101101",
  56812=>"001100010",
  56813=>"011011110",
  56814=>"111000101",
  56815=>"100000011",
  56816=>"000001011",
  56817=>"101000110",
  56818=>"011001010",
  56819=>"010110000",
  56820=>"001001000",
  56821=>"110000000",
  56822=>"000111111",
  56823=>"001000110",
  56824=>"101111001",
  56825=>"011100110",
  56826=>"001000000",
  56827=>"110000110",
  56828=>"001110100",
  56829=>"101011000",
  56830=>"111100100",
  56831=>"110110111",
  56832=>"100100111",
  56833=>"101010000",
  56834=>"010110001",
  56835=>"000011011",
  56836=>"000001001",
  56837=>"001101101",
  56838=>"100110000",
  56839=>"100000000",
  56840=>"100110001",
  56841=>"010011010",
  56842=>"111110000",
  56843=>"001100111",
  56844=>"000100100",
  56845=>"100010001",
  56846=>"000011100",
  56847=>"110110010",
  56848=>"111101101",
  56849=>"110100101",
  56850=>"111111111",
  56851=>"010011000",
  56852=>"000100010",
  56853=>"010010000",
  56854=>"001100111",
  56855=>"100100010",
  56856=>"100111000",
  56857=>"001111000",
  56858=>"000010010",
  56859=>"000110101",
  56860=>"100111110",
  56861=>"010101111",
  56862=>"111001110",
  56863=>"110101101",
  56864=>"011001101",
  56865=>"010010101",
  56866=>"010001010",
  56867=>"011100101",
  56868=>"001011111",
  56869=>"101000000",
  56870=>"010110110",
  56871=>"001011110",
  56872=>"101001100",
  56873=>"111010100",
  56874=>"101111010",
  56875=>"100010101",
  56876=>"111111001",
  56877=>"111100001",
  56878=>"000100100",
  56879=>"010110001",
  56880=>"011100101",
  56881=>"101011000",
  56882=>"110110001",
  56883=>"011110111",
  56884=>"001110101",
  56885=>"110100000",
  56886=>"001000101",
  56887=>"101001101",
  56888=>"011000000",
  56889=>"000101011",
  56890=>"110010111",
  56891=>"011011100",
  56892=>"100010101",
  56893=>"010000000",
  56894=>"111100000",
  56895=>"100101000",
  56896=>"000000010",
  56897=>"000111001",
  56898=>"110110100",
  56899=>"101011110",
  56900=>"011000110",
  56901=>"000111000",
  56902=>"011110010",
  56903=>"111011001",
  56904=>"011010111",
  56905=>"001101110",
  56906=>"100111100",
  56907=>"101000000",
  56908=>"111001101",
  56909=>"011111111",
  56910=>"111100110",
  56911=>"001101001",
  56912=>"100110001",
  56913=>"001010011",
  56914=>"000010001",
  56915=>"010000000",
  56916=>"111100010",
  56917=>"111010000",
  56918=>"101100101",
  56919=>"000111100",
  56920=>"011000011",
  56921=>"100101000",
  56922=>"110101111",
  56923=>"110111101",
  56924=>"100111111",
  56925=>"011110000",
  56926=>"100101001",
  56927=>"011001111",
  56928=>"010110010",
  56929=>"000001001",
  56930=>"011100001",
  56931=>"010100010",
  56932=>"000000110",
  56933=>"100000000",
  56934=>"110000100",
  56935=>"100111100",
  56936=>"001110101",
  56937=>"110101000",
  56938=>"010100000",
  56939=>"000101100",
  56940=>"101111110",
  56941=>"101110111",
  56942=>"011101010",
  56943=>"100000010",
  56944=>"110011110",
  56945=>"111100110",
  56946=>"111100010",
  56947=>"000010100",
  56948=>"011010110",
  56949=>"111111100",
  56950=>"111010001",
  56951=>"110111000",
  56952=>"110010010",
  56953=>"100111101",
  56954=>"100110101",
  56955=>"110011110",
  56956=>"011011101",
  56957=>"101000010",
  56958=>"011101100",
  56959=>"011111000",
  56960=>"011100110",
  56961=>"101010101",
  56962=>"110100111",
  56963=>"010101100",
  56964=>"110010110",
  56965=>"010000010",
  56966=>"001011011",
  56967=>"011001000",
  56968=>"100110011",
  56969=>"111110100",
  56970=>"001000111",
  56971=>"000011110",
  56972=>"100011001",
  56973=>"000000101",
  56974=>"000011111",
  56975=>"001001011",
  56976=>"010000001",
  56977=>"101010111",
  56978=>"001100000",
  56979=>"010101000",
  56980=>"010000010",
  56981=>"001011110",
  56982=>"101000001",
  56983=>"001011000",
  56984=>"101110111",
  56985=>"110100001",
  56986=>"001111110",
  56987=>"101100100",
  56988=>"011000111",
  56989=>"101110001",
  56990=>"101011011",
  56991=>"001101110",
  56992=>"110100011",
  56993=>"101010000",
  56994=>"100111000",
  56995=>"010111111",
  56996=>"111111001",
  56997=>"101110111",
  56998=>"110110100",
  56999=>"011011100",
  57000=>"010000000",
  57001=>"110100101",
  57002=>"010000100",
  57003=>"000110001",
  57004=>"110000001",
  57005=>"111111101",
  57006=>"101111011",
  57007=>"110110001",
  57008=>"100111101",
  57009=>"001100001",
  57010=>"100100111",
  57011=>"010000000",
  57012=>"011010010",
  57013=>"000111001",
  57014=>"011001000",
  57015=>"110010110",
  57016=>"001001011",
  57017=>"111101101",
  57018=>"110101101",
  57019=>"000000111",
  57020=>"111111011",
  57021=>"000111001",
  57022=>"100001000",
  57023=>"111101000",
  57024=>"000110100",
  57025=>"000001110",
  57026=>"101000010",
  57027=>"001110101",
  57028=>"001010101",
  57029=>"000110101",
  57030=>"000001100",
  57031=>"110001000",
  57032=>"111011111",
  57033=>"001110011",
  57034=>"100010100",
  57035=>"000101001",
  57036=>"011101110",
  57037=>"110111100",
  57038=>"110100111",
  57039=>"000000110",
  57040=>"111111101",
  57041=>"101111011",
  57042=>"101011110",
  57043=>"000101110",
  57044=>"010000110",
  57045=>"001101000",
  57046=>"001011001",
  57047=>"111010001",
  57048=>"111001100",
  57049=>"011110101",
  57050=>"011101011",
  57051=>"101001001",
  57052=>"100001110",
  57053=>"001100000",
  57054=>"011100110",
  57055=>"010010011",
  57056=>"001100111",
  57057=>"111110110",
  57058=>"100011011",
  57059=>"110110111",
  57060=>"100110010",
  57061=>"001100101",
  57062=>"111010001",
  57063=>"111011000",
  57064=>"111010110",
  57065=>"011100001",
  57066=>"110100010",
  57067=>"100000101",
  57068=>"101000100",
  57069=>"010000000",
  57070=>"000000101",
  57071=>"100101000",
  57072=>"111110011",
  57073=>"011100011",
  57074=>"000000111",
  57075=>"000111011",
  57076=>"110000001",
  57077=>"110001001",
  57078=>"101010110",
  57079=>"101011100",
  57080=>"001111001",
  57081=>"100100001",
  57082=>"101111011",
  57083=>"101100001",
  57084=>"010100110",
  57085=>"001010100",
  57086=>"000001100",
  57087=>"100101110",
  57088=>"000001000",
  57089=>"011001110",
  57090=>"100101010",
  57091=>"000010101",
  57092=>"010000011",
  57093=>"100001011",
  57094=>"001000110",
  57095=>"001000011",
  57096=>"010111000",
  57097=>"111010010",
  57098=>"011110111",
  57099=>"001101101",
  57100=>"101100111",
  57101=>"111010010",
  57102=>"000100011",
  57103=>"010110001",
  57104=>"000011001",
  57105=>"100011000",
  57106=>"100001010",
  57107=>"001110000",
  57108=>"110011111",
  57109=>"001011001",
  57110=>"110000111",
  57111=>"010011010",
  57112=>"110100000",
  57113=>"110010010",
  57114=>"111111111",
  57115=>"101111001",
  57116=>"000111001",
  57117=>"000000100",
  57118=>"101110001",
  57119=>"010110010",
  57120=>"011111101",
  57121=>"110111101",
  57122=>"111111100",
  57123=>"010011111",
  57124=>"101011000",
  57125=>"001101110",
  57126=>"000111101",
  57127=>"111111110",
  57128=>"001110110",
  57129=>"000111000",
  57130=>"000100010",
  57131=>"001110111",
  57132=>"110010000",
  57133=>"111010000",
  57134=>"000011111",
  57135=>"001100101",
  57136=>"000011111",
  57137=>"010110010",
  57138=>"010111101",
  57139=>"111100101",
  57140=>"100001000",
  57141=>"001100001",
  57142=>"110110000",
  57143=>"100000110",
  57144=>"001110001",
  57145=>"001001010",
  57146=>"100111001",
  57147=>"001111101",
  57148=>"101010101",
  57149=>"000101011",
  57150=>"100010010",
  57151=>"000100000",
  57152=>"000111111",
  57153=>"011011101",
  57154=>"100101011",
  57155=>"001100000",
  57156=>"111100000",
  57157=>"010111011",
  57158=>"111000001",
  57159=>"001101011",
  57160=>"100100001",
  57161=>"100100100",
  57162=>"111011001",
  57163=>"000100011",
  57164=>"100011101",
  57165=>"110011011",
  57166=>"111111011",
  57167=>"001111000",
  57168=>"111011000",
  57169=>"011101001",
  57170=>"011111111",
  57171=>"001101110",
  57172=>"001100111",
  57173=>"001100101",
  57174=>"100001000",
  57175=>"110001011",
  57176=>"010101100",
  57177=>"111111110",
  57178=>"101010001",
  57179=>"100010110",
  57180=>"100000000",
  57181=>"011111101",
  57182=>"001100010",
  57183=>"011010111",
  57184=>"101001101",
  57185=>"001110001",
  57186=>"101110001",
  57187=>"011011001",
  57188=>"110111110",
  57189=>"010100001",
  57190=>"111111101",
  57191=>"001001111",
  57192=>"010010110",
  57193=>"011101111",
  57194=>"101001011",
  57195=>"100000011",
  57196=>"110011110",
  57197=>"011011100",
  57198=>"011000001",
  57199=>"111001101",
  57200=>"000000011",
  57201=>"001011011",
  57202=>"010100010",
  57203=>"111011110",
  57204=>"111010111",
  57205=>"111100011",
  57206=>"000110100",
  57207=>"011110000",
  57208=>"010010110",
  57209=>"110000010",
  57210=>"001011010",
  57211=>"010110110",
  57212=>"011101111",
  57213=>"001100010",
  57214=>"011011100",
  57215=>"000001010",
  57216=>"110111010",
  57217=>"111000110",
  57218=>"110100100",
  57219=>"110111001",
  57220=>"110100100",
  57221=>"001010110",
  57222=>"110001100",
  57223=>"000000110",
  57224=>"011110101",
  57225=>"011010010",
  57226=>"001111001",
  57227=>"001110000",
  57228=>"100100111",
  57229=>"111000110",
  57230=>"111101011",
  57231=>"000000011",
  57232=>"000011100",
  57233=>"101111101",
  57234=>"001110010",
  57235=>"010000000",
  57236=>"001101000",
  57237=>"011101111",
  57238=>"100010010",
  57239=>"101010110",
  57240=>"000100000",
  57241=>"010110011",
  57242=>"010111010",
  57243=>"100110001",
  57244=>"001011110",
  57245=>"111001000",
  57246=>"111100101",
  57247=>"001100100",
  57248=>"001001000",
  57249=>"101110111",
  57250=>"111011010",
  57251=>"101100111",
  57252=>"101111101",
  57253=>"011000010",
  57254=>"111100001",
  57255=>"111111110",
  57256=>"110011110",
  57257=>"101101111",
  57258=>"111000110",
  57259=>"101010010",
  57260=>"010111111",
  57261=>"100111000",
  57262=>"100110100",
  57263=>"100010101",
  57264=>"010110100",
  57265=>"111101001",
  57266=>"101010000",
  57267=>"000110001",
  57268=>"100001101",
  57269=>"000000000",
  57270=>"101111100",
  57271=>"011100110",
  57272=>"100111111",
  57273=>"011000111",
  57274=>"010111000",
  57275=>"101011100",
  57276=>"001001100",
  57277=>"100011100",
  57278=>"111110110",
  57279=>"000101110",
  57280=>"001111010",
  57281=>"010100101",
  57282=>"111100101",
  57283=>"011100011",
  57284=>"100011000",
  57285=>"110101100",
  57286=>"110101011",
  57287=>"101010111",
  57288=>"000000110",
  57289=>"001111110",
  57290=>"010000100",
  57291=>"110000111",
  57292=>"110100010",
  57293=>"001000011",
  57294=>"010000111",
  57295=>"011110110",
  57296=>"000000000",
  57297=>"011000111",
  57298=>"101000101",
  57299=>"001110101",
  57300=>"000011011",
  57301=>"000010001",
  57302=>"110111110",
  57303=>"101111110",
  57304=>"010010111",
  57305=>"001111011",
  57306=>"111001110",
  57307=>"100010011",
  57308=>"101101101",
  57309=>"010001111",
  57310=>"000100100",
  57311=>"101101010",
  57312=>"000100000",
  57313=>"000011101",
  57314=>"001001111",
  57315=>"110000101",
  57316=>"011111110",
  57317=>"000000010",
  57318=>"110010110",
  57319=>"010011001",
  57320=>"000011110",
  57321=>"001111000",
  57322=>"000111111",
  57323=>"010001010",
  57324=>"000010011",
  57325=>"111000111",
  57326=>"000010000",
  57327=>"111000110",
  57328=>"011111111",
  57329=>"110000100",
  57330=>"111000110",
  57331=>"001111100",
  57332=>"011011001",
  57333=>"110011110",
  57334=>"011010101",
  57335=>"111001000",
  57336=>"100100111",
  57337=>"011000010",
  57338=>"011001011",
  57339=>"111000101",
  57340=>"110101110",
  57341=>"110001110",
  57342=>"011010111",
  57343=>"000000100",
  57344=>"010111010",
  57345=>"101111110",
  57346=>"110101000",
  57347=>"011000100",
  57348=>"001100100",
  57349=>"111010110",
  57350=>"111111100",
  57351=>"011001000",
  57352=>"001011011",
  57353=>"100010110",
  57354=>"111111111",
  57355=>"110000011",
  57356=>"111000001",
  57357=>"101110000",
  57358=>"100101100",
  57359=>"101100011",
  57360=>"001001001",
  57361=>"011000110",
  57362=>"111010000",
  57363=>"110100011",
  57364=>"111111101",
  57365=>"010000011",
  57366=>"010111100",
  57367=>"011010011",
  57368=>"010110000",
  57369=>"000000001",
  57370=>"010001100",
  57371=>"010011011",
  57372=>"001111100",
  57373=>"110010011",
  57374=>"010111111",
  57375=>"110001001",
  57376=>"101110111",
  57377=>"001100011",
  57378=>"100000110",
  57379=>"101001000",
  57380=>"000001101",
  57381=>"100110001",
  57382=>"001101100",
  57383=>"111011111",
  57384=>"011100011",
  57385=>"000111001",
  57386=>"001010000",
  57387=>"110111100",
  57388=>"101111111",
  57389=>"011100110",
  57390=>"010111100",
  57391=>"111100111",
  57392=>"110010010",
  57393=>"111101010",
  57394=>"010011101",
  57395=>"100110010",
  57396=>"000101111",
  57397=>"001101110",
  57398=>"111111000",
  57399=>"100110101",
  57400=>"101000000",
  57401=>"010010001",
  57402=>"100010000",
  57403=>"100110001",
  57404=>"010111010",
  57405=>"010011011",
  57406=>"000011100",
  57407=>"110000010",
  57408=>"001100000",
  57409=>"001011001",
  57410=>"000010100",
  57411=>"101110000",
  57412=>"111100100",
  57413=>"110111100",
  57414=>"111001110",
  57415=>"011010000",
  57416=>"001111010",
  57417=>"101000100",
  57418=>"000000011",
  57419=>"100010100",
  57420=>"001110111",
  57421=>"100001011",
  57422=>"001111110",
  57423=>"010100001",
  57424=>"111011010",
  57425=>"110100011",
  57426=>"111101011",
  57427=>"011011100",
  57428=>"001101101",
  57429=>"001100100",
  57430=>"101001001",
  57431=>"001110001",
  57432=>"000101101",
  57433=>"100110011",
  57434=>"000100011",
  57435=>"101110111",
  57436=>"000001000",
  57437=>"110001000",
  57438=>"111000001",
  57439=>"000010011",
  57440=>"100011000",
  57441=>"000010000",
  57442=>"001000111",
  57443=>"101101101",
  57444=>"111111110",
  57445=>"010100101",
  57446=>"111011001",
  57447=>"010100101",
  57448=>"011101111",
  57449=>"010001011",
  57450=>"111111110",
  57451=>"100100000",
  57452=>"000111011",
  57453=>"110110110",
  57454=>"011110001",
  57455=>"011001000",
  57456=>"000100010",
  57457=>"101010001",
  57458=>"110010010",
  57459=>"000101001",
  57460=>"110111110",
  57461=>"011100010",
  57462=>"111110011",
  57463=>"111011100",
  57464=>"100101100",
  57465=>"001010010",
  57466=>"010101111",
  57467=>"001101100",
  57468=>"110111010",
  57469=>"001101100",
  57470=>"011111100",
  57471=>"100111101",
  57472=>"011011001",
  57473=>"010001101",
  57474=>"100110110",
  57475=>"111111010",
  57476=>"101111100",
  57477=>"100010010",
  57478=>"100101010",
  57479=>"110010010",
  57480=>"110100010",
  57481=>"111011010",
  57482=>"111011010",
  57483=>"110111010",
  57484=>"011011110",
  57485=>"101001100",
  57486=>"010100001",
  57487=>"100110101",
  57488=>"001110010",
  57489=>"010100001",
  57490=>"000010010",
  57491=>"000010001",
  57492=>"010010110",
  57493=>"110100100",
  57494=>"010001000",
  57495=>"100011111",
  57496=>"111011101",
  57497=>"010111010",
  57498=>"101010011",
  57499=>"011010111",
  57500=>"011100010",
  57501=>"100011010",
  57502=>"100010111",
  57503=>"001101001",
  57504=>"001001100",
  57505=>"010101010",
  57506=>"011110000",
  57507=>"111011100",
  57508=>"010100001",
  57509=>"000001000",
  57510=>"011001110",
  57511=>"101010001",
  57512=>"011111100",
  57513=>"110001000",
  57514=>"101000101",
  57515=>"010111011",
  57516=>"011000010",
  57517=>"011001000",
  57518=>"000111001",
  57519=>"100001011",
  57520=>"000101000",
  57521=>"111110111",
  57522=>"111001110",
  57523=>"011001010",
  57524=>"101110101",
  57525=>"000010000",
  57526=>"110111000",
  57527=>"011000110",
  57528=>"100111011",
  57529=>"001011101",
  57530=>"111100100",
  57531=>"101110001",
  57532=>"001101111",
  57533=>"011101111",
  57534=>"110110100",
  57535=>"011010011",
  57536=>"101110101",
  57537=>"010000001",
  57538=>"001001111",
  57539=>"100000111",
  57540=>"001100011",
  57541=>"010100000",
  57542=>"001100100",
  57543=>"010111100",
  57544=>"001101111",
  57545=>"001011000",
  57546=>"000000100",
  57547=>"110110111",
  57548=>"011010101",
  57549=>"000101110",
  57550=>"011001011",
  57551=>"001110001",
  57552=>"010010110",
  57553=>"000010100",
  57554=>"011110001",
  57555=>"011000010",
  57556=>"100011111",
  57557=>"111110010",
  57558=>"001011001",
  57559=>"110000000",
  57560=>"011000000",
  57561=>"110101110",
  57562=>"001100101",
  57563=>"010110101",
  57564=>"011000100",
  57565=>"011111001",
  57566=>"100011001",
  57567=>"110111001",
  57568=>"101011000",
  57569=>"011001001",
  57570=>"010001011",
  57571=>"110110010",
  57572=>"010110011",
  57573=>"001110001",
  57574=>"001110010",
  57575=>"101111100",
  57576=>"100101101",
  57577=>"001011101",
  57578=>"010001101",
  57579=>"111010011",
  57580=>"001110011",
  57581=>"100011111",
  57582=>"111001001",
  57583=>"000011100",
  57584=>"010100010",
  57585=>"011100111",
  57586=>"110001010",
  57587=>"001001000",
  57588=>"110111100",
  57589=>"011111101",
  57590=>"101110111",
  57591=>"001100101",
  57592=>"111100110",
  57593=>"110001000",
  57594=>"010000000",
  57595=>"001101001",
  57596=>"111100101",
  57597=>"101111100",
  57598=>"001111110",
  57599=>"000111001",
  57600=>"000001110",
  57601=>"110111010",
  57602=>"100110001",
  57603=>"111101001",
  57604=>"101010110",
  57605=>"000111110",
  57606=>"110111010",
  57607=>"011011110",
  57608=>"010110110",
  57609=>"000010101",
  57610=>"111110010",
  57611=>"100010110",
  57612=>"001011001",
  57613=>"100011011",
  57614=>"011110100",
  57615=>"001000000",
  57616=>"110000110",
  57617=>"110000011",
  57618=>"000000010",
  57619=>"101100011",
  57620=>"100111000",
  57621=>"001110000",
  57622=>"010101101",
  57623=>"000110110",
  57624=>"111010110",
  57625=>"101010111",
  57626=>"001001011",
  57627=>"111011111",
  57628=>"110100010",
  57629=>"101010110",
  57630=>"100000011",
  57631=>"001010011",
  57632=>"001011011",
  57633=>"011101110",
  57634=>"110101000",
  57635=>"110010100",
  57636=>"100001010",
  57637=>"001010110",
  57638=>"110000010",
  57639=>"010110100",
  57640=>"000111001",
  57641=>"110011110",
  57642=>"010010000",
  57643=>"100010111",
  57644=>"000010010",
  57645=>"001001110",
  57646=>"101111001",
  57647=>"010000101",
  57648=>"101101110",
  57649=>"101101101",
  57650=>"001110000",
  57651=>"011011110",
  57652=>"111100100",
  57653=>"111001011",
  57654=>"101001111",
  57655=>"000111010",
  57656=>"000101011",
  57657=>"111101100",
  57658=>"011101111",
  57659=>"100111000",
  57660=>"001001011",
  57661=>"100010101",
  57662=>"010011110",
  57663=>"101000101",
  57664=>"010011110",
  57665=>"110000111",
  57666=>"011101100",
  57667=>"100111110",
  57668=>"001010101",
  57669=>"110101100",
  57670=>"011010101",
  57671=>"100000011",
  57672=>"111001101",
  57673=>"110000010",
  57674=>"010111111",
  57675=>"101110101",
  57676=>"100010001",
  57677=>"000000101",
  57678=>"110101000",
  57679=>"111101001",
  57680=>"011011000",
  57681=>"000110011",
  57682=>"000000000",
  57683=>"001111111",
  57684=>"111000000",
  57685=>"001000100",
  57686=>"010011010",
  57687=>"111001000",
  57688=>"000101000",
  57689=>"100011011",
  57690=>"110011010",
  57691=>"100110000",
  57692=>"011110011",
  57693=>"001101000",
  57694=>"101100001",
  57695=>"100100101",
  57696=>"100100001",
  57697=>"101110110",
  57698=>"000111010",
  57699=>"010101001",
  57700=>"110010110",
  57701=>"011010110",
  57702=>"011100010",
  57703=>"101110110",
  57704=>"111011000",
  57705=>"010000010",
  57706=>"110010100",
  57707=>"001001001",
  57708=>"101001111",
  57709=>"100000001",
  57710=>"010111001",
  57711=>"001000111",
  57712=>"000001001",
  57713=>"110100010",
  57714=>"100011011",
  57715=>"000111011",
  57716=>"101100111",
  57717=>"100110001",
  57718=>"101111001",
  57719=>"111111001",
  57720=>"101011110",
  57721=>"011010100",
  57722=>"101101001",
  57723=>"110110100",
  57724=>"000101101",
  57725=>"100010000",
  57726=>"101101101",
  57727=>"111001000",
  57728=>"001111111",
  57729=>"000011001",
  57730=>"000100101",
  57731=>"001001001",
  57732=>"111001010",
  57733=>"001001010",
  57734=>"100010001",
  57735=>"000101010",
  57736=>"001101001",
  57737=>"011001100",
  57738=>"011011010",
  57739=>"001000110",
  57740=>"000000100",
  57741=>"101010010",
  57742=>"110000101",
  57743=>"110011010",
  57744=>"110011111",
  57745=>"001111101",
  57746=>"011111000",
  57747=>"100101001",
  57748=>"101011101",
  57749=>"001000110",
  57750=>"000110011",
  57751=>"000100001",
  57752=>"111000000",
  57753=>"101111010",
  57754=>"110110110",
  57755=>"010110101",
  57756=>"100000110",
  57757=>"000000011",
  57758=>"011110010",
  57759=>"110010110",
  57760=>"111010010",
  57761=>"000011101",
  57762=>"000100000",
  57763=>"010010000",
  57764=>"101101010",
  57765=>"110101011",
  57766=>"000100010",
  57767=>"100111111",
  57768=>"011110111",
  57769=>"010000100",
  57770=>"001000001",
  57771=>"110100011",
  57772=>"011100010",
  57773=>"100101010",
  57774=>"010010111",
  57775=>"000000111",
  57776=>"110011100",
  57777=>"011101011",
  57778=>"001000100",
  57779=>"110111110",
  57780=>"011000011",
  57781=>"110001011",
  57782=>"000000010",
  57783=>"000111101",
  57784=>"001110101",
  57785=>"000010101",
  57786=>"100011010",
  57787=>"110110000",
  57788=>"000011010",
  57789=>"110011011",
  57790=>"011001100",
  57791=>"001000101",
  57792=>"011100100",
  57793=>"111010101",
  57794=>"110000011",
  57795=>"001011111",
  57796=>"010110011",
  57797=>"100100110",
  57798=>"101011011",
  57799=>"110111100",
  57800=>"101111111",
  57801=>"101011010",
  57802=>"001111111",
  57803=>"101101111",
  57804=>"111111010",
  57805=>"010100100",
  57806=>"011100011",
  57807=>"001000100",
  57808=>"010100110",
  57809=>"111110101",
  57810=>"011111110",
  57811=>"101110001",
  57812=>"010111010",
  57813=>"011010110",
  57814=>"101000100",
  57815=>"001100001",
  57816=>"011101000",
  57817=>"000111101",
  57818=>"011001010",
  57819=>"001000110",
  57820=>"001111101",
  57821=>"011100001",
  57822=>"011111000",
  57823=>"100100000",
  57824=>"001010100",
  57825=>"001011101",
  57826=>"011101110",
  57827=>"000011110",
  57828=>"101011011",
  57829=>"111000011",
  57830=>"010011100",
  57831=>"010011101",
  57832=>"101000010",
  57833=>"110000101",
  57834=>"000101000",
  57835=>"101101010",
  57836=>"111001011",
  57837=>"010010000",
  57838=>"011100011",
  57839=>"000010111",
  57840=>"100011010",
  57841=>"011010011",
  57842=>"111010111",
  57843=>"001100001",
  57844=>"100010000",
  57845=>"101100000",
  57846=>"000001001",
  57847=>"011100011",
  57848=>"110111111",
  57849=>"000011010",
  57850=>"100101100",
  57851=>"111101100",
  57852=>"011110001",
  57853=>"111111000",
  57854=>"011011011",
  57855=>"000001001",
  57856=>"000111011",
  57857=>"011011010",
  57858=>"101101100",
  57859=>"000010010",
  57860=>"111010001",
  57861=>"111100010",
  57862=>"011000101",
  57863=>"111111010",
  57864=>"111110001",
  57865=>"110111101",
  57866=>"100101010",
  57867=>"100001110",
  57868=>"001010110",
  57869=>"101011110",
  57870=>"010001011",
  57871=>"001110111",
  57872=>"111001011",
  57873=>"000000111",
  57874=>"000000100",
  57875=>"111110101",
  57876=>"000000001",
  57877=>"100000011",
  57878=>"000000001",
  57879=>"110010110",
  57880=>"101011100",
  57881=>"001000100",
  57882=>"100100100",
  57883=>"110010000",
  57884=>"000001010",
  57885=>"001000110",
  57886=>"100100110",
  57887=>"010100101",
  57888=>"010000001",
  57889=>"010011110",
  57890=>"000010100",
  57891=>"111100001",
  57892=>"111011101",
  57893=>"101000010",
  57894=>"000100000",
  57895=>"000011011",
  57896=>"011100000",
  57897=>"010001011",
  57898=>"101111000",
  57899=>"111110001",
  57900=>"010110100",
  57901=>"110001001",
  57902=>"001111100",
  57903=>"111101111",
  57904=>"111000010",
  57905=>"110101100",
  57906=>"011100000",
  57907=>"110000010",
  57908=>"011111000",
  57909=>"110010100",
  57910=>"000101110",
  57911=>"101011011",
  57912=>"010011011",
  57913=>"110011010",
  57914=>"000100011",
  57915=>"010110100",
  57916=>"101100100",
  57917=>"001110100",
  57918=>"010101011",
  57919=>"111110100",
  57920=>"101110110",
  57921=>"101010010",
  57922=>"010011000",
  57923=>"101101100",
  57924=>"001000101",
  57925=>"010100100",
  57926=>"001010110",
  57927=>"001101110",
  57928=>"111100010",
  57929=>"000101010",
  57930=>"000110010",
  57931=>"001001111",
  57932=>"111101110",
  57933=>"001110000",
  57934=>"011110100",
  57935=>"010011000",
  57936=>"010100100",
  57937=>"101010000",
  57938=>"010110110",
  57939=>"100111100",
  57940=>"100011000",
  57941=>"101010001",
  57942=>"111100111",
  57943=>"100010110",
  57944=>"010111110",
  57945=>"100010011",
  57946=>"011000011",
  57947=>"100000001",
  57948=>"001101111",
  57949=>"000100010",
  57950=>"100010010",
  57951=>"001001111",
  57952=>"111011110",
  57953=>"001010001",
  57954=>"101110111",
  57955=>"110100010",
  57956=>"011010000",
  57957=>"000011011",
  57958=>"001000111",
  57959=>"100100110",
  57960=>"011011110",
  57961=>"100000100",
  57962=>"000010011",
  57963=>"011110000",
  57964=>"010000010",
  57965=>"111010000",
  57966=>"101011000",
  57967=>"010010101",
  57968=>"110001010",
  57969=>"001000001",
  57970=>"100110001",
  57971=>"000111010",
  57972=>"101100010",
  57973=>"010001000",
  57974=>"101011101",
  57975=>"011001010",
  57976=>"001001101",
  57977=>"111100111",
  57978=>"110101000",
  57979=>"100010000",
  57980=>"011000000",
  57981=>"101011000",
  57982=>"000101111",
  57983=>"111101011",
  57984=>"100010000",
  57985=>"010011010",
  57986=>"011100101",
  57987=>"010000100",
  57988=>"100001010",
  57989=>"001001000",
  57990=>"100101010",
  57991=>"000001000",
  57992=>"010110101",
  57993=>"011100000",
  57994=>"100111011",
  57995=>"000110101",
  57996=>"100011100",
  57997=>"000100001",
  57998=>"101100111",
  57999=>"010110001",
  58000=>"010101110",
  58001=>"000010111",
  58002=>"101110110",
  58003=>"110111101",
  58004=>"101101100",
  58005=>"000011110",
  58006=>"001000110",
  58007=>"010001100",
  58008=>"110000000",
  58009=>"101010100",
  58010=>"011010101",
  58011=>"111101000",
  58012=>"000111110",
  58013=>"100010111",
  58014=>"010011000",
  58015=>"000011000",
  58016=>"000001100",
  58017=>"100110111",
  58018=>"011111101",
  58019=>"111111100",
  58020=>"010000001",
  58021=>"001011001",
  58022=>"011010100",
  58023=>"100010011",
  58024=>"100110101",
  58025=>"001111000",
  58026=>"000000101",
  58027=>"101100100",
  58028=>"000100000",
  58029=>"010001101",
  58030=>"111110011",
  58031=>"100101101",
  58032=>"010110001",
  58033=>"101001010",
  58034=>"101010101",
  58035=>"001111011",
  58036=>"001001000",
  58037=>"101010000",
  58038=>"011100101",
  58039=>"000111000",
  58040=>"100101101",
  58041=>"101101101",
  58042=>"001110010",
  58043=>"101111001",
  58044=>"011100101",
  58045=>"011000011",
  58046=>"101011010",
  58047=>"101000001",
  58048=>"111000001",
  58049=>"001011111",
  58050=>"111010101",
  58051=>"011101101",
  58052=>"010010000",
  58053=>"000111100",
  58054=>"010110111",
  58055=>"000011001",
  58056=>"000100100",
  58057=>"100100111",
  58058=>"111010111",
  58059=>"000111001",
  58060=>"010100101",
  58061=>"111101111",
  58062=>"101101100",
  58063=>"001010000",
  58064=>"101010110",
  58065=>"100010000",
  58066=>"010001000",
  58067=>"111101011",
  58068=>"101111110",
  58069=>"010110000",
  58070=>"101000101",
  58071=>"101110010",
  58072=>"111010100",
  58073=>"001100000",
  58074=>"100001011",
  58075=>"010111011",
  58076=>"110001101",
  58077=>"010000000",
  58078=>"000110000",
  58079=>"111010011",
  58080=>"110011110",
  58081=>"000111110",
  58082=>"001010011",
  58083=>"011010001",
  58084=>"011010100",
  58085=>"001001110",
  58086=>"010001100",
  58087=>"010000001",
  58088=>"100010011",
  58089=>"010010100",
  58090=>"011101001",
  58091=>"010111100",
  58092=>"000101011",
  58093=>"001110001",
  58094=>"011110000",
  58095=>"100001101",
  58096=>"110001110",
  58097=>"001000001",
  58098=>"000000111",
  58099=>"100110001",
  58100=>"111000001",
  58101=>"001110000",
  58102=>"110111000",
  58103=>"000000111",
  58104=>"111000000",
  58105=>"000111100",
  58106=>"100011110",
  58107=>"101101010",
  58108=>"110110010",
  58109=>"110100100",
  58110=>"011010001",
  58111=>"011011001",
  58112=>"110111001",
  58113=>"010111100",
  58114=>"111111110",
  58115=>"000010001",
  58116=>"001000010",
  58117=>"001100101",
  58118=>"111101010",
  58119=>"000011101",
  58120=>"010110011",
  58121=>"111111010",
  58122=>"111100101",
  58123=>"001110100",
  58124=>"011101010",
  58125=>"011010101",
  58126=>"111100011",
  58127=>"111010111",
  58128=>"111111000",
  58129=>"111011001",
  58130=>"011111111",
  58131=>"010101011",
  58132=>"101001011",
  58133=>"010101011",
  58134=>"000010000",
  58135=>"010001011",
  58136=>"110010000",
  58137=>"000111011",
  58138=>"001100111",
  58139=>"111000110",
  58140=>"001100001",
  58141=>"011100110",
  58142=>"111100011",
  58143=>"110111111",
  58144=>"110111111",
  58145=>"111010001",
  58146=>"110011101",
  58147=>"010010011",
  58148=>"110100001",
  58149=>"100000000",
  58150=>"001001001",
  58151=>"010011100",
  58152=>"111010100",
  58153=>"100111111",
  58154=>"000010111",
  58155=>"111100000",
  58156=>"100001110",
  58157=>"000011010",
  58158=>"100011001",
  58159=>"000000001",
  58160=>"000011110",
  58161=>"110100000",
  58162=>"101010100",
  58163=>"010111001",
  58164=>"101010000",
  58165=>"100101111",
  58166=>"001000111",
  58167=>"100010100",
  58168=>"101000100",
  58169=>"001000110",
  58170=>"011100000",
  58171=>"100100100",
  58172=>"110000001",
  58173=>"001100100",
  58174=>"101111111",
  58175=>"001101011",
  58176=>"000010100",
  58177=>"000011011",
  58178=>"101111000",
  58179=>"100111101",
  58180=>"101000011",
  58181=>"011111001",
  58182=>"010010100",
  58183=>"101001010",
  58184=>"010011011",
  58185=>"111011000",
  58186=>"111011010",
  58187=>"101010000",
  58188=>"100101001",
  58189=>"010010001",
  58190=>"001001100",
  58191=>"001101111",
  58192=>"110110110",
  58193=>"110010001",
  58194=>"011101010",
  58195=>"010110001",
  58196=>"010010100",
  58197=>"100000011",
  58198=>"100000010",
  58199=>"011000000",
  58200=>"111111011",
  58201=>"101011001",
  58202=>"101011101",
  58203=>"000101100",
  58204=>"111001100",
  58205=>"111100011",
  58206=>"001110001",
  58207=>"000111000",
  58208=>"110011000",
  58209=>"010011100",
  58210=>"001000101",
  58211=>"101101110",
  58212=>"110110001",
  58213=>"010111100",
  58214=>"110011000",
  58215=>"001101001",
  58216=>"011111100",
  58217=>"110110001",
  58218=>"100100111",
  58219=>"011000110",
  58220=>"011000100",
  58221=>"100010011",
  58222=>"111001001",
  58223=>"101101000",
  58224=>"010101110",
  58225=>"000101100",
  58226=>"110000011",
  58227=>"111001010",
  58228=>"101010010",
  58229=>"000110100",
  58230=>"010010110",
  58231=>"100101001",
  58232=>"111100011",
  58233=>"010101000",
  58234=>"000111101",
  58235=>"111111001",
  58236=>"001011111",
  58237=>"000100010",
  58238=>"110010000",
  58239=>"111111101",
  58240=>"011001000",
  58241=>"101101000",
  58242=>"000100011",
  58243=>"001001101",
  58244=>"100111101",
  58245=>"010001111",
  58246=>"000100101",
  58247=>"000101101",
  58248=>"010011001",
  58249=>"101000000",
  58250=>"101100100",
  58251=>"111000000",
  58252=>"000001111",
  58253=>"001111010",
  58254=>"100010011",
  58255=>"001101010",
  58256=>"101001011",
  58257=>"011001101",
  58258=>"000010111",
  58259=>"010101000",
  58260=>"000000011",
  58261=>"001000110",
  58262=>"001011110",
  58263=>"000101101",
  58264=>"010101100",
  58265=>"001011000",
  58266=>"111101010",
  58267=>"101111011",
  58268=>"100011001",
  58269=>"001010010",
  58270=>"010111101",
  58271=>"111110111",
  58272=>"111001111",
  58273=>"000111100",
  58274=>"001111001",
  58275=>"001011001",
  58276=>"011111000",
  58277=>"011001100",
  58278=>"101010000",
  58279=>"100100100",
  58280=>"011110100",
  58281=>"010111011",
  58282=>"101010110",
  58283=>"111010010",
  58284=>"100010101",
  58285=>"111011011",
  58286=>"101000100",
  58287=>"010000110",
  58288=>"010000111",
  58289=>"101110110",
  58290=>"011110101",
  58291=>"101100001",
  58292=>"100100001",
  58293=>"011111111",
  58294=>"011111111",
  58295=>"110100010",
  58296=>"010110000",
  58297=>"000100110",
  58298=>"001010011",
  58299=>"111001010",
  58300=>"101111001",
  58301=>"011000011",
  58302=>"101011011",
  58303=>"100011010",
  58304=>"110100100",
  58305=>"100110010",
  58306=>"010111111",
  58307=>"011011111",
  58308=>"101110100",
  58309=>"011111110",
  58310=>"010000001",
  58311=>"101011010",
  58312=>"111000100",
  58313=>"100100100",
  58314=>"110101011",
  58315=>"101110010",
  58316=>"111001110",
  58317=>"000000111",
  58318=>"100010100",
  58319=>"111010001",
  58320=>"110001110",
  58321=>"110010101",
  58322=>"010011011",
  58323=>"101010110",
  58324=>"100000000",
  58325=>"111010001",
  58326=>"010000111",
  58327=>"011111111",
  58328=>"110011110",
  58329=>"101111111",
  58330=>"111110001",
  58331=>"100001010",
  58332=>"100101010",
  58333=>"010111110",
  58334=>"111111001",
  58335=>"110011100",
  58336=>"111111110",
  58337=>"000101000",
  58338=>"001111100",
  58339=>"100110111",
  58340=>"001010000",
  58341=>"011111101",
  58342=>"101010011",
  58343=>"100101000",
  58344=>"011110001",
  58345=>"111010110",
  58346=>"101101111",
  58347=>"011100000",
  58348=>"000100101",
  58349=>"111011101",
  58350=>"101110101",
  58351=>"011101100",
  58352=>"110010010",
  58353=>"110101000",
  58354=>"111101111",
  58355=>"111001110",
  58356=>"110110010",
  58357=>"100000111",
  58358=>"110001111",
  58359=>"011101001",
  58360=>"111101101",
  58361=>"010101001",
  58362=>"100100001",
  58363=>"010111111",
  58364=>"011111011",
  58365=>"110100001",
  58366=>"000111101",
  58367=>"000111111",
  58368=>"000011110",
  58369=>"010111010",
  58370=>"011100011",
  58371=>"011011011",
  58372=>"010010010",
  58373=>"001001001",
  58374=>"011110110",
  58375=>"001101000",
  58376=>"111101111",
  58377=>"011110011",
  58378=>"001011111",
  58379=>"110000001",
  58380=>"110101001",
  58381=>"110011000",
  58382=>"111101010",
  58383=>"110010010",
  58384=>"010101011",
  58385=>"111011001",
  58386=>"110000000",
  58387=>"111101110",
  58388=>"001101100",
  58389=>"011000100",
  58390=>"011001011",
  58391=>"101001110",
  58392=>"100101100",
  58393=>"010010101",
  58394=>"100000011",
  58395=>"100100010",
  58396=>"011001000",
  58397=>"101010110",
  58398=>"111110110",
  58399=>"010101011",
  58400=>"010010000",
  58401=>"111111101",
  58402=>"110000011",
  58403=>"000000011",
  58404=>"110101110",
  58405=>"110000010",
  58406=>"110010111",
  58407=>"100110110",
  58408=>"100110011",
  58409=>"101011001",
  58410=>"010011000",
  58411=>"110100001",
  58412=>"001101101",
  58413=>"110010111",
  58414=>"000111011",
  58415=>"111101000",
  58416=>"110101100",
  58417=>"100100101",
  58418=>"101010001",
  58419=>"101100001",
  58420=>"110011111",
  58421=>"110100000",
  58422=>"111011101",
  58423=>"011011001",
  58424=>"100000111",
  58425=>"000111001",
  58426=>"100111111",
  58427=>"001010111",
  58428=>"101001000",
  58429=>"001101010",
  58430=>"101011011",
  58431=>"101100001",
  58432=>"001100000",
  58433=>"000010110",
  58434=>"101000000",
  58435=>"000011110",
  58436=>"000000101",
  58437=>"001100111",
  58438=>"111100000",
  58439=>"101111100",
  58440=>"010001011",
  58441=>"000010011",
  58442=>"000110010",
  58443=>"110010110",
  58444=>"110100110",
  58445=>"010111111",
  58446=>"011100110",
  58447=>"111001011",
  58448=>"010111101",
  58449=>"100110101",
  58450=>"110111110",
  58451=>"011010110",
  58452=>"111011000",
  58453=>"110010101",
  58454=>"001000111",
  58455=>"110011100",
  58456=>"101110011",
  58457=>"100100101",
  58458=>"011111101",
  58459=>"111000111",
  58460=>"011010000",
  58461=>"010011110",
  58462=>"000000001",
  58463=>"000010011",
  58464=>"011100110",
  58465=>"001110001",
  58466=>"100101011",
  58467=>"010111111",
  58468=>"101101000",
  58469=>"101101011",
  58470=>"110010011",
  58471=>"000010101",
  58472=>"111010100",
  58473=>"000001111",
  58474=>"111101000",
  58475=>"001001001",
  58476=>"100011011",
  58477=>"010010100",
  58478=>"000101111",
  58479=>"000000011",
  58480=>"011001111",
  58481=>"101110110",
  58482=>"001011010",
  58483=>"010111011",
  58484=>"111100101",
  58485=>"011000001",
  58486=>"111011000",
  58487=>"000101000",
  58488=>"011010100",
  58489=>"111111011",
  58490=>"100111000",
  58491=>"000010010",
  58492=>"111110101",
  58493=>"001011110",
  58494=>"110101110",
  58495=>"010001010",
  58496=>"101011001",
  58497=>"110010000",
  58498=>"001000101",
  58499=>"011111001",
  58500=>"000000000",
  58501=>"000010110",
  58502=>"000110000",
  58503=>"010000000",
  58504=>"111100001",
  58505=>"011100001",
  58506=>"110011001",
  58507=>"000100000",
  58508=>"101111111",
  58509=>"110010011",
  58510=>"000001000",
  58511=>"111001011",
  58512=>"110101111",
  58513=>"001010001",
  58514=>"010010101",
  58515=>"100010001",
  58516=>"000100101",
  58517=>"010111111",
  58518=>"001011010",
  58519=>"111010110",
  58520=>"001110000",
  58521=>"001111011",
  58522=>"000110000",
  58523=>"001100101",
  58524=>"100011000",
  58525=>"010110011",
  58526=>"000011000",
  58527=>"100101011",
  58528=>"101000000",
  58529=>"101010101",
  58530=>"111100000",
  58531=>"001110001",
  58532=>"111101100",
  58533=>"101110111",
  58534=>"011111001",
  58535=>"011100010",
  58536=>"001100000",
  58537=>"101101111",
  58538=>"000001100",
  58539=>"011110110",
  58540=>"111101100",
  58541=>"001010011",
  58542=>"011110000",
  58543=>"101010111",
  58544=>"001110110",
  58545=>"101001111",
  58546=>"001101001",
  58547=>"100111101",
  58548=>"110100111",
  58549=>"011000000",
  58550=>"011111011",
  58551=>"101011110",
  58552=>"000110110",
  58553=>"111001100",
  58554=>"101001111",
  58555=>"101001111",
  58556=>"110101000",
  58557=>"100011011",
  58558=>"010110110",
  58559=>"100011000",
  58560=>"011011011",
  58561=>"101101100",
  58562=>"010101000",
  58563=>"011011010",
  58564=>"100100010",
  58565=>"100010110",
  58566=>"001100110",
  58567=>"010010000",
  58568=>"011110000",
  58569=>"010110111",
  58570=>"001101010",
  58571=>"101011000",
  58572=>"110000100",
  58573=>"101100010",
  58574=>"110000010",
  58575=>"111110111",
  58576=>"001001010",
  58577=>"000101010",
  58578=>"111111011",
  58579=>"000001101",
  58580=>"101001000",
  58581=>"001011001",
  58582=>"011111110",
  58583=>"110011100",
  58584=>"110111111",
  58585=>"010101111",
  58586=>"110100010",
  58587=>"110011111",
  58588=>"101011100",
  58589=>"001111010",
  58590=>"101100110",
  58591=>"100011010",
  58592=>"100000100",
  58593=>"111100101",
  58594=>"000010111",
  58595=>"011010111",
  58596=>"011001001",
  58597=>"000000111",
  58598=>"100111110",
  58599=>"100011001",
  58600=>"100111110",
  58601=>"001100000",
  58602=>"111010001",
  58603=>"101101010",
  58604=>"110101000",
  58605=>"100000101",
  58606=>"111110000",
  58607=>"000000010",
  58608=>"110001100",
  58609=>"001000010",
  58610=>"100001011",
  58611=>"001100101",
  58612=>"101100000",
  58613=>"000110110",
  58614=>"100110000",
  58615=>"100011011",
  58616=>"011111101",
  58617=>"110111000",
  58618=>"000100000",
  58619=>"001100011",
  58620=>"011101111",
  58621=>"000000100",
  58622=>"111111000",
  58623=>"000101111",
  58624=>"111001110",
  58625=>"101010111",
  58626=>"001111101",
  58627=>"100111101",
  58628=>"010111111",
  58629=>"101111001",
  58630=>"101010100",
  58631=>"110101000",
  58632=>"100000111",
  58633=>"100000010",
  58634=>"010010001",
  58635=>"011110111",
  58636=>"110111111",
  58637=>"111100101",
  58638=>"110011000",
  58639=>"000100011",
  58640=>"111100001",
  58641=>"111010000",
  58642=>"001011111",
  58643=>"001100111",
  58644=>"100001011",
  58645=>"111010100",
  58646=>"001001001",
  58647=>"111001010",
  58648=>"001101101",
  58649=>"100110101",
  58650=>"111100001",
  58651=>"001011000",
  58652=>"110010111",
  58653=>"100110010",
  58654=>"001000101",
  58655=>"100100011",
  58656=>"000001101",
  58657=>"110110010",
  58658=>"111010111",
  58659=>"110111110",
  58660=>"110001001",
  58661=>"011101110",
  58662=>"111100010",
  58663=>"110100001",
  58664=>"001000111",
  58665=>"101100110",
  58666=>"010010010",
  58667=>"111101001",
  58668=>"110101000",
  58669=>"000100001",
  58670=>"101010101",
  58671=>"010010000",
  58672=>"010100101",
  58673=>"011101001",
  58674=>"100010011",
  58675=>"100111000",
  58676=>"000000100",
  58677=>"111110111",
  58678=>"111000001",
  58679=>"100110011",
  58680=>"001100111",
  58681=>"011111100",
  58682=>"110100110",
  58683=>"000111110",
  58684=>"000101110",
  58685=>"001010001",
  58686=>"100000011",
  58687=>"011111110",
  58688=>"111111011",
  58689=>"000100110",
  58690=>"010101011",
  58691=>"011010001",
  58692=>"001010010",
  58693=>"001111111",
  58694=>"111001011",
  58695=>"101011010",
  58696=>"010000000",
  58697=>"100111010",
  58698=>"101111110",
  58699=>"011101010",
  58700=>"100101010",
  58701=>"010010111",
  58702=>"110000111",
  58703=>"110101001",
  58704=>"100001111",
  58705=>"111100000",
  58706=>"001001110",
  58707=>"010111010",
  58708=>"001110001",
  58709=>"000101111",
  58710=>"010010001",
  58711=>"011011010",
  58712=>"111000110",
  58713=>"111000101",
  58714=>"111111001",
  58715=>"110001111",
  58716=>"000010100",
  58717=>"011001001",
  58718=>"001000000",
  58719=>"000001111",
  58720=>"011110011",
  58721=>"111110000",
  58722=>"001111010",
  58723=>"101000000",
  58724=>"010100110",
  58725=>"001100100",
  58726=>"101000001",
  58727=>"100110010",
  58728=>"000000111",
  58729=>"010010011",
  58730=>"011001100",
  58731=>"000100101",
  58732=>"101100101",
  58733=>"010101110",
  58734=>"011000000",
  58735=>"100110011",
  58736=>"100011101",
  58737=>"010100010",
  58738=>"001001111",
  58739=>"000111100",
  58740=>"011110000",
  58741=>"000110001",
  58742=>"001111011",
  58743=>"100011111",
  58744=>"011101011",
  58745=>"101111000",
  58746=>"010111011",
  58747=>"000110101",
  58748=>"011111000",
  58749=>"001111100",
  58750=>"101001100",
  58751=>"111100011",
  58752=>"100011010",
  58753=>"101101100",
  58754=>"000100010",
  58755=>"111110010",
  58756=>"101001100",
  58757=>"110101001",
  58758=>"000001001",
  58759=>"100101011",
  58760=>"000111111",
  58761=>"010101010",
  58762=>"001111000",
  58763=>"011001001",
  58764=>"000000000",
  58765=>"100010000",
  58766=>"111100011",
  58767=>"111111110",
  58768=>"010111110",
  58769=>"001001000",
  58770=>"100000011",
  58771=>"111011010",
  58772=>"001010011",
  58773=>"010011100",
  58774=>"100101111",
  58775=>"110111110",
  58776=>"111101000",
  58777=>"101001010",
  58778=>"100110100",
  58779=>"000010011",
  58780=>"110010111",
  58781=>"010110010",
  58782=>"001011100",
  58783=>"000111000",
  58784=>"001011110",
  58785=>"001000101",
  58786=>"000000000",
  58787=>"000111100",
  58788=>"011111000",
  58789=>"010000001",
  58790=>"010101001",
  58791=>"111001100",
  58792=>"110000101",
  58793=>"110000100",
  58794=>"000110010",
  58795=>"011011001",
  58796=>"000010100",
  58797=>"010110100",
  58798=>"110000010",
  58799=>"110101000",
  58800=>"001010110",
  58801=>"001010101",
  58802=>"101000001",
  58803=>"010110111",
  58804=>"110010110",
  58805=>"011110011",
  58806=>"100000100",
  58807=>"101100101",
  58808=>"111101000",
  58809=>"001010000",
  58810=>"100011000",
  58811=>"111111100",
  58812=>"010101101",
  58813=>"101011001",
  58814=>"010011010",
  58815=>"001011001",
  58816=>"000100000",
  58817=>"101001101",
  58818=>"000001010",
  58819=>"110110110",
  58820=>"010011011",
  58821=>"111100100",
  58822=>"011100111",
  58823=>"011100001",
  58824=>"001101111",
  58825=>"110001011",
  58826=>"011001001",
  58827=>"110001000",
  58828=>"110111001",
  58829=>"011011110",
  58830=>"001010101",
  58831=>"101100111",
  58832=>"100100101",
  58833=>"001101001",
  58834=>"111011110",
  58835=>"010100010",
  58836=>"000111110",
  58837=>"000110101",
  58838=>"000101101",
  58839=>"101010110",
  58840=>"001010111",
  58841=>"111001010",
  58842=>"110101010",
  58843=>"101000100",
  58844=>"111101110",
  58845=>"110111010",
  58846=>"101010000",
  58847=>"011111110",
  58848=>"100110110",
  58849=>"111111101",
  58850=>"101001011",
  58851=>"110001111",
  58852=>"111011100",
  58853=>"000010001",
  58854=>"101100001",
  58855=>"010110001",
  58856=>"110000110",
  58857=>"010111010",
  58858=>"111011011",
  58859=>"101101101",
  58860=>"000100000",
  58861=>"001001111",
  58862=>"000111011",
  58863=>"001010110",
  58864=>"001001010",
  58865=>"000110011",
  58866=>"111100110",
  58867=>"100100011",
  58868=>"010011110",
  58869=>"001001001",
  58870=>"101111101",
  58871=>"110010100",
  58872=>"001110110",
  58873=>"001010110",
  58874=>"011010111",
  58875=>"111111100",
  58876=>"110010100",
  58877=>"011000000",
  58878=>"001111010",
  58879=>"010011111",
  58880=>"011111001",
  58881=>"100101110",
  58882=>"000000011",
  58883=>"111010000",
  58884=>"110111010",
  58885=>"110011101",
  58886=>"111101111",
  58887=>"001001100",
  58888=>"010111001",
  58889=>"111000000",
  58890=>"111000001",
  58891=>"100110101",
  58892=>"010001000",
  58893=>"011111011",
  58894=>"111000111",
  58895=>"000001001",
  58896=>"100011100",
  58897=>"011000011",
  58898=>"010111110",
  58899=>"010001010",
  58900=>"001110011",
  58901=>"111110011",
  58902=>"001110100",
  58903=>"011100110",
  58904=>"100100001",
  58905=>"000110010",
  58906=>"100101101",
  58907=>"111011010",
  58908=>"010010110",
  58909=>"111101000",
  58910=>"111110111",
  58911=>"111100100",
  58912=>"010111110",
  58913=>"110010100",
  58914=>"101101000",
  58915=>"000110001",
  58916=>"100000101",
  58917=>"110010011",
  58918=>"110010000",
  58919=>"001000100",
  58920=>"101000100",
  58921=>"101101100",
  58922=>"001010000",
  58923=>"101001100",
  58924=>"000111011",
  58925=>"111010100",
  58926=>"001001000",
  58927=>"000011000",
  58928=>"000101100",
  58929=>"011110101",
  58930=>"000011000",
  58931=>"110011110",
  58932=>"001100101",
  58933=>"001100010",
  58934=>"110000110",
  58935=>"111110111",
  58936=>"110111010",
  58937=>"001100001",
  58938=>"001010000",
  58939=>"000101111",
  58940=>"100111111",
  58941=>"110100110",
  58942=>"111110110",
  58943=>"110000000",
  58944=>"101001100",
  58945=>"111011100",
  58946=>"001000001",
  58947=>"011000111",
  58948=>"101101110",
  58949=>"101101111",
  58950=>"000111101",
  58951=>"110001011",
  58952=>"010010111",
  58953=>"110110011",
  58954=>"100111001",
  58955=>"000110011",
  58956=>"111011111",
  58957=>"100000010",
  58958=>"001000001",
  58959=>"101111011",
  58960=>"001110100",
  58961=>"000100010",
  58962=>"101111111",
  58963=>"010110110",
  58964=>"011101110",
  58965=>"001101001",
  58966=>"011100110",
  58967=>"111010001",
  58968=>"000000100",
  58969=>"110110000",
  58970=>"001101000",
  58971=>"110111100",
  58972=>"010010101",
  58973=>"111111111",
  58974=>"000111001",
  58975=>"111001000",
  58976=>"001000111",
  58977=>"011011001",
  58978=>"111101011",
  58979=>"000100110",
  58980=>"110011010",
  58981=>"101011110",
  58982=>"011001010",
  58983=>"100001011",
  58984=>"011101000",
  58985=>"000000100",
  58986=>"100101111",
  58987=>"110000111",
  58988=>"100000100",
  58989=>"100010011",
  58990=>"010110010",
  58991=>"110001111",
  58992=>"100101001",
  58993=>"100110000",
  58994=>"111010011",
  58995=>"111100100",
  58996=>"101000000",
  58997=>"101001100",
  58998=>"000111111",
  58999=>"101110000",
  59000=>"111100110",
  59001=>"010111011",
  59002=>"000010010",
  59003=>"100110111",
  59004=>"111110011",
  59005=>"101011011",
  59006=>"110000000",
  59007=>"110001101",
  59008=>"000001110",
  59009=>"111011111",
  59010=>"000001000",
  59011=>"001000000",
  59012=>"001011011",
  59013=>"111011011",
  59014=>"000111011",
  59015=>"000111110",
  59016=>"110001110",
  59017=>"000011101",
  59018=>"000001110",
  59019=>"101111111",
  59020=>"000101101",
  59021=>"001000101",
  59022=>"110100110",
  59023=>"000111000",
  59024=>"111001011",
  59025=>"110001000",
  59026=>"101000110",
  59027=>"110110010",
  59028=>"110001000",
  59029=>"101001001",
  59030=>"001011110",
  59031=>"010110101",
  59032=>"110000100",
  59033=>"011011101",
  59034=>"000100111",
  59035=>"111000101",
  59036=>"110001010",
  59037=>"101111001",
  59038=>"011100010",
  59039=>"101001100",
  59040=>"000101000",
  59041=>"000100001",
  59042=>"111010001",
  59043=>"110101110",
  59044=>"001001000",
  59045=>"010011111",
  59046=>"111001001",
  59047=>"101100010",
  59048=>"011000011",
  59049=>"001110001",
  59050=>"110100000",
  59051=>"000100000",
  59052=>"111000001",
  59053=>"110110111",
  59054=>"011100101",
  59055=>"011101100",
  59056=>"000001010",
  59057=>"001010101",
  59058=>"001000101",
  59059=>"000000000",
  59060=>"011100000",
  59061=>"100000001",
  59062=>"100010011",
  59063=>"100000011",
  59064=>"111110100",
  59065=>"011110000",
  59066=>"111101010",
  59067=>"011001100",
  59068=>"111011011",
  59069=>"000000011",
  59070=>"000010010",
  59071=>"010110110",
  59072=>"000110100",
  59073=>"000110000",
  59074=>"001111000",
  59075=>"010110101",
  59076=>"101010011",
  59077=>"101010001",
  59078=>"111110010",
  59079=>"100000011",
  59080=>"011000100",
  59081=>"010111111",
  59082=>"101110101",
  59083=>"100000000",
  59084=>"110110011",
  59085=>"010110101",
  59086=>"100111101",
  59087=>"100001011",
  59088=>"001000001",
  59089=>"011011001",
  59090=>"001000000",
  59091=>"110001100",
  59092=>"100100000",
  59093=>"110001011",
  59094=>"010111010",
  59095=>"000000111",
  59096=>"110101011",
  59097=>"110101101",
  59098=>"111111011",
  59099=>"100010010",
  59100=>"111101101",
  59101=>"101000101",
  59102=>"101111001",
  59103=>"010110100",
  59104=>"011101111",
  59105=>"100110001",
  59106=>"001100010",
  59107=>"001001000",
  59108=>"101100110",
  59109=>"100101100",
  59110=>"000111100",
  59111=>"001101011",
  59112=>"001001000",
  59113=>"111001011",
  59114=>"001000010",
  59115=>"101100011",
  59116=>"001111111",
  59117=>"100001010",
  59118=>"000010001",
  59119=>"100010000",
  59120=>"010011110",
  59121=>"100010101",
  59122=>"100001010",
  59123=>"101010011",
  59124=>"011011010",
  59125=>"100000010",
  59126=>"101001000",
  59127=>"010010101",
  59128=>"111010111",
  59129=>"000101010",
  59130=>"011110010",
  59131=>"010010011",
  59132=>"110010000",
  59133=>"111011100",
  59134=>"000000011",
  59135=>"011001101",
  59136=>"111101110",
  59137=>"111111011",
  59138=>"110110110",
  59139=>"001000011",
  59140=>"011110010",
  59141=>"011101011",
  59142=>"000101000",
  59143=>"111010111",
  59144=>"010011000",
  59145=>"111010000",
  59146=>"110000100",
  59147=>"000010010",
  59148=>"001100000",
  59149=>"111000111",
  59150=>"111100000",
  59151=>"111010110",
  59152=>"000001110",
  59153=>"000111011",
  59154=>"101101100",
  59155=>"100110011",
  59156=>"011011111",
  59157=>"010010001",
  59158=>"001001000",
  59159=>"110011111",
  59160=>"110010101",
  59161=>"000110100",
  59162=>"001011111",
  59163=>"111111101",
  59164=>"111100110",
  59165=>"000100011",
  59166=>"001111001",
  59167=>"010111100",
  59168=>"111001010",
  59169=>"100111100",
  59170=>"100111100",
  59171=>"001101001",
  59172=>"011000011",
  59173=>"101000011",
  59174=>"000101011",
  59175=>"010001111",
  59176=>"101110010",
  59177=>"000001001",
  59178=>"010110010",
  59179=>"111110001",
  59180=>"111001010",
  59181=>"101101111",
  59182=>"000000011",
  59183=>"001000001",
  59184=>"010010100",
  59185=>"111111101",
  59186=>"111101111",
  59187=>"011111001",
  59188=>"000100011",
  59189=>"010010001",
  59190=>"101000101",
  59191=>"010111011",
  59192=>"111110001",
  59193=>"000010101",
  59194=>"110000110",
  59195=>"000000111",
  59196=>"001011110",
  59197=>"111100110",
  59198=>"010110001",
  59199=>"010001001",
  59200=>"011111101",
  59201=>"011010011",
  59202=>"011101101",
  59203=>"011000110",
  59204=>"000011101",
  59205=>"001110100",
  59206=>"100000011",
  59207=>"010011010",
  59208=>"010011111",
  59209=>"011101010",
  59210=>"000000011",
  59211=>"110001101",
  59212=>"100001111",
  59213=>"101111010",
  59214=>"011011001",
  59215=>"010110001",
  59216=>"111111010",
  59217=>"011001000",
  59218=>"110010010",
  59219=>"100010111",
  59220=>"100100110",
  59221=>"011100100",
  59222=>"010000010",
  59223=>"110000001",
  59224=>"010000111",
  59225=>"011101101",
  59226=>"010100110",
  59227=>"110100111",
  59228=>"000110000",
  59229=>"001000101",
  59230=>"110111001",
  59231=>"001000011",
  59232=>"100110011",
  59233=>"001101100",
  59234=>"100011011",
  59235=>"101010001",
  59236=>"101010010",
  59237=>"110101011",
  59238=>"001000101",
  59239=>"000111000",
  59240=>"100011110",
  59241=>"100010010",
  59242=>"110011111",
  59243=>"101101101",
  59244=>"101001010",
  59245=>"110100000",
  59246=>"101000100",
  59247=>"101111010",
  59248=>"100110111",
  59249=>"011100110",
  59250=>"100000100",
  59251=>"101110111",
  59252=>"011110101",
  59253=>"011110011",
  59254=>"100111111",
  59255=>"010111101",
  59256=>"010000101",
  59257=>"100001101",
  59258=>"010011011",
  59259=>"011110101",
  59260=>"101000100",
  59261=>"110000000",
  59262=>"000111101",
  59263=>"000110110",
  59264=>"101110010",
  59265=>"001000001",
  59266=>"010110110",
  59267=>"001000101",
  59268=>"101011110",
  59269=>"000001001",
  59270=>"000000101",
  59271=>"100101010",
  59272=>"010011111",
  59273=>"100010111",
  59274=>"111111101",
  59275=>"010100101",
  59276=>"101011111",
  59277=>"001100101",
  59278=>"000010110",
  59279=>"111101010",
  59280=>"000001111",
  59281=>"110101001",
  59282=>"111111001",
  59283=>"010011111",
  59284=>"001110011",
  59285=>"111101000",
  59286=>"110111001",
  59287=>"001110101",
  59288=>"100001000",
  59289=>"100000101",
  59290=>"101000001",
  59291=>"000001010",
  59292=>"010010101",
  59293=>"011110111",
  59294=>"100100011",
  59295=>"111111001",
  59296=>"101000101",
  59297=>"111111010",
  59298=>"011100100",
  59299=>"001101000",
  59300=>"110110001",
  59301=>"000011011",
  59302=>"111001101",
  59303=>"111101001",
  59304=>"110011001",
  59305=>"001110101",
  59306=>"011111101",
  59307=>"110010111",
  59308=>"101000100",
  59309=>"010101010",
  59310=>"111110100",
  59311=>"010000101",
  59312=>"001001011",
  59313=>"001100110",
  59314=>"010000000",
  59315=>"101001110",
  59316=>"111101110",
  59317=>"110011010",
  59318=>"100011111",
  59319=>"110100101",
  59320=>"110100110",
  59321=>"100111010",
  59322=>"111110101",
  59323=>"011111100",
  59324=>"101000011",
  59325=>"000010101",
  59326=>"010110111",
  59327=>"010000000",
  59328=>"010010001",
  59329=>"110011010",
  59330=>"001101110",
  59331=>"010001111",
  59332=>"010010111",
  59333=>"000001101",
  59334=>"111100000",
  59335=>"111110110",
  59336=>"110110011",
  59337=>"110110100",
  59338=>"001000011",
  59339=>"001000100",
  59340=>"111011100",
  59341=>"010101101",
  59342=>"001010000",
  59343=>"011010001",
  59344=>"011001101",
  59345=>"011000101",
  59346=>"010010000",
  59347=>"010110111",
  59348=>"001111111",
  59349=>"110110000",
  59350=>"000010111",
  59351=>"111110001",
  59352=>"101110000",
  59353=>"001011100",
  59354=>"101111001",
  59355=>"000000101",
  59356=>"110100111",
  59357=>"110110000",
  59358=>"001111100",
  59359=>"100100010",
  59360=>"001010111",
  59361=>"011100010",
  59362=>"000111010",
  59363=>"011010011",
  59364=>"000110111",
  59365=>"100010001",
  59366=>"000011111",
  59367=>"010001101",
  59368=>"011011011",
  59369=>"111010001",
  59370=>"001000010",
  59371=>"001010110",
  59372=>"101100111",
  59373=>"100110011",
  59374=>"100111011",
  59375=>"111111101",
  59376=>"000101000",
  59377=>"000001000",
  59378=>"000100111",
  59379=>"001000101",
  59380=>"010111110",
  59381=>"110111011",
  59382=>"000111110",
  59383=>"011010010",
  59384=>"110101000",
  59385=>"101000101",
  59386=>"001111111",
  59387=>"101001001",
  59388=>"001110010",
  59389=>"101011100",
  59390=>"110110001",
  59391=>"101111101",
  59392=>"011101000",
  59393=>"000000111",
  59394=>"111000000",
  59395=>"000101010",
  59396=>"001100110",
  59397=>"101101100",
  59398=>"010001011",
  59399=>"001100101",
  59400=>"000101111",
  59401=>"110010010",
  59402=>"000110111",
  59403=>"100100111",
  59404=>"101010000",
  59405=>"000100000",
  59406=>"101100011",
  59407=>"010000000",
  59408=>"011001000",
  59409=>"111010010",
  59410=>"110001110",
  59411=>"001111000",
  59412=>"010110001",
  59413=>"100110100",
  59414=>"111100011",
  59415=>"100010011",
  59416=>"000000110",
  59417=>"110110100",
  59418=>"111110110",
  59419=>"111100110",
  59420=>"000111110",
  59421=>"101111110",
  59422=>"000010010",
  59423=>"011001011",
  59424=>"010100000",
  59425=>"001001111",
  59426=>"111000111",
  59427=>"110101110",
  59428=>"000001110",
  59429=>"100100100",
  59430=>"001101011",
  59431=>"111001100",
  59432=>"100111011",
  59433=>"010010001",
  59434=>"000101100",
  59435=>"110100000",
  59436=>"100100000",
  59437=>"010010010",
  59438=>"011100101",
  59439=>"000000010",
  59440=>"010000111",
  59441=>"101010100",
  59442=>"010111101",
  59443=>"011011110",
  59444=>"111111100",
  59445=>"010000100",
  59446=>"011000110",
  59447=>"110100101",
  59448=>"101001111",
  59449=>"001011000",
  59450=>"101111111",
  59451=>"100100101",
  59452=>"100101001",
  59453=>"000110111",
  59454=>"011111000",
  59455=>"101011100",
  59456=>"110100100",
  59457=>"011110010",
  59458=>"010110000",
  59459=>"111010011",
  59460=>"111011011",
  59461=>"100111001",
  59462=>"101001101",
  59463=>"010101101",
  59464=>"000100111",
  59465=>"101010101",
  59466=>"111010011",
  59467=>"011100110",
  59468=>"110000010",
  59469=>"010101001",
  59470=>"110010000",
  59471=>"001101011",
  59472=>"001000100",
  59473=>"101001100",
  59474=>"101111110",
  59475=>"011000111",
  59476=>"001110100",
  59477=>"110111100",
  59478=>"000110110",
  59479=>"011000010",
  59480=>"000110011",
  59481=>"000111100",
  59482=>"110010110",
  59483=>"000000000",
  59484=>"001000001",
  59485=>"000000101",
  59486=>"101101100",
  59487=>"010011000",
  59488=>"000010110",
  59489=>"001001101",
  59490=>"100001101",
  59491=>"110100011",
  59492=>"111011111",
  59493=>"111111000",
  59494=>"011001100",
  59495=>"011001000",
  59496=>"000011100",
  59497=>"110110001",
  59498=>"000001011",
  59499=>"111000001",
  59500=>"010101000",
  59501=>"001010011",
  59502=>"100010000",
  59503=>"001000000",
  59504=>"000001010",
  59505=>"111011101",
  59506=>"101010111",
  59507=>"011110101",
  59508=>"110100011",
  59509=>"101100001",
  59510=>"100000010",
  59511=>"010110001",
  59512=>"010100110",
  59513=>"101111110",
  59514=>"000011101",
  59515=>"010011110",
  59516=>"001000011",
  59517=>"111111000",
  59518=>"000101011",
  59519=>"000011011",
  59520=>"010110011",
  59521=>"010110110",
  59522=>"110011101",
  59523=>"001001101",
  59524=>"011011010",
  59525=>"110100010",
  59526=>"100011010",
  59527=>"010110111",
  59528=>"101000101",
  59529=>"100000001",
  59530=>"011001010",
  59531=>"100100011",
  59532=>"110001001",
  59533=>"110110101",
  59534=>"111101010",
  59535=>"100111101",
  59536=>"110111001",
  59537=>"101011111",
  59538=>"011101101",
  59539=>"001010010",
  59540=>"011101110",
  59541=>"000010111",
  59542=>"101110111",
  59543=>"011010011",
  59544=>"010111100",
  59545=>"101101110",
  59546=>"101111011",
  59547=>"000001111",
  59548=>"010110100",
  59549=>"001110101",
  59550=>"000100000",
  59551=>"000010011",
  59552=>"000110010",
  59553=>"110000010",
  59554=>"100111011",
  59555=>"010000000",
  59556=>"111101011",
  59557=>"011001100",
  59558=>"001001000",
  59559=>"110101111",
  59560=>"000000101",
  59561=>"001100011",
  59562=>"110010000",
  59563=>"100110011",
  59564=>"101011001",
  59565=>"100000000",
  59566=>"110100001",
  59567=>"101000011",
  59568=>"001111110",
  59569=>"010101100",
  59570=>"000101101",
  59571=>"111011100",
  59572=>"100001000",
  59573=>"010111011",
  59574=>"000101100",
  59575=>"000001100",
  59576=>"110101101",
  59577=>"010001000",
  59578=>"011001110",
  59579=>"101111010",
  59580=>"100111010",
  59581=>"000000101",
  59582=>"100011111",
  59583=>"010111110",
  59584=>"110110000",
  59585=>"101000100",
  59586=>"001011000",
  59587=>"111111100",
  59588=>"011100110",
  59589=>"110100001",
  59590=>"001001000",
  59591=>"111001010",
  59592=>"000011011",
  59593=>"100000010",
  59594=>"111011011",
  59595=>"110010010",
  59596=>"001011000",
  59597=>"101100111",
  59598=>"110010010",
  59599=>"100100100",
  59600=>"100111111",
  59601=>"001000110",
  59602=>"010000001",
  59603=>"100001000",
  59604=>"111110010",
  59605=>"100001110",
  59606=>"011000010",
  59607=>"110011111",
  59608=>"000001000",
  59609=>"100111110",
  59610=>"100010111",
  59611=>"111011101",
  59612=>"100110011",
  59613=>"110000110",
  59614=>"000000000",
  59615=>"101110110",
  59616=>"101100001",
  59617=>"111000100",
  59618=>"000000110",
  59619=>"111101111",
  59620=>"001111001",
  59621=>"110010001",
  59622=>"110011010",
  59623=>"101101001",
  59624=>"101111001",
  59625=>"001001101",
  59626=>"000000010",
  59627=>"000100000",
  59628=>"000111001",
  59629=>"011100100",
  59630=>"110100001",
  59631=>"101001100",
  59632=>"010110110",
  59633=>"111000110",
  59634=>"000110000",
  59635=>"110110010",
  59636=>"111010101",
  59637=>"110101111",
  59638=>"101010110",
  59639=>"000011111",
  59640=>"011000001",
  59641=>"010011101",
  59642=>"011001100",
  59643=>"100000101",
  59644=>"101001110",
  59645=>"101000110",
  59646=>"111001010",
  59647=>"010000111",
  59648=>"000101010",
  59649=>"100001100",
  59650=>"111100101",
  59651=>"010100001",
  59652=>"010101101",
  59653=>"001111011",
  59654=>"101000011",
  59655=>"110101101",
  59656=>"100000001",
  59657=>"000011100",
  59658=>"001001011",
  59659=>"010100011",
  59660=>"001010011",
  59661=>"011100011",
  59662=>"110000011",
  59663=>"101101000",
  59664=>"010011011",
  59665=>"100000010",
  59666=>"100100010",
  59667=>"101000010",
  59668=>"001110000",
  59669=>"000010000",
  59670=>"111011110",
  59671=>"000010001",
  59672=>"001111101",
  59673=>"001001000",
  59674=>"000000110",
  59675=>"011000100",
  59676=>"000101111",
  59677=>"010110100",
  59678=>"000110010",
  59679=>"101011111",
  59680=>"000001011",
  59681=>"100001010",
  59682=>"110011100",
  59683=>"111001000",
  59684=>"010011101",
  59685=>"010000101",
  59686=>"001001011",
  59687=>"100010010",
  59688=>"100011101",
  59689=>"111111100",
  59690=>"000011110",
  59691=>"110111010",
  59692=>"100000001",
  59693=>"011101100",
  59694=>"011010010",
  59695=>"010111110",
  59696=>"000001010",
  59697=>"110100000",
  59698=>"110101110",
  59699=>"110110100",
  59700=>"100101011",
  59701=>"000111111",
  59702=>"111001011",
  59703=>"111111101",
  59704=>"100010010",
  59705=>"000011000",
  59706=>"000111000",
  59707=>"001011101",
  59708=>"100111011",
  59709=>"011010011",
  59710=>"011100001",
  59711=>"010000001",
  59712=>"001100100",
  59713=>"100010000",
  59714=>"110110110",
  59715=>"000101001",
  59716=>"001101101",
  59717=>"111001110",
  59718=>"110010010",
  59719=>"011111101",
  59720=>"100010011",
  59721=>"100010001",
  59722=>"010011111",
  59723=>"100110010",
  59724=>"001111011",
  59725=>"000001110",
  59726=>"100001111",
  59727=>"011001100",
  59728=>"110111100",
  59729=>"011110001",
  59730=>"001111001",
  59731=>"101010010",
  59732=>"011010010",
  59733=>"000001111",
  59734=>"101011001",
  59735=>"111010101",
  59736=>"001000010",
  59737=>"000110100",
  59738=>"100000001",
  59739=>"010010001",
  59740=>"001010000",
  59741=>"100010110",
  59742=>"110010010",
  59743=>"110100000",
  59744=>"101111111",
  59745=>"000101111",
  59746=>"001001110",
  59747=>"001010011",
  59748=>"001110000",
  59749=>"001100010",
  59750=>"101000010",
  59751=>"001000001",
  59752=>"000100000",
  59753=>"010000010",
  59754=>"110000110",
  59755=>"011011010",
  59756=>"001110000",
  59757=>"100110101",
  59758=>"011000000",
  59759=>"001111001",
  59760=>"001101011",
  59761=>"011111100",
  59762=>"000111110",
  59763=>"001001001",
  59764=>"001111111",
  59765=>"100101010",
  59766=>"000110010",
  59767=>"011010010",
  59768=>"111111110",
  59769=>"010001001",
  59770=>"101011000",
  59771=>"000000011",
  59772=>"100001011",
  59773=>"001110010",
  59774=>"111101011",
  59775=>"011110111",
  59776=>"111001011",
  59777=>"110010111",
  59778=>"011011110",
  59779=>"011100010",
  59780=>"010110111",
  59781=>"000101100",
  59782=>"000000001",
  59783=>"100110100",
  59784=>"111011010",
  59785=>"000111000",
  59786=>"100111010",
  59787=>"011000000",
  59788=>"110111010",
  59789=>"001100110",
  59790=>"011001010",
  59791=>"110001001",
  59792=>"011110000",
  59793=>"101101101",
  59794=>"000101100",
  59795=>"110100000",
  59796=>"010101000",
  59797=>"100101111",
  59798=>"011100000",
  59799=>"011100011",
  59800=>"101001010",
  59801=>"010101010",
  59802=>"001100000",
  59803=>"000000100",
  59804=>"110011001",
  59805=>"010110000",
  59806=>"110100101",
  59807=>"011110010",
  59808=>"110000110",
  59809=>"000000010",
  59810=>"111011110",
  59811=>"011001101",
  59812=>"101110100",
  59813=>"101001110",
  59814=>"001100110",
  59815=>"001000011",
  59816=>"011100011",
  59817=>"000010010",
  59818=>"101001101",
  59819=>"001110101",
  59820=>"001100010",
  59821=>"101111111",
  59822=>"011010111",
  59823=>"010110000",
  59824=>"000000010",
  59825=>"001100000",
  59826=>"100001101",
  59827=>"110011100",
  59828=>"011010000",
  59829=>"111011101",
  59830=>"110001111",
  59831=>"110101111",
  59832=>"111100010",
  59833=>"010101100",
  59834=>"111001001",
  59835=>"111011110",
  59836=>"000000001",
  59837=>"001011010",
  59838=>"110110001",
  59839=>"110100101",
  59840=>"011111110",
  59841=>"110110001",
  59842=>"110111000",
  59843=>"100110111",
  59844=>"111101000",
  59845=>"000010000",
  59846=>"110010100",
  59847=>"111100000",
  59848=>"000011001",
  59849=>"000110111",
  59850=>"011011001",
  59851=>"101010111",
  59852=>"001000101",
  59853=>"101000010",
  59854=>"101011011",
  59855=>"001011000",
  59856=>"110000011",
  59857=>"111101111",
  59858=>"001000010",
  59859=>"100011000",
  59860=>"101101011",
  59861=>"001111000",
  59862=>"100111100",
  59863=>"111001001",
  59864=>"111110111",
  59865=>"001111111",
  59866=>"011111111",
  59867=>"111011000",
  59868=>"100000010",
  59869=>"011010000",
  59870=>"010010011",
  59871=>"110000011",
  59872=>"010000001",
  59873=>"000110111",
  59874=>"100000100",
  59875=>"000100000",
  59876=>"010011000",
  59877=>"100111011",
  59878=>"001101101",
  59879=>"100011010",
  59880=>"101011001",
  59881=>"100000001",
  59882=>"000100001",
  59883=>"111001110",
  59884=>"111100111",
  59885=>"000011011",
  59886=>"110010111",
  59887=>"100100100",
  59888=>"101110010",
  59889=>"100110001",
  59890=>"000111010",
  59891=>"010001001",
  59892=>"100111011",
  59893=>"001010101",
  59894=>"111110001",
  59895=>"001000100",
  59896=>"001100110",
  59897=>"101110000",
  59898=>"110011000",
  59899=>"000000001",
  59900=>"010110001",
  59901=>"110111000",
  59902=>"100111101",
  59903=>"000011001",
  59904=>"011001100",
  59905=>"000011110",
  59906=>"011001001",
  59907=>"001111100",
  59908=>"110100010",
  59909=>"010110000",
  59910=>"000111110",
  59911=>"000010011",
  59912=>"100001011",
  59913=>"011000110",
  59914=>"011110000",
  59915=>"111001110",
  59916=>"101111001",
  59917=>"110101000",
  59918=>"011010000",
  59919=>"001010110",
  59920=>"110010000",
  59921=>"110101111",
  59922=>"011100101",
  59923=>"101110111",
  59924=>"000011000",
  59925=>"001011101",
  59926=>"100110011",
  59927=>"111111000",
  59928=>"010011010",
  59929=>"110101100",
  59930=>"110111101",
  59931=>"101011010",
  59932=>"111110001",
  59933=>"010011010",
  59934=>"001010111",
  59935=>"111110111",
  59936=>"001101101",
  59937=>"100101000",
  59938=>"010000111",
  59939=>"010111101",
  59940=>"101000001",
  59941=>"011001001",
  59942=>"101000100",
  59943=>"001011010",
  59944=>"000000010",
  59945=>"101101110",
  59946=>"111111101",
  59947=>"001010100",
  59948=>"100011101",
  59949=>"010101000",
  59950=>"010001101",
  59951=>"101000101",
  59952=>"110101100",
  59953=>"111101101",
  59954=>"010001100",
  59955=>"011000011",
  59956=>"001010010",
  59957=>"001010110",
  59958=>"110100010",
  59959=>"110000110",
  59960=>"000001111",
  59961=>"001111011",
  59962=>"010100101",
  59963=>"101011110",
  59964=>"001110000",
  59965=>"001011111",
  59966=>"111101100",
  59967=>"111110110",
  59968=>"001010011",
  59969=>"100011001",
  59970=>"000101101",
  59971=>"110011100",
  59972=>"101101011",
  59973=>"000011001",
  59974=>"111011111",
  59975=>"011000100",
  59976=>"001100110",
  59977=>"111000001",
  59978=>"111110001",
  59979=>"011000011",
  59980=>"010010111",
  59981=>"100100011",
  59982=>"110011001",
  59983=>"111001000",
  59984=>"111111111",
  59985=>"000010000",
  59986=>"100110101",
  59987=>"101101000",
  59988=>"010111011",
  59989=>"111111011",
  59990=>"100001010",
  59991=>"100111101",
  59992=>"110000110",
  59993=>"100001011",
  59994=>"111111000",
  59995=>"000101011",
  59996=>"001100010",
  59997=>"111001000",
  59998=>"001011100",
  59999=>"110100101",
  60000=>"101101110",
  60001=>"111110001",
  60002=>"010110100",
  60003=>"011011110",
  60004=>"101110011",
  60005=>"001101100",
  60006=>"001011111",
  60007=>"111100010",
  60008=>"001001000",
  60009=>"111001110",
  60010=>"100111110",
  60011=>"011000110",
  60012=>"110010010",
  60013=>"011001001",
  60014=>"000001010",
  60015=>"010111100",
  60016=>"000100011",
  60017=>"011100000",
  60018=>"000001010",
  60019=>"001101001",
  60020=>"100010100",
  60021=>"111010100",
  60022=>"000110000",
  60023=>"100111010",
  60024=>"110111011",
  60025=>"111110111",
  60026=>"010010110",
  60027=>"001010001",
  60028=>"010101011",
  60029=>"011010110",
  60030=>"101111011",
  60031=>"000100010",
  60032=>"001010100",
  60033=>"101110111",
  60034=>"011001001",
  60035=>"101100100",
  60036=>"101010001",
  60037=>"010100000",
  60038=>"000011001",
  60039=>"011101010",
  60040=>"010010111",
  60041=>"000110111",
  60042=>"100010001",
  60043=>"111010000",
  60044=>"100000010",
  60045=>"010000111",
  60046=>"101110010",
  60047=>"001100101",
  60048=>"010100010",
  60049=>"001000011",
  60050=>"111001110",
  60051=>"011001111",
  60052=>"110000011",
  60053=>"010010010",
  60054=>"110110110",
  60055=>"000101000",
  60056=>"101011100",
  60057=>"110011011",
  60058=>"100100100",
  60059=>"111100111",
  60060=>"110111011",
  60061=>"000111010",
  60062=>"000110010",
  60063=>"110001010",
  60064=>"000100110",
  60065=>"011001101",
  60066=>"111000111",
  60067=>"000000011",
  60068=>"110110101",
  60069=>"011001010",
  60070=>"101000000",
  60071=>"110000100",
  60072=>"010100111",
  60073=>"001011010",
  60074=>"001101100",
  60075=>"100100011",
  60076=>"111111000",
  60077=>"000010011",
  60078=>"100100000",
  60079=>"110101001",
  60080=>"010101011",
  60081=>"110001101",
  60082=>"101000001",
  60083=>"111111101",
  60084=>"010100001",
  60085=>"110100000",
  60086=>"101011000",
  60087=>"010001110",
  60088=>"010111100",
  60089=>"111110101",
  60090=>"010110110",
  60091=>"100010011",
  60092=>"010101010",
  60093=>"111111111",
  60094=>"011101100",
  60095=>"011001111",
  60096=>"000011111",
  60097=>"111011000",
  60098=>"101101100",
  60099=>"011110000",
  60100=>"011000110",
  60101=>"110101001",
  60102=>"010010010",
  60103=>"010111011",
  60104=>"111100111",
  60105=>"100101011",
  60106=>"111101010",
  60107=>"000100100",
  60108=>"010000001",
  60109=>"010100101",
  60110=>"111011110",
  60111=>"100111111",
  60112=>"000101000",
  60113=>"111000111",
  60114=>"101110111",
  60115=>"111101110",
  60116=>"100100001",
  60117=>"000000010",
  60118=>"011011111",
  60119=>"111000100",
  60120=>"000000011",
  60121=>"101101010",
  60122=>"010111110",
  60123=>"111100001",
  60124=>"111101010",
  60125=>"000011011",
  60126=>"000110000",
  60127=>"110001110",
  60128=>"100000011",
  60129=>"011001110",
  60130=>"111100011",
  60131=>"110101111",
  60132=>"010000100",
  60133=>"001111101",
  60134=>"011100001",
  60135=>"110100010",
  60136=>"011010011",
  60137=>"000001111",
  60138=>"101011110",
  60139=>"101000001",
  60140=>"010011000",
  60141=>"001001011",
  60142=>"010110010",
  60143=>"000000110",
  60144=>"100110101",
  60145=>"101000111",
  60146=>"001001011",
  60147=>"111001001",
  60148=>"011010010",
  60149=>"110000001",
  60150=>"000100011",
  60151=>"011000111",
  60152=>"111001101",
  60153=>"110011101",
  60154=>"111000101",
  60155=>"011000100",
  60156=>"000000010",
  60157=>"010100010",
  60158=>"110000001",
  60159=>"111000011",
  60160=>"100101000",
  60161=>"010001000",
  60162=>"110110000",
  60163=>"000110011",
  60164=>"011101111",
  60165=>"100110100",
  60166=>"111011111",
  60167=>"111101011",
  60168=>"100010000",
  60169=>"001101011",
  60170=>"001000110",
  60171=>"011010111",
  60172=>"000000010",
  60173=>"000100001",
  60174=>"100010011",
  60175=>"011110001",
  60176=>"111111010",
  60177=>"001101000",
  60178=>"010001001",
  60179=>"100011111",
  60180=>"010100010",
  60181=>"101011111",
  60182=>"000100101",
  60183=>"110000010",
  60184=>"000010010",
  60185=>"111111110",
  60186=>"000001110",
  60187=>"100000010",
  60188=>"011011010",
  60189=>"010011010",
  60190=>"100001000",
  60191=>"000100001",
  60192=>"100000111",
  60193=>"011010110",
  60194=>"101000010",
  60195=>"111011111",
  60196=>"001101111",
  60197=>"101101111",
  60198=>"111110111",
  60199=>"111110011",
  60200=>"100101011",
  60201=>"000110001",
  60202=>"100111101",
  60203=>"111000010",
  60204=>"110110100",
  60205=>"000111101",
  60206=>"111100101",
  60207=>"101001000",
  60208=>"000000110",
  60209=>"111000100",
  60210=>"100101100",
  60211=>"000010101",
  60212=>"000100100",
  60213=>"000101111",
  60214=>"111010111",
  60215=>"110101101",
  60216=>"010010000",
  60217=>"100101100",
  60218=>"011000101",
  60219=>"001111011",
  60220=>"011010101",
  60221=>"011001010",
  60222=>"110011011",
  60223=>"110010001",
  60224=>"010000101",
  60225=>"100101111",
  60226=>"110111011",
  60227=>"000001000",
  60228=>"110001100",
  60229=>"110001101",
  60230=>"000010010",
  60231=>"011010110",
  60232=>"000100110",
  60233=>"111001111",
  60234=>"000011110",
  60235=>"100011101",
  60236=>"100010101",
  60237=>"111011110",
  60238=>"001100011",
  60239=>"100000000",
  60240=>"000001000",
  60241=>"100111111",
  60242=>"110101111",
  60243=>"100111011",
  60244=>"110011111",
  60245=>"100010111",
  60246=>"100001101",
  60247=>"101011100",
  60248=>"111101111",
  60249=>"000111101",
  60250=>"001111111",
  60251=>"000000001",
  60252=>"101100000",
  60253=>"111011010",
  60254=>"001010011",
  60255=>"011110111",
  60256=>"010100010",
  60257=>"110110110",
  60258=>"000101101",
  60259=>"000011100",
  60260=>"101100110",
  60261=>"010110111",
  60262=>"110010100",
  60263=>"110111010",
  60264=>"110001011",
  60265=>"111000110",
  60266=>"000110001",
  60267=>"011011111",
  60268=>"001110000",
  60269=>"111100011",
  60270=>"000010111",
  60271=>"101001100",
  60272=>"000000000",
  60273=>"000011110",
  60274=>"111100000",
  60275=>"111101011",
  60276=>"011000000",
  60277=>"000000010",
  60278=>"001010111",
  60279=>"101001011",
  60280=>"101011111",
  60281=>"111001011",
  60282=>"111001110",
  60283=>"010000110",
  60284=>"000000100",
  60285=>"111100010",
  60286=>"110110110",
  60287=>"000111111",
  60288=>"010010001",
  60289=>"110001011",
  60290=>"111100001",
  60291=>"001001100",
  60292=>"011000011",
  60293=>"000100000",
  60294=>"110101011",
  60295=>"111001110",
  60296=>"010100011",
  60297=>"010011111",
  60298=>"000101110",
  60299=>"000110110",
  60300=>"010110000",
  60301=>"111000011",
  60302=>"000110110",
  60303=>"111111100",
  60304=>"000111001",
  60305=>"011010100",
  60306=>"001010010",
  60307=>"111010010",
  60308=>"110111001",
  60309=>"011010110",
  60310=>"001011000",
  60311=>"100111000",
  60312=>"101001011",
  60313=>"111111001",
  60314=>"010000100",
  60315=>"001111100",
  60316=>"110011000",
  60317=>"110010100",
  60318=>"110000100",
  60319=>"110000000",
  60320=>"111111000",
  60321=>"010110001",
  60322=>"001101000",
  60323=>"100010110",
  60324=>"001011100",
  60325=>"111000011",
  60326=>"001010010",
  60327=>"010000111",
  60328=>"001000010",
  60329=>"100000001",
  60330=>"001001000",
  60331=>"111110000",
  60332=>"010000110",
  60333=>"110111101",
  60334=>"110101111",
  60335=>"110011000",
  60336=>"011010110",
  60337=>"001000101",
  60338=>"010010010",
  60339=>"100000110",
  60340=>"011100110",
  60341=>"000111010",
  60342=>"100100101",
  60343=>"011000001",
  60344=>"011011111",
  60345=>"010100010",
  60346=>"111011001",
  60347=>"001000000",
  60348=>"010100000",
  60349=>"100011111",
  60350=>"001110000",
  60351=>"010000000",
  60352=>"111111111",
  60353=>"001000110",
  60354=>"000111110",
  60355=>"110001101",
  60356=>"110100111",
  60357=>"000101101",
  60358=>"100010001",
  60359=>"001011001",
  60360=>"110000101",
  60361=>"100010110",
  60362=>"000110010",
  60363=>"100110100",
  60364=>"011011111",
  60365=>"110011110",
  60366=>"000010110",
  60367=>"110010101",
  60368=>"111000010",
  60369=>"000011001",
  60370=>"100011101",
  60371=>"101010011",
  60372=>"001010100",
  60373=>"111001011",
  60374=>"010110100",
  60375=>"100001010",
  60376=>"111110000",
  60377=>"101001100",
  60378=>"000011111",
  60379=>"100101011",
  60380=>"001110111",
  60381=>"001011100",
  60382=>"011101000",
  60383=>"011101110",
  60384=>"111010001",
  60385=>"111010010",
  60386=>"100000100",
  60387=>"000011010",
  60388=>"111010100",
  60389=>"110111010",
  60390=>"000010000",
  60391=>"000000100",
  60392=>"001010111",
  60393=>"110101101",
  60394=>"011100111",
  60395=>"111110000",
  60396=>"101001111",
  60397=>"010001110",
  60398=>"000101001",
  60399=>"001100111",
  60400=>"011000001",
  60401=>"000001101",
  60402=>"110001000",
  60403=>"001110111",
  60404=>"001100110",
  60405=>"101101000",
  60406=>"010010011",
  60407=>"101101101",
  60408=>"111111011",
  60409=>"100101011",
  60410=>"111000001",
  60411=>"100110000",
  60412=>"011100001",
  60413=>"000010100",
  60414=>"001101011",
  60415=>"110011010",
  60416=>"001001000",
  60417=>"100001100",
  60418=>"010000100",
  60419=>"000100011",
  60420=>"010001100",
  60421=>"000100110",
  60422=>"101000011",
  60423=>"001000111",
  60424=>"100110001",
  60425=>"101100101",
  60426=>"000111111",
  60427=>"001101000",
  60428=>"111011011",
  60429=>"000001100",
  60430=>"110100000",
  60431=>"100101011",
  60432=>"001111010",
  60433=>"001100011",
  60434=>"001100001",
  60435=>"000000100",
  60436=>"111101111",
  60437=>"001100100",
  60438=>"100111010",
  60439=>"101111110",
  60440=>"000010010",
  60441=>"111001110",
  60442=>"011011111",
  60443=>"111101011",
  60444=>"000000001",
  60445=>"111001110",
  60446=>"110101011",
  60447=>"101011000",
  60448=>"000110100",
  60449=>"011110101",
  60450=>"000001111",
  60451=>"100101011",
  60452=>"001111101",
  60453=>"011100010",
  60454=>"101000110",
  60455=>"010100000",
  60456=>"000111111",
  60457=>"100001100",
  60458=>"100011001",
  60459=>"100000101",
  60460=>"110101010",
  60461=>"001101100",
  60462=>"110101100",
  60463=>"010011000",
  60464=>"011101010",
  60465=>"100000101",
  60466=>"111101001",
  60467=>"110001110",
  60468=>"111110000",
  60469=>"110010011",
  60470=>"101000100",
  60471=>"100111011",
  60472=>"000000110",
  60473=>"111011000",
  60474=>"101010011",
  60475=>"001101010",
  60476=>"000000101",
  60477=>"110011101",
  60478=>"000011100",
  60479=>"001100111",
  60480=>"111101000",
  60481=>"001001100",
  60482=>"111100010",
  60483=>"100010001",
  60484=>"110001111",
  60485=>"110100100",
  60486=>"110100100",
  60487=>"111000010",
  60488=>"110111001",
  60489=>"101010011",
  60490=>"111100001",
  60491=>"010011111",
  60492=>"111000110",
  60493=>"111001011",
  60494=>"011000011",
  60495=>"000110001",
  60496=>"000000010",
  60497=>"111111011",
  60498=>"010000110",
  60499=>"000110101",
  60500=>"010110110",
  60501=>"111001000",
  60502=>"100011101",
  60503=>"101101001",
  60504=>"111110111",
  60505=>"000011110",
  60506=>"110010011",
  60507=>"010101000",
  60508=>"010100011",
  60509=>"111100011",
  60510=>"110000111",
  60511=>"001101101",
  60512=>"100100110",
  60513=>"100110110",
  60514=>"001111101",
  60515=>"000111011",
  60516=>"001111101",
  60517=>"000000111",
  60518=>"101101111",
  60519=>"110000000",
  60520=>"000101001",
  60521=>"101001011",
  60522=>"011101001",
  60523=>"111101001",
  60524=>"000101111",
  60525=>"000010000",
  60526=>"100000010",
  60527=>"101001101",
  60528=>"011000010",
  60529=>"010000000",
  60530=>"110101101",
  60531=>"001011000",
  60532=>"001111101",
  60533=>"011101011",
  60534=>"110011000",
  60535=>"101101010",
  60536=>"111010110",
  60537=>"110101100",
  60538=>"111101011",
  60539=>"111100100",
  60540=>"001111101",
  60541=>"000010110",
  60542=>"101011101",
  60543=>"111001101",
  60544=>"000010111",
  60545=>"101111011",
  60546=>"111101001",
  60547=>"100010010",
  60548=>"101010001",
  60549=>"011000001",
  60550=>"010101010",
  60551=>"101101001",
  60552=>"100111100",
  60553=>"000110011",
  60554=>"011001001",
  60555=>"110101100",
  60556=>"111000111",
  60557=>"000110010",
  60558=>"011110001",
  60559=>"100000100",
  60560=>"101000101",
  60561=>"111010110",
  60562=>"011110110",
  60563=>"111101111",
  60564=>"110001111",
  60565=>"011011100",
  60566=>"101000111",
  60567=>"000010011",
  60568=>"110011000",
  60569=>"101100101",
  60570=>"010101111",
  60571=>"000001011",
  60572=>"111110100",
  60573=>"100100111",
  60574=>"101110010",
  60575=>"001011100",
  60576=>"110010111",
  60577=>"110000001",
  60578=>"101101011",
  60579=>"101101000",
  60580=>"110111111",
  60581=>"011100001",
  60582=>"000111100",
  60583=>"011100110",
  60584=>"101001011",
  60585=>"001010000",
  60586=>"011010011",
  60587=>"001100100",
  60588=>"111010100",
  60589=>"101010110",
  60590=>"011010001",
  60591=>"011011011",
  60592=>"001011010",
  60593=>"110100111",
  60594=>"011101101",
  60595=>"011110011",
  60596=>"011110101",
  60597=>"011111111",
  60598=>"100111101",
  60599=>"000000000",
  60600=>"001001001",
  60601=>"100101101",
  60602=>"010000010",
  60603=>"110000001",
  60604=>"101101011",
  60605=>"001010011",
  60606=>"000000111",
  60607=>"111110100",
  60608=>"100110110",
  60609=>"000101001",
  60610=>"110101010",
  60611=>"000101001",
  60612=>"111110111",
  60613=>"001110111",
  60614=>"101111010",
  60615=>"110101111",
  60616=>"101010111",
  60617=>"010100101",
  60618=>"010000110",
  60619=>"010001100",
  60620=>"001110100",
  60621=>"111100111",
  60622=>"011001001",
  60623=>"010001101",
  60624=>"000100011",
  60625=>"010110100",
  60626=>"011110000",
  60627=>"101101110",
  60628=>"011100010",
  60629=>"010000100",
  60630=>"000010001",
  60631=>"100010010",
  60632=>"111101011",
  60633=>"011110100",
  60634=>"000101000",
  60635=>"111100100",
  60636=>"000011011",
  60637=>"000011110",
  60638=>"011101101",
  60639=>"001000001",
  60640=>"000111000",
  60641=>"111101111",
  60642=>"001001111",
  60643=>"111111111",
  60644=>"111111111",
  60645=>"111010110",
  60646=>"111111101",
  60647=>"111111010",
  60648=>"001100101",
  60649=>"101011000",
  60650=>"101010000",
  60651=>"111110100",
  60652=>"101111111",
  60653=>"000011001",
  60654=>"001011011",
  60655=>"000100000",
  60656=>"001001110",
  60657=>"001111101",
  60658=>"000100011",
  60659=>"101011110",
  60660=>"100001101",
  60661=>"011100101",
  60662=>"000110111",
  60663=>"101000011",
  60664=>"101000001",
  60665=>"101001011",
  60666=>"111111110",
  60667=>"111110101",
  60668=>"001010010",
  60669=>"111101100",
  60670=>"111101100",
  60671=>"010111100",
  60672=>"110111011",
  60673=>"100000101",
  60674=>"001100111",
  60675=>"011111000",
  60676=>"100100101",
  60677=>"100010001",
  60678=>"001010111",
  60679=>"011010010",
  60680=>"111001101",
  60681=>"110100110",
  60682=>"101101111",
  60683=>"100110110",
  60684=>"100000001",
  60685=>"111000000",
  60686=>"110100100",
  60687=>"110000111",
  60688=>"011101011",
  60689=>"011011001",
  60690=>"100001011",
  60691=>"100101111",
  60692=>"001110100",
  60693=>"000000001",
  60694=>"010100010",
  60695=>"110100000",
  60696=>"100111000",
  60697=>"111000101",
  60698=>"100101010",
  60699=>"000101011",
  60700=>"001111011",
  60701=>"111010100",
  60702=>"110100010",
  60703=>"000100110",
  60704=>"000110101",
  60705=>"110110100",
  60706=>"010110111",
  60707=>"001011101",
  60708=>"010110001",
  60709=>"100111001",
  60710=>"000001101",
  60711=>"100100001",
  60712=>"110001100",
  60713=>"100000111",
  60714=>"000010010",
  60715=>"010111010",
  60716=>"110100011",
  60717=>"100001000",
  60718=>"000000011",
  60719=>"011010011",
  60720=>"110011100",
  60721=>"001110010",
  60722=>"010010000",
  60723=>"011001100",
  60724=>"010101111",
  60725=>"011101000",
  60726=>"111000110",
  60727=>"101111001",
  60728=>"111000001",
  60729=>"011110010",
  60730=>"111101010",
  60731=>"001111011",
  60732=>"100111011",
  60733=>"100111001",
  60734=>"111011111",
  60735=>"011100000",
  60736=>"100010001",
  60737=>"111111010",
  60738=>"101001010",
  60739=>"111100110",
  60740=>"011110101",
  60741=>"011101110",
  60742=>"001100100",
  60743=>"111101111",
  60744=>"000011110",
  60745=>"111101101",
  60746=>"011111011",
  60747=>"100111101",
  60748=>"001010010",
  60749=>"110010000",
  60750=>"100000110",
  60751=>"100110001",
  60752=>"000000011",
  60753=>"010101100",
  60754=>"111010011",
  60755=>"010001000",
  60756=>"000000001",
  60757=>"001101000",
  60758=>"010000110",
  60759=>"010110011",
  60760=>"000101000",
  60761=>"110010000",
  60762=>"010100001",
  60763=>"101000011",
  60764=>"000001101",
  60765=>"111001101",
  60766=>"001000000",
  60767=>"010000000",
  60768=>"011000010",
  60769=>"101010000",
  60770=>"111111101",
  60771=>"001010011",
  60772=>"010011000",
  60773=>"010011111",
  60774=>"001100110",
  60775=>"111111011",
  60776=>"111111001",
  60777=>"000100101",
  60778=>"111101111",
  60779=>"000000100",
  60780=>"110010011",
  60781=>"101110010",
  60782=>"110111100",
  60783=>"111100000",
  60784=>"011111001",
  60785=>"110101011",
  60786=>"101011111",
  60787=>"010001111",
  60788=>"100100101",
  60789=>"100110010",
  60790=>"010010010",
  60791=>"010011101",
  60792=>"111111101",
  60793=>"001110001",
  60794=>"001111110",
  60795=>"000100011",
  60796=>"111000100",
  60797=>"111011011",
  60798=>"101100001",
  60799=>"010000110",
  60800=>"011010101",
  60801=>"100010010",
  60802=>"011101000",
  60803=>"001101001",
  60804=>"011010010",
  60805=>"110010000",
  60806=>"111011010",
  60807=>"110100001",
  60808=>"010101111",
  60809=>"110011100",
  60810=>"110100010",
  60811=>"001000111",
  60812=>"011000000",
  60813=>"000101110",
  60814=>"110001101",
  60815=>"111111010",
  60816=>"101100010",
  60817=>"011001111",
  60818=>"001111111",
  60819=>"110100111",
  60820=>"100000011",
  60821=>"101101111",
  60822=>"101100000",
  60823=>"110011111",
  60824=>"000100101",
  60825=>"111001100",
  60826=>"111000011",
  60827=>"111111000",
  60828=>"010000100",
  60829=>"101110000",
  60830=>"001100101",
  60831=>"101110010",
  60832=>"001100000",
  60833=>"000100001",
  60834=>"100110111",
  60835=>"010100111",
  60836=>"110100011",
  60837=>"110000100",
  60838=>"101011001",
  60839=>"101010011",
  60840=>"111110101",
  60841=>"010000010",
  60842=>"001011000",
  60843=>"000100010",
  60844=>"001011000",
  60845=>"001110011",
  60846=>"101000000",
  60847=>"001010000",
  60848=>"100010001",
  60849=>"101000100",
  60850=>"010001011",
  60851=>"111101111",
  60852=>"100111111",
  60853=>"100010011",
  60854=>"010001110",
  60855=>"001000001",
  60856=>"110111010",
  60857=>"010100100",
  60858=>"100101100",
  60859=>"010110011",
  60860=>"110010101",
  60861=>"101000100",
  60862=>"011011110",
  60863=>"011010010",
  60864=>"111000100",
  60865=>"010000010",
  60866=>"011000000",
  60867=>"110001101",
  60868=>"111001110",
  60869=>"000100010",
  60870=>"001010011",
  60871=>"111001110",
  60872=>"000110111",
  60873=>"001101011",
  60874=>"101000100",
  60875=>"111001011",
  60876=>"110110111",
  60877=>"101111011",
  60878=>"110110110",
  60879=>"000000000",
  60880=>"111101000",
  60881=>"010010101",
  60882=>"110101001",
  60883=>"000001010",
  60884=>"111000101",
  60885=>"001011111",
  60886=>"100000011",
  60887=>"110110010",
  60888=>"110001101",
  60889=>"001111110",
  60890=>"000001011",
  60891=>"111100000",
  60892=>"011111111",
  60893=>"000001101",
  60894=>"001000000",
  60895=>"000110010",
  60896=>"100101010",
  60897=>"110111111",
  60898=>"011101110",
  60899=>"111010001",
  60900=>"011010110",
  60901=>"000101101",
  60902=>"001001100",
  60903=>"111110001",
  60904=>"010111101",
  60905=>"001010110",
  60906=>"100010100",
  60907=>"010001010",
  60908=>"111101000",
  60909=>"100001101",
  60910=>"000001001",
  60911=>"011001110",
  60912=>"111001011",
  60913=>"111110101",
  60914=>"011010001",
  60915=>"111110111",
  60916=>"000110100",
  60917=>"100100111",
  60918=>"111011001",
  60919=>"000101101",
  60920=>"000100000",
  60921=>"110001010",
  60922=>"011101000",
  60923=>"110000100",
  60924=>"110101110",
  60925=>"011111000",
  60926=>"010010100",
  60927=>"111000011",
  60928=>"000010000",
  60929=>"011011100",
  60930=>"110001000",
  60931=>"111011000",
  60932=>"101110111",
  60933=>"100101111",
  60934=>"011000011",
  60935=>"001010000",
  60936=>"010000001",
  60937=>"011110001",
  60938=>"001101110",
  60939=>"001000000",
  60940=>"111100011",
  60941=>"011000111",
  60942=>"000100001",
  60943=>"011111001",
  60944=>"010010000",
  60945=>"110001110",
  60946=>"011011110",
  60947=>"001110100",
  60948=>"110010001",
  60949=>"010000001",
  60950=>"111011101",
  60951=>"001100110",
  60952=>"010110010",
  60953=>"001011111",
  60954=>"110001010",
  60955=>"011010100",
  60956=>"101001101",
  60957=>"001010001",
  60958=>"001010110",
  60959=>"010011010",
  60960=>"000100000",
  60961=>"111000001",
  60962=>"001100011",
  60963=>"000110011",
  60964=>"100011000",
  60965=>"000001010",
  60966=>"001010000",
  60967=>"111100010",
  60968=>"000111000",
  60969=>"110110111",
  60970=>"111011000",
  60971=>"010000011",
  60972=>"010011011",
  60973=>"010010101",
  60974=>"001000111",
  60975=>"000100010",
  60976=>"011101000",
  60977=>"011001100",
  60978=>"001100100",
  60979=>"101001010",
  60980=>"100010011",
  60981=>"000000010",
  60982=>"110111111",
  60983=>"010000101",
  60984=>"000000010",
  60985=>"001110101",
  60986=>"010000011",
  60987=>"110010111",
  60988=>"111010111",
  60989=>"100011100",
  60990=>"101000010",
  60991=>"110101111",
  60992=>"110101010",
  60993=>"000111100",
  60994=>"011010001",
  60995=>"000010100",
  60996=>"011000101",
  60997=>"111110011",
  60998=>"101111011",
  60999=>"001110101",
  61000=>"010011100",
  61001=>"110110000",
  61002=>"110000010",
  61003=>"000110001",
  61004=>"010010001",
  61005=>"110101010",
  61006=>"101100000",
  61007=>"010010000",
  61008=>"111000111",
  61009=>"000001010",
  61010=>"101000101",
  61011=>"010001110",
  61012=>"101110000",
  61013=>"100110100",
  61014=>"001000001",
  61015=>"011111001",
  61016=>"001000111",
  61017=>"110010111",
  61018=>"001101101",
  61019=>"111010101",
  61020=>"110111110",
  61021=>"000101101",
  61022=>"100011001",
  61023=>"101001010",
  61024=>"111000000",
  61025=>"111001100",
  61026=>"111101001",
  61027=>"010000011",
  61028=>"101100111",
  61029=>"111011101",
  61030=>"010101110",
  61031=>"100010010",
  61032=>"010100000",
  61033=>"111111111",
  61034=>"100001011",
  61035=>"100011111",
  61036=>"111101011",
  61037=>"110001110",
  61038=>"010110100",
  61039=>"101110001",
  61040=>"000111000",
  61041=>"011000010",
  61042=>"010010001",
  61043=>"001100100",
  61044=>"100000100",
  61045=>"110000011",
  61046=>"111101110",
  61047=>"110000111",
  61048=>"110001100",
  61049=>"110111101",
  61050=>"011010111",
  61051=>"000100111",
  61052=>"100001000",
  61053=>"010000100",
  61054=>"101101111",
  61055=>"011111110",
  61056=>"100100010",
  61057=>"111111100",
  61058=>"001101000",
  61059=>"010001010",
  61060=>"010111001",
  61061=>"111001010",
  61062=>"000110011",
  61063=>"100000001",
  61064=>"000110100",
  61065=>"110110000",
  61066=>"000100011",
  61067=>"100001111",
  61068=>"010001100",
  61069=>"000100100",
  61070=>"011001010",
  61071=>"010111000",
  61072=>"110001110",
  61073=>"101011011",
  61074=>"011011010",
  61075=>"000010100",
  61076=>"000100100",
  61077=>"011010010",
  61078=>"000101011",
  61079=>"011101100",
  61080=>"011011001",
  61081=>"101011010",
  61082=>"100011000",
  61083=>"100101011",
  61084=>"000110110",
  61085=>"101101110",
  61086=>"111111110",
  61087=>"110100100",
  61088=>"111100110",
  61089=>"111110001",
  61090=>"010110110",
  61091=>"000000000",
  61092=>"110111011",
  61093=>"100000101",
  61094=>"100101000",
  61095=>"000100011",
  61096=>"101011000",
  61097=>"000111010",
  61098=>"001111110",
  61099=>"011000110",
  61100=>"000110100",
  61101=>"100100010",
  61102=>"011000010",
  61103=>"000110000",
  61104=>"101010010",
  61105=>"110101100",
  61106=>"011000010",
  61107=>"111111001",
  61108=>"011011011",
  61109=>"000111011",
  61110=>"000110000",
  61111=>"011011110",
  61112=>"101100111",
  61113=>"111111001",
  61114=>"111010110",
  61115=>"011000000",
  61116=>"111101000",
  61117=>"111000001",
  61118=>"000100111",
  61119=>"100101110",
  61120=>"101010100",
  61121=>"101111001",
  61122=>"111000110",
  61123=>"010100010",
  61124=>"010111011",
  61125=>"111100000",
  61126=>"100101110",
  61127=>"011000011",
  61128=>"011111001",
  61129=>"100110011",
  61130=>"011011011",
  61131=>"100110000",
  61132=>"101111110",
  61133=>"010110001",
  61134=>"101100010",
  61135=>"011011101",
  61136=>"110011111",
  61137=>"111110000",
  61138=>"000110101",
  61139=>"001011001",
  61140=>"010100010",
  61141=>"011011111",
  61142=>"101000000",
  61143=>"010110000",
  61144=>"100101010",
  61145=>"011001010",
  61146=>"001000100",
  61147=>"000001010",
  61148=>"000101111",
  61149=>"011101101",
  61150=>"000010110",
  61151=>"001011000",
  61152=>"001011111",
  61153=>"100010111",
  61154=>"110001110",
  61155=>"010001001",
  61156=>"101110101",
  61157=>"011110110",
  61158=>"001011001",
  61159=>"010000100",
  61160=>"101100001",
  61161=>"001010000",
  61162=>"110111100",
  61163=>"111111000",
  61164=>"000000001",
  61165=>"000101001",
  61166=>"001011000",
  61167=>"000000010",
  61168=>"110000001",
  61169=>"100100110",
  61170=>"010000100",
  61171=>"000000000",
  61172=>"001001000",
  61173=>"011111101",
  61174=>"010100100",
  61175=>"100001000",
  61176=>"010011001",
  61177=>"101101111",
  61178=>"010110010",
  61179=>"001001101",
  61180=>"101000000",
  61181=>"110000011",
  61182=>"001101001",
  61183=>"001010000",
  61184=>"011110001",
  61185=>"110100100",
  61186=>"000100100",
  61187=>"010101101",
  61188=>"000111011",
  61189=>"101000001",
  61190=>"110111000",
  61191=>"000011011",
  61192=>"010101000",
  61193=>"101010010",
  61194=>"000101100",
  61195=>"101010001",
  61196=>"010100101",
  61197=>"110110001",
  61198=>"110101010",
  61199=>"101010000",
  61200=>"101100000",
  61201=>"100110011",
  61202=>"000010110",
  61203=>"000101111",
  61204=>"101000001",
  61205=>"101000010",
  61206=>"010010001",
  61207=>"110010000",
  61208=>"001010101",
  61209=>"010011000",
  61210=>"001101011",
  61211=>"010000100",
  61212=>"100000000",
  61213=>"010111100",
  61214=>"110011100",
  61215=>"011010111",
  61216=>"101100010",
  61217=>"100011001",
  61218=>"000101011",
  61219=>"000001101",
  61220=>"001000100",
  61221=>"100110101",
  61222=>"100011111",
  61223=>"010110110",
  61224=>"111000111",
  61225=>"011000100",
  61226=>"011010111",
  61227=>"111010111",
  61228=>"100010010",
  61229=>"000010100",
  61230=>"011111010",
  61231=>"001000101",
  61232=>"011010010",
  61233=>"100100011",
  61234=>"001011001",
  61235=>"000000100",
  61236=>"110101000",
  61237=>"011010011",
  61238=>"111001100",
  61239=>"101000011",
  61240=>"000000001",
  61241=>"011101101",
  61242=>"100110010",
  61243=>"000100101",
  61244=>"000000000",
  61245=>"101111111",
  61246=>"111001010",
  61247=>"111010101",
  61248=>"110000110",
  61249=>"001000110",
  61250=>"100111101",
  61251=>"110011010",
  61252=>"110100111",
  61253=>"000100100",
  61254=>"011000111",
  61255=>"101111111",
  61256=>"000001100",
  61257=>"010011110",
  61258=>"011101111",
  61259=>"010110011",
  61260=>"001110010",
  61261=>"110011111",
  61262=>"000100001",
  61263=>"011000001",
  61264=>"101000111",
  61265=>"011100000",
  61266=>"001001010",
  61267=>"010000100",
  61268=>"110111110",
  61269=>"100010111",
  61270=>"010101001",
  61271=>"010111111",
  61272=>"101111110",
  61273=>"011001101",
  61274=>"011001110",
  61275=>"001000001",
  61276=>"111010110",
  61277=>"101010010",
  61278=>"100011111",
  61279=>"101101101",
  61280=>"100010101",
  61281=>"111101100",
  61282=>"001101111",
  61283=>"111101101",
  61284=>"011011101",
  61285=>"010010010",
  61286=>"110100111",
  61287=>"110001101",
  61288=>"100001010",
  61289=>"110111010",
  61290=>"001010010",
  61291=>"011001010",
  61292=>"011101101",
  61293=>"100011000",
  61294=>"000100000",
  61295=>"010011110",
  61296=>"001000011",
  61297=>"001100110",
  61298=>"101010110",
  61299=>"100011111",
  61300=>"101100110",
  61301=>"110000010",
  61302=>"111100000",
  61303=>"010100001",
  61304=>"101011000",
  61305=>"101110101",
  61306=>"000000101",
  61307=>"010010010",
  61308=>"100100111",
  61309=>"011111100",
  61310=>"000100010",
  61311=>"001000110",
  61312=>"101011101",
  61313=>"100100001",
  61314=>"101100010",
  61315=>"110100101",
  61316=>"001111010",
  61317=>"000111110",
  61318=>"110100000",
  61319=>"100011011",
  61320=>"001001101",
  61321=>"010000001",
  61322=>"000010100",
  61323=>"101001010",
  61324=>"001001011",
  61325=>"010110110",
  61326=>"101101010",
  61327=>"100011110",
  61328=>"011100101",
  61329=>"010001111",
  61330=>"101100001",
  61331=>"000000101",
  61332=>"100000110",
  61333=>"000101100",
  61334=>"111011100",
  61335=>"000110011",
  61336=>"111101101",
  61337=>"010001011",
  61338=>"010011111",
  61339=>"001111110",
  61340=>"000000001",
  61341=>"001000010",
  61342=>"100101000",
  61343=>"000010010",
  61344=>"100011100",
  61345=>"011010101",
  61346=>"011011000",
  61347=>"110001000",
  61348=>"000100101",
  61349=>"100011011",
  61350=>"110011101",
  61351=>"010101111",
  61352=>"000110101",
  61353=>"101111111",
  61354=>"001011101",
  61355=>"010110110",
  61356=>"011001110",
  61357=>"110010111",
  61358=>"001101001",
  61359=>"101001111",
  61360=>"101110111",
  61361=>"011010011",
  61362=>"010110111",
  61363=>"100110000",
  61364=>"000011111",
  61365=>"110110111",
  61366=>"011011001",
  61367=>"110111000",
  61368=>"110011011",
  61369=>"001010111",
  61370=>"101010110",
  61371=>"010000110",
  61372=>"100011001",
  61373=>"111011101",
  61374=>"010000110",
  61375=>"110000111",
  61376=>"111101001",
  61377=>"101001001",
  61378=>"000111001",
  61379=>"000000010",
  61380=>"001111101",
  61381=>"100010110",
  61382=>"111100111",
  61383=>"110000010",
  61384=>"000000111",
  61385=>"010100110",
  61386=>"110101110",
  61387=>"001001110",
  61388=>"101010101",
  61389=>"010001000",
  61390=>"001010100",
  61391=>"111010100",
  61392=>"011011110",
  61393=>"010110110",
  61394=>"110011111",
  61395=>"101111000",
  61396=>"001000111",
  61397=>"011111000",
  61398=>"001110000",
  61399=>"010101011",
  61400=>"000000001",
  61401=>"100101110",
  61402=>"001101001",
  61403=>"000000100",
  61404=>"000110111",
  61405=>"001110010",
  61406=>"011100010",
  61407=>"010110000",
  61408=>"101110111",
  61409=>"001000000",
  61410=>"000101100",
  61411=>"000100111",
  61412=>"111011001",
  61413=>"001001110",
  61414=>"011000001",
  61415=>"000011010",
  61416=>"011111101",
  61417=>"101010111",
  61418=>"010000110",
  61419=>"101100100",
  61420=>"011101101",
  61421=>"101101111",
  61422=>"010010111",
  61423=>"111011111",
  61424=>"111111011",
  61425=>"110111011",
  61426=>"101100111",
  61427=>"000000010",
  61428=>"100011101",
  61429=>"010001010",
  61430=>"001000101",
  61431=>"010000010",
  61432=>"001010000",
  61433=>"100111111",
  61434=>"100100001",
  61435=>"111000000",
  61436=>"111001010",
  61437=>"100100011",
  61438=>"000011010",
  61439=>"010000100",
  61440=>"110011001",
  61441=>"111001001",
  61442=>"111010111",
  61443=>"001001000",
  61444=>"001110101",
  61445=>"011001110",
  61446=>"111010000",
  61447=>"110011111",
  61448=>"001101011",
  61449=>"001100111",
  61450=>"111010010",
  61451=>"010111111",
  61452=>"001000110",
  61453=>"000101001",
  61454=>"011100110",
  61455=>"001000100",
  61456=>"100000000",
  61457=>"011010100",
  61458=>"000010011",
  61459=>"010111100",
  61460=>"000000001",
  61461=>"111011110",
  61462=>"010001011",
  61463=>"011000011",
  61464=>"101001111",
  61465=>"101101101",
  61466=>"111111001",
  61467=>"011101010",
  61468=>"101110110",
  61469=>"001000010",
  61470=>"110010010",
  61471=>"000000010",
  61472=>"011010010",
  61473=>"101111111",
  61474=>"011011001",
  61475=>"101011111",
  61476=>"110101110",
  61477=>"011011100",
  61478=>"001001100",
  61479=>"111011111",
  61480=>"010001001",
  61481=>"111000000",
  61482=>"110100110",
  61483=>"000101101",
  61484=>"101001010",
  61485=>"000110111",
  61486=>"000011010",
  61487=>"000101111",
  61488=>"001011101",
  61489=>"110001110",
  61490=>"000001100",
  61491=>"011000101",
  61492=>"100000110",
  61493=>"011000000",
  61494=>"100101101",
  61495=>"100001111",
  61496=>"101011011",
  61497=>"001011010",
  61498=>"110111101",
  61499=>"110111011",
  61500=>"110001001",
  61501=>"010000110",
  61502=>"011001111",
  61503=>"000101011",
  61504=>"011111000",
  61505=>"000001100",
  61506=>"100000001",
  61507=>"110010000",
  61508=>"110001001",
  61509=>"000001010",
  61510=>"111100111",
  61511=>"111110000",
  61512=>"011011001",
  61513=>"110111000",
  61514=>"010010110",
  61515=>"010011001",
  61516=>"101110101",
  61517=>"111101011",
  61518=>"100110010",
  61519=>"110110001",
  61520=>"110100010",
  61521=>"000111100",
  61522=>"001001010",
  61523=>"100110101",
  61524=>"111011000",
  61525=>"001000000",
  61526=>"001011101",
  61527=>"000000101",
  61528=>"110011000",
  61529=>"001011111",
  61530=>"011000100",
  61531=>"010010101",
  61532=>"000010011",
  61533=>"001110110",
  61534=>"101111001",
  61535=>"011011001",
  61536=>"100100000",
  61537=>"100010110",
  61538=>"000000110",
  61539=>"011000001",
  61540=>"100010010",
  61541=>"000000111",
  61542=>"010100000",
  61543=>"000101000",
  61544=>"110101110",
  61545=>"011110000",
  61546=>"010111010",
  61547=>"110000100",
  61548=>"000011000",
  61549=>"001100010",
  61550=>"110111011",
  61551=>"101010101",
  61552=>"000111100",
  61553=>"100000001",
  61554=>"011100110",
  61555=>"110101000",
  61556=>"111010011",
  61557=>"010001110",
  61558=>"100000000",
  61559=>"000101101",
  61560=>"110110110",
  61561=>"111010110",
  61562=>"000101010",
  61563=>"001100011",
  61564=>"001100101",
  61565=>"110000100",
  61566=>"110110000",
  61567=>"100000011",
  61568=>"101001111",
  61569=>"100101101",
  61570=>"010101111",
  61571=>"010001101",
  61572=>"100101110",
  61573=>"000010110",
  61574=>"100110001",
  61575=>"000110100",
  61576=>"000011010",
  61577=>"101000010",
  61578=>"000101100",
  61579=>"011111110",
  61580=>"001110000",
  61581=>"100110000",
  61582=>"100101010",
  61583=>"111110101",
  61584=>"000000011",
  61585=>"001110110",
  61586=>"000001000",
  61587=>"000001000",
  61588=>"011000000",
  61589=>"010100111",
  61590=>"111101001",
  61591=>"011010001",
  61592=>"001101110",
  61593=>"111001001",
  61594=>"100111010",
  61595=>"101111100",
  61596=>"010111100",
  61597=>"100101100",
  61598=>"110000111",
  61599=>"100101000",
  61600=>"100001111",
  61601=>"011000110",
  61602=>"100100101",
  61603=>"100101001",
  61604=>"101011111",
  61605=>"110011011",
  61606=>"110000000",
  61607=>"001101100",
  61608=>"001111001",
  61609=>"001010101",
  61610=>"011110110",
  61611=>"111111101",
  61612=>"101011111",
  61613=>"010111111",
  61614=>"110001101",
  61615=>"010000111",
  61616=>"101010001",
  61617=>"000110010",
  61618=>"100100110",
  61619=>"010101110",
  61620=>"101011000",
  61621=>"110110010",
  61622=>"110010011",
  61623=>"101010100",
  61624=>"110000101",
  61625=>"111100000",
  61626=>"010011010",
  61627=>"010100010",
  61628=>"010010110",
  61629=>"011100110",
  61630=>"011101011",
  61631=>"011001100",
  61632=>"100010100",
  61633=>"000010000",
  61634=>"000011000",
  61635=>"110000000",
  61636=>"001100010",
  61637=>"011011001",
  61638=>"001101100",
  61639=>"110101010",
  61640=>"010000011",
  61641=>"010000011",
  61642=>"011010111",
  61643=>"110100010",
  61644=>"011101001",
  61645=>"010010001",
  61646=>"010000100",
  61647=>"001011001",
  61648=>"100111011",
  61649=>"000111000",
  61650=>"001100011",
  61651=>"111000010",
  61652=>"010010010",
  61653=>"000101010",
  61654=>"011010111",
  61655=>"000000011",
  61656=>"111001100",
  61657=>"110101001",
  61658=>"000000011",
  61659=>"001010001",
  61660=>"111000000",
  61661=>"011111010",
  61662=>"101011101",
  61663=>"001010101",
  61664=>"101100110",
  61665=>"010000110",
  61666=>"010000100",
  61667=>"000000000",
  61668=>"010110100",
  61669=>"110101100",
  61670=>"000100101",
  61671=>"100011000",
  61672=>"101011011",
  61673=>"010010101",
  61674=>"011010001",
  61675=>"010111011",
  61676=>"100101110",
  61677=>"000000000",
  61678=>"010010011",
  61679=>"100000110",
  61680=>"010101010",
  61681=>"101111011",
  61682=>"100110001",
  61683=>"000000001",
  61684=>"100010011",
  61685=>"110000100",
  61686=>"011111000",
  61687=>"110001111",
  61688=>"110110001",
  61689=>"111001110",
  61690=>"100101000",
  61691=>"111010111",
  61692=>"011111101",
  61693=>"011100110",
  61694=>"111110101",
  61695=>"010000001",
  61696=>"000010110",
  61697=>"010100001",
  61698=>"101011100",
  61699=>"100100111",
  61700=>"101111001",
  61701=>"001100111",
  61702=>"001010111",
  61703=>"110101100",
  61704=>"000001010",
  61705=>"001010000",
  61706=>"001000000",
  61707=>"110110010",
  61708=>"000100100",
  61709=>"011100101",
  61710=>"100101011",
  61711=>"011111010",
  61712=>"011110000",
  61713=>"011111011",
  61714=>"110101100",
  61715=>"100111010",
  61716=>"000100000",
  61717=>"000000100",
  61718=>"010100100",
  61719=>"000101000",
  61720=>"110111010",
  61721=>"010100111",
  61722=>"111110000",
  61723=>"111110111",
  61724=>"011000000",
  61725=>"100010001",
  61726=>"011111110",
  61727=>"011001000",
  61728=>"010010111",
  61729=>"110001000",
  61730=>"001001011",
  61731=>"110100111",
  61732=>"001101110",
  61733=>"000101111",
  61734=>"110100100",
  61735=>"101100011",
  61736=>"001011010",
  61737=>"001110001",
  61738=>"101100110",
  61739=>"001110010",
  61740=>"011000100",
  61741=>"010001001",
  61742=>"011010010",
  61743=>"111000101",
  61744=>"000001110",
  61745=>"010010000",
  61746=>"111111111",
  61747=>"110110101",
  61748=>"110000100",
  61749=>"000110100",
  61750=>"011111101",
  61751=>"001100001",
  61752=>"011000100",
  61753=>"111010110",
  61754=>"111110010",
  61755=>"111101100",
  61756=>"111110011",
  61757=>"110111101",
  61758=>"100010110",
  61759=>"101001101",
  61760=>"000100110",
  61761=>"110100000",
  61762=>"101100100",
  61763=>"001111001",
  61764=>"101000010",
  61765=>"101111110",
  61766=>"100010110",
  61767=>"100101000",
  61768=>"000100110",
  61769=>"011010101",
  61770=>"011011101",
  61771=>"101100100",
  61772=>"010011000",
  61773=>"010000100",
  61774=>"100110011",
  61775=>"010001101",
  61776=>"010110000",
  61777=>"101111101",
  61778=>"001000000",
  61779=>"001100110",
  61780=>"001111000",
  61781=>"101111000",
  61782=>"110010010",
  61783=>"010111100",
  61784=>"101110011",
  61785=>"000010100",
  61786=>"001010110",
  61787=>"010010010",
  61788=>"001010000",
  61789=>"100101101",
  61790=>"100101001",
  61791=>"011010001",
  61792=>"011010000",
  61793=>"011111111",
  61794=>"110000000",
  61795=>"001010011",
  61796=>"000001101",
  61797=>"000000010",
  61798=>"111000001",
  61799=>"100000011",
  61800=>"001010110",
  61801=>"001111101",
  61802=>"100010111",
  61803=>"000011110",
  61804=>"100010000",
  61805=>"111100111",
  61806=>"001000111",
  61807=>"100011010",
  61808=>"000100000",
  61809=>"100001010",
  61810=>"001110001",
  61811=>"010100000",
  61812=>"011101110",
  61813=>"101101101",
  61814=>"111110001",
  61815=>"000111000",
  61816=>"100100101",
  61817=>"110011001",
  61818=>"101100111",
  61819=>"010110010",
  61820=>"111100101",
  61821=>"011110100",
  61822=>"110000001",
  61823=>"111000110",
  61824=>"001101100",
  61825=>"110000001",
  61826=>"111111011",
  61827=>"000110111",
  61828=>"000001111",
  61829=>"001110001",
  61830=>"010000011",
  61831=>"110111001",
  61832=>"010110000",
  61833=>"101000100",
  61834=>"110110111",
  61835=>"110110011",
  61836=>"110111010",
  61837=>"111111001",
  61838=>"000010000",
  61839=>"011011100",
  61840=>"100100111",
  61841=>"010000100",
  61842=>"101110100",
  61843=>"101010111",
  61844=>"100110100",
  61845=>"100100101",
  61846=>"010000001",
  61847=>"001110010",
  61848=>"000111111",
  61849=>"001100110",
  61850=>"110101001",
  61851=>"000011110",
  61852=>"101110001",
  61853=>"110110001",
  61854=>"001010011",
  61855=>"101101111",
  61856=>"011111111",
  61857=>"100100101",
  61858=>"011000000",
  61859=>"110000111",
  61860=>"000000011",
  61861=>"100111000",
  61862=>"000000000",
  61863=>"000100001",
  61864=>"111101111",
  61865=>"001000100",
  61866=>"101000000",
  61867=>"110100011",
  61868=>"000101111",
  61869=>"001100011",
  61870=>"110111000",
  61871=>"111011110",
  61872=>"000010001",
  61873=>"000110111",
  61874=>"110101011",
  61875=>"000000000",
  61876=>"111111001",
  61877=>"001001111",
  61878=>"010011000",
  61879=>"000100000",
  61880=>"011010100",
  61881=>"001010100",
  61882=>"000010001",
  61883=>"100111111",
  61884=>"111000100",
  61885=>"101011101",
  61886=>"000000001",
  61887=>"111110010",
  61888=>"011000111",
  61889=>"001010011",
  61890=>"111110100",
  61891=>"001110001",
  61892=>"000110101",
  61893=>"011101010",
  61894=>"110111101",
  61895=>"010010100",
  61896=>"100101000",
  61897=>"101000100",
  61898=>"110001000",
  61899=>"101010010",
  61900=>"010011100",
  61901=>"011100110",
  61902=>"100110100",
  61903=>"100000111",
  61904=>"111111001",
  61905=>"000110100",
  61906=>"001111010",
  61907=>"001110110",
  61908=>"010001110",
  61909=>"011101000",
  61910=>"100100100",
  61911=>"000000110",
  61912=>"000011010",
  61913=>"110000001",
  61914=>"111011010",
  61915=>"001010101",
  61916=>"111100001",
  61917=>"111110111",
  61918=>"001001011",
  61919=>"001010001",
  61920=>"101111000",
  61921=>"111111000",
  61922=>"110111010",
  61923=>"001101111",
  61924=>"100110100",
  61925=>"110111000",
  61926=>"001100101",
  61927=>"101111001",
  61928=>"011001111",
  61929=>"011101000",
  61930=>"000010110",
  61931=>"010100110",
  61932=>"110010100",
  61933=>"110100010",
  61934=>"000000100",
  61935=>"100010010",
  61936=>"100110010",
  61937=>"111101011",
  61938=>"001100101",
  61939=>"111010001",
  61940=>"001110010",
  61941=>"001100110",
  61942=>"011001110",
  61943=>"101111001",
  61944=>"101101001",
  61945=>"111100001",
  61946=>"001011110",
  61947=>"100001000",
  61948=>"101100000",
  61949=>"100100010",
  61950=>"110110011",
  61951=>"100000010",
  61952=>"000000111",
  61953=>"010010111",
  61954=>"111011101",
  61955=>"001100100",
  61956=>"100000111",
  61957=>"001110000",
  61958=>"011111110",
  61959=>"011101110",
  61960=>"010010100",
  61961=>"011000111",
  61962=>"110110000",
  61963=>"000101101",
  61964=>"000110110",
  61965=>"010101011",
  61966=>"100100000",
  61967=>"110000101",
  61968=>"101100110",
  61969=>"110000011",
  61970=>"101001111",
  61971=>"010100000",
  61972=>"000110000",
  61973=>"001000100",
  61974=>"101101100",
  61975=>"101001001",
  61976=>"001110010",
  61977=>"110010000",
  61978=>"101000100",
  61979=>"110000010",
  61980=>"000100101",
  61981=>"001101101",
  61982=>"100111110",
  61983=>"001100100",
  61984=>"101110100",
  61985=>"111101101",
  61986=>"010100111",
  61987=>"110010101",
  61988=>"100111000",
  61989=>"000110011",
  61990=>"000100001",
  61991=>"110100100",
  61992=>"110100000",
  61993=>"011110000",
  61994=>"111000111",
  61995=>"100101000",
  61996=>"100111100",
  61997=>"110010100",
  61998=>"011101100",
  61999=>"110100101",
  62000=>"110111010",
  62001=>"011011100",
  62002=>"100010111",
  62003=>"111001011",
  62004=>"010110101",
  62005=>"111110011",
  62006=>"101100101",
  62007=>"010000011",
  62008=>"101001001",
  62009=>"010011100",
  62010=>"010100000",
  62011=>"000011010",
  62012=>"010010010",
  62013=>"110000001",
  62014=>"110100110",
  62015=>"011100000",
  62016=>"010100010",
  62017=>"000011100",
  62018=>"100010111",
  62019=>"010101110",
  62020=>"011000101",
  62021=>"100101011",
  62022=>"101110101",
  62023=>"110010000",
  62024=>"001010011",
  62025=>"000101010",
  62026=>"100110100",
  62027=>"000110000",
  62028=>"110011111",
  62029=>"000100111",
  62030=>"010110111",
  62031=>"110000011",
  62032=>"100001110",
  62033=>"011111101",
  62034=>"000111000",
  62035=>"101111000",
  62036=>"001000000",
  62037=>"101101101",
  62038=>"011010101",
  62039=>"110111111",
  62040=>"011111100",
  62041=>"111111110",
  62042=>"111110111",
  62043=>"101011000",
  62044=>"000100011",
  62045=>"100110100",
  62046=>"111101000",
  62047=>"101100000",
  62048=>"101100001",
  62049=>"010100010",
  62050=>"000111110",
  62051=>"100010111",
  62052=>"111100101",
  62053=>"011100001",
  62054=>"111111001",
  62055=>"010111010",
  62056=>"000101110",
  62057=>"110100000",
  62058=>"011110010",
  62059=>"000001011",
  62060=>"010001100",
  62061=>"010011111",
  62062=>"000010010",
  62063=>"100111100",
  62064=>"100100001",
  62065=>"000100011",
  62066=>"011110101",
  62067=>"100010110",
  62068=>"100110101",
  62069=>"010110010",
  62070=>"101101001",
  62071=>"001110101",
  62072=>"010011011",
  62073=>"100101100",
  62074=>"101011011",
  62075=>"000111111",
  62076=>"100100100",
  62077=>"110101010",
  62078=>"011110110",
  62079=>"100000011",
  62080=>"111110110",
  62081=>"110011110",
  62082=>"111100100",
  62083=>"111101100",
  62084=>"000110110",
  62085=>"100101101",
  62086=>"000110011",
  62087=>"101100000",
  62088=>"111000001",
  62089=>"011000111",
  62090=>"100011111",
  62091=>"011011000",
  62092=>"011100100",
  62093=>"110001100",
  62094=>"111011001",
  62095=>"001011001",
  62096=>"000011000",
  62097=>"001100010",
  62098=>"010101100",
  62099=>"011001101",
  62100=>"010100001",
  62101=>"010010110",
  62102=>"101100010",
  62103=>"001011001",
  62104=>"110001111",
  62105=>"000110011",
  62106=>"101111111",
  62107=>"001110100",
  62108=>"111000000",
  62109=>"111001100",
  62110=>"010111100",
  62111=>"101111111",
  62112=>"100010111",
  62113=>"101001101",
  62114=>"010100000",
  62115=>"000100000",
  62116=>"011100111",
  62117=>"111001100",
  62118=>"110010000",
  62119=>"110010011",
  62120=>"001001001",
  62121=>"011010010",
  62122=>"001110000",
  62123=>"001010000",
  62124=>"101011010",
  62125=>"100000000",
  62126=>"001011011",
  62127=>"101010001",
  62128=>"010011000",
  62129=>"100100111",
  62130=>"111000000",
  62131=>"000100000",
  62132=>"000000101",
  62133=>"101110100",
  62134=>"101100000",
  62135=>"111111000",
  62136=>"010000100",
  62137=>"110010111",
  62138=>"001011111",
  62139=>"111100000",
  62140=>"101101110",
  62141=>"101010001",
  62142=>"110000101",
  62143=>"010111101",
  62144=>"011010011",
  62145=>"001011101",
  62146=>"000100010",
  62147=>"100100001",
  62148=>"011001111",
  62149=>"100100100",
  62150=>"110000100",
  62151=>"000011110",
  62152=>"111101110",
  62153=>"000000000",
  62154=>"110001000",
  62155=>"010111010",
  62156=>"110011101",
  62157=>"110100110",
  62158=>"000100101",
  62159=>"000100101",
  62160=>"110111110",
  62161=>"111101011",
  62162=>"000011101",
  62163=>"010000011",
  62164=>"111101101",
  62165=>"000101011",
  62166=>"010111010",
  62167=>"001110111",
  62168=>"000010010",
  62169=>"011100000",
  62170=>"000000100",
  62171=>"011000010",
  62172=>"101101001",
  62173=>"101001111",
  62174=>"101110101",
  62175=>"001001110",
  62176=>"100000001",
  62177=>"010101001",
  62178=>"011000000",
  62179=>"000010101",
  62180=>"000000011",
  62181=>"110100110",
  62182=>"110000110",
  62183=>"100000101",
  62184=>"010010010",
  62185=>"101111101",
  62186=>"000001111",
  62187=>"110110101",
  62188=>"100001000",
  62189=>"100110000",
  62190=>"011011001",
  62191=>"101000100",
  62192=>"000100010",
  62193=>"110100010",
  62194=>"000010001",
  62195=>"110001011",
  62196=>"101011110",
  62197=>"111100000",
  62198=>"000000100",
  62199=>"110100011",
  62200=>"101101111",
  62201=>"000011001",
  62202=>"010100101",
  62203=>"001001101",
  62204=>"011011000",
  62205=>"111100101",
  62206=>"010001101",
  62207=>"001011111",
  62208=>"010111111",
  62209=>"101110011",
  62210=>"110101110",
  62211=>"101001101",
  62212=>"110111110",
  62213=>"010000100",
  62214=>"001101001",
  62215=>"011011110",
  62216=>"001101010",
  62217=>"010101111",
  62218=>"110001101",
  62219=>"110101110",
  62220=>"001001101",
  62221=>"010000001",
  62222=>"011001001",
  62223=>"111101110",
  62224=>"000011011",
  62225=>"100100100",
  62226=>"000010110",
  62227=>"110101110",
  62228=>"110010001",
  62229=>"101011110",
  62230=>"100000011",
  62231=>"000010101",
  62232=>"010011011",
  62233=>"001101001",
  62234=>"010010001",
  62235=>"110010111",
  62236=>"100011001",
  62237=>"110101011",
  62238=>"111100100",
  62239=>"010100010",
  62240=>"110110110",
  62241=>"001011001",
  62242=>"111110110",
  62243=>"000000110",
  62244=>"100010001",
  62245=>"101110100",
  62246=>"100000110",
  62247=>"000100110",
  62248=>"100100111",
  62249=>"111110011",
  62250=>"010100111",
  62251=>"011110100",
  62252=>"110101000",
  62253=>"100010100",
  62254=>"000000011",
  62255=>"000101000",
  62256=>"000100111",
  62257=>"110001000",
  62258=>"000001100",
  62259=>"101100111",
  62260=>"110111110",
  62261=>"101111100",
  62262=>"010100000",
  62263=>"110001011",
  62264=>"011111101",
  62265=>"001111100",
  62266=>"011001000",
  62267=>"000101000",
  62268=>"000111010",
  62269=>"010011001",
  62270=>"111100101",
  62271=>"011100010",
  62272=>"010000000",
  62273=>"000011010",
  62274=>"001011011",
  62275=>"100100100",
  62276=>"111100001",
  62277=>"111011101",
  62278=>"011000001",
  62279=>"100000000",
  62280=>"000000101",
  62281=>"100011000",
  62282=>"000111111",
  62283=>"001110110",
  62284=>"111101010",
  62285=>"111011010",
  62286=>"011111100",
  62287=>"101000111",
  62288=>"000111001",
  62289=>"111010110",
  62290=>"100100000",
  62291=>"101111100",
  62292=>"101010000",
  62293=>"100011100",
  62294=>"011100001",
  62295=>"110010000",
  62296=>"011101100",
  62297=>"111110110",
  62298=>"110110001",
  62299=>"000111000",
  62300=>"100010011",
  62301=>"101100100",
  62302=>"000010001",
  62303=>"001000110",
  62304=>"111001110",
  62305=>"111001000",
  62306=>"000000000",
  62307=>"010001010",
  62308=>"010000110",
  62309=>"111110010",
  62310=>"111101110",
  62311=>"111111100",
  62312=>"000000100",
  62313=>"011101101",
  62314=>"011010100",
  62315=>"111111010",
  62316=>"111010101",
  62317=>"011011010",
  62318=>"111111100",
  62319=>"010011010",
  62320=>"001000100",
  62321=>"010001010",
  62322=>"001011000",
  62323=>"001010101",
  62324=>"010001001",
  62325=>"011110000",
  62326=>"111010010",
  62327=>"010011001",
  62328=>"010010111",
  62329=>"000110001",
  62330=>"100110110",
  62331=>"100111111",
  62332=>"100010000",
  62333=>"110001110",
  62334=>"010001110",
  62335=>"011011111",
  62336=>"011001110",
  62337=>"110011101",
  62338=>"001100100",
  62339=>"010100111",
  62340=>"011000000",
  62341=>"010001111",
  62342=>"000100000",
  62343=>"101010100",
  62344=>"101001001",
  62345=>"111111100",
  62346=>"000001001",
  62347=>"000101100",
  62348=>"011100001",
  62349=>"111100010",
  62350=>"111001110",
  62351=>"110011000",
  62352=>"010100100",
  62353=>"101000110",
  62354=>"110001000",
  62355=>"111110111",
  62356=>"101000000",
  62357=>"001000101",
  62358=>"110101011",
  62359=>"011101101",
  62360=>"000000001",
  62361=>"100111100",
  62362=>"101110110",
  62363=>"111111101",
  62364=>"100000010",
  62365=>"011010000",
  62366=>"001110000",
  62367=>"001101010",
  62368=>"001101110",
  62369=>"000011000",
  62370=>"011111010",
  62371=>"100110111",
  62372=>"011011100",
  62373=>"001010100",
  62374=>"001011000",
  62375=>"110011001",
  62376=>"011111000",
  62377=>"110010001",
  62378=>"111001110",
  62379=>"101001011",
  62380=>"001111110",
  62381=>"101110001",
  62382=>"101111000",
  62383=>"110010111",
  62384=>"110010000",
  62385=>"111111001",
  62386=>"001101110",
  62387=>"110011101",
  62388=>"011100010",
  62389=>"000100011",
  62390=>"100000111",
  62391=>"001110100",
  62392=>"001001000",
  62393=>"110110110",
  62394=>"101010011",
  62395=>"111110111",
  62396=>"001101111",
  62397=>"001110100",
  62398=>"111100100",
  62399=>"111110110",
  62400=>"101111111",
  62401=>"101011011",
  62402=>"000000001",
  62403=>"111011001",
  62404=>"011111111",
  62405=>"010001111",
  62406=>"100101001",
  62407=>"101011000",
  62408=>"000100110",
  62409=>"010111000",
  62410=>"000001000",
  62411=>"101101010",
  62412=>"011000101",
  62413=>"001100110",
  62414=>"110001101",
  62415=>"110001101",
  62416=>"111001011",
  62417=>"011000011",
  62418=>"101101111",
  62419=>"101011000",
  62420=>"000001100",
  62421=>"010111100",
  62422=>"001101111",
  62423=>"000100010",
  62424=>"011111000",
  62425=>"001001001",
  62426=>"010101011",
  62427=>"000101101",
  62428=>"110110010",
  62429=>"011111011",
  62430=>"111001100",
  62431=>"111100111",
  62432=>"101001100",
  62433=>"000101000",
  62434=>"000000010",
  62435=>"000100001",
  62436=>"101100000",
  62437=>"010011001",
  62438=>"101110001",
  62439=>"111111100",
  62440=>"000010110",
  62441=>"001010111",
  62442=>"010111101",
  62443=>"110111000",
  62444=>"010001000",
  62445=>"010111101",
  62446=>"101010010",
  62447=>"000000111",
  62448=>"000101000",
  62449=>"001110001",
  62450=>"111010101",
  62451=>"011101101",
  62452=>"100100110",
  62453=>"000010001",
  62454=>"111011100",
  62455=>"000000011",
  62456=>"111101011",
  62457=>"001010010",
  62458=>"011000000",
  62459=>"100001000",
  62460=>"111101000",
  62461=>"100110111",
  62462=>"000100011",
  62463=>"010011001",
  62464=>"000101101",
  62465=>"110101001",
  62466=>"011001010",
  62467=>"011010001",
  62468=>"000101010",
  62469=>"011100101",
  62470=>"000000011",
  62471=>"100100101",
  62472=>"000100000",
  62473=>"101000111",
  62474=>"110100101",
  62475=>"011100001",
  62476=>"000100001",
  62477=>"000000111",
  62478=>"111101111",
  62479=>"000111001",
  62480=>"100010110",
  62481=>"100101101",
  62482=>"111110111",
  62483=>"001010001",
  62484=>"111010011",
  62485=>"111001011",
  62486=>"001111111",
  62487=>"100100100",
  62488=>"010101110",
  62489=>"110011011",
  62490=>"001001010",
  62491=>"010110101",
  62492=>"100100100",
  62493=>"011010110",
  62494=>"100110001",
  62495=>"000101001",
  62496=>"001110011",
  62497=>"101001100",
  62498=>"111011110",
  62499=>"001011100",
  62500=>"110110001",
  62501=>"011100110",
  62502=>"110000001",
  62503=>"100010010",
  62504=>"100001000",
  62505=>"000111000",
  62506=>"001001101",
  62507=>"100100101",
  62508=>"100100010",
  62509=>"011001011",
  62510=>"100101001",
  62511=>"100011111",
  62512=>"110010101",
  62513=>"101011111",
  62514=>"011101111",
  62515=>"000101001",
  62516=>"101001011",
  62517=>"000000001",
  62518=>"001000000",
  62519=>"011010101",
  62520=>"101110011",
  62521=>"100000001",
  62522=>"111000101",
  62523=>"001111001",
  62524=>"110000011",
  62525=>"100110010",
  62526=>"011111111",
  62527=>"010011110",
  62528=>"001110011",
  62529=>"001100000",
  62530=>"011001010",
  62531=>"000110111",
  62532=>"111100001",
  62533=>"110100111",
  62534=>"100010001",
  62535=>"010000110",
  62536=>"101111110",
  62537=>"000100000",
  62538=>"000000010",
  62539=>"000101110",
  62540=>"011110111",
  62541=>"001011000",
  62542=>"110000110",
  62543=>"010100001",
  62544=>"111001100",
  62545=>"100011010",
  62546=>"010111001",
  62547=>"001001000",
  62548=>"010001101",
  62549=>"101100111",
  62550=>"100111111",
  62551=>"000000011",
  62552=>"010111001",
  62553=>"001010011",
  62554=>"101011100",
  62555=>"110111000",
  62556=>"101111111",
  62557=>"111001001",
  62558=>"001000000",
  62559=>"001000011",
  62560=>"111100011",
  62561=>"101001000",
  62562=>"110010101",
  62563=>"000101000",
  62564=>"100000000",
  62565=>"011010100",
  62566=>"101100111",
  62567=>"000111001",
  62568=>"000000111",
  62569=>"101000110",
  62570=>"100000101",
  62571=>"101000100",
  62572=>"111011000",
  62573=>"111111101",
  62574=>"111110010",
  62575=>"111101111",
  62576=>"100110001",
  62577=>"001101111",
  62578=>"100011001",
  62579=>"000010101",
  62580=>"110110110",
  62581=>"110010110",
  62582=>"001011111",
  62583=>"110100001",
  62584=>"001110100",
  62585=>"111000001",
  62586=>"011010011",
  62587=>"010000100",
  62588=>"000100110",
  62589=>"111100000",
  62590=>"100011100",
  62591=>"000011101",
  62592=>"100000010",
  62593=>"001110100",
  62594=>"011001100",
  62595=>"101010111",
  62596=>"011111000",
  62597=>"011001011",
  62598=>"110000110",
  62599=>"101000100",
  62600=>"111010100",
  62601=>"000001001",
  62602=>"101111100",
  62603=>"010111111",
  62604=>"001100100",
  62605=>"100110000",
  62606=>"101101000",
  62607=>"011110110",
  62608=>"001001111",
  62609=>"100110110",
  62610=>"001001000",
  62611=>"000101000",
  62612=>"111010011",
  62613=>"011110100",
  62614=>"001101111",
  62615=>"000010010",
  62616=>"000001001",
  62617=>"011111000",
  62618=>"110001010",
  62619=>"100000011",
  62620=>"001100110",
  62621=>"101111011",
  62622=>"101011110",
  62623=>"101001000",
  62624=>"110101000",
  62625=>"100000110",
  62626=>"000001010",
  62627=>"010100111",
  62628=>"001110111",
  62629=>"000010100",
  62630=>"110111100",
  62631=>"010010011",
  62632=>"100110011",
  62633=>"110001011",
  62634=>"010001111",
  62635=>"111101000",
  62636=>"010001000",
  62637=>"010100010",
  62638=>"000001110",
  62639=>"001000100",
  62640=>"001100001",
  62641=>"100011011",
  62642=>"001001010",
  62643=>"000011010",
  62644=>"001110011",
  62645=>"110110101",
  62646=>"000101110",
  62647=>"110000010",
  62648=>"010100001",
  62649=>"111010000",
  62650=>"100001011",
  62651=>"011011110",
  62652=>"111001001",
  62653=>"000101111",
  62654=>"001011001",
  62655=>"010001110",
  62656=>"110001110",
  62657=>"000011000",
  62658=>"000000010",
  62659=>"001001001",
  62660=>"000101100",
  62661=>"010100001",
  62662=>"010001011",
  62663=>"000000001",
  62664=>"011001110",
  62665=>"011101011",
  62666=>"101101111",
  62667=>"011110100",
  62668=>"010101010",
  62669=>"101101010",
  62670=>"001000001",
  62671=>"111101011",
  62672=>"011011101",
  62673=>"111110001",
  62674=>"100000000",
  62675=>"000100101",
  62676=>"100111111",
  62677=>"110011000",
  62678=>"010111111",
  62679=>"000001001",
  62680=>"000110101",
  62681=>"111100100",
  62682=>"001000001",
  62683=>"011100100",
  62684=>"011000001",
  62685=>"001101111",
  62686=>"100111100",
  62687=>"010010000",
  62688=>"111010011",
  62689=>"110111100",
  62690=>"100100011",
  62691=>"000011000",
  62692=>"000101110",
  62693=>"011001110",
  62694=>"110100000",
  62695=>"010110100",
  62696=>"100111101",
  62697=>"111111101",
  62698=>"010010010",
  62699=>"000001000",
  62700=>"010011101",
  62701=>"101010010",
  62702=>"101101001",
  62703=>"110101000",
  62704=>"101010001",
  62705=>"101000000",
  62706=>"011000000",
  62707=>"001101111",
  62708=>"001010101",
  62709=>"001000111",
  62710=>"111100110",
  62711=>"001101001",
  62712=>"001001010",
  62713=>"110000000",
  62714=>"010001010",
  62715=>"001100101",
  62716=>"110000100",
  62717=>"101000010",
  62718=>"000001001",
  62719=>"010111001",
  62720=>"110011111",
  62721=>"101001001",
  62722=>"011111011",
  62723=>"101101010",
  62724=>"100100001",
  62725=>"000011011",
  62726=>"110111110",
  62727=>"011001101",
  62728=>"110111111",
  62729=>"110110001",
  62730=>"111100001",
  62731=>"011011000",
  62732=>"000101011",
  62733=>"000010110",
  62734=>"101100110",
  62735=>"000101111",
  62736=>"101001000",
  62737=>"011011110",
  62738=>"011011110",
  62739=>"000110110",
  62740=>"001001011",
  62741=>"010101100",
  62742=>"111110111",
  62743=>"001101010",
  62744=>"100000100",
  62745=>"011100100",
  62746=>"100000111",
  62747=>"110110101",
  62748=>"111011111",
  62749=>"111001010",
  62750=>"111101110",
  62751=>"011010010",
  62752=>"011100101",
  62753=>"110010100",
  62754=>"000100001",
  62755=>"001000000",
  62756=>"101001101",
  62757=>"111001001",
  62758=>"111001110",
  62759=>"101011000",
  62760=>"110110000",
  62761=>"011100101",
  62762=>"001101100",
  62763=>"001000111",
  62764=>"100010000",
  62765=>"011000100",
  62766=>"010000011",
  62767=>"111100011",
  62768=>"011101110",
  62769=>"100001010",
  62770=>"000001111",
  62771=>"111001001",
  62772=>"011010010",
  62773=>"000100111",
  62774=>"001000111",
  62775=>"101001001",
  62776=>"010101011",
  62777=>"100011110",
  62778=>"011000110",
  62779=>"101010111",
  62780=>"110001010",
  62781=>"110110110",
  62782=>"110110111",
  62783=>"110011110",
  62784=>"011000000",
  62785=>"011111000",
  62786=>"011011000",
  62787=>"110111000",
  62788=>"000111100",
  62789=>"001011001",
  62790=>"111000000",
  62791=>"010011000",
  62792=>"010111101",
  62793=>"001100010",
  62794=>"101001110",
  62795=>"010001111",
  62796=>"110011101",
  62797=>"111001010",
  62798=>"101000011",
  62799=>"001010001",
  62800=>"110111100",
  62801=>"001001000",
  62802=>"111100001",
  62803=>"100000100",
  62804=>"010010000",
  62805=>"011001111",
  62806=>"101110101",
  62807=>"010001111",
  62808=>"100101001",
  62809=>"101111010",
  62810=>"100110011",
  62811=>"100100110",
  62812=>"001001111",
  62813=>"000101101",
  62814=>"101010011",
  62815=>"100011100",
  62816=>"001010100",
  62817=>"111001101",
  62818=>"000101000",
  62819=>"101011000",
  62820=>"011100001",
  62821=>"101000010",
  62822=>"101000101",
  62823=>"100001001",
  62824=>"100000101",
  62825=>"011111101",
  62826=>"100110101",
  62827=>"101010110",
  62828=>"111000010",
  62829=>"000001001",
  62830=>"000011000",
  62831=>"110111000",
  62832=>"101010011",
  62833=>"000110100",
  62834=>"110101110",
  62835=>"100111110",
  62836=>"000000011",
  62837=>"010000101",
  62838=>"100100000",
  62839=>"100000001",
  62840=>"001111100",
  62841=>"101011110",
  62842=>"110110111",
  62843=>"011010111",
  62844=>"110100000",
  62845=>"011111100",
  62846=>"001110100",
  62847=>"101111111",
  62848=>"000111001",
  62849=>"000001001",
  62850=>"011111001",
  62851=>"000111100",
  62852=>"110010101",
  62853=>"001101101",
  62854=>"110010110",
  62855=>"011010010",
  62856=>"100000101",
  62857=>"010110111",
  62858=>"001000111",
  62859=>"001001000",
  62860=>"110100110",
  62861=>"110101101",
  62862=>"100000110",
  62863=>"100101110",
  62864=>"000101001",
  62865=>"010101000",
  62866=>"100010000",
  62867=>"000111110",
  62868=>"011000100",
  62869=>"100010001",
  62870=>"110001110",
  62871=>"101111111",
  62872=>"001000000",
  62873=>"110100010",
  62874=>"101110000",
  62875=>"100101001",
  62876=>"010011100",
  62877=>"110001110",
  62878=>"001000110",
  62879=>"111100111",
  62880=>"100101101",
  62881=>"001100100",
  62882=>"111100011",
  62883=>"100111101",
  62884=>"101011010",
  62885=>"000000001",
  62886=>"110000011",
  62887=>"110001010",
  62888=>"111010000",
  62889=>"100001100",
  62890=>"011100010",
  62891=>"011110110",
  62892=>"101000110",
  62893=>"001100001",
  62894=>"100000000",
  62895=>"110111111",
  62896=>"000000011",
  62897=>"100101101",
  62898=>"001111110",
  62899=>"010111000",
  62900=>"101100000",
  62901=>"110000001",
  62902=>"111000110",
  62903=>"000110011",
  62904=>"110001110",
  62905=>"100101101",
  62906=>"001001001",
  62907=>"110101110",
  62908=>"100110100",
  62909=>"111111101",
  62910=>"111010101",
  62911=>"101011000",
  62912=>"000101111",
  62913=>"101000000",
  62914=>"000010100",
  62915=>"000111011",
  62916=>"101000110",
  62917=>"011100110",
  62918=>"000010100",
  62919=>"111000001",
  62920=>"000111100",
  62921=>"101101111",
  62922=>"001010001",
  62923=>"101011111",
  62924=>"100110111",
  62925=>"010000010",
  62926=>"010001110",
  62927=>"101100110",
  62928=>"001110110",
  62929=>"000001010",
  62930=>"010111100",
  62931=>"101110101",
  62932=>"010110101",
  62933=>"010001010",
  62934=>"001100101",
  62935=>"101101011",
  62936=>"001101001",
  62937=>"011100111",
  62938=>"100100011",
  62939=>"110101001",
  62940=>"100101010",
  62941=>"111000110",
  62942=>"001101010",
  62943=>"101111011",
  62944=>"101110101",
  62945=>"111101111",
  62946=>"111010010",
  62947=>"010110101",
  62948=>"001111011",
  62949=>"101111000",
  62950=>"110010010",
  62951=>"101001001",
  62952=>"010011000",
  62953=>"111001111",
  62954=>"000011000",
  62955=>"011000001",
  62956=>"010101010",
  62957=>"011100001",
  62958=>"100000010",
  62959=>"101011101",
  62960=>"111111111",
  62961=>"101100011",
  62962=>"000011000",
  62963=>"011000100",
  62964=>"001110101",
  62965=>"011011111",
  62966=>"011001000",
  62967=>"100110010",
  62968=>"101010100",
  62969=>"101101111",
  62970=>"110110101",
  62971=>"110101110",
  62972=>"000000010",
  62973=>"110110111",
  62974=>"110111010",
  62975=>"100011010",
  62976=>"111010000",
  62977=>"101000000",
  62978=>"001100111",
  62979=>"000011100",
  62980=>"010001111",
  62981=>"010001011",
  62982=>"111011110",
  62983=>"000101111",
  62984=>"000110000",
  62985=>"100110111",
  62986=>"001110001",
  62987=>"100100001",
  62988=>"001100010",
  62989=>"010100110",
  62990=>"011111000",
  62991=>"110001001",
  62992=>"001110101",
  62993=>"011011110",
  62994=>"101101101",
  62995=>"100010111",
  62996=>"001001111",
  62997=>"011101100",
  62998=>"001011001",
  62999=>"000011010",
  63000=>"001101000",
  63001=>"011001101",
  63002=>"101001000",
  63003=>"000000011",
  63004=>"100001111",
  63005=>"110011011",
  63006=>"000100110",
  63007=>"011011011",
  63008=>"011000001",
  63009=>"011110100",
  63010=>"000100001",
  63011=>"111000001",
  63012=>"110111011",
  63013=>"011011010",
  63014=>"010011100",
  63015=>"011111101",
  63016=>"110001001",
  63017=>"000011111",
  63018=>"111101110",
  63019=>"010001110",
  63020=>"110011111",
  63021=>"101010111",
  63022=>"000001010",
  63023=>"101110100",
  63024=>"110011110",
  63025=>"101010001",
  63026=>"011101101",
  63027=>"001010011",
  63028=>"000001011",
  63029=>"001011100",
  63030=>"011001100",
  63031=>"000001110",
  63032=>"011001110",
  63033=>"111001101",
  63034=>"000100110",
  63035=>"001011110",
  63036=>"110001101",
  63037=>"000100010",
  63038=>"100111111",
  63039=>"111110111",
  63040=>"110111011",
  63041=>"100001001",
  63042=>"011001100",
  63043=>"100011100",
  63044=>"110011111",
  63045=>"100110011",
  63046=>"101001010",
  63047=>"111001111",
  63048=>"011010101",
  63049=>"101010111",
  63050=>"101011101",
  63051=>"100100011",
  63052=>"101010101",
  63053=>"001101011",
  63054=>"010100111",
  63055=>"110001001",
  63056=>"001011000",
  63057=>"000100000",
  63058=>"010010000",
  63059=>"100011101",
  63060=>"100110010",
  63061=>"011010111",
  63062=>"101001101",
  63063=>"100000011",
  63064=>"100101111",
  63065=>"101001000",
  63066=>"101010101",
  63067=>"101010011",
  63068=>"000101011",
  63069=>"000110001",
  63070=>"101000000",
  63071=>"110100110",
  63072=>"101010010",
  63073=>"000010010",
  63074=>"000100110",
  63075=>"110001000",
  63076=>"011001101",
  63077=>"111000110",
  63078=>"100001000",
  63079=>"101001001",
  63080=>"000110010",
  63081=>"100000010",
  63082=>"000010000",
  63083=>"100100000",
  63084=>"000111110",
  63085=>"001101101",
  63086=>"101100011",
  63087=>"100001000",
  63088=>"010010100",
  63089=>"001000000",
  63090=>"111100000",
  63091=>"100010010",
  63092=>"011100010",
  63093=>"001110110",
  63094=>"110011110",
  63095=>"110000001",
  63096=>"001111011",
  63097=>"001101000",
  63098=>"011011000",
  63099=>"000101001",
  63100=>"110001111",
  63101=>"011011011",
  63102=>"001010111",
  63103=>"000110100",
  63104=>"100010010",
  63105=>"101100001",
  63106=>"111010011",
  63107=>"110010011",
  63108=>"010011101",
  63109=>"010000100",
  63110=>"111110111",
  63111=>"010101011",
  63112=>"110111110",
  63113=>"000000101",
  63114=>"011110110",
  63115=>"011000001",
  63116=>"011010110",
  63117=>"011010000",
  63118=>"100101111",
  63119=>"101100011",
  63120=>"010100000",
  63121=>"011100100",
  63122=>"110000100",
  63123=>"011110100",
  63124=>"110111110",
  63125=>"100011010",
  63126=>"011111001",
  63127=>"001010000",
  63128=>"111111011",
  63129=>"000110000",
  63130=>"011111101",
  63131=>"100110001",
  63132=>"100000101",
  63133=>"110110100",
  63134=>"011011000",
  63135=>"001010111",
  63136=>"111100110",
  63137=>"000010111",
  63138=>"110100101",
  63139=>"101111001",
  63140=>"101101000",
  63141=>"010100100",
  63142=>"011011101",
  63143=>"011001100",
  63144=>"111010000",
  63145=>"111000000",
  63146=>"011000001",
  63147=>"000011111",
  63148=>"001101000",
  63149=>"100000100",
  63150=>"011011010",
  63151=>"110101011",
  63152=>"000001110",
  63153=>"110111001",
  63154=>"001000011",
  63155=>"101010100",
  63156=>"110011110",
  63157=>"100001100",
  63158=>"111000111",
  63159=>"110011010",
  63160=>"111001111",
  63161=>"010001000",
  63162=>"010011010",
  63163=>"100011010",
  63164=>"101101101",
  63165=>"110101001",
  63166=>"100001000",
  63167=>"001101110",
  63168=>"010011001",
  63169=>"001100000",
  63170=>"010101000",
  63171=>"110001000",
  63172=>"001000001",
  63173=>"001001001",
  63174=>"100000010",
  63175=>"011101001",
  63176=>"101000011",
  63177=>"011010000",
  63178=>"100110000",
  63179=>"001100101",
  63180=>"010100100",
  63181=>"000101000",
  63182=>"000101100",
  63183=>"100110110",
  63184=>"000011011",
  63185=>"011000001",
  63186=>"010010111",
  63187=>"111101001",
  63188=>"110100001",
  63189=>"011001010",
  63190=>"010100100",
  63191=>"111111001",
  63192=>"000110110",
  63193=>"010101010",
  63194=>"011110101",
  63195=>"001010111",
  63196=>"011011111",
  63197=>"111111010",
  63198=>"100011010",
  63199=>"011110100",
  63200=>"001011101",
  63201=>"010100011",
  63202=>"111010010",
  63203=>"000111110",
  63204=>"011101100",
  63205=>"000011111",
  63206=>"011000111",
  63207=>"001011000",
  63208=>"000000101",
  63209=>"101101011",
  63210=>"001000001",
  63211=>"100010011",
  63212=>"010000011",
  63213=>"110111011",
  63214=>"001010010",
  63215=>"100100110",
  63216=>"111111100",
  63217=>"000000000",
  63218=>"110100001",
  63219=>"010110100",
  63220=>"000100111",
  63221=>"000011010",
  63222=>"010000111",
  63223=>"010010001",
  63224=>"111011001",
  63225=>"001111011",
  63226=>"001000111",
  63227=>"000010110",
  63228=>"100001100",
  63229=>"000010101",
  63230=>"110110110",
  63231=>"010000001",
  63232=>"000010000",
  63233=>"100101010",
  63234=>"011111100",
  63235=>"101101100",
  63236=>"011110100",
  63237=>"101001101",
  63238=>"011110000",
  63239=>"100111100",
  63240=>"100100101",
  63241=>"101010100",
  63242=>"001011011",
  63243=>"011000000",
  63244=>"101001000",
  63245=>"001101011",
  63246=>"000100100",
  63247=>"111001110",
  63248=>"111100001",
  63249=>"000110001",
  63250=>"001110001",
  63251=>"110000101",
  63252=>"011110000",
  63253=>"001011011",
  63254=>"101001000",
  63255=>"000001100",
  63256=>"011000101",
  63257=>"111101111",
  63258=>"000001100",
  63259=>"001100110",
  63260=>"101000001",
  63261=>"011111001",
  63262=>"100110011",
  63263=>"110011100",
  63264=>"011010111",
  63265=>"111000100",
  63266=>"010011110",
  63267=>"001110001",
  63268=>"010010001",
  63269=>"100010001",
  63270=>"011110101",
  63271=>"000111000",
  63272=>"111100000",
  63273=>"000001010",
  63274=>"111000001",
  63275=>"100001111",
  63276=>"110011000",
  63277=>"000100000",
  63278=>"000011011",
  63279=>"000110010",
  63280=>"000011111",
  63281=>"110000101",
  63282=>"011010111",
  63283=>"111010001",
  63284=>"101110100",
  63285=>"011100100",
  63286=>"110010010",
  63287=>"111011111",
  63288=>"001001001",
  63289=>"111111001",
  63290=>"110010001",
  63291=>"110011000",
  63292=>"010110100",
  63293=>"111001011",
  63294=>"011000110",
  63295=>"001000111",
  63296=>"100001000",
  63297=>"010101110",
  63298=>"100011110",
  63299=>"101100011",
  63300=>"011011010",
  63301=>"001011000",
  63302=>"001001010",
  63303=>"011111101",
  63304=>"111110000",
  63305=>"011101101",
  63306=>"100000000",
  63307=>"011101000",
  63308=>"101011101",
  63309=>"101100011",
  63310=>"111010011",
  63311=>"111010010",
  63312=>"111000010",
  63313=>"011010010",
  63314=>"101010101",
  63315=>"101010101",
  63316=>"100010001",
  63317=>"011101011",
  63318=>"011001000",
  63319=>"110101011",
  63320=>"010000011",
  63321=>"000110010",
  63322=>"010101100",
  63323=>"100101100",
  63324=>"110100011",
  63325=>"011011111",
  63326=>"100010001",
  63327=>"000000000",
  63328=>"010000001",
  63329=>"001000000",
  63330=>"000011101",
  63331=>"111100100",
  63332=>"111101001",
  63333=>"000111001",
  63334=>"101110010",
  63335=>"001100111",
  63336=>"000011111",
  63337=>"110111001",
  63338=>"101011000",
  63339=>"111001110",
  63340=>"101010101",
  63341=>"111000101",
  63342=>"100111010",
  63343=>"011100110",
  63344=>"000010110",
  63345=>"001100110",
  63346=>"100111110",
  63347=>"011000001",
  63348=>"001000010",
  63349=>"100101000",
  63350=>"100100110",
  63351=>"100100011",
  63352=>"101000100",
  63353=>"000111011",
  63354=>"110001000",
  63355=>"111110010",
  63356=>"000000000",
  63357=>"000000011",
  63358=>"110111100",
  63359=>"111110100",
  63360=>"000001110",
  63361=>"110101101",
  63362=>"000010000",
  63363=>"001110010",
  63364=>"101000000",
  63365=>"001101101",
  63366=>"000111010",
  63367=>"011010110",
  63368=>"001101101",
  63369=>"010001110",
  63370=>"100100110",
  63371=>"100100100",
  63372=>"010000111",
  63373=>"011101011",
  63374=>"000101111",
  63375=>"101010001",
  63376=>"111110011",
  63377=>"101001110",
  63378=>"001000000",
  63379=>"111110010",
  63380=>"111101010",
  63381=>"000011011",
  63382=>"111110000",
  63383=>"001001010",
  63384=>"011010111",
  63385=>"010000100",
  63386=>"110110001",
  63387=>"000110000",
  63388=>"111001110",
  63389=>"001001011",
  63390=>"000111000",
  63391=>"001001011",
  63392=>"111111011",
  63393=>"001101100",
  63394=>"100101110",
  63395=>"001110001",
  63396=>"010110011",
  63397=>"011100100",
  63398=>"110111111",
  63399=>"000100001",
  63400=>"100100100",
  63401=>"101010010",
  63402=>"110011110",
  63403=>"100101010",
  63404=>"100100100",
  63405=>"011101110",
  63406=>"001101100",
  63407=>"101110010",
  63408=>"011000010",
  63409=>"100001010",
  63410=>"010000100",
  63411=>"001011101",
  63412=>"010001111",
  63413=>"111111010",
  63414=>"111011100",
  63415=>"001000101",
  63416=>"000011011",
  63417=>"100000101",
  63418=>"000010110",
  63419=>"011101000",
  63420=>"001111011",
  63421=>"010000011",
  63422=>"011010000",
  63423=>"011111000",
  63424=>"010111111",
  63425=>"110101011",
  63426=>"100101111",
  63427=>"110111110",
  63428=>"010001110",
  63429=>"100010010",
  63430=>"110001010",
  63431=>"100011000",
  63432=>"010000011",
  63433=>"101110010",
  63434=>"101100110",
  63435=>"010111110",
  63436=>"110100000",
  63437=>"100110111",
  63438=>"010001010",
  63439=>"000111011",
  63440=>"001111011",
  63441=>"101000011",
  63442=>"100010000",
  63443=>"101100111",
  63444=>"010001000",
  63445=>"100010001",
  63446=>"100001011",
  63447=>"000010011",
  63448=>"000100110",
  63449=>"101101110",
  63450=>"111010111",
  63451=>"000111001",
  63452=>"111010100",
  63453=>"101100011",
  63454=>"101000011",
  63455=>"110010101",
  63456=>"110010101",
  63457=>"110100111",
  63458=>"001101011",
  63459=>"001001000",
  63460=>"001010010",
  63461=>"111010110",
  63462=>"111000000",
  63463=>"101011111",
  63464=>"111010010",
  63465=>"011001111",
  63466=>"010111010",
  63467=>"010110001",
  63468=>"111110100",
  63469=>"001001000",
  63470=>"100000001",
  63471=>"001110011",
  63472=>"010110101",
  63473=>"011100111",
  63474=>"010110010",
  63475=>"110000010",
  63476=>"101000000",
  63477=>"010011011",
  63478=>"100010010",
  63479=>"100001101",
  63480=>"010101101",
  63481=>"000000000",
  63482=>"111101101",
  63483=>"001000010",
  63484=>"010001000",
  63485=>"100010100",
  63486=>"101110010",
  63487=>"000101001",
  63488=>"111111111",
  63489=>"111110111",
  63490=>"100111001",
  63491=>"111100101",
  63492=>"011010111",
  63493=>"101111011",
  63494=>"010000101",
  63495=>"010110000",
  63496=>"000100011",
  63497=>"111111000",
  63498=>"001000010",
  63499=>"001011000",
  63500=>"001001010",
  63501=>"000111111",
  63502=>"111100001",
  63503=>"110101010",
  63504=>"100001110",
  63505=>"000100011",
  63506=>"000001001",
  63507=>"111111111",
  63508=>"101101000",
  63509=>"010000011",
  63510=>"111110011",
  63511=>"010110111",
  63512=>"111111111",
  63513=>"000001111",
  63514=>"000101101",
  63515=>"110111001",
  63516=>"101111001",
  63517=>"011111000",
  63518=>"011011010",
  63519=>"011100001",
  63520=>"000101101",
  63521=>"101101001",
  63522=>"111011010",
  63523=>"110011101",
  63524=>"101011010",
  63525=>"101000110",
  63526=>"110110101",
  63527=>"000111001",
  63528=>"000011011",
  63529=>"100010011",
  63530=>"110100011",
  63531=>"101110101",
  63532=>"000001101",
  63533=>"000100000",
  63534=>"010000011",
  63535=>"011100100",
  63536=>"110100010",
  63537=>"001001100",
  63538=>"010001001",
  63539=>"011101011",
  63540=>"011101110",
  63541=>"111111111",
  63542=>"011001111",
  63543=>"011001000",
  63544=>"100001100",
  63545=>"010010110",
  63546=>"011011001",
  63547=>"001011110",
  63548=>"011101100",
  63549=>"100000111",
  63550=>"101001011",
  63551=>"101000110",
  63552=>"011001110",
  63553=>"010100110",
  63554=>"010010001",
  63555=>"100000000",
  63556=>"110010011",
  63557=>"101011110",
  63558=>"111001100",
  63559=>"000101111",
  63560=>"111000111",
  63561=>"010111001",
  63562=>"110101010",
  63563=>"111101110",
  63564=>"111001110",
  63565=>"001001101",
  63566=>"001000111",
  63567=>"111111101",
  63568=>"011111010",
  63569=>"000000000",
  63570=>"101000111",
  63571=>"000010101",
  63572=>"110101010",
  63573=>"110010010",
  63574=>"011000000",
  63575=>"010010100",
  63576=>"111101100",
  63577=>"100110110",
  63578=>"110000101",
  63579=>"111010011",
  63580=>"101100101",
  63581=>"000000111",
  63582=>"000001111",
  63583=>"010001001",
  63584=>"011011100",
  63585=>"101001000",
  63586=>"001100011",
  63587=>"101111111",
  63588=>"001010010",
  63589=>"111101010",
  63590=>"110110110",
  63591=>"110011000",
  63592=>"000110110",
  63593=>"101101101",
  63594=>"010001111",
  63595=>"111111001",
  63596=>"011010010",
  63597=>"100000001",
  63598=>"100001001",
  63599=>"000101100",
  63600=>"001100001",
  63601=>"100110100",
  63602=>"100000000",
  63603=>"111001010",
  63604=>"000001001",
  63605=>"101110100",
  63606=>"011011011",
  63607=>"100001100",
  63608=>"110000000",
  63609=>"001101010",
  63610=>"110110111",
  63611=>"111101010",
  63612=>"001111000",
  63613=>"011001001",
  63614=>"001100101",
  63615=>"111011111",
  63616=>"110111110",
  63617=>"101010011",
  63618=>"111100000",
  63619=>"000111100",
  63620=>"100011000",
  63621=>"010100111",
  63622=>"001011010",
  63623=>"001101001",
  63624=>"001100111",
  63625=>"111111010",
  63626=>"000011001",
  63627=>"010000011",
  63628=>"001110000",
  63629=>"011011000",
  63630=>"001101101",
  63631=>"011100011",
  63632=>"000000010",
  63633=>"101101101",
  63634=>"110000010",
  63635=>"010000101",
  63636=>"010001101",
  63637=>"000011110",
  63638=>"101101101",
  63639=>"000100001",
  63640=>"101111101",
  63641=>"111111101",
  63642=>"000010100",
  63643=>"101001000",
  63644=>"011110101",
  63645=>"010101011",
  63646=>"000111000",
  63647=>"000110001",
  63648=>"110100010",
  63649=>"001101110",
  63650=>"001110101",
  63651=>"010100000",
  63652=>"000000001",
  63653=>"111111000",
  63654=>"010101010",
  63655=>"110101111",
  63656=>"101001110",
  63657=>"010100000",
  63658=>"010010000",
  63659=>"000000010",
  63660=>"010000101",
  63661=>"101010000",
  63662=>"000011101",
  63663=>"101010110",
  63664=>"010001001",
  63665=>"010000010",
  63666=>"110111000",
  63667=>"010011000",
  63668=>"011111100",
  63669=>"001000000",
  63670=>"000011001",
  63671=>"000010001",
  63672=>"100101111",
  63673=>"001001111",
  63674=>"011000101",
  63675=>"000000001",
  63676=>"100000100",
  63677=>"110100100",
  63678=>"110101100",
  63679=>"000101001",
  63680=>"000000010",
  63681=>"000000000",
  63682=>"111001111",
  63683=>"110101001",
  63684=>"011100010",
  63685=>"000100010",
  63686=>"010001110",
  63687=>"000000110",
  63688=>"110001101",
  63689=>"010000011",
  63690=>"111111011",
  63691=>"111010011",
  63692=>"011111101",
  63693=>"001110001",
  63694=>"011000111",
  63695=>"011111100",
  63696=>"101110001",
  63697=>"010001101",
  63698=>"000000000",
  63699=>"111001111",
  63700=>"100100100",
  63701=>"001001111",
  63702=>"001001110",
  63703=>"110000001",
  63704=>"011000111",
  63705=>"000010010",
  63706=>"101000001",
  63707=>"001101100",
  63708=>"101010100",
  63709=>"001001001",
  63710=>"101011000",
  63711=>"010011000",
  63712=>"111101111",
  63713=>"010000001",
  63714=>"110100001",
  63715=>"010100000",
  63716=>"000011010",
  63717=>"111101101",
  63718=>"110101110",
  63719=>"000111111",
  63720=>"000110001",
  63721=>"010111000",
  63722=>"101010101",
  63723=>"000000100",
  63724=>"010010011",
  63725=>"010011010",
  63726=>"101001110",
  63727=>"010100000",
  63728=>"111000101",
  63729=>"010100110",
  63730=>"000001111",
  63731=>"100111101",
  63732=>"110111100",
  63733=>"011110000",
  63734=>"010010010",
  63735=>"001011001",
  63736=>"010001001",
  63737=>"011101011",
  63738=>"100101000",
  63739=>"110010000",
  63740=>"010000101",
  63741=>"100110111",
  63742=>"010001101",
  63743=>"110101000",
  63744=>"000110000",
  63745=>"101011000",
  63746=>"011001011",
  63747=>"010000001",
  63748=>"100001000",
  63749=>"110000000",
  63750=>"010010000",
  63751=>"010001001",
  63752=>"110110010",
  63753=>"001100100",
  63754=>"100110011",
  63755=>"100101100",
  63756=>"111110100",
  63757=>"110101100",
  63758=>"110010100",
  63759=>"011110110",
  63760=>"010100001",
  63761=>"110011000",
  63762=>"011101011",
  63763=>"011110101",
  63764=>"000001001",
  63765=>"001111001",
  63766=>"111110001",
  63767=>"101100110",
  63768=>"101000001",
  63769=>"010001111",
  63770=>"001111111",
  63771=>"000000011",
  63772=>"000101001",
  63773=>"101100010",
  63774=>"011101100",
  63775=>"000111010",
  63776=>"010000000",
  63777=>"111100001",
  63778=>"111000100",
  63779=>"000010101",
  63780=>"011111100",
  63781=>"100000000",
  63782=>"100000000",
  63783=>"110000001",
  63784=>"010011110",
  63785=>"101001101",
  63786=>"110110011",
  63787=>"101101110",
  63788=>"001000000",
  63789=>"111001111",
  63790=>"101001000",
  63791=>"111100110",
  63792=>"110111000",
  63793=>"111011000",
  63794=>"111000101",
  63795=>"010010100",
  63796=>"110100111",
  63797=>"001010111",
  63798=>"111111100",
  63799=>"001010011",
  63800=>"101010011",
  63801=>"100101011",
  63802=>"111010111",
  63803=>"000010000",
  63804=>"110001110",
  63805=>"111010011",
  63806=>"011000100",
  63807=>"010111111",
  63808=>"111100110",
  63809=>"000010100",
  63810=>"111110001",
  63811=>"101100101",
  63812=>"001000101",
  63813=>"100001001",
  63814=>"111001101",
  63815=>"001011000",
  63816=>"001001001",
  63817=>"011100101",
  63818=>"001110110",
  63819=>"000001111",
  63820=>"101000010",
  63821=>"111011100",
  63822=>"000110101",
  63823=>"001111011",
  63824=>"001111110",
  63825=>"011101100",
  63826=>"000000001",
  63827=>"111001011",
  63828=>"100110000",
  63829=>"101101011",
  63830=>"001011001",
  63831=>"000111001",
  63832=>"010110000",
  63833=>"101110001",
  63834=>"000000110",
  63835=>"110000000",
  63836=>"011101001",
  63837=>"000011000",
  63838=>"101111001",
  63839=>"000111000",
  63840=>"010110100",
  63841=>"100110100",
  63842=>"100111100",
  63843=>"101000110",
  63844=>"101101011",
  63845=>"111000000",
  63846=>"001100001",
  63847=>"110000101",
  63848=>"010100110",
  63849=>"111011101",
  63850=>"010101100",
  63851=>"101010110",
  63852=>"101110000",
  63853=>"000001111",
  63854=>"011110111",
  63855=>"000011001",
  63856=>"110100100",
  63857=>"011110011",
  63858=>"111111101",
  63859=>"100000110",
  63860=>"001101010",
  63861=>"100110001",
  63862=>"000111111",
  63863=>"001000010",
  63864=>"100100000",
  63865=>"011011011",
  63866=>"111111011",
  63867=>"000111111",
  63868=>"111110010",
  63869=>"010011100",
  63870=>"000110010",
  63871=>"000111111",
  63872=>"000010111",
  63873=>"100000000",
  63874=>"010111110",
  63875=>"110110000",
  63876=>"011010011",
  63877=>"010100111",
  63878=>"001110010",
  63879=>"100111111",
  63880=>"101100000",
  63881=>"001000100",
  63882=>"101111100",
  63883=>"110011111",
  63884=>"011010001",
  63885=>"011010001",
  63886=>"000100110",
  63887=>"011111010",
  63888=>"010000111",
  63889=>"110111000",
  63890=>"101000001",
  63891=>"101000111",
  63892=>"110011101",
  63893=>"110101110",
  63894=>"011101111",
  63895=>"010001110",
  63896=>"101100111",
  63897=>"110101110",
  63898=>"001101111",
  63899=>"000101111",
  63900=>"011100101",
  63901=>"001111000",
  63902=>"001110111",
  63903=>"101011111",
  63904=>"101110001",
  63905=>"001000011",
  63906=>"111010001",
  63907=>"101000111",
  63908=>"100001110",
  63909=>"100011011",
  63910=>"001100000",
  63911=>"001001010",
  63912=>"110000011",
  63913=>"100100100",
  63914=>"111101000",
  63915=>"111100101",
  63916=>"111101010",
  63917=>"000111011",
  63918=>"000011100",
  63919=>"101000001",
  63920=>"111110100",
  63921=>"111000111",
  63922=>"000111101",
  63923=>"001010111",
  63924=>"010001011",
  63925=>"100011110",
  63926=>"011011111",
  63927=>"111110101",
  63928=>"100111100",
  63929=>"110001111",
  63930=>"100101011",
  63931=>"111010101",
  63932=>"010010000",
  63933=>"001011001",
  63934=>"011111110",
  63935=>"100100111",
  63936=>"100000110",
  63937=>"111101010",
  63938=>"101110101",
  63939=>"110011001",
  63940=>"000110100",
  63941=>"000001001",
  63942=>"011111100",
  63943=>"100001111",
  63944=>"111010101",
  63945=>"101001101",
  63946=>"101010111",
  63947=>"100101110",
  63948=>"000001000",
  63949=>"101110011",
  63950=>"001110101",
  63951=>"000111010",
  63952=>"010110101",
  63953=>"101111101",
  63954=>"011100000",
  63955=>"101111000",
  63956=>"010011010",
  63957=>"000101000",
  63958=>"000011111",
  63959=>"001010110",
  63960=>"001011101",
  63961=>"011100101",
  63962=>"110101111",
  63963=>"110011001",
  63964=>"011101101",
  63965=>"010101010",
  63966=>"100101101",
  63967=>"100011000",
  63968=>"010100111",
  63969=>"100000111",
  63970=>"111101111",
  63971=>"100110010",
  63972=>"100100110",
  63973=>"000101110",
  63974=>"100110011",
  63975=>"000011100",
  63976=>"010111111",
  63977=>"000101001",
  63978=>"000100100",
  63979=>"111010101",
  63980=>"001111010",
  63981=>"110001111",
  63982=>"110101111",
  63983=>"100111011",
  63984=>"000000110",
  63985=>"010001000",
  63986=>"110111101",
  63987=>"011111000",
  63988=>"011000001",
  63989=>"000000110",
  63990=>"111100000",
  63991=>"101001111",
  63992=>"111101100",
  63993=>"010111001",
  63994=>"100000100",
  63995=>"001101000",
  63996=>"100100111",
  63997=>"101110010",
  63998=>"000000100",
  63999=>"110000111",
  64000=>"110101010",
  64001=>"000111010",
  64002=>"111110101",
  64003=>"111101011",
  64004=>"110101110",
  64005=>"010100010",
  64006=>"000111011",
  64007=>"000010111",
  64008=>"010110001",
  64009=>"010101100",
  64010=>"001010111",
  64011=>"111111101",
  64012=>"100010110",
  64013=>"010101100",
  64014=>"111010101",
  64015=>"110101111",
  64016=>"101001010",
  64017=>"000010010",
  64018=>"111000110",
  64019=>"001100111",
  64020=>"111001010",
  64021=>"100011001",
  64022=>"011001010",
  64023=>"111010110",
  64024=>"000100000",
  64025=>"010111001",
  64026=>"011101100",
  64027=>"000010000",
  64028=>"111111111",
  64029=>"111101101",
  64030=>"000111110",
  64031=>"001011010",
  64032=>"101001011",
  64033=>"100110101",
  64034=>"001101111",
  64035=>"110010100",
  64036=>"100100110",
  64037=>"000000111",
  64038=>"010011111",
  64039=>"111110100",
  64040=>"010011101",
  64041=>"000100100",
  64042=>"110001000",
  64043=>"000110011",
  64044=>"110110111",
  64045=>"111100111",
  64046=>"110100011",
  64047=>"011000010",
  64048=>"111100011",
  64049=>"111011011",
  64050=>"011110011",
  64051=>"101001001",
  64052=>"111100111",
  64053=>"001010100",
  64054=>"111011110",
  64055=>"001000111",
  64056=>"100110100",
  64057=>"101100111",
  64058=>"111001010",
  64059=>"001000001",
  64060=>"100110001",
  64061=>"000000100",
  64062=>"001010010",
  64063=>"000011000",
  64064=>"011001101",
  64065=>"100011101",
  64066=>"101001001",
  64067=>"000011011",
  64068=>"010101101",
  64069=>"101001101",
  64070=>"010111000",
  64071=>"010011011",
  64072=>"110000011",
  64073=>"101101100",
  64074=>"111110011",
  64075=>"101110100",
  64076=>"011101010",
  64077=>"010000001",
  64078=>"000011000",
  64079=>"001000110",
  64080=>"001110001",
  64081=>"001100001",
  64082=>"110011011",
  64083=>"001000011",
  64084=>"111110111",
  64085=>"101101010",
  64086=>"110101111",
  64087=>"110110110",
  64088=>"001000100",
  64089=>"100000010",
  64090=>"111101111",
  64091=>"101100101",
  64092=>"001000100",
  64093=>"111000011",
  64094=>"100110110",
  64095=>"000111101",
  64096=>"000111001",
  64097=>"101000100",
  64098=>"111010101",
  64099=>"011010011",
  64100=>"100110111",
  64101=>"001000101",
  64102=>"110100100",
  64103=>"001101100",
  64104=>"110010001",
  64105=>"001000011",
  64106=>"100011011",
  64107=>"100001011",
  64108=>"111011011",
  64109=>"101111101",
  64110=>"100100010",
  64111=>"011100011",
  64112=>"011010100",
  64113=>"101111100",
  64114=>"111010001",
  64115=>"000000011",
  64116=>"010000111",
  64117=>"101100110",
  64118=>"011101101",
  64119=>"100111000",
  64120=>"011000100",
  64121=>"010110010",
  64122=>"101100001",
  64123=>"101111110",
  64124=>"110000011",
  64125=>"001011000",
  64126=>"010100101",
  64127=>"010000100",
  64128=>"111111001",
  64129=>"000011000",
  64130=>"111100001",
  64131=>"011000011",
  64132=>"000101100",
  64133=>"101010110",
  64134=>"111000101",
  64135=>"000000001",
  64136=>"110100010",
  64137=>"101001111",
  64138=>"101100000",
  64139=>"011011010",
  64140=>"000111010",
  64141=>"111001010",
  64142=>"001111110",
  64143=>"001011001",
  64144=>"010111111",
  64145=>"111000111",
  64146=>"011010000",
  64147=>"011100000",
  64148=>"100100100",
  64149=>"110111101",
  64150=>"110110110",
  64151=>"011001001",
  64152=>"101001011",
  64153=>"000100000",
  64154=>"010100111",
  64155=>"001001001",
  64156=>"001101101",
  64157=>"101111001",
  64158=>"010101111",
  64159=>"101100011",
  64160=>"101110011",
  64161=>"000100011",
  64162=>"010100100",
  64163=>"010111000",
  64164=>"100110000",
  64165=>"000110001",
  64166=>"001100111",
  64167=>"000000011",
  64168=>"010000011",
  64169=>"111101111",
  64170=>"001000000",
  64171=>"001001101",
  64172=>"111111111",
  64173=>"000001001",
  64174=>"011101000",
  64175=>"001101110",
  64176=>"101100100",
  64177=>"101110000",
  64178=>"111110010",
  64179=>"100101111",
  64180=>"111000010",
  64181=>"000111001",
  64182=>"111101111",
  64183=>"011111110",
  64184=>"000000011",
  64185=>"000001110",
  64186=>"011010010",
  64187=>"101101100",
  64188=>"100000101",
  64189=>"111100001",
  64190=>"100101110",
  64191=>"011101110",
  64192=>"100000010",
  64193=>"111000100",
  64194=>"100000001",
  64195=>"010011100",
  64196=>"000001000",
  64197=>"001101100",
  64198=>"110110011",
  64199=>"100001001",
  64200=>"000111001",
  64201=>"000111100",
  64202=>"001101001",
  64203=>"110111010",
  64204=>"111000111",
  64205=>"011011010",
  64206=>"110010110",
  64207=>"110000110",
  64208=>"110111110",
  64209=>"101110001",
  64210=>"011010110",
  64211=>"010011110",
  64212=>"001000111",
  64213=>"000001111",
  64214=>"100110110",
  64215=>"001101011",
  64216=>"111011010",
  64217=>"011100000",
  64218=>"000011100",
  64219=>"111101110",
  64220=>"010011010",
  64221=>"000110001",
  64222=>"111011001",
  64223=>"010000110",
  64224=>"001010000",
  64225=>"110000001",
  64226=>"110100110",
  64227=>"010001111",
  64228=>"011010001",
  64229=>"010000001",
  64230=>"100100100",
  64231=>"101001001",
  64232=>"111000101",
  64233=>"111001100",
  64234=>"100001001",
  64235=>"100000010",
  64236=>"000001110",
  64237=>"101100001",
  64238=>"101100111",
  64239=>"011100101",
  64240=>"101011111",
  64241=>"000110111",
  64242=>"110010000",
  64243=>"010000000",
  64244=>"010011001",
  64245=>"111011010",
  64246=>"011100000",
  64247=>"110100100",
  64248=>"000010001",
  64249=>"111011110",
  64250=>"011111001",
  64251=>"101110101",
  64252=>"001000110",
  64253=>"111011111",
  64254=>"010101110",
  64255=>"110111111",
  64256=>"111010011",
  64257=>"011110010",
  64258=>"100111101",
  64259=>"111010010",
  64260=>"001000110",
  64261=>"101010010",
  64262=>"100000111",
  64263=>"011100000",
  64264=>"110010011",
  64265=>"010000010",
  64266=>"111110101",
  64267=>"111101100",
  64268=>"011010111",
  64269=>"000100101",
  64270=>"110101000",
  64271=>"001000000",
  64272=>"110101001",
  64273=>"111011001",
  64274=>"110000100",
  64275=>"011010001",
  64276=>"010001000",
  64277=>"111110110",
  64278=>"101011111",
  64279=>"000010010",
  64280=>"111001101",
  64281=>"011110111",
  64282=>"010000001",
  64283=>"000100001",
  64284=>"101111100",
  64285=>"000010110",
  64286=>"100011101",
  64287=>"100011010",
  64288=>"111011110",
  64289=>"111010111",
  64290=>"000100000",
  64291=>"110011110",
  64292=>"010001011",
  64293=>"010010010",
  64294=>"101110100",
  64295=>"011101110",
  64296=>"000110100",
  64297=>"110111011",
  64298=>"101000011",
  64299=>"101110000",
  64300=>"100010111",
  64301=>"000100000",
  64302=>"000110101",
  64303=>"111011000",
  64304=>"111001111",
  64305=>"100100100",
  64306=>"011011010",
  64307=>"111100010",
  64308=>"000001001",
  64309=>"100001111",
  64310=>"101010011",
  64311=>"000000011",
  64312=>"111111110",
  64313=>"110110010",
  64314=>"001111010",
  64315=>"111001101",
  64316=>"010101110",
  64317=>"000000110",
  64318=>"110001000",
  64319=>"000110011",
  64320=>"101001110",
  64321=>"001101011",
  64322=>"000000000",
  64323=>"001100111",
  64324=>"100011000",
  64325=>"111110000",
  64326=>"100110011",
  64327=>"000101000",
  64328=>"111110100",
  64329=>"110001100",
  64330=>"110010110",
  64331=>"011110000",
  64332=>"101000010",
  64333=>"010000111",
  64334=>"011101111",
  64335=>"001010001",
  64336=>"001100011",
  64337=>"011001011",
  64338=>"011101011",
  64339=>"111100010",
  64340=>"100010000",
  64341=>"110011000",
  64342=>"011110001",
  64343=>"111101011",
  64344=>"010001100",
  64345=>"101101001",
  64346=>"110110011",
  64347=>"001100111",
  64348=>"000000110",
  64349=>"101000111",
  64350=>"101101100",
  64351=>"000000010",
  64352=>"110011111",
  64353=>"101101110",
  64354=>"110100001",
  64355=>"111110100",
  64356=>"000001100",
  64357=>"111011010",
  64358=>"111001010",
  64359=>"101101111",
  64360=>"001101000",
  64361=>"011101001",
  64362=>"110100111",
  64363=>"010001010",
  64364=>"101000010",
  64365=>"111111101",
  64366=>"111000000",
  64367=>"000000111",
  64368=>"110010011",
  64369=>"100000000",
  64370=>"001101110",
  64371=>"101001000",
  64372=>"110001110",
  64373=>"011001010",
  64374=>"011011000",
  64375=>"100011000",
  64376=>"001001111",
  64377=>"111110011",
  64378=>"100100100",
  64379=>"110011111",
  64380=>"110001011",
  64381=>"111011001",
  64382=>"000001100",
  64383=>"000111001",
  64384=>"100001101",
  64385=>"111100110",
  64386=>"000111110",
  64387=>"010111011",
  64388=>"011110101",
  64389=>"111000011",
  64390=>"000110000",
  64391=>"111001110",
  64392=>"010111001",
  64393=>"111000100",
  64394=>"000110100",
  64395=>"010011000",
  64396=>"010000111",
  64397=>"100110100",
  64398=>"100001011",
  64399=>"101011111",
  64400=>"110101110",
  64401=>"011011010",
  64402=>"001001100",
  64403=>"011110001",
  64404=>"001100111",
  64405=>"001001001",
  64406=>"001101000",
  64407=>"101011100",
  64408=>"011001110",
  64409=>"101101110",
  64410=>"001100011",
  64411=>"010011010",
  64412=>"011010101",
  64413=>"100001100",
  64414=>"110110001",
  64415=>"100010111",
  64416=>"111011110",
  64417=>"111100000",
  64418=>"100001100",
  64419=>"100000011",
  64420=>"001100101",
  64421=>"101110010",
  64422=>"010000101",
  64423=>"110111110",
  64424=>"010111111",
  64425=>"010111111",
  64426=>"101010110",
  64427=>"111110110",
  64428=>"101111011",
  64429=>"111101011",
  64430=>"111100001",
  64431=>"100110101",
  64432=>"001101001",
  64433=>"001010111",
  64434=>"111100111",
  64435=>"000000101",
  64436=>"011000100",
  64437=>"101000010",
  64438=>"000001000",
  64439=>"100100100",
  64440=>"011011011",
  64441=>"101111010",
  64442=>"111011100",
  64443=>"001011111",
  64444=>"100101000",
  64445=>"000000110",
  64446=>"110100011",
  64447=>"111101001",
  64448=>"111110011",
  64449=>"011101111",
  64450=>"000000001",
  64451=>"000101011",
  64452=>"000000100",
  64453=>"101010110",
  64454=>"100000110",
  64455=>"100010111",
  64456=>"101010101",
  64457=>"011101100",
  64458=>"110010001",
  64459=>"101000000",
  64460=>"000011100",
  64461=>"110110101",
  64462=>"010000111",
  64463=>"000010010",
  64464=>"000000010",
  64465=>"000011111",
  64466=>"010011010",
  64467=>"100100000",
  64468=>"000011101",
  64469=>"111000100",
  64470=>"110111010",
  64471=>"111000011",
  64472=>"011011100",
  64473=>"011010010",
  64474=>"011001101",
  64475=>"111100100",
  64476=>"101000101",
  64477=>"011010011",
  64478=>"111100100",
  64479=>"001010111",
  64480=>"011010111",
  64481=>"000010111",
  64482=>"001101001",
  64483=>"101000010",
  64484=>"110110100",
  64485=>"111010011",
  64486=>"001101110",
  64487=>"000001001",
  64488=>"111100100",
  64489=>"110110010",
  64490=>"001100100",
  64491=>"111000100",
  64492=>"011100100",
  64493=>"011111111",
  64494=>"100000111",
  64495=>"000010001",
  64496=>"000010100",
  64497=>"010000010",
  64498=>"001010000",
  64499=>"111110111",
  64500=>"010001110",
  64501=>"110101111",
  64502=>"110111110",
  64503=>"110101101",
  64504=>"101010000",
  64505=>"111010011",
  64506=>"001101111",
  64507=>"110110011",
  64508=>"010100011",
  64509=>"100111001",
  64510=>"001111000",
  64511=>"101110101",
  64512=>"110011100",
  64513=>"111111010",
  64514=>"011001111",
  64515=>"000010101",
  64516=>"000111011",
  64517=>"000100010",
  64518=>"011110010",
  64519=>"000011001",
  64520=>"010000001",
  64521=>"110010010",
  64522=>"000010100",
  64523=>"111001001",
  64524=>"101100001",
  64525=>"000001011",
  64526=>"101011111",
  64527=>"100110011",
  64528=>"001010011",
  64529=>"000011001",
  64530=>"101111111",
  64531=>"010001010",
  64532=>"100010111",
  64533=>"111001110",
  64534=>"010001000",
  64535=>"101010001",
  64536=>"100001110",
  64537=>"100001001",
  64538=>"010100100",
  64539=>"100001100",
  64540=>"111111111",
  64541=>"101010001",
  64542=>"111000000",
  64543=>"001010011",
  64544=>"101011000",
  64545=>"010000110",
  64546=>"101110111",
  64547=>"101011101",
  64548=>"100011110",
  64549=>"111001010",
  64550=>"000010100",
  64551=>"100011001",
  64552=>"010110000",
  64553=>"100011111",
  64554=>"111101000",
  64555=>"011100110",
  64556=>"100001100",
  64557=>"000101000",
  64558=>"011110010",
  64559=>"110100011",
  64560=>"111010000",
  64561=>"010011000",
  64562=>"011101000",
  64563=>"111110000",
  64564=>"011001111",
  64565=>"110001100",
  64566=>"011010010",
  64567=>"100101100",
  64568=>"001111111",
  64569=>"110000111",
  64570=>"000111110",
  64571=>"100100000",
  64572=>"110110000",
  64573=>"011101011",
  64574=>"110000011",
  64575=>"110010010",
  64576=>"010010010",
  64577=>"010111011",
  64578=>"100110000",
  64579=>"101011001",
  64580=>"100010011",
  64581=>"001110010",
  64582=>"110100001",
  64583=>"111000011",
  64584=>"100001011",
  64585=>"001010110",
  64586=>"110100101",
  64587=>"010100011",
  64588=>"000001110",
  64589=>"001001100",
  64590=>"010011010",
  64591=>"111001100",
  64592=>"001100111",
  64593=>"101110010",
  64594=>"001001110",
  64595=>"001111110",
  64596=>"001110011",
  64597=>"110111110",
  64598=>"111001111",
  64599=>"100001001",
  64600=>"001100000",
  64601=>"100001001",
  64602=>"111110011",
  64603=>"010011001",
  64604=>"110000000",
  64605=>"100100101",
  64606=>"100111011",
  64607=>"100101101",
  64608=>"010001100",
  64609=>"110110111",
  64610=>"100001011",
  64611=>"011010001",
  64612=>"111100000",
  64613=>"011011100",
  64614=>"000111101",
  64615=>"001101001",
  64616=>"100110001",
  64617=>"010101101",
  64618=>"101101010",
  64619=>"100100100",
  64620=>"100110010",
  64621=>"011001111",
  64622=>"101101011",
  64623=>"011010101",
  64624=>"110001000",
  64625=>"011000100",
  64626=>"100111100",
  64627=>"001110100",
  64628=>"011010001",
  64629=>"110110000",
  64630=>"100001110",
  64631=>"001111011",
  64632=>"100010110",
  64633=>"100001111",
  64634=>"011110100",
  64635=>"000010100",
  64636=>"010010101",
  64637=>"010011000",
  64638=>"001100111",
  64639=>"100110011",
  64640=>"010001111",
  64641=>"110010001",
  64642=>"001010001",
  64643=>"101101111",
  64644=>"000101000",
  64645=>"011101000",
  64646=>"010001101",
  64647=>"011000111",
  64648=>"000100000",
  64649=>"010111010",
  64650=>"110100000",
  64651=>"010100000",
  64652=>"000000001",
  64653=>"101110011",
  64654=>"011001000",
  64655=>"000111010",
  64656=>"100111001",
  64657=>"000111000",
  64658=>"010101100",
  64659=>"000010101",
  64660=>"000110100",
  64661=>"111000011",
  64662=>"001000000",
  64663=>"010001001",
  64664=>"101011010",
  64665=>"001000110",
  64666=>"100110111",
  64667=>"001101101",
  64668=>"101111110",
  64669=>"001001100",
  64670=>"110000000",
  64671=>"101010010",
  64672=>"010011000",
  64673=>"011111001",
  64674=>"101101111",
  64675=>"001000111",
  64676=>"110101111",
  64677=>"100111001",
  64678=>"000000011",
  64679=>"100110110",
  64680=>"110010100",
  64681=>"010001000",
  64682=>"010100000",
  64683=>"011001111",
  64684=>"000011011",
  64685=>"000001111",
  64686=>"011100111",
  64687=>"001010001",
  64688=>"111111001",
  64689=>"011001111",
  64690=>"000011011",
  64691=>"010011001",
  64692=>"001101111",
  64693=>"011101011",
  64694=>"010110011",
  64695=>"000111110",
  64696=>"100100000",
  64697=>"010111011",
  64698=>"011100011",
  64699=>"110100000",
  64700=>"001110101",
  64701=>"111000111",
  64702=>"011110111",
  64703=>"011100111",
  64704=>"010000110",
  64705=>"000110001",
  64706=>"111110111",
  64707=>"100001000",
  64708=>"000101010",
  64709=>"011000111",
  64710=>"010000111",
  64711=>"110101011",
  64712=>"011001001",
  64713=>"011000011",
  64714=>"100000110",
  64715=>"100001010",
  64716=>"110100100",
  64717=>"100001111",
  64718=>"111101110",
  64719=>"101111011",
  64720=>"100010000",
  64721=>"111100011",
  64722=>"010010010",
  64723=>"111101111",
  64724=>"011100010",
  64725=>"000100011",
  64726=>"110100100",
  64727=>"011011000",
  64728=>"011100001",
  64729=>"000001010",
  64730=>"010101111",
  64731=>"010000010",
  64732=>"001010010",
  64733=>"001001101",
  64734=>"110000110",
  64735=>"011101010",
  64736=>"001011000",
  64737=>"101111101",
  64738=>"101000111",
  64739=>"010001000",
  64740=>"011101001",
  64741=>"110100111",
  64742=>"000010000",
  64743=>"011111100",
  64744=>"100000011",
  64745=>"110010101",
  64746=>"101100001",
  64747=>"000011000",
  64748=>"111101011",
  64749=>"101001110",
  64750=>"101101011",
  64751=>"011010001",
  64752=>"101110000",
  64753=>"010110001",
  64754=>"000111001",
  64755=>"110110001",
  64756=>"111011000",
  64757=>"101011000",
  64758=>"101111000",
  64759=>"000010011",
  64760=>"110111000",
  64761=>"110110110",
  64762=>"000110111",
  64763=>"110000010",
  64764=>"010011001",
  64765=>"111001110",
  64766=>"000011100",
  64767=>"111010110",
  64768=>"000000000",
  64769=>"010110100",
  64770=>"100001010",
  64771=>"100110011",
  64772=>"000101111",
  64773=>"000000001",
  64774=>"111011101",
  64775=>"001011011",
  64776=>"010010000",
  64777=>"111111000",
  64778=>"000001000",
  64779=>"001000100",
  64780=>"100011011",
  64781=>"111000110",
  64782=>"011100111",
  64783=>"111011101",
  64784=>"000000000",
  64785=>"011111010",
  64786=>"000100000",
  64787=>"110000110",
  64788=>"111100110",
  64789=>"101101001",
  64790=>"100100111",
  64791=>"000010111",
  64792=>"011000101",
  64793=>"101000110",
  64794=>"001000010",
  64795=>"001011011",
  64796=>"110001011",
  64797=>"000000010",
  64798=>"000111111",
  64799=>"000100111",
  64800=>"000000001",
  64801=>"111001011",
  64802=>"001101100",
  64803=>"000011000",
  64804=>"111100100",
  64805=>"011110000",
  64806=>"000111100",
  64807=>"011000101",
  64808=>"111001001",
  64809=>"011100011",
  64810=>"000101010",
  64811=>"000000011",
  64812=>"111001011",
  64813=>"110000010",
  64814=>"000010111",
  64815=>"011111111",
  64816=>"000110000",
  64817=>"110010011",
  64818=>"111111110",
  64819=>"000100011",
  64820=>"001100011",
  64821=>"111010010",
  64822=>"110000011",
  64823=>"011000000",
  64824=>"001111110",
  64825=>"001111111",
  64826=>"010100011",
  64827=>"100111100",
  64828=>"110110101",
  64829=>"101100010",
  64830=>"101110100",
  64831=>"001010000",
  64832=>"001011100",
  64833=>"100110101",
  64834=>"000001110",
  64835=>"011001001",
  64836=>"011010000",
  64837=>"000001110",
  64838=>"001100010",
  64839=>"010111110",
  64840=>"000001110",
  64841=>"001010000",
  64842=>"010101011",
  64843=>"111011110",
  64844=>"110101111",
  64845=>"111001011",
  64846=>"011010010",
  64847=>"110001100",
  64848=>"011010011",
  64849=>"100010010",
  64850=>"110011001",
  64851=>"111001100",
  64852=>"110100111",
  64853=>"110100010",
  64854=>"110110100",
  64855=>"001101100",
  64856=>"101100001",
  64857=>"000011111",
  64858=>"101101111",
  64859=>"101000010",
  64860=>"101011011",
  64861=>"110000000",
  64862=>"010001010",
  64863=>"001100011",
  64864=>"111111100",
  64865=>"100011000",
  64866=>"111110111",
  64867=>"111010101",
  64868=>"110010110",
  64869=>"011010010",
  64870=>"001111011",
  64871=>"010010011",
  64872=>"100100011",
  64873=>"010100011",
  64874=>"001101110",
  64875=>"100001101",
  64876=>"111100001",
  64877=>"110011001",
  64878=>"100000100",
  64879=>"000010111",
  64880=>"001110001",
  64881=>"100010101",
  64882=>"110010100",
  64883=>"011101011",
  64884=>"110001010",
  64885=>"101001111",
  64886=>"101001101",
  64887=>"110001110",
  64888=>"101000110",
  64889=>"001101000",
  64890=>"100011100",
  64891=>"011001100",
  64892=>"100011100",
  64893=>"011111111",
  64894=>"101001100",
  64895=>"101100101",
  64896=>"110001100",
  64897=>"100110011",
  64898=>"010111001",
  64899=>"000100001",
  64900=>"101001010",
  64901=>"100000000",
  64902=>"001011011",
  64903=>"110001111",
  64904=>"010001000",
  64905=>"111000111",
  64906=>"111100111",
  64907=>"000010001",
  64908=>"101011011",
  64909=>"110100011",
  64910=>"010001011",
  64911=>"101000100",
  64912=>"001010001",
  64913=>"000101011",
  64914=>"100101110",
  64915=>"100011101",
  64916=>"100001111",
  64917=>"000011111",
  64918=>"011110111",
  64919=>"010000000",
  64920=>"110000100",
  64921=>"111101011",
  64922=>"010110011",
  64923=>"000100100",
  64924=>"001111001",
  64925=>"000100101",
  64926=>"101001101",
  64927=>"110100011",
  64928=>"001100000",
  64929=>"111001110",
  64930=>"000000000",
  64931=>"110010011",
  64932=>"010101010",
  64933=>"010101110",
  64934=>"010010100",
  64935=>"001011001",
  64936=>"111010110",
  64937=>"010110111",
  64938=>"000000111",
  64939=>"010010110",
  64940=>"011010100",
  64941=>"100101100",
  64942=>"000011100",
  64943=>"001001011",
  64944=>"001001100",
  64945=>"110101111",
  64946=>"011100000",
  64947=>"000110001",
  64948=>"101111001",
  64949=>"110110011",
  64950=>"011000101",
  64951=>"111111100",
  64952=>"001000110",
  64953=>"110110001",
  64954=>"100001110",
  64955=>"111010000",
  64956=>"110111011",
  64957=>"010110110",
  64958=>"100100000",
  64959=>"100011001",
  64960=>"010110011",
  64961=>"110011001",
  64962=>"110100010",
  64963=>"010101001",
  64964=>"000101101",
  64965=>"111000001",
  64966=>"110110010",
  64967=>"011111101",
  64968=>"100011001",
  64969=>"110001100",
  64970=>"100001100",
  64971=>"011010010",
  64972=>"110101110",
  64973=>"000100101",
  64974=>"000001110",
  64975=>"010010000",
  64976=>"000110111",
  64977=>"001110011",
  64978=>"010010110",
  64979=>"101011011",
  64980=>"110011010",
  64981=>"010111001",
  64982=>"011011110",
  64983=>"010000001",
  64984=>"111110100",
  64985=>"111001000",
  64986=>"100000001",
  64987=>"110001001",
  64988=>"100001110",
  64989=>"110011000",
  64990=>"011101010",
  64991=>"010111011",
  64992=>"001000100",
  64993=>"000111100",
  64994=>"011011100",
  64995=>"001010110",
  64996=>"001111110",
  64997=>"101010111",
  64998=>"100011111",
  64999=>"010011001",
  65000=>"001100101",
  65001=>"111101000",
  65002=>"010101011",
  65003=>"010100111",
  65004=>"100010110",
  65005=>"011010100",
  65006=>"000100100",
  65007=>"001110100",
  65008=>"011111010",
  65009=>"101100101",
  65010=>"000000000",
  65011=>"000101001",
  65012=>"100010111",
  65013=>"001111110",
  65014=>"000010001",
  65015=>"011110011",
  65016=>"010111111",
  65017=>"010011100",
  65018=>"010011111",
  65019=>"010100010",
  65020=>"010111011",
  65021=>"101000000",
  65022=>"100001101",
  65023=>"101000001",
  65024=>"010110110",
  65025=>"001111111",
  65026=>"011010111",
  65027=>"100101101",
  65028=>"010100000",
  65029=>"000001011",
  65030=>"000000011",
  65031=>"011001110",
  65032=>"100101100",
  65033=>"101011011",
  65034=>"111001011",
  65035=>"100111111",
  65036=>"101100011",
  65037=>"010110100",
  65038=>"000111011",
  65039=>"111010001",
  65040=>"010111110",
  65041=>"000110000",
  65042=>"100101101",
  65043=>"111011101",
  65044=>"001000100",
  65045=>"011000110",
  65046=>"010111100",
  65047=>"101111000",
  65048=>"011101110",
  65049=>"111100001",
  65050=>"000100110",
  65051=>"010100010",
  65052=>"001011110",
  65053=>"100101001",
  65054=>"010000111",
  65055=>"100001111",
  65056=>"111111101",
  65057=>"100011100",
  65058=>"010110010",
  65059=>"011100010",
  65060=>"110100110",
  65061=>"111101101",
  65062=>"010010010",
  65063=>"010010001",
  65064=>"001111001",
  65065=>"100001111",
  65066=>"100000101",
  65067=>"100111010",
  65068=>"011011000",
  65069=>"011110110",
  65070=>"110011101",
  65071=>"010010011",
  65072=>"100101000",
  65073=>"101110001",
  65074=>"110001001",
  65075=>"110110111",
  65076=>"100010110",
  65077=>"000100011",
  65078=>"001110001",
  65079=>"101011101",
  65080=>"110010110",
  65081=>"101001111",
  65082=>"100110000",
  65083=>"010110100",
  65084=>"010110110",
  65085=>"100001010",
  65086=>"101111100",
  65087=>"001011000",
  65088=>"101111001",
  65089=>"111000011",
  65090=>"110000000",
  65091=>"110001001",
  65092=>"001100111",
  65093=>"110111101",
  65094=>"000011110",
  65095=>"110001010",
  65096=>"011011101",
  65097=>"001101011",
  65098=>"110010110",
  65099=>"010111110",
  65100=>"001010111",
  65101=>"110010110",
  65102=>"000110101",
  65103=>"011000100",
  65104=>"000110110",
  65105=>"000110011",
  65106=>"000110011",
  65107=>"010110011",
  65108=>"000011001",
  65109=>"100110000",
  65110=>"000110110",
  65111=>"011100011",
  65112=>"110011011",
  65113=>"111000000",
  65114=>"101101011",
  65115=>"010010000",
  65116=>"111110010",
  65117=>"100100110",
  65118=>"000110101",
  65119=>"110111001",
  65120=>"100001111",
  65121=>"111000000",
  65122=>"000010111",
  65123=>"001100010",
  65124=>"100101001",
  65125=>"100111000",
  65126=>"010101100",
  65127=>"111110111",
  65128=>"111001101",
  65129=>"101111001",
  65130=>"010011011",
  65131=>"110101110",
  65132=>"111000111",
  65133=>"000000101",
  65134=>"110001010",
  65135=>"011100010",
  65136=>"000011000",
  65137=>"010001101",
  65138=>"001100011",
  65139=>"100011110",
  65140=>"100101000",
  65141=>"110101010",
  65142=>"100100110",
  65143=>"000110110",
  65144=>"111110111",
  65145=>"010010001",
  65146=>"100010000",
  65147=>"001101000",
  65148=>"101011111",
  65149=>"000100100",
  65150=>"011011111",
  65151=>"011110011",
  65152=>"101111100",
  65153=>"101000100",
  65154=>"001101010",
  65155=>"100101011",
  65156=>"000000011",
  65157=>"011101110",
  65158=>"000101111",
  65159=>"011001011",
  65160=>"000110010",
  65161=>"000100001",
  65162=>"111100101",
  65163=>"110011100",
  65164=>"101110100",
  65165=>"000100010",
  65166=>"101001010",
  65167=>"101111100",
  65168=>"111100010",
  65169=>"101111001",
  65170=>"110010011",
  65171=>"000110110",
  65172=>"010101010",
  65173=>"100100111",
  65174=>"011001001",
  65175=>"110101110",
  65176=>"001000110",
  65177=>"110110000",
  65178=>"000111111",
  65179=>"111000110",
  65180=>"000100110",
  65181=>"100001000",
  65182=>"110011010",
  65183=>"010100010",
  65184=>"010010110",
  65185=>"000110111",
  65186=>"010110110",
  65187=>"010010001",
  65188=>"011111000",
  65189=>"000111101",
  65190=>"001100110",
  65191=>"110100000",
  65192=>"101010011",
  65193=>"000011101",
  65194=>"111110001",
  65195=>"000000000",
  65196=>"001000110",
  65197=>"000010110",
  65198=>"000101101",
  65199=>"000011011",
  65200=>"100111011",
  65201=>"000100101",
  65202=>"100110101",
  65203=>"011100001",
  65204=>"101010100",
  65205=>"001010000",
  65206=>"101101000",
  65207=>"100110110",
  65208=>"010101100",
  65209=>"011001111",
  65210=>"011000001",
  65211=>"100100011",
  65212=>"011111101",
  65213=>"111000111",
  65214=>"111000100",
  65215=>"000110110",
  65216=>"100111100",
  65217=>"100000001",
  65218=>"100100000",
  65219=>"011010100",
  65220=>"100111001",
  65221=>"101100111",
  65222=>"001001000",
  65223=>"011001001",
  65224=>"000100111",
  65225=>"001101100",
  65226=>"010110101",
  65227=>"110011110",
  65228=>"010011110",
  65229=>"101011111",
  65230=>"101010100",
  65231=>"100111001",
  65232=>"110110110",
  65233=>"001111101",
  65234=>"100011110",
  65235=>"010010101",
  65236=>"100000010",
  65237=>"101001111",
  65238=>"010000111",
  65239=>"100000110",
  65240=>"010111100",
  65241=>"001000011",
  65242=>"100010001",
  65243=>"001111000",
  65244=>"101111110",
  65245=>"001111000",
  65246=>"011011111",
  65247=>"111000101",
  65248=>"101101001",
  65249=>"011100101",
  65250=>"100010111",
  65251=>"010100001",
  65252=>"001001101",
  65253=>"011010100",
  65254=>"101011000",
  65255=>"100000000",
  65256=>"000000011",
  65257=>"001000101",
  65258=>"010000111",
  65259=>"010001110",
  65260=>"101100010",
  65261=>"111110111",
  65262=>"100001100",
  65263=>"101101000",
  65264=>"110001110",
  65265=>"101101110",
  65266=>"101111100",
  65267=>"100001101",
  65268=>"010111001",
  65269=>"101110011",
  65270=>"101001001",
  65271=>"011011110",
  65272=>"011001001",
  65273=>"111101111",
  65274=>"101001100",
  65275=>"110101100",
  65276=>"111001111",
  65277=>"010000011",
  65278=>"111001101",
  65279=>"111100000",
  65280=>"000010010",
  65281=>"101011101",
  65282=>"011001100",
  65283=>"111000001",
  65284=>"111111111",
  65285=>"001000001",
  65286=>"111111111",
  65287=>"110101100",
  65288=>"001110110",
  65289=>"101100001",
  65290=>"111111011",
  65291=>"111001110",
  65292=>"001101011",
  65293=>"101101111",
  65294=>"011111111",
  65295=>"111001110",
  65296=>"100110100",
  65297=>"100100111",
  65298=>"011001011",
  65299=>"011100100",
  65300=>"111101001",
  65301=>"011001101",
  65302=>"011000011",
  65303=>"001010011",
  65304=>"101101100",
  65305=>"000000111",
  65306=>"100010010",
  65307=>"000010011",
  65308=>"001001111",
  65309=>"010010101",
  65310=>"100010111",
  65311=>"101101000",
  65312=>"000100010",
  65313=>"000000011",
  65314=>"101000101",
  65315=>"111100010",
  65316=>"111100100",
  65317=>"011100000",
  65318=>"101010011",
  65319=>"101110110",
  65320=>"111111100",
  65321=>"110101101",
  65322=>"011101110",
  65323=>"011011010",
  65324=>"111111000",
  65325=>"000000110",
  65326=>"110110100",
  65327=>"000000000",
  65328=>"000110001",
  65329=>"011100000",
  65330=>"100011011",
  65331=>"101111001",
  65332=>"100010011",
  65333=>"110110011",
  65334=>"100110110",
  65335=>"001100010",
  65336=>"111101110",
  65337=>"000000110",
  65338=>"011000110",
  65339=>"101010101",
  65340=>"110011011",
  65341=>"000000010",
  65342=>"000000000",
  65343=>"101001101",
  65344=>"001110000",
  65345=>"010111111",
  65346=>"100111111",
  65347=>"000110110",
  65348=>"111000110",
  65349=>"011101011",
  65350=>"100111110",
  65351=>"000100110",
  65352=>"100001101",
  65353=>"101100001",
  65354=>"111100110",
  65355=>"100101001",
  65356=>"100011010",
  65357=>"000010110",
  65358=>"100010010",
  65359=>"111111001",
  65360=>"100110110",
  65361=>"101001001",
  65362=>"010000111",
  65363=>"001111110",
  65364=>"101000100",
  65365=>"101111010",
  65366=>"011010111",
  65367=>"000110000",
  65368=>"100101111",
  65369=>"011000100",
  65370=>"011111111",
  65371=>"110110010",
  65372=>"101100000",
  65373=>"011011010",
  65374=>"001001010",
  65375=>"001000011",
  65376=>"110000010",
  65377=>"110000101",
  65378=>"111101111",
  65379=>"110101000",
  65380=>"001001001",
  65381=>"010100000",
  65382=>"101010111",
  65383=>"100101110",
  65384=>"011000001",
  65385=>"101000010",
  65386=>"110100101",
  65387=>"111000101",
  65388=>"011011110",
  65389=>"010001000",
  65390=>"101100000",
  65391=>"011000001",
  65392=>"001001111",
  65393=>"011101011",
  65394=>"011111001",
  65395=>"110100011",
  65396=>"100010100",
  65397=>"011111111",
  65398=>"011100111",
  65399=>"001110001",
  65400=>"110001001",
  65401=>"000010011",
  65402=>"001001101",
  65403=>"001111000",
  65404=>"000110000",
  65405=>"101010101",
  65406=>"110010110",
  65407=>"101101101",
  65408=>"000101011",
  65409=>"000001001",
  65410=>"101011100",
  65411=>"000110010",
  65412=>"111110010",
  65413=>"110010000",
  65414=>"100010111",
  65415=>"110100001",
  65416=>"100111010",
  65417=>"110110100",
  65418=>"000000101",
  65419=>"001000011",
  65420=>"111001011",
  65421=>"101110001",
  65422=>"001000010",
  65423=>"101001001",
  65424=>"111100011",
  65425=>"100000111",
  65426=>"000001011",
  65427=>"110110101",
  65428=>"100110101",
  65429=>"010111100",
  65430=>"000110111",
  65431=>"001000110",
  65432=>"110010110",
  65433=>"100110100",
  65434=>"111110011",
  65435=>"100011101",
  65436=>"000011110",
  65437=>"000110001",
  65438=>"011100110",
  65439=>"111111111",
  65440=>"001111001",
  65441=>"001111000",
  65442=>"110111110",
  65443=>"110011000",
  65444=>"101010000",
  65445=>"000111010",
  65446=>"100001001",
  65447=>"000101111",
  65448=>"000011011",
  65449=>"010000111",
  65450=>"100011110",
  65451=>"100101010",
  65452=>"110011001",
  65453=>"010101010",
  65454=>"111100101",
  65455=>"101111001",
  65456=>"111110111",
  65457=>"101110110",
  65458=>"111101001",
  65459=>"001001011",
  65460=>"111001101",
  65461=>"100010100",
  65462=>"001101100",
  65463=>"011101111",
  65464=>"100100111",
  65465=>"110001001",
  65466=>"111001010",
  65467=>"101100111",
  65468=>"000000110",
  65469=>"000101010",
  65470=>"010010001",
  65471=>"010100010",
  65472=>"010000011",
  65473=>"001010000",
  65474=>"010111100",
  65475=>"000000110",
  65476=>"111000111",
  65477=>"100101110",
  65478=>"111001000",
  65479=>"011001101",
  65480=>"100111001",
  65481=>"011111011",
  65482=>"010001001",
  65483=>"100111110",
  65484=>"010010001",
  65485=>"000100111",
  65486=>"100010100",
  65487=>"101111001",
  65488=>"100111010",
  65489=>"100010000",
  65490=>"101111011",
  65491=>"010111110",
  65492=>"010001000",
  65493=>"111111001",
  65494=>"110000101",
  65495=>"111101011",
  65496=>"101100011",
  65497=>"000100000",
  65498=>"111000011",
  65499=>"101100110",
  65500=>"110110010",
  65501=>"110010111",
  65502=>"010001101",
  65503=>"100100111",
  65504=>"011001100",
  65505=>"100010111",
  65506=>"011011111",
  65507=>"101100010",
  65508=>"101100011",
  65509=>"001110100",
  65510=>"111010101",
  65511=>"001000000",
  65512=>"001000010",
  65513=>"000000001",
  65514=>"001000110",
  65515=>"110100111",
  65516=>"000000011",
  65517=>"110010010",
  65518=>"000001100",
  65519=>"010111101",
  65520=>"010100010",
  65521=>"000101111",
  65522=>"110011011",
  65523=>"100111001",
  65524=>"011111110",
  65525=>"001011011",
  65526=>"001010001",
  65527=>"000100000",
  65528=>"011001011",
  65529=>"111111111",
  65530=>"101010111",
  65531=>"011011010",
  65532=>"000111101",
  65533=>"011101111",
  65534=>"101001111",
  65535=>"011101011");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;