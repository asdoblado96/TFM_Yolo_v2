LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_2_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_2_WROM;

ARCHITECTURE RTL OF L8_2_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"111000000",
  1=>"000011111",
  2=>"101010011",
  3=>"010100100",
  4=>"010010111",
  5=>"110001010",
  6=>"000001101",
  7=>"101100010",
  8=>"000001110",
  9=>"010000111",
  10=>"001101100",
  11=>"101000010",
  12=>"110011000",
  13=>"001110100",
  14=>"110110011",
  15=>"111010010",
  16=>"000000001",
  17=>"001011111",
  18=>"101111110",
  19=>"000100011",
  20=>"000000011",
  21=>"000101100",
  22=>"110000010",
  23=>"111001010",
  24=>"101001100",
  25=>"110011011",
  26=>"111101110",
  27=>"110110111",
  28=>"001000001",
  29=>"010000101",
  30=>"101111010",
  31=>"000101010",
  32=>"100110111",
  33=>"000001100",
  34=>"101011100",
  35=>"110101011",
  36=>"010001000",
  37=>"100001110",
  38=>"110110100",
  39=>"100010101",
  40=>"000111010",
  41=>"100001000",
  42=>"010011000",
  43=>"001110001",
  44=>"111111011",
  45=>"101011110",
  46=>"011111010",
  47=>"011010011",
  48=>"011101010",
  49=>"111010111",
  50=>"101110000",
  51=>"111101010",
  52=>"000000000",
  53=>"110001001",
  54=>"111101111",
  55=>"011111110",
  56=>"000010101",
  57=>"001110110",
  58=>"000100011",
  59=>"000001101",
  60=>"000011111",
  61=>"010100111",
  62=>"101010001",
  63=>"001110111",
  64=>"110000100",
  65=>"000001010",
  66=>"000000110",
  67=>"110110010",
  68=>"000010110",
  69=>"010000010",
  70=>"100100101",
  71=>"010001101",
  72=>"111001000",
  73=>"101110000",
  74=>"001100000",
  75=>"011100001",
  76=>"001011110",
  77=>"111010001",
  78=>"000111111",
  79=>"111000001",
  80=>"100010101",
  81=>"111111000",
  82=>"111010001",
  83=>"001100001",
  84=>"000000000",
  85=>"011000100",
  86=>"011110000",
  87=>"110100111",
  88=>"000001101",
  89=>"001100101",
  90=>"110000111",
  91=>"011011000",
  92=>"000000000",
  93=>"010111011",
  94=>"100010010",
  95=>"010000000",
  96=>"100100100",
  97=>"111011000",
  98=>"001011000",
  99=>"100100111",
  100=>"110100100",
  101=>"000001011",
  102=>"011000100",
  103=>"000001010",
  104=>"011001111",
  105=>"010110100",
  106=>"110001010",
  107=>"000101011",
  108=>"000110010",
  109=>"000100001",
  110=>"010000111",
  111=>"000101001",
  112=>"000001000",
  113=>"001110100",
  114=>"010110000",
  115=>"001101111",
  116=>"001111110",
  117=>"101001010",
  118=>"100000001",
  119=>"110110111",
  120=>"010010111",
  121=>"100111101",
  122=>"101000110",
  123=>"101001110",
  124=>"010101011",
  125=>"000001011",
  126=>"100101110",
  127=>"011110010",
  128=>"001110011",
  129=>"000111111",
  130=>"001010010",
  131=>"101100001",
  132=>"111001100",
  133=>"011010100",
  134=>"000000011",
  135=>"001100011",
  136=>"101110110",
  137=>"111010001",
  138=>"000000001",
  139=>"000110110",
  140=>"000101101",
  141=>"011000011",
  142=>"101110000",
  143=>"101011011",
  144=>"100010011",
  145=>"101001010",
  146=>"001111110",
  147=>"100111011",
  148=>"000010110",
  149=>"000100011",
  150=>"100100110",
  151=>"101011010",
  152=>"010000011",
  153=>"110011110",
  154=>"000010000",
  155=>"001101011",
  156=>"100111010",
  157=>"011000011",
  158=>"100000000",
  159=>"110001100",
  160=>"011111100",
  161=>"111101100",
  162=>"010101011",
  163=>"001010100",
  164=>"101110111",
  165=>"111001101",
  166=>"000101111",
  167=>"000000100",
  168=>"101011011",
  169=>"101110111",
  170=>"100011110",
  171=>"100100110",
  172=>"000001010",
  173=>"010100110",
  174=>"101100010",
  175=>"110001110",
  176=>"011010001",
  177=>"000001001",
  178=>"101111100",
  179=>"001110110",
  180=>"001010100",
  181=>"010000000",
  182=>"010000000",
  183=>"101111111",
  184=>"001100111",
  185=>"001011000",
  186=>"100001011",
  187=>"000111011",
  188=>"010010011",
  189=>"110011011",
  190=>"000100111",
  191=>"101011001",
  192=>"000101011",
  193=>"011001110",
  194=>"011000000",
  195=>"110011110",
  196=>"111101011",
  197=>"100101100",
  198=>"101001111",
  199=>"010001110",
  200=>"000101000",
  201=>"111010101",
  202=>"001100111",
  203=>"100101100",
  204=>"011011110",
  205=>"110011110",
  206=>"101000001",
  207=>"010010101",
  208=>"000111001",
  209=>"100111001",
  210=>"011000000",
  211=>"000010010",
  212=>"001001111",
  213=>"101110111",
  214=>"001011110",
  215=>"001101010",
  216=>"000100001",
  217=>"111111100",
  218=>"010100111",
  219=>"110110111",
  220=>"010010101",
  221=>"011011111",
  222=>"101010110",
  223=>"101000111",
  224=>"000001011",
  225=>"011001111",
  226=>"010101010",
  227=>"111100111",
  228=>"110111111",
  229=>"010110100",
  230=>"010000000",
  231=>"101011000",
  232=>"011101011",
  233=>"111001010",
  234=>"101001011",
  235=>"111101100",
  236=>"000111110",
  237=>"000110001",
  238=>"100001010",
  239=>"111111100",
  240=>"110101111",
  241=>"111001001",
  242=>"000000011",
  243=>"000000100",
  244=>"101111010",
  245=>"010111100",
  246=>"011000010",
  247=>"100110100",
  248=>"010011010",
  249=>"011011011",
  250=>"010001100",
  251=>"011100000",
  252=>"001000111",
  253=>"100011010",
  254=>"110000110",
  255=>"000110010",
  256=>"011110111",
  257=>"111111101",
  258=>"110001000",
  259=>"000110110",
  260=>"111101101",
  261=>"001101001",
  262=>"110111111",
  263=>"100010010",
  264=>"101100100",
  265=>"000000001",
  266=>"000110000",
  267=>"001100011",
  268=>"011101000",
  269=>"111000111",
  270=>"001000000",
  271=>"011111000",
  272=>"111011101",
  273=>"101101100",
  274=>"111101010",
  275=>"000010101",
  276=>"100100111",
  277=>"011110101",
  278=>"101011011",
  279=>"011010000",
  280=>"110111100",
  281=>"001010101",
  282=>"100000001",
  283=>"010001100",
  284=>"110101100",
  285=>"111011000",
  286=>"111101101",
  287=>"100100000",
  288=>"100101110",
  289=>"001101011",
  290=>"111001111",
  291=>"000111000",
  292=>"110010110",
  293=>"010011010",
  294=>"000010101",
  295=>"110011001",
  296=>"000101110",
  297=>"110111100",
  298=>"100111101",
  299=>"001010000",
  300=>"000010100",
  301=>"011111011",
  302=>"101011010",
  303=>"100010000",
  304=>"000111011",
  305=>"011111011",
  306=>"111111111",
  307=>"001000111",
  308=>"101100001",
  309=>"011100001",
  310=>"001100111",
  311=>"010000111",
  312=>"110100110",
  313=>"100100101",
  314=>"100001000",
  315=>"111111011",
  316=>"000000101",
  317=>"000100010",
  318=>"100010001",
  319=>"101111011",
  320=>"010110001",
  321=>"101101111",
  322=>"111110001",
  323=>"100001100",
  324=>"010000010",
  325=>"001011100",
  326=>"010100100",
  327=>"111000100",
  328=>"100000000",
  329=>"101000010",
  330=>"110100010",
  331=>"110100011",
  332=>"111100101",
  333=>"000000010",
  334=>"001000111",
  335=>"000001000",
  336=>"010010111",
  337=>"000110101",
  338=>"000000010",
  339=>"000010000",
  340=>"100000000",
  341=>"110111111",
  342=>"111111111",
  343=>"111100101",
  344=>"000001111",
  345=>"001010111",
  346=>"001110011",
  347=>"110110110",
  348=>"000011101",
  349=>"111110000",
  350=>"101010100",
  351=>"101110011",
  352=>"110111111",
  353=>"010011101",
  354=>"010010011",
  355=>"011000000",
  356=>"000000100",
  357=>"011010001",
  358=>"000010011",
  359=>"101111001",
  360=>"111001101",
  361=>"101010001",
  362=>"001101010",
  363=>"010110000",
  364=>"001101101",
  365=>"010011111",
  366=>"110110010",
  367=>"000110011",
  368=>"001100000",
  369=>"110001101",
  370=>"000111000",
  371=>"010110010",
  372=>"111011101",
  373=>"001000101",
  374=>"010011001",
  375=>"110100110",
  376=>"000000011",
  377=>"001011100",
  378=>"101001110",
  379=>"111100111",
  380=>"000011001",
  381=>"111101011",
  382=>"010001111",
  383=>"111001111",
  384=>"101111011",
  385=>"100100000",
  386=>"100101110",
  387=>"010111011",
  388=>"110011100",
  389=>"100011000",
  390=>"111100100",
  391=>"000000001",
  392=>"000001000",
  393=>"101111101",
  394=>"110010101",
  395=>"100100111",
  396=>"110100011",
  397=>"001011011",
  398=>"111001010",
  399=>"111100100",
  400=>"010101100",
  401=>"000000000",
  402=>"110110101",
  403=>"111001111",
  404=>"001100001",
  405=>"011100000",
  406=>"100110000",
  407=>"010101100",
  408=>"000010111",
  409=>"000010000",
  410=>"110100010",
  411=>"111101001",
  412=>"111011001",
  413=>"000100000",
  414=>"000001101",
  415=>"000101101",
  416=>"111000001",
  417=>"100111000",
  418=>"101110110",
  419=>"001000100",
  420=>"101010101",
  421=>"010000110",
  422=>"111000100",
  423=>"000111000",
  424=>"001110100",
  425=>"001011001",
  426=>"110000001",
  427=>"010111101",
  428=>"110100000",
  429=>"110111101",
  430=>"011000011",
  431=>"010110100",
  432=>"100100000",
  433=>"010000010",
  434=>"010010001",
  435=>"111101110",
  436=>"000100010",
  437=>"111100010",
  438=>"111000101",
  439=>"110101010",
  440=>"001111110",
  441=>"110000011",
  442=>"100000000",
  443=>"110111100",
  444=>"001101110",
  445=>"011100111",
  446=>"000001000",
  447=>"111111000",
  448=>"011010011",
  449=>"011100001",
  450=>"010001100",
  451=>"111110000",
  452=>"000000010",
  453=>"101101111",
  454=>"101111011",
  455=>"000001010",
  456=>"000100000",
  457=>"101011011",
  458=>"011111010",
  459=>"001010101",
  460=>"101001110",
  461=>"100100011",
  462=>"011011001",
  463=>"011110111",
  464=>"111011001",
  465=>"001001111",
  466=>"101011000",
  467=>"001111000",
  468=>"111100001",
  469=>"000110101",
  470=>"000010011",
  471=>"100010100",
  472=>"111000000",
  473=>"011010000",
  474=>"100100000",
  475=>"111001100",
  476=>"001100100",
  477=>"011001010",
  478=>"000111110",
  479=>"111011111",
  480=>"001010001",
  481=>"111100011",
  482=>"011010010",
  483=>"010001001",
  484=>"110111110",
  485=>"110111101",
  486=>"000110110",
  487=>"111100100",
  488=>"111110000",
  489=>"101101011",
  490=>"010001001",
  491=>"101111110",
  492=>"010110001",
  493=>"000110001",
  494=>"000000001",
  495=>"011000100",
  496=>"011000101",
  497=>"000011000",
  498=>"111010011",
  499=>"110110000",
  500=>"110101100",
  501=>"111100011",
  502=>"011100101",
  503=>"111011111",
  504=>"000001010",
  505=>"110000001",
  506=>"010010011",
  507=>"110101001",
  508=>"101011100",
  509=>"010010001",
  510=>"001111011",
  511=>"010110111",
  512=>"111110010",
  513=>"001001001",
  514=>"100100101",
  515=>"010100100",
  516=>"100100010",
  517=>"000111001",
  518=>"100010001",
  519=>"001111000",
  520=>"001100000",
  521=>"100110101",
  522=>"010101010",
  523=>"001001100",
  524=>"011101111",
  525=>"111110010",
  526=>"010110010",
  527=>"010011101",
  528=>"011000000",
  529=>"000111111",
  530=>"100101011",
  531=>"101010011",
  532=>"010001001",
  533=>"110111011",
  534=>"010110100",
  535=>"101111010",
  536=>"111010100",
  537=>"011110110",
  538=>"110111000",
  539=>"000001111",
  540=>"000011000",
  541=>"101001100",
  542=>"011110101",
  543=>"100000111",
  544=>"000100111",
  545=>"110011111",
  546=>"000111101",
  547=>"011100101",
  548=>"110110111",
  549=>"111111101",
  550=>"001101011",
  551=>"111010000",
  552=>"001010001",
  553=>"000100111",
  554=>"100100010",
  555=>"010010010",
  556=>"001011011",
  557=>"000001110",
  558=>"011010010",
  559=>"000101001",
  560=>"000111001",
  561=>"011011100",
  562=>"101101001",
  563=>"011111000",
  564=>"101110100",
  565=>"100101111",
  566=>"100011011",
  567=>"110111001",
  568=>"100110010",
  569=>"110110100",
  570=>"110111101",
  571=>"100111111",
  572=>"110010010",
  573=>"111010011",
  574=>"111001011",
  575=>"100000001",
  576=>"110101100",
  577=>"001001011",
  578=>"001100010",
  579=>"101111001",
  580=>"101100110",
  581=>"011000000",
  582=>"010001100",
  583=>"100000000",
  584=>"000110100",
  585=>"110111010",
  586=>"000001100",
  587=>"000110011",
  588=>"000010000",
  589=>"001010100",
  590=>"101101101",
  591=>"010011001",
  592=>"110000000",
  593=>"100101111",
  594=>"110011010",
  595=>"101000010",
  596=>"111010010",
  597=>"101110100",
  598=>"011100010",
  599=>"010110010",
  600=>"100010100",
  601=>"000010001",
  602=>"010100101",
  603=>"110111110",
  604=>"100110110",
  605=>"001100100",
  606=>"100110101",
  607=>"010001100",
  608=>"110110001",
  609=>"101100011",
  610=>"010101010",
  611=>"100110010",
  612=>"001010010",
  613=>"000111010",
  614=>"111001001",
  615=>"001010011",
  616=>"011111111",
  617=>"110111110",
  618=>"000001110",
  619=>"111101010",
  620=>"101110011",
  621=>"110101011",
  622=>"111101101",
  623=>"101001101",
  624=>"101001100",
  625=>"111010011",
  626=>"011100001",
  627=>"011100110",
  628=>"100111101",
  629=>"011110011",
  630=>"101001100",
  631=>"111010100",
  632=>"101000110",
  633=>"000010011",
  634=>"011011000",
  635=>"111100110",
  636=>"100101000",
  637=>"111110100",
  638=>"010101010",
  639=>"101000111",
  640=>"000000100",
  641=>"111001001",
  642=>"010001011",
  643=>"001000001",
  644=>"111010011",
  645=>"110101110",
  646=>"110101011",
  647=>"100101011",
  648=>"100000100",
  649=>"001100010",
  650=>"101101101",
  651=>"101001101",
  652=>"110011101",
  653=>"001001111",
  654=>"010001110",
  655=>"100010101",
  656=>"110101001",
  657=>"011101000",
  658=>"001001111",
  659=>"001101011",
  660=>"101001101",
  661=>"100101011",
  662=>"010111101",
  663=>"001001110",
  664=>"111111100",
  665=>"001110001",
  666=>"100111101",
  667=>"100100000",
  668=>"110001100",
  669=>"011010001",
  670=>"000011010",
  671=>"010110000",
  672=>"001000001",
  673=>"100110111",
  674=>"111000101",
  675=>"100001101",
  676=>"000101111",
  677=>"110110101",
  678=>"000001010",
  679=>"000001101",
  680=>"100001000",
  681=>"010010001",
  682=>"000000111",
  683=>"110001100",
  684=>"101010100",
  685=>"011010010",
  686=>"010001111",
  687=>"010100001",
  688=>"011010100",
  689=>"001010011",
  690=>"000010011",
  691=>"100001111",
  692=>"111010111",
  693=>"000111010",
  694=>"011010000",
  695=>"110011001",
  696=>"111000101",
  697=>"100110110",
  698=>"100010111",
  699=>"100011100",
  700=>"110010110",
  701=>"000000000",
  702=>"111001011",
  703=>"001000000",
  704=>"100001011",
  705=>"101111000",
  706=>"111000111",
  707=>"001110100",
  708=>"001100000",
  709=>"101011101",
  710=>"010110000",
  711=>"000100111",
  712=>"110000001",
  713=>"111010100",
  714=>"101011100",
  715=>"101100100",
  716=>"011111001",
  717=>"110010001",
  718=>"110010111",
  719=>"000001001",
  720=>"101101111",
  721=>"001000100",
  722=>"101000111",
  723=>"010010110",
  724=>"001111011",
  725=>"000000000",
  726=>"100110011",
  727=>"000011100",
  728=>"010101110",
  729=>"101010101",
  730=>"110101000",
  731=>"111000001",
  732=>"110011111",
  733=>"000001010",
  734=>"000001010",
  735=>"101100011",
  736=>"011111111",
  737=>"101000011",
  738=>"011110100",
  739=>"100111011",
  740=>"011010100",
  741=>"110110001",
  742=>"000101111",
  743=>"010000100",
  744=>"110010000",
  745=>"011001010",
  746=>"011111100",
  747=>"010010101",
  748=>"000111001",
  749=>"111110100",
  750=>"100100011",
  751=>"011000010",
  752=>"010100101",
  753=>"000010111",
  754=>"100100100",
  755=>"001000100",
  756=>"000101001",
  757=>"000010011",
  758=>"100101010",
  759=>"111101111",
  760=>"000010111",
  761=>"101110111",
  762=>"011001101",
  763=>"111011100",
  764=>"010111100",
  765=>"001110111",
  766=>"011000011",
  767=>"011100111",
  768=>"010011111",
  769=>"000110001",
  770=>"101000110",
  771=>"000011000",
  772=>"011000000",
  773=>"110001110",
  774=>"001010110",
  775=>"110010011",
  776=>"011110111",
  777=>"110111111",
  778=>"100000101",
  779=>"101010001",
  780=>"001110001",
  781=>"111011101",
  782=>"110101010",
  783=>"011001100",
  784=>"101001001",
  785=>"101110001",
  786=>"100011100",
  787=>"110010000",
  788=>"101011110",
  789=>"111000111",
  790=>"010111111",
  791=>"011101111",
  792=>"000000011",
  793=>"001001000",
  794=>"000000100",
  795=>"001010111",
  796=>"100110100",
  797=>"011011010",
  798=>"110100100",
  799=>"010110101",
  800=>"010000101",
  801=>"011010111",
  802=>"001111000",
  803=>"001000111",
  804=>"101110000",
  805=>"101010001",
  806=>"110010101",
  807=>"000101010",
  808=>"101011111",
  809=>"000010000",
  810=>"111111110",
  811=>"011101011",
  812=>"011110110",
  813=>"010100010",
  814=>"110110100",
  815=>"110000110",
  816=>"010101011",
  817=>"000101011",
  818=>"011101101",
  819=>"111111111",
  820=>"110010101",
  821=>"111011010",
  822=>"111111111",
  823=>"010100001",
  824=>"000010110",
  825=>"011010000",
  826=>"101100101",
  827=>"101111111",
  828=>"000110001",
  829=>"110100111",
  830=>"111011100",
  831=>"101110111",
  832=>"010111011",
  833=>"101011000",
  834=>"101010001",
  835=>"111011000",
  836=>"011001011",
  837=>"101001111",
  838=>"001111110",
  839=>"000100111",
  840=>"100001000",
  841=>"111101101",
  842=>"011101000",
  843=>"011110110",
  844=>"001101010",
  845=>"011000110",
  846=>"010110101",
  847=>"101011101",
  848=>"111110010",
  849=>"010001101",
  850=>"000110110",
  851=>"111010010",
  852=>"010111100",
  853=>"101001111",
  854=>"011000010",
  855=>"011011000",
  856=>"001011001",
  857=>"101000111",
  858=>"010001011",
  859=>"110010100",
  860=>"110010011",
  861=>"111101101",
  862=>"000101110",
  863=>"010001101",
  864=>"101011101",
  865=>"011000000",
  866=>"001000100",
  867=>"100010110",
  868=>"000010010",
  869=>"011110101",
  870=>"000011110",
  871=>"111110101",
  872=>"111010010",
  873=>"010011101",
  874=>"011111111",
  875=>"111000000",
  876=>"001011100",
  877=>"010000001",
  878=>"010001110",
  879=>"111111100",
  880=>"010000101",
  881=>"111000101",
  882=>"100110010",
  883=>"110100111",
  884=>"111100111",
  885=>"000110010",
  886=>"010101001",
  887=>"010101101",
  888=>"010100100",
  889=>"011001010",
  890=>"100101000",
  891=>"101010001",
  892=>"000001010",
  893=>"100100011",
  894=>"001110110",
  895=>"011100001",
  896=>"011001001",
  897=>"101001001",
  898=>"000001000",
  899=>"100000010",
  900=>"101111001",
  901=>"011111011",
  902=>"110100010",
  903=>"011110010",
  904=>"000100000",
  905=>"011011111",
  906=>"000110110",
  907=>"000010101",
  908=>"010000000",
  909=>"010011100",
  910=>"101100001",
  911=>"111110110",
  912=>"111000001",
  913=>"001000010",
  914=>"001010101",
  915=>"001101011",
  916=>"100001010",
  917=>"110110100",
  918=>"101000000",
  919=>"011010001",
  920=>"011001101",
  921=>"000010110",
  922=>"100001001",
  923=>"001111110",
  924=>"000100101",
  925=>"010010101",
  926=>"001010111",
  927=>"000111011",
  928=>"101001101",
  929=>"111000010",
  930=>"001001100",
  931=>"001011010",
  932=>"101011000",
  933=>"000011000",
  934=>"010100000",
  935=>"000001000",
  936=>"110101001",
  937=>"001000101",
  938=>"011010000",
  939=>"001101101",
  940=>"110100001",
  941=>"000101111",
  942=>"011101011",
  943=>"101001111",
  944=>"101000101",
  945=>"101000010",
  946=>"001000110",
  947=>"010110001",
  948=>"110110100",
  949=>"001010010",
  950=>"001000000",
  951=>"111111101",
  952=>"110010100",
  953=>"001010101",
  954=>"110101110",
  955=>"000100000",
  956=>"000001001",
  957=>"111110000",
  958=>"100111111",
  959=>"011100010",
  960=>"101110011",
  961=>"001010011",
  962=>"100111001",
  963=>"000100010",
  964=>"111110000",
  965=>"000000010",
  966=>"101101000",
  967=>"001101111",
  968=>"001010110",
  969=>"111011100",
  970=>"000110110",
  971=>"010011101",
  972=>"111110111",
  973=>"110101011",
  974=>"010000000",
  975=>"111110000",
  976=>"000011011",
  977=>"001110011",
  978=>"101110101",
  979=>"010011010",
  980=>"111101001",
  981=>"101001111",
  982=>"010010110",
  983=>"000111011",
  984=>"101010101",
  985=>"100000001",
  986=>"101001011",
  987=>"101111101",
  988=>"001010000",
  989=>"010011011",
  990=>"101100010",
  991=>"011111101",
  992=>"101000001",
  993=>"011110010",
  994=>"100101111",
  995=>"011010011",
  996=>"000000001",
  997=>"110000011",
  998=>"111010001",
  999=>"100000111",
  1000=>"001011111",
  1001=>"011110000",
  1002=>"000110000",
  1003=>"110000110",
  1004=>"111111011",
  1005=>"011010100",
  1006=>"010101011",
  1007=>"001100001",
  1008=>"010000011",
  1009=>"000010000",
  1010=>"101110000",
  1011=>"011010101",
  1012=>"100111100",
  1013=>"011110011",
  1014=>"111101000",
  1015=>"100101011",
  1016=>"011110000",
  1017=>"011001001",
  1018=>"111111001",
  1019=>"000000110",
  1020=>"001001000",
  1021=>"000101000",
  1022=>"110001100",
  1023=>"001000000",
  1024=>"100101000",
  1025=>"111111001",
  1026=>"111000101",
  1027=>"001100100",
  1028=>"001111110",
  1029=>"010111110",
  1030=>"111110111",
  1031=>"000110110",
  1032=>"111111001",
  1033=>"011011000",
  1034=>"101100110",
  1035=>"101000101",
  1036=>"101101010",
  1037=>"001000011",
  1038=>"011011010",
  1039=>"000001010",
  1040=>"111010010",
  1041=>"010001100",
  1042=>"101111000",
  1043=>"101101111",
  1044=>"010000010",
  1045=>"001010110",
  1046=>"010100101",
  1047=>"001100011",
  1048=>"001100111",
  1049=>"001000011",
  1050=>"100111011",
  1051=>"111101101",
  1052=>"000001101",
  1053=>"011010110",
  1054=>"011111100",
  1055=>"111001001",
  1056=>"001011100",
  1057=>"000110110",
  1058=>"000110111",
  1059=>"011010110",
  1060=>"110101010",
  1061=>"101110011",
  1062=>"010000000",
  1063=>"100110100",
  1064=>"000000111",
  1065=>"001110000",
  1066=>"111100001",
  1067=>"000111111",
  1068=>"011110000",
  1069=>"011100101",
  1070=>"100010100",
  1071=>"001001001",
  1072=>"100101110",
  1073=>"001011000",
  1074=>"100010001",
  1075=>"000000100",
  1076=>"100100000",
  1077=>"001010001",
  1078=>"000000001",
  1079=>"010100100",
  1080=>"011101111",
  1081=>"001010001",
  1082=>"100011100",
  1083=>"101001001",
  1084=>"000011001",
  1085=>"000110100",
  1086=>"001101011",
  1087=>"100010000",
  1088=>"000011000",
  1089=>"100101010",
  1090=>"011001011",
  1091=>"101100100",
  1092=>"001111010",
  1093=>"100001101",
  1094=>"110100011",
  1095=>"111010110",
  1096=>"111111110",
  1097=>"011110000",
  1098=>"111010011",
  1099=>"001010000",
  1100=>"001001110",
  1101=>"011100011",
  1102=>"010001111",
  1103=>"101100110",
  1104=>"100001100",
  1105=>"100001100",
  1106=>"101111110",
  1107=>"111010011",
  1108=>"001110110",
  1109=>"101111111",
  1110=>"001100101",
  1111=>"100101101",
  1112=>"110000010",
  1113=>"100011000",
  1114=>"111111001",
  1115=>"001000000",
  1116=>"001001010",
  1117=>"001010100",
  1118=>"100001001",
  1119=>"000101101",
  1120=>"001011111",
  1121=>"010000110",
  1122=>"111001011",
  1123=>"110101110",
  1124=>"111110110",
  1125=>"100011010",
  1126=>"001001100",
  1127=>"011100011",
  1128=>"010110110",
  1129=>"110110100",
  1130=>"100100100",
  1131=>"011110010",
  1132=>"110011001",
  1133=>"000110100",
  1134=>"001000100",
  1135=>"000001111",
  1136=>"001110101",
  1137=>"100000001",
  1138=>"101001011",
  1139=>"001101100",
  1140=>"101100011",
  1141=>"111101110",
  1142=>"111000001",
  1143=>"110010000",
  1144=>"111001000",
  1145=>"111111100",
  1146=>"110111110",
  1147=>"001111110",
  1148=>"000100001",
  1149=>"111111011",
  1150=>"001100010",
  1151=>"001011100",
  1152=>"000010100",
  1153=>"001110100",
  1154=>"010001000",
  1155=>"101000110",
  1156=>"110111000",
  1157=>"100010110",
  1158=>"111010111",
  1159=>"000100011",
  1160=>"100101000",
  1161=>"000110000",
  1162=>"101100010",
  1163=>"000011011",
  1164=>"010100111",
  1165=>"000000011",
  1166=>"111101000",
  1167=>"111110100",
  1168=>"010111001",
  1169=>"111001101",
  1170=>"000001011",
  1171=>"000010100",
  1172=>"000000100",
  1173=>"010111101",
  1174=>"101011101",
  1175=>"101000110",
  1176=>"101000110",
  1177=>"011001110",
  1178=>"001001000",
  1179=>"011110010",
  1180=>"110110111",
  1181=>"100100100",
  1182=>"001101101",
  1183=>"111101011",
  1184=>"010101010",
  1185=>"110010010",
  1186=>"101100000",
  1187=>"000101101",
  1188=>"101110100",
  1189=>"001000110",
  1190=>"100000011",
  1191=>"011100100",
  1192=>"010001011",
  1193=>"000011111",
  1194=>"101100101",
  1195=>"011001110",
  1196=>"011010100",
  1197=>"101001000",
  1198=>"100100110",
  1199=>"101110110",
  1200=>"011101011",
  1201=>"010010001",
  1202=>"000111110",
  1203=>"110001110",
  1204=>"011011100",
  1205=>"101110011",
  1206=>"101001100",
  1207=>"100001010",
  1208=>"101101101",
  1209=>"101101100",
  1210=>"001011100",
  1211=>"111100110",
  1212=>"110101011",
  1213=>"110010101",
  1214=>"000011100",
  1215=>"011100010",
  1216=>"010111011",
  1217=>"100100110",
  1218=>"101010100",
  1219=>"111011010",
  1220=>"111000110",
  1221=>"101111111",
  1222=>"001101101",
  1223=>"011000010",
  1224=>"111001001",
  1225=>"010110001",
  1226=>"110110101",
  1227=>"111000001",
  1228=>"001111010",
  1229=>"111110100",
  1230=>"110011000",
  1231=>"000100100",
  1232=>"111100000",
  1233=>"110110000",
  1234=>"000000001",
  1235=>"100101001",
  1236=>"110001000",
  1237=>"001111110",
  1238=>"100110010",
  1239=>"110110110",
  1240=>"110011100",
  1241=>"111111001",
  1242=>"000100001",
  1243=>"000111001",
  1244=>"001011000",
  1245=>"001110001",
  1246=>"011000000",
  1247=>"000011000",
  1248=>"100000011",
  1249=>"100010010",
  1250=>"111100011",
  1251=>"110111111",
  1252=>"001011000",
  1253=>"000111000",
  1254=>"110011100",
  1255=>"100111110",
  1256=>"010110100",
  1257=>"111100010",
  1258=>"001110011",
  1259=>"000010101",
  1260=>"000111010",
  1261=>"110001110",
  1262=>"110001100",
  1263=>"011111011",
  1264=>"111000001",
  1265=>"001101100",
  1266=>"000101111",
  1267=>"010011110",
  1268=>"001101110",
  1269=>"010000111",
  1270=>"011001111",
  1271=>"110101000",
  1272=>"001011010",
  1273=>"000010010",
  1274=>"001110000",
  1275=>"101110100",
  1276=>"110110001",
  1277=>"011100011",
  1278=>"000111111",
  1279=>"101001011",
  1280=>"111100000",
  1281=>"010011100",
  1282=>"010111101",
  1283=>"000110000",
  1284=>"111010101",
  1285=>"010100111",
  1286=>"011100010",
  1287=>"110000110",
  1288=>"000111000",
  1289=>"010011110",
  1290=>"011011111",
  1291=>"011000000",
  1292=>"000010111",
  1293=>"110011001",
  1294=>"101100100",
  1295=>"010000011",
  1296=>"101110001",
  1297=>"010110100",
  1298=>"011001101",
  1299=>"110111011",
  1300=>"001001000",
  1301=>"010111010",
  1302=>"110000101",
  1303=>"001111110",
  1304=>"100010100",
  1305=>"110111110",
  1306=>"010101100",
  1307=>"101101011",
  1308=>"001001000",
  1309=>"000001100",
  1310=>"010000001",
  1311=>"001110101",
  1312=>"011011001",
  1313=>"011101010",
  1314=>"111001001",
  1315=>"011001111",
  1316=>"001011011",
  1317=>"110000010",
  1318=>"010100001",
  1319=>"100110010",
  1320=>"101101101",
  1321=>"100000101",
  1322=>"100000000",
  1323=>"110010100",
  1324=>"010111000",
  1325=>"110011100",
  1326=>"010011110",
  1327=>"110000000",
  1328=>"000000011",
  1329=>"000010101",
  1330=>"011001111",
  1331=>"001100100",
  1332=>"110100010",
  1333=>"000011111",
  1334=>"100010110",
  1335=>"001000111",
  1336=>"010000101",
  1337=>"101111011",
  1338=>"010111101",
  1339=>"011011111",
  1340=>"000110111",
  1341=>"100000111",
  1342=>"000011111",
  1343=>"101001001",
  1344=>"011011010",
  1345=>"000011010",
  1346=>"110100011",
  1347=>"001011010",
  1348=>"000001111",
  1349=>"000010100",
  1350=>"100010001",
  1351=>"100000011",
  1352=>"001110101",
  1353=>"100001111",
  1354=>"111110010",
  1355=>"101111010",
  1356=>"000000001",
  1357=>"101111011",
  1358=>"010100010",
  1359=>"101001101",
  1360=>"000100010",
  1361=>"101111000",
  1362=>"111101010",
  1363=>"110100110",
  1364=>"001010011",
  1365=>"100001110",
  1366=>"110110000",
  1367=>"100000000",
  1368=>"000000110",
  1369=>"001001110",
  1370=>"001111111",
  1371=>"010000110",
  1372=>"101000100",
  1373=>"101101001",
  1374=>"110010001",
  1375=>"111111011",
  1376=>"110010110",
  1377=>"110011100",
  1378=>"010100011",
  1379=>"111010010",
  1380=>"111101111",
  1381=>"010110010",
  1382=>"001001011",
  1383=>"010100110",
  1384=>"010011010",
  1385=>"010001001",
  1386=>"100010100",
  1387=>"101100100",
  1388=>"101000010",
  1389=>"111110011",
  1390=>"010101001",
  1391=>"011000011",
  1392=>"110111001",
  1393=>"110011011",
  1394=>"001111101",
  1395=>"100010010",
  1396=>"001110001",
  1397=>"011011010",
  1398=>"011100011",
  1399=>"111101000",
  1400=>"000010111",
  1401=>"010111101",
  1402=>"110010100",
  1403=>"001000101",
  1404=>"101110101",
  1405=>"110001100",
  1406=>"101000111",
  1407=>"000100010",
  1408=>"100010101",
  1409=>"011110100",
  1410=>"001000000",
  1411=>"101100010",
  1412=>"000110110",
  1413=>"100011011",
  1414=>"110111111",
  1415=>"110100101",
  1416=>"000001011",
  1417=>"000010101",
  1418=>"011110011",
  1419=>"011000111",
  1420=>"111001010",
  1421=>"001011000",
  1422=>"101000001",
  1423=>"001110011",
  1424=>"001101000",
  1425=>"011000000",
  1426=>"000101011",
  1427=>"011001111",
  1428=>"010110001",
  1429=>"000000101",
  1430=>"101001111",
  1431=>"100101111",
  1432=>"000111101",
  1433=>"000111001",
  1434=>"100011101",
  1435=>"001011101",
  1436=>"000001000",
  1437=>"111011100",
  1438=>"111100000",
  1439=>"011110010",
  1440=>"000101000",
  1441=>"111000010",
  1442=>"010101111",
  1443=>"110011000",
  1444=>"011111011",
  1445=>"001101001",
  1446=>"010010100",
  1447=>"101000101",
  1448=>"111011100",
  1449=>"000100011",
  1450=>"000000000",
  1451=>"001000000",
  1452=>"000011011",
  1453=>"011000001",
  1454=>"000111101",
  1455=>"101100010",
  1456=>"101110000",
  1457=>"111010010",
  1458=>"101101111",
  1459=>"011010010",
  1460=>"110011011",
  1461=>"111111011",
  1462=>"101110100",
  1463=>"011011110",
  1464=>"101011101",
  1465=>"111101001",
  1466=>"110101000",
  1467=>"010011010",
  1468=>"011111001",
  1469=>"011111001",
  1470=>"110110101",
  1471=>"010100110",
  1472=>"100100100",
  1473=>"001001010",
  1474=>"011001111",
  1475=>"001000110",
  1476=>"000110111",
  1477=>"000110110",
  1478=>"010001011",
  1479=>"000101100",
  1480=>"011000111",
  1481=>"011110100",
  1482=>"101000001",
  1483=>"000100110",
  1484=>"000001111",
  1485=>"011110001",
  1486=>"100110101",
  1487=>"010000001",
  1488=>"101001010",
  1489=>"010011000",
  1490=>"100100110",
  1491=>"010111011",
  1492=>"100101100",
  1493=>"010111011",
  1494=>"010110001",
  1495=>"111011000",
  1496=>"111001100",
  1497=>"110011101",
  1498=>"000011011",
  1499=>"010011001",
  1500=>"111100101",
  1501=>"111110101",
  1502=>"101100110",
  1503=>"111010001",
  1504=>"011001111",
  1505=>"011010111",
  1506=>"100110010",
  1507=>"100000100",
  1508=>"000000000",
  1509=>"101111001",
  1510=>"111001101",
  1511=>"110000111",
  1512=>"110000100",
  1513=>"101110011",
  1514=>"100000110",
  1515=>"000101001",
  1516=>"101110000",
  1517=>"001010011",
  1518=>"000111101",
  1519=>"100100111",
  1520=>"100000100",
  1521=>"011010111",
  1522=>"000011011",
  1523=>"101001100",
  1524=>"101010111",
  1525=>"100000001",
  1526=>"010100111",
  1527=>"000100000",
  1528=>"110010101",
  1529=>"010110010",
  1530=>"110101011",
  1531=>"100010101",
  1532=>"100101101",
  1533=>"010100110",
  1534=>"101011000",
  1535=>"111101100",
  1536=>"100100010",
  1537=>"000110001",
  1538=>"010001110",
  1539=>"111101110",
  1540=>"101011100",
  1541=>"110100100",
  1542=>"000111010",
  1543=>"000010001",
  1544=>"001000000",
  1545=>"010001110",
  1546=>"001001001",
  1547=>"011011111",
  1548=>"010011000",
  1549=>"110010000",
  1550=>"000100100",
  1551=>"111111101",
  1552=>"110101101",
  1553=>"111011010",
  1554=>"001110101",
  1555=>"011100110",
  1556=>"110000111",
  1557=>"110001110",
  1558=>"001101001",
  1559=>"101110001",
  1560=>"001011101",
  1561=>"011101110",
  1562=>"001101101",
  1563=>"111111010",
  1564=>"001000100",
  1565=>"110010111",
  1566=>"011101010",
  1567=>"000101001",
  1568=>"100011111",
  1569=>"010011011",
  1570=>"101000010",
  1571=>"100111101",
  1572=>"000000000",
  1573=>"011010010",
  1574=>"000000100",
  1575=>"101111110",
  1576=>"101010011",
  1577=>"011111001",
  1578=>"111010111",
  1579=>"101101000",
  1580=>"100111011",
  1581=>"111101100",
  1582=>"100100001",
  1583=>"010001001",
  1584=>"100000001",
  1585=>"100111110",
  1586=>"010010100",
  1587=>"101111100",
  1588=>"001101011",
  1589=>"010011101",
  1590=>"010000110",
  1591=>"110010111",
  1592=>"000100100",
  1593=>"100111101",
  1594=>"110111010",
  1595=>"110010100",
  1596=>"000000110",
  1597=>"100101001",
  1598=>"100011001",
  1599=>"000111100",
  1600=>"011000000",
  1601=>"000100000",
  1602=>"000111010",
  1603=>"100111111",
  1604=>"101000100",
  1605=>"001111101",
  1606=>"001000001",
  1607=>"111100111",
  1608=>"111001101",
  1609=>"011000001",
  1610=>"000111110",
  1611=>"111101001",
  1612=>"011101110",
  1613=>"110001110",
  1614=>"101111110",
  1615=>"010100100",
  1616=>"100111100",
  1617=>"011000001",
  1618=>"110110000",
  1619=>"101001011",
  1620=>"010010010",
  1621=>"011000000",
  1622=>"010110100",
  1623=>"100111101",
  1624=>"100011011",
  1625=>"101111101",
  1626=>"000101001",
  1627=>"001010001",
  1628=>"001110100",
  1629=>"001010101",
  1630=>"010010100",
  1631=>"110101101",
  1632=>"110011011",
  1633=>"001110010",
  1634=>"001000011",
  1635=>"001100100",
  1636=>"101010011",
  1637=>"110011101",
  1638=>"011110000",
  1639=>"111010010",
  1640=>"000100000",
  1641=>"100110100",
  1642=>"100001001",
  1643=>"100110000",
  1644=>"011100000",
  1645=>"000001100",
  1646=>"011000101",
  1647=>"110010001",
  1648=>"000110001",
  1649=>"010010010",
  1650=>"011010111",
  1651=>"101000101",
  1652=>"101001010",
  1653=>"000111000",
  1654=>"000000111",
  1655=>"011000100",
  1656=>"110111011",
  1657=>"111100000",
  1658=>"000001101",
  1659=>"100001010",
  1660=>"000110100",
  1661=>"100010111",
  1662=>"111110010",
  1663=>"100100101",
  1664=>"110111110",
  1665=>"001110111",
  1666=>"101000010",
  1667=>"000100111",
  1668=>"011001011",
  1669=>"111110010",
  1670=>"000111011",
  1671=>"111101001",
  1672=>"011000101",
  1673=>"101001001",
  1674=>"011110100",
  1675=>"011100001",
  1676=>"101100001",
  1677=>"000101000",
  1678=>"011101001",
  1679=>"111111101",
  1680=>"110011010",
  1681=>"000010001",
  1682=>"111100111",
  1683=>"100001001",
  1684=>"000001110",
  1685=>"010101010",
  1686=>"111000010",
  1687=>"001001110",
  1688=>"001110001",
  1689=>"010010001",
  1690=>"111101100",
  1691=>"111100011",
  1692=>"100100001",
  1693=>"110101000",
  1694=>"011111001",
  1695=>"111011111",
  1696=>"010010000",
  1697=>"000100011",
  1698=>"100111101",
  1699=>"011101110",
  1700=>"100001000",
  1701=>"111010000",
  1702=>"110000111",
  1703=>"000100100",
  1704=>"011010011",
  1705=>"111101100",
  1706=>"011000001",
  1707=>"000010101",
  1708=>"100001010",
  1709=>"010010010",
  1710=>"001010111",
  1711=>"110011111",
  1712=>"000000111",
  1713=>"100011101",
  1714=>"011011011",
  1715=>"101110001",
  1716=>"010110000",
  1717=>"000001101",
  1718=>"100001010",
  1719=>"000000010",
  1720=>"100101001",
  1721=>"100010101",
  1722=>"001111001",
  1723=>"101001100",
  1724=>"001000010",
  1725=>"111011111",
  1726=>"101000001",
  1727=>"000111110",
  1728=>"010111011",
  1729=>"010010000",
  1730=>"011001110",
  1731=>"100110111",
  1732=>"010000110",
  1733=>"000000010",
  1734=>"100000010",
  1735=>"011011111",
  1736=>"000101011",
  1737=>"000111101",
  1738=>"111001111",
  1739=>"000001100",
  1740=>"010000010",
  1741=>"010010011",
  1742=>"010100110",
  1743=>"111111001",
  1744=>"011110001",
  1745=>"100001010",
  1746=>"111000100",
  1747=>"000011111",
  1748=>"101111110",
  1749=>"101100100",
  1750=>"101110011",
  1751=>"111001001",
  1752=>"101101111",
  1753=>"100000101",
  1754=>"101110101",
  1755=>"110001001",
  1756=>"010011001",
  1757=>"001111111",
  1758=>"110101100",
  1759=>"000100000",
  1760=>"100010011",
  1761=>"100101110",
  1762=>"111101001",
  1763=>"101010100",
  1764=>"001100010",
  1765=>"010000101",
  1766=>"000100100",
  1767=>"010010000",
  1768=>"010110101",
  1769=>"011110101",
  1770=>"001101011",
  1771=>"110000111",
  1772=>"111011001",
  1773=>"100110111",
  1774=>"010011011",
  1775=>"111001011",
  1776=>"110100000",
  1777=>"011101100",
  1778=>"101010000",
  1779=>"001110101",
  1780=>"001001011",
  1781=>"010011101",
  1782=>"111011011",
  1783=>"000010100",
  1784=>"010001000",
  1785=>"011110010",
  1786=>"011100000",
  1787=>"100111010",
  1788=>"101010011",
  1789=>"010100100",
  1790=>"001011110",
  1791=>"011010001",
  1792=>"000110010",
  1793=>"000001001",
  1794=>"100110101",
  1795=>"100110110",
  1796=>"101010000",
  1797=>"000111011",
  1798=>"000001011",
  1799=>"010011010",
  1800=>"000000001",
  1801=>"010111111",
  1802=>"000110000",
  1803=>"101100111",
  1804=>"010010110",
  1805=>"001010110",
  1806=>"100110101",
  1807=>"001110111",
  1808=>"000001001",
  1809=>"100101110",
  1810=>"111010011",
  1811=>"010000001",
  1812=>"010100010",
  1813=>"110101111",
  1814=>"001110010",
  1815=>"101001011",
  1816=>"001000111",
  1817=>"000010011",
  1818=>"111011011",
  1819=>"001111101",
  1820=>"110101100",
  1821=>"101101100",
  1822=>"110111000",
  1823=>"010000101",
  1824=>"101100110",
  1825=>"111110001",
  1826=>"101111000",
  1827=>"101011011",
  1828=>"001110000",
  1829=>"000010001",
  1830=>"100000100",
  1831=>"111111011",
  1832=>"011100000",
  1833=>"101111101",
  1834=>"010100000",
  1835=>"000111111",
  1836=>"110010010",
  1837=>"010000011",
  1838=>"101101111",
  1839=>"000001100",
  1840=>"000100100",
  1841=>"110000001",
  1842=>"100101110",
  1843=>"000110010",
  1844=>"111100011",
  1845=>"111011101",
  1846=>"111101101",
  1847=>"111100000",
  1848=>"000010101",
  1849=>"110111111",
  1850=>"110100000",
  1851=>"001101001",
  1852=>"001011000",
  1853=>"001111010",
  1854=>"110001101",
  1855=>"100110110",
  1856=>"000100110",
  1857=>"000110110",
  1858=>"111101110",
  1859=>"000000101",
  1860=>"011111100",
  1861=>"101110110",
  1862=>"101100101",
  1863=>"011100000",
  1864=>"111011000",
  1865=>"010110101",
  1866=>"100000000",
  1867=>"110000110",
  1868=>"110000011",
  1869=>"101100101",
  1870=>"111011010",
  1871=>"111111011",
  1872=>"111100110",
  1873=>"110001111",
  1874=>"101101110",
  1875=>"000000100",
  1876=>"110100111",
  1877=>"101011010",
  1878=>"111101100",
  1879=>"010011110",
  1880=>"000000110",
  1881=>"101111101",
  1882=>"101101110",
  1883=>"100111110",
  1884=>"111101111",
  1885=>"001011110",
  1886=>"101011010",
  1887=>"101100101",
  1888=>"110001000",
  1889=>"101011010",
  1890=>"001000000",
  1891=>"010110001",
  1892=>"111010101",
  1893=>"001101101",
  1894=>"111111000",
  1895=>"001101100",
  1896=>"110100101",
  1897=>"011010010",
  1898=>"010101011",
  1899=>"111101010",
  1900=>"000100001",
  1901=>"011011011",
  1902=>"000111110",
  1903=>"011000100",
  1904=>"111101100",
  1905=>"111011011",
  1906=>"101111111",
  1907=>"001101111",
  1908=>"000101000",
  1909=>"011000110",
  1910=>"010000100",
  1911=>"110010000",
  1912=>"011100100",
  1913=>"101001000",
  1914=>"101100110",
  1915=>"111111111",
  1916=>"101011010",
  1917=>"101011101",
  1918=>"101110011",
  1919=>"110010010",
  1920=>"010110010",
  1921=>"011000110",
  1922=>"111111100",
  1923=>"010011111",
  1924=>"111100100",
  1925=>"101001110",
  1926=>"111100111",
  1927=>"100010010",
  1928=>"011011010",
  1929=>"110000100",
  1930=>"001111001",
  1931=>"101100010",
  1932=>"001000011",
  1933=>"111111110",
  1934=>"101010010",
  1935=>"101111101",
  1936=>"111100001",
  1937=>"100010100",
  1938=>"101111000",
  1939=>"100100011",
  1940=>"011011011",
  1941=>"111111101",
  1942=>"001000110",
  1943=>"110010011",
  1944=>"001100101",
  1945=>"111101000",
  1946=>"011011100",
  1947=>"100011111",
  1948=>"001111011",
  1949=>"110101000",
  1950=>"111101001",
  1951=>"100110100",
  1952=>"001101101",
  1953=>"110001111",
  1954=>"111010101",
  1955=>"010100011",
  1956=>"110111100",
  1957=>"001101111",
  1958=>"000011110",
  1959=>"010110101",
  1960=>"100101101",
  1961=>"101000011",
  1962=>"011010010",
  1963=>"011011010",
  1964=>"001110100",
  1965=>"100101011",
  1966=>"011101000",
  1967=>"011000010",
  1968=>"011111100",
  1969=>"111111111",
  1970=>"010000010",
  1971=>"110001110",
  1972=>"010111111",
  1973=>"010000000",
  1974=>"111111011",
  1975=>"000000111",
  1976=>"000110110",
  1977=>"010010111",
  1978=>"011011100",
  1979=>"010101010",
  1980=>"011011100",
  1981=>"001011110",
  1982=>"111111011",
  1983=>"110000000",
  1984=>"100000111",
  1985=>"111010101",
  1986=>"000111001",
  1987=>"111011011",
  1988=>"110001100",
  1989=>"000101001",
  1990=>"010110111",
  1991=>"101011011",
  1992=>"010000001",
  1993=>"000110011",
  1994=>"001001000",
  1995=>"110101111",
  1996=>"011011011",
  1997=>"001010000",
  1998=>"110000110",
  1999=>"011111011",
  2000=>"001111110",
  2001=>"001110000",
  2002=>"000100000",
  2003=>"001110001",
  2004=>"100001001",
  2005=>"000000111",
  2006=>"101100101",
  2007=>"000100010",
  2008=>"011101100",
  2009=>"001111010",
  2010=>"010000001",
  2011=>"011110011",
  2012=>"010000011",
  2013=>"010000001",
  2014=>"100011111",
  2015=>"111001001",
  2016=>"000000110",
  2017=>"001111011",
  2018=>"100110010",
  2019=>"101000011",
  2020=>"111001011",
  2021=>"111111001",
  2022=>"000101011",
  2023=>"011001110",
  2024=>"101011010",
  2025=>"010100011",
  2026=>"111101101",
  2027=>"001110011",
  2028=>"100110000",
  2029=>"001101101",
  2030=>"010010101",
  2031=>"111101010",
  2032=>"001010011",
  2033=>"111110110",
  2034=>"011010110",
  2035=>"111000011",
  2036=>"011111111",
  2037=>"111111000",
  2038=>"001111101",
  2039=>"100100001",
  2040=>"110001001",
  2041=>"011101101",
  2042=>"111001100",
  2043=>"101000111",
  2044=>"110010101",
  2045=>"100000001",
  2046=>"001110000",
  2047=>"111011010",
  2048=>"001100010",
  2049=>"111111101",
  2050=>"111111010",
  2051=>"001010011",
  2052=>"000100010",
  2053=>"001110100",
  2054=>"110110100",
  2055=>"001100000",
  2056=>"111111111",
  2057=>"001000010",
  2058=>"010111000",
  2059=>"110101001",
  2060=>"010110100",
  2061=>"000010001",
  2062=>"110111011",
  2063=>"110010110",
  2064=>"110000010",
  2065=>"100010111",
  2066=>"010010000",
  2067=>"011010011",
  2068=>"100011101",
  2069=>"110000101",
  2070=>"011001011",
  2071=>"001011100",
  2072=>"100011101",
  2073=>"100001001",
  2074=>"000110010",
  2075=>"000011111",
  2076=>"100110110",
  2077=>"101101101",
  2078=>"000111010",
  2079=>"111101111",
  2080=>"100001100",
  2081=>"100011100",
  2082=>"100101110",
  2083=>"111000110",
  2084=>"111100111",
  2085=>"111100100",
  2086=>"010001010",
  2087=>"111001001",
  2088=>"011100111",
  2089=>"101001001",
  2090=>"010010110",
  2091=>"100100001",
  2092=>"010011110",
  2093=>"100000011",
  2094=>"011111010",
  2095=>"111000000",
  2096=>"100100001",
  2097=>"010100101",
  2098=>"000100000",
  2099=>"000100100",
  2100=>"101011111",
  2101=>"101110000",
  2102=>"111000010",
  2103=>"111111000",
  2104=>"110100100",
  2105=>"011100110",
  2106=>"000010000",
  2107=>"000110101",
  2108=>"100110111",
  2109=>"100100100",
  2110=>"001000011",
  2111=>"010111101",
  2112=>"110111000",
  2113=>"000100001",
  2114=>"101110111",
  2115=>"010010100",
  2116=>"111111111",
  2117=>"000000010",
  2118=>"000011011",
  2119=>"101100000",
  2120=>"000111111",
  2121=>"001010111",
  2122=>"101111110",
  2123=>"110110111",
  2124=>"001111010",
  2125=>"101110011",
  2126=>"101100000",
  2127=>"011011111",
  2128=>"100110100",
  2129=>"101100111",
  2130=>"100100001",
  2131=>"001010011",
  2132=>"111101111",
  2133=>"111011110",
  2134=>"001010010",
  2135=>"001011011",
  2136=>"000000111",
  2137=>"000111110",
  2138=>"110000110",
  2139=>"001100001",
  2140=>"000001100",
  2141=>"010110110",
  2142=>"011000110",
  2143=>"001100010",
  2144=>"010010001",
  2145=>"101101101",
  2146=>"101001000",
  2147=>"100011010",
  2148=>"101111000",
  2149=>"000110000",
  2150=>"101001001",
  2151=>"010111100",
  2152=>"010011000",
  2153=>"111110011",
  2154=>"001001100",
  2155=>"010010111",
  2156=>"001110101",
  2157=>"011110001",
  2158=>"000011000",
  2159=>"001011101",
  2160=>"000001011",
  2161=>"000001010",
  2162=>"101010001",
  2163=>"000111011",
  2164=>"011100011",
  2165=>"111011011",
  2166=>"000001100",
  2167=>"010010011",
  2168=>"011010001",
  2169=>"001011000",
  2170=>"000111110",
  2171=>"001001000",
  2172=>"000001000",
  2173=>"110111011",
  2174=>"011111000",
  2175=>"011001101",
  2176=>"001101000",
  2177=>"000111100",
  2178=>"010100010",
  2179=>"111100110",
  2180=>"001100100",
  2181=>"111100111",
  2182=>"100100110",
  2183=>"100010110",
  2184=>"000011101",
  2185=>"001110010",
  2186=>"000111100",
  2187=>"111000001",
  2188=>"000001101",
  2189=>"010100100",
  2190=>"110010110",
  2191=>"101101000",
  2192=>"111100111",
  2193=>"011001100",
  2194=>"000100010",
  2195=>"001011111",
  2196=>"001010001",
  2197=>"110101011",
  2198=>"000100110",
  2199=>"001000111",
  2200=>"110111111",
  2201=>"111111101",
  2202=>"000011111",
  2203=>"000001010",
  2204=>"110100010",
  2205=>"101101110",
  2206=>"010111101",
  2207=>"111100110",
  2208=>"100100011",
  2209=>"111110010",
  2210=>"100010111",
  2211=>"010001001",
  2212=>"111010110",
  2213=>"001011001",
  2214=>"101000101",
  2215=>"000000111",
  2216=>"110010110",
  2217=>"101110111",
  2218=>"111011101",
  2219=>"100011101",
  2220=>"010011000",
  2221=>"110101101",
  2222=>"011001111",
  2223=>"001100011",
  2224=>"000011001",
  2225=>"101010000",
  2226=>"111110010",
  2227=>"100000111",
  2228=>"000000010",
  2229=>"111110010",
  2230=>"010100111",
  2231=>"101011010",
  2232=>"101010001",
  2233=>"101111110",
  2234=>"000000100",
  2235=>"111111111",
  2236=>"101110100",
  2237=>"101111111",
  2238=>"010001011",
  2239=>"100000100",
  2240=>"011000111",
  2241=>"001011011",
  2242=>"001101010",
  2243=>"010111010",
  2244=>"101110011",
  2245=>"001010100",
  2246=>"110111100",
  2247=>"101110011",
  2248=>"111110001",
  2249=>"110001000",
  2250=>"111100111",
  2251=>"101111001",
  2252=>"111000011",
  2253=>"111000001",
  2254=>"011011101",
  2255=>"110000111",
  2256=>"000100101",
  2257=>"011111000",
  2258=>"010000011",
  2259=>"101000100",
  2260=>"011011111",
  2261=>"111111000",
  2262=>"001001000",
  2263=>"010000001",
  2264=>"001110010",
  2265=>"111100000",
  2266=>"000010100",
  2267=>"100110000",
  2268=>"110001101",
  2269=>"011001011",
  2270=>"101001010",
  2271=>"100011010",
  2272=>"011011101",
  2273=>"111000000",
  2274=>"110111010",
  2275=>"000100010",
  2276=>"000011000",
  2277=>"101101100",
  2278=>"110011110",
  2279=>"111100000",
  2280=>"011010100",
  2281=>"010011011",
  2282=>"100100100",
  2283=>"000010110",
  2284=>"111011000",
  2285=>"010100101",
  2286=>"100101010",
  2287=>"000101101",
  2288=>"010011100",
  2289=>"010000111",
  2290=>"110101001",
  2291=>"110101110",
  2292=>"001000000",
  2293=>"111001111",
  2294=>"111101111",
  2295=>"001011101",
  2296=>"001101000",
  2297=>"011000111",
  2298=>"101111011",
  2299=>"000010001",
  2300=>"010101101",
  2301=>"100011011",
  2302=>"111101100",
  2303=>"000101111",
  2304=>"001000011",
  2305=>"011110111",
  2306=>"001110010",
  2307=>"010101101",
  2308=>"101110010",
  2309=>"101000011",
  2310=>"000100100",
  2311=>"000001110",
  2312=>"100111101",
  2313=>"101101010",
  2314=>"110101100",
  2315=>"100011011",
  2316=>"100011011",
  2317=>"000110000",
  2318=>"101000000",
  2319=>"000001100",
  2320=>"010000101",
  2321=>"000000000",
  2322=>"111110000",
  2323=>"011100101",
  2324=>"001010110",
  2325=>"001110000",
  2326=>"111011111",
  2327=>"010011011",
  2328=>"001010100",
  2329=>"001110110",
  2330=>"000011100",
  2331=>"000001011",
  2332=>"010100001",
  2333=>"110010001",
  2334=>"101000011",
  2335=>"000110100",
  2336=>"100110011",
  2337=>"100110001",
  2338=>"000111010",
  2339=>"010110000",
  2340=>"010001110",
  2341=>"111101101",
  2342=>"001000110",
  2343=>"000000101",
  2344=>"011111011",
  2345=>"001110010",
  2346=>"100110001",
  2347=>"110010111",
  2348=>"111111110",
  2349=>"100001110",
  2350=>"000010000",
  2351=>"011010100",
  2352=>"110011001",
  2353=>"001110111",
  2354=>"011011110",
  2355=>"011010100",
  2356=>"111110001",
  2357=>"001000011",
  2358=>"001111011",
  2359=>"111110011",
  2360=>"110110011",
  2361=>"110110000",
  2362=>"010010101",
  2363=>"110100000",
  2364=>"000111101",
  2365=>"110100000",
  2366=>"000011110",
  2367=>"101001000",
  2368=>"111101001",
  2369=>"100000110",
  2370=>"101110010",
  2371=>"111010011",
  2372=>"101111100",
  2373=>"010010010",
  2374=>"011011101",
  2375=>"001111010",
  2376=>"111111110",
  2377=>"110100100",
  2378=>"100010000",
  2379=>"110000100",
  2380=>"010010110",
  2381=>"011000001",
  2382=>"100000001",
  2383=>"101001000",
  2384=>"010011100",
  2385=>"010111001",
  2386=>"010100100",
  2387=>"000110100",
  2388=>"101000111",
  2389=>"001100101",
  2390=>"010011000",
  2391=>"000100101",
  2392=>"111001000",
  2393=>"100111101",
  2394=>"010100011",
  2395=>"000001000",
  2396=>"100101100",
  2397=>"101011000",
  2398=>"110001011",
  2399=>"110110100",
  2400=>"000010100",
  2401=>"101000111",
  2402=>"001101000",
  2403=>"111001001",
  2404=>"110111001",
  2405=>"111101010",
  2406=>"110000111",
  2407=>"100100100",
  2408=>"110010000",
  2409=>"101001100",
  2410=>"001100100",
  2411=>"101111001",
  2412=>"001000000",
  2413=>"000001010",
  2414=>"010111110",
  2415=>"101000110",
  2416=>"001101110",
  2417=>"001011101",
  2418=>"000111111",
  2419=>"111011001",
  2420=>"010011001",
  2421=>"110000100",
  2422=>"001110000",
  2423=>"110111011",
  2424=>"000000111",
  2425=>"011011001",
  2426=>"110111110",
  2427=>"111110110",
  2428=>"001101111",
  2429=>"010001011",
  2430=>"111000101",
  2431=>"100001110",
  2432=>"100010010",
  2433=>"000101000",
  2434=>"011111100",
  2435=>"110111110",
  2436=>"010001011",
  2437=>"000100001",
  2438=>"010000011",
  2439=>"111111011",
  2440=>"011011001",
  2441=>"010000000",
  2442=>"011100000",
  2443=>"110001100",
  2444=>"011001011",
  2445=>"110100101",
  2446=>"000001000",
  2447=>"010100000",
  2448=>"011101010",
  2449=>"010100000",
  2450=>"001001111",
  2451=>"101000110",
  2452=>"010101111",
  2453=>"000100011",
  2454=>"100000001",
  2455=>"000110100",
  2456=>"110110001",
  2457=>"101001100",
  2458=>"000111000",
  2459=>"000000101",
  2460=>"110101011",
  2461=>"110111011",
  2462=>"111110001",
  2463=>"111011000",
  2464=>"100101101",
  2465=>"011100010",
  2466=>"001110111",
  2467=>"100110101",
  2468=>"101100010",
  2469=>"000100001",
  2470=>"011011111",
  2471=>"101011000",
  2472=>"110101110",
  2473=>"010000111",
  2474=>"100001011",
  2475=>"001000001",
  2476=>"000010001",
  2477=>"011010110",
  2478=>"000101001",
  2479=>"001100001",
  2480=>"110110001",
  2481=>"011000111",
  2482=>"111111001",
  2483=>"010011000",
  2484=>"111011101",
  2485=>"001100011",
  2486=>"111000100",
  2487=>"011100111",
  2488=>"100011010",
  2489=>"000010011",
  2490=>"001101000",
  2491=>"101011100",
  2492=>"010000110",
  2493=>"111101111",
  2494=>"001011000",
  2495=>"101011010",
  2496=>"101011101",
  2497=>"111010101",
  2498=>"110110101",
  2499=>"011001000",
  2500=>"101000000",
  2501=>"011011100",
  2502=>"100111010",
  2503=>"001110000",
  2504=>"000100000",
  2505=>"101101011",
  2506=>"000111010",
  2507=>"000110110",
  2508=>"100011000",
  2509=>"010110001",
  2510=>"111011000",
  2511=>"010000000",
  2512=>"101100100",
  2513=>"000001100",
  2514=>"111101000",
  2515=>"010100001",
  2516=>"111000100",
  2517=>"101010100",
  2518=>"010001010",
  2519=>"100100100",
  2520=>"000110010",
  2521=>"001110110",
  2522=>"110110001",
  2523=>"000100011",
  2524=>"001001010",
  2525=>"010101101",
  2526=>"001110100",
  2527=>"010110001",
  2528=>"010111010",
  2529=>"010111010",
  2530=>"111110000",
  2531=>"011100000",
  2532=>"100101011",
  2533=>"100011111",
  2534=>"011011010",
  2535=>"110110100",
  2536=>"100001001",
  2537=>"101000010",
  2538=>"101010010",
  2539=>"111001001",
  2540=>"101000100",
  2541=>"100000000",
  2542=>"101110010",
  2543=>"011011010",
  2544=>"010000101",
  2545=>"001000001",
  2546=>"111010001",
  2547=>"001000011",
  2548=>"110011000",
  2549=>"011100110",
  2550=>"110111111",
  2551=>"001101000",
  2552=>"111110111",
  2553=>"000010011",
  2554=>"101110000",
  2555=>"111010001",
  2556=>"101001101",
  2557=>"000001110",
  2558=>"101111111",
  2559=>"101001101",
  2560=>"101010101",
  2561=>"010000100",
  2562=>"110011101",
  2563=>"000100101",
  2564=>"101111101",
  2565=>"000010111",
  2566=>"000001001",
  2567=>"000100111",
  2568=>"000000011",
  2569=>"011100011",
  2570=>"100000010",
  2571=>"001000000",
  2572=>"110101001",
  2573=>"000010110",
  2574=>"000000101",
  2575=>"110111000",
  2576=>"110100111",
  2577=>"111000110",
  2578=>"100110111",
  2579=>"111100011",
  2580=>"000000110",
  2581=>"001011000",
  2582=>"100001000",
  2583=>"010111100",
  2584=>"101100100",
  2585=>"011101110",
  2586=>"111101001",
  2587=>"101011010",
  2588=>"000010100",
  2589=>"000111011",
  2590=>"111011011",
  2591=>"111101001",
  2592=>"110100000",
  2593=>"000100000",
  2594=>"010110010",
  2595=>"000011010",
  2596=>"111001011",
  2597=>"100110101",
  2598=>"110101001",
  2599=>"001001101",
  2600=>"011001010",
  2601=>"101100110",
  2602=>"100101000",
  2603=>"100111011",
  2604=>"000001010",
  2605=>"001101010",
  2606=>"000000110",
  2607=>"111000110",
  2608=>"110101110",
  2609=>"100100010",
  2610=>"100101000",
  2611=>"111110010",
  2612=>"110110001",
  2613=>"110110101",
  2614=>"101111011",
  2615=>"100010011",
  2616=>"100001100",
  2617=>"100111111",
  2618=>"110111110",
  2619=>"010100111",
  2620=>"110110100",
  2621=>"000110000",
  2622=>"111001011",
  2623=>"111111110",
  2624=>"101111111",
  2625=>"011010010",
  2626=>"101111100",
  2627=>"010001100",
  2628=>"011101000",
  2629=>"110101010",
  2630=>"000000111",
  2631=>"111101001",
  2632=>"010001101",
  2633=>"001000101",
  2634=>"011101111",
  2635=>"111001011",
  2636=>"101100000",
  2637=>"100001101",
  2638=>"000010000",
  2639=>"101000000",
  2640=>"011101110",
  2641=>"101011111",
  2642=>"111000011",
  2643=>"110101001",
  2644=>"010001000",
  2645=>"100100111",
  2646=>"111001011",
  2647=>"001101010",
  2648=>"011110100",
  2649=>"111101011",
  2650=>"101101100",
  2651=>"111111101",
  2652=>"110011100",
  2653=>"100100101",
  2654=>"010001001",
  2655=>"101010010",
  2656=>"011100101",
  2657=>"011011000",
  2658=>"101011100",
  2659=>"110000111",
  2660=>"010111001",
  2661=>"000010110",
  2662=>"111010110",
  2663=>"000001001",
  2664=>"001001010",
  2665=>"111101011",
  2666=>"000101101",
  2667=>"001010110",
  2668=>"100111100",
  2669=>"001111011",
  2670=>"000011010",
  2671=>"010111000",
  2672=>"110101001",
  2673=>"000010000",
  2674=>"000100011",
  2675=>"001111010",
  2676=>"100101100",
  2677=>"010010101",
  2678=>"101101111",
  2679=>"010110001",
  2680=>"110101001",
  2681=>"110111001",
  2682=>"111001000",
  2683=>"101111111",
  2684=>"100010101",
  2685=>"010001100",
  2686=>"000111010",
  2687=>"001011001",
  2688=>"010001001",
  2689=>"000111110",
  2690=>"010000010",
  2691=>"001001010",
  2692=>"111111000",
  2693=>"100000111",
  2694=>"101001100",
  2695=>"000101001",
  2696=>"010100001",
  2697=>"111100001",
  2698=>"000111100",
  2699=>"110011011",
  2700=>"110001110",
  2701=>"011010001",
  2702=>"000011101",
  2703=>"110100100",
  2704=>"001101110",
  2705=>"101001111",
  2706=>"111010101",
  2707=>"110000001",
  2708=>"110000001",
  2709=>"011101010",
  2710=>"110111111",
  2711=>"001101000",
  2712=>"111111001",
  2713=>"011010000",
  2714=>"001000010",
  2715=>"101010101",
  2716=>"011011101",
  2717=>"001011011",
  2718=>"111111110",
  2719=>"001000010",
  2720=>"100011100",
  2721=>"000001101",
  2722=>"000111000",
  2723=>"101110100",
  2724=>"010101110",
  2725=>"100111111",
  2726=>"011001011",
  2727=>"000111011",
  2728=>"000001001",
  2729=>"000100000",
  2730=>"010011100",
  2731=>"011101000",
  2732=>"110001110",
  2733=>"101001010",
  2734=>"101111101",
  2735=>"111101011",
  2736=>"010010011",
  2737=>"101011011",
  2738=>"101110000",
  2739=>"000100110",
  2740=>"011010111",
  2741=>"101011101",
  2742=>"000011010",
  2743=>"011011011",
  2744=>"011101000",
  2745=>"100001011",
  2746=>"000000101",
  2747=>"111110011",
  2748=>"101010001",
  2749=>"001101011",
  2750=>"011000010",
  2751=>"001111111",
  2752=>"001110111",
  2753=>"011100000",
  2754=>"010001001",
  2755=>"011101001",
  2756=>"110100010",
  2757=>"010111101",
  2758=>"101111000",
  2759=>"010101010",
  2760=>"001101101",
  2761=>"001000000",
  2762=>"011101101",
  2763=>"001111000",
  2764=>"010100000",
  2765=>"011111100",
  2766=>"010101110",
  2767=>"000101110",
  2768=>"001100100",
  2769=>"001101101",
  2770=>"010110101",
  2771=>"100100011",
  2772=>"000111111",
  2773=>"111111100",
  2774=>"010111001",
  2775=>"001001100",
  2776=>"011100000",
  2777=>"011000110",
  2778=>"010001110",
  2779=>"100101110",
  2780=>"001101110",
  2781=>"000101010",
  2782=>"000001100",
  2783=>"010110011",
  2784=>"111100111",
  2785=>"100101001",
  2786=>"011101100",
  2787=>"100010010",
  2788=>"110111011",
  2789=>"010000000",
  2790=>"011000001",
  2791=>"001100000",
  2792=>"111000011",
  2793=>"000000001",
  2794=>"101111111",
  2795=>"010001100",
  2796=>"001100001",
  2797=>"001111010",
  2798=>"011110101",
  2799=>"111000101",
  2800=>"000100010",
  2801=>"101111011",
  2802=>"001101111",
  2803=>"010010110",
  2804=>"110000100",
  2805=>"100011110",
  2806=>"000011010",
  2807=>"110011010",
  2808=>"100110000",
  2809=>"010101010",
  2810=>"000001000",
  2811=>"011001001",
  2812=>"111111000",
  2813=>"110001110",
  2814=>"000001100",
  2815=>"110101100",
  2816=>"001101000",
  2817=>"111001100",
  2818=>"000100010",
  2819=>"110101011",
  2820=>"001011001",
  2821=>"010010100",
  2822=>"110110000",
  2823=>"101011011",
  2824=>"101100110",
  2825=>"001110001",
  2826=>"010001010",
  2827=>"010010000",
  2828=>"000100101",
  2829=>"000000000",
  2830=>"110101101",
  2831=>"001111000",
  2832=>"110011111",
  2833=>"000010001",
  2834=>"000101110",
  2835=>"110001010",
  2836=>"100111110",
  2837=>"011100100",
  2838=>"010111110",
  2839=>"000000001",
  2840=>"110010110",
  2841=>"111001111",
  2842=>"110001001",
  2843=>"010011111",
  2844=>"011111101",
  2845=>"111011010",
  2846=>"001001011",
  2847=>"000011110",
  2848=>"100100101",
  2849=>"010111001",
  2850=>"111011011",
  2851=>"000001111",
  2852=>"100111101",
  2853=>"111110011",
  2854=>"110010100",
  2855=>"110111111",
  2856=>"101101010",
  2857=>"000110001",
  2858=>"001101111",
  2859=>"010110100",
  2860=>"000101110",
  2861=>"111010010",
  2862=>"000111111",
  2863=>"001110100",
  2864=>"001100111",
  2865=>"100100100",
  2866=>"111000100",
  2867=>"100010100",
  2868=>"100010001",
  2869=>"001111101",
  2870=>"110011100",
  2871=>"101111111",
  2872=>"100110000",
  2873=>"001110001",
  2874=>"110001010",
  2875=>"011101000",
  2876=>"101101001",
  2877=>"001001000",
  2878=>"000111000",
  2879=>"100111111",
  2880=>"010000011",
  2881=>"111111001",
  2882=>"110001101",
  2883=>"010000011",
  2884=>"110001001",
  2885=>"100001100",
  2886=>"110110011",
  2887=>"000011011",
  2888=>"101110100",
  2889=>"011000100",
  2890=>"100110111",
  2891=>"011011001",
  2892=>"111100011",
  2893=>"101101110",
  2894=>"110110111",
  2895=>"110001100",
  2896=>"000011110",
  2897=>"101010110",
  2898=>"100010101",
  2899=>"001000000",
  2900=>"111111001",
  2901=>"010101011",
  2902=>"001011000",
  2903=>"011000010",
  2904=>"110100010",
  2905=>"010110110",
  2906=>"111001111",
  2907=>"100001001",
  2908=>"011110111",
  2909=>"010000110",
  2910=>"101100011",
  2911=>"110101011",
  2912=>"111001100",
  2913=>"100010101",
  2914=>"010010000",
  2915=>"010010010",
  2916=>"011011010",
  2917=>"110111001",
  2918=>"000111110",
  2919=>"110011100",
  2920=>"000110000",
  2921=>"100111110",
  2922=>"011101111",
  2923=>"101101000",
  2924=>"110001110",
  2925=>"000011101",
  2926=>"001000110",
  2927=>"000110111",
  2928=>"001100101",
  2929=>"100000001",
  2930=>"001101110",
  2931=>"011001110",
  2932=>"110001101",
  2933=>"000110000",
  2934=>"100101101",
  2935=>"101100001",
  2936=>"000101110",
  2937=>"101011110",
  2938=>"111100000",
  2939=>"110001011",
  2940=>"001001101",
  2941=>"100011001",
  2942=>"011001101",
  2943=>"111011110",
  2944=>"000111101",
  2945=>"101001010",
  2946=>"100110001",
  2947=>"010000101",
  2948=>"001110100",
  2949=>"000101101",
  2950=>"011111110",
  2951=>"110001001",
  2952=>"001110001",
  2953=>"101010000",
  2954=>"111101011",
  2955=>"010100001",
  2956=>"000000001",
  2957=>"010001000",
  2958=>"111111111",
  2959=>"111110110",
  2960=>"111100001",
  2961=>"110010110",
  2962=>"000000100",
  2963=>"110011110",
  2964=>"011011111",
  2965=>"101110011",
  2966=>"111011010",
  2967=>"010001000",
  2968=>"111110001",
  2969=>"011001111",
  2970=>"101011011",
  2971=>"110110101",
  2972=>"110011010",
  2973=>"011000101",
  2974=>"011001001",
  2975=>"000111000",
  2976=>"100000111",
  2977=>"000010110",
  2978=>"010001001",
  2979=>"100000100",
  2980=>"000010110",
  2981=>"000100100",
  2982=>"001101111",
  2983=>"110010011",
  2984=>"001010110",
  2985=>"100001110",
  2986=>"111110100",
  2987=>"101000010",
  2988=>"000000100",
  2989=>"111111000",
  2990=>"000111101",
  2991=>"011111110",
  2992=>"110000111",
  2993=>"000111000",
  2994=>"111100101",
  2995=>"010000010",
  2996=>"110000111",
  2997=>"000000000",
  2998=>"011110001",
  2999=>"011001111",
  3000=>"111110100",
  3001=>"100000101",
  3002=>"100101111",
  3003=>"000000010",
  3004=>"001110010",
  3005=>"000001000",
  3006=>"111100001",
  3007=>"110111110",
  3008=>"111111010",
  3009=>"110100100",
  3010=>"010101001",
  3011=>"100011100",
  3012=>"001101001",
  3013=>"000010100",
  3014=>"101001001",
  3015=>"100111111",
  3016=>"110000111",
  3017=>"100010111",
  3018=>"100110011",
  3019=>"110111011",
  3020=>"001001101",
  3021=>"000101011",
  3022=>"000000110",
  3023=>"110101011",
  3024=>"111111011",
  3025=>"111001100",
  3026=>"100010001",
  3027=>"001101011",
  3028=>"000000110",
  3029=>"111110111",
  3030=>"101000000",
  3031=>"000011100",
  3032=>"111000101",
  3033=>"101101000",
  3034=>"110011110",
  3035=>"011000000",
  3036=>"111111010",
  3037=>"000110000",
  3038=>"111111101",
  3039=>"111101111",
  3040=>"000000100",
  3041=>"100110110",
  3042=>"110010000",
  3043=>"100111111",
  3044=>"000000000",
  3045=>"110100111",
  3046=>"010101000",
  3047=>"110100111",
  3048=>"010011111",
  3049=>"100101100",
  3050=>"000100011",
  3051=>"000100110",
  3052=>"101001110",
  3053=>"111100010",
  3054=>"101000100",
  3055=>"000010100",
  3056=>"010101011",
  3057=>"101111011",
  3058=>"001110111",
  3059=>"010100010",
  3060=>"100110100",
  3061=>"100011111",
  3062=>"100110100",
  3063=>"110111101",
  3064=>"111000001",
  3065=>"100001111",
  3066=>"000101010",
  3067=>"101001100",
  3068=>"101001111",
  3069=>"110110111",
  3070=>"110101100",
  3071=>"010000011",
  3072=>"011000100",
  3073=>"111101001",
  3074=>"010000001",
  3075=>"111100001",
  3076=>"110101110",
  3077=>"010010101",
  3078=>"101111010",
  3079=>"011100000",
  3080=>"001011101",
  3081=>"101000100",
  3082=>"001011111",
  3083=>"100100110",
  3084=>"110010011",
  3085=>"111101000",
  3086=>"100101110",
  3087=>"111101011",
  3088=>"001100000",
  3089=>"001010111",
  3090=>"110111110",
  3091=>"001111100",
  3092=>"111011011",
  3093=>"000000101",
  3094=>"010011011",
  3095=>"101001010",
  3096=>"010001010",
  3097=>"000011111",
  3098=>"000000010",
  3099=>"110000100",
  3100=>"110100000",
  3101=>"100011101",
  3102=>"100100110",
  3103=>"000111100",
  3104=>"010100100",
  3105=>"100001111",
  3106=>"011001111",
  3107=>"111100000",
  3108=>"011100110",
  3109=>"111110010",
  3110=>"110000010",
  3111=>"111001001",
  3112=>"010110001",
  3113=>"101010111",
  3114=>"010100101",
  3115=>"011101011",
  3116=>"011011100",
  3117=>"011100101",
  3118=>"110100101",
  3119=>"110101001",
  3120=>"001001000",
  3121=>"110110111",
  3122=>"111010000",
  3123=>"000111000",
  3124=>"001000100",
  3125=>"010111010",
  3126=>"100001100",
  3127=>"010110110",
  3128=>"000110110",
  3129=>"001010101",
  3130=>"010000100",
  3131=>"011010100",
  3132=>"001011000",
  3133=>"011111101",
  3134=>"111101000",
  3135=>"101100001",
  3136=>"001010110",
  3137=>"011001011",
  3138=>"100000011",
  3139=>"010010011",
  3140=>"101000110",
  3141=>"011110111",
  3142=>"011000011",
  3143=>"111111011",
  3144=>"001111010",
  3145=>"101111010",
  3146=>"001101010",
  3147=>"111100011",
  3148=>"100101100",
  3149=>"100100100",
  3150=>"110000001",
  3151=>"110111101",
  3152=>"001110011",
  3153=>"011111001",
  3154=>"110011111",
  3155=>"000000111",
  3156=>"010000101",
  3157=>"110100110",
  3158=>"001100000",
  3159=>"111110111",
  3160=>"101110000",
  3161=>"110000111",
  3162=>"011101011",
  3163=>"000001001",
  3164=>"010011011",
  3165=>"110000111",
  3166=>"010100010",
  3167=>"010001011",
  3168=>"001111111",
  3169=>"111010111",
  3170=>"000010011",
  3171=>"111010000",
  3172=>"010000100",
  3173=>"011110001",
  3174=>"011011111",
  3175=>"000110101",
  3176=>"000000000",
  3177=>"101100010",
  3178=>"010111000",
  3179=>"001100111",
  3180=>"001001000",
  3181=>"011010000",
  3182=>"001011100",
  3183=>"010111111",
  3184=>"010000000",
  3185=>"000011101",
  3186=>"110001000",
  3187=>"111101100",
  3188=>"100111110",
  3189=>"010100010",
  3190=>"111010010",
  3191=>"101100111",
  3192=>"010001000",
  3193=>"001111101",
  3194=>"110011111",
  3195=>"101011001",
  3196=>"000110110",
  3197=>"100011000",
  3198=>"000100111",
  3199=>"001000000",
  3200=>"001111001",
  3201=>"110111010",
  3202=>"010010100",
  3203=>"000010000",
  3204=>"000100001",
  3205=>"101000000",
  3206=>"000111000",
  3207=>"000011100",
  3208=>"110111111",
  3209=>"110000111",
  3210=>"001010100",
  3211=>"111111010",
  3212=>"001001011",
  3213=>"101000111",
  3214=>"000010111",
  3215=>"010001111",
  3216=>"100110110",
  3217=>"000001000",
  3218=>"110110111",
  3219=>"000000111",
  3220=>"001011101",
  3221=>"010100110",
  3222=>"100111110",
  3223=>"001101110",
  3224=>"000000100",
  3225=>"111110101",
  3226=>"101001001",
  3227=>"001000011",
  3228=>"001001111",
  3229=>"000011000",
  3230=>"011011011",
  3231=>"110011111",
  3232=>"010111001",
  3233=>"111101101",
  3234=>"110001000",
  3235=>"111001111",
  3236=>"001001001",
  3237=>"010101101",
  3238=>"111011011",
  3239=>"101110010",
  3240=>"001001001",
  3241=>"010010000",
  3242=>"111111100",
  3243=>"100010101",
  3244=>"001011010",
  3245=>"010100001",
  3246=>"010110100",
  3247=>"101001100",
  3248=>"010101000",
  3249=>"010110100",
  3250=>"010100011",
  3251=>"110001010",
  3252=>"001011111",
  3253=>"001010001",
  3254=>"111010111",
  3255=>"100101010",
  3256=>"000101100",
  3257=>"010110111",
  3258=>"100001100",
  3259=>"011010010",
  3260=>"101011100",
  3261=>"001001111",
  3262=>"100011111",
  3263=>"111010111",
  3264=>"100110110",
  3265=>"001000011",
  3266=>"001100110",
  3267=>"101110110",
  3268=>"101110010",
  3269=>"101101000",
  3270=>"100101101",
  3271=>"010101000",
  3272=>"011101111",
  3273=>"101110010",
  3274=>"010110000",
  3275=>"101010111",
  3276=>"111101111",
  3277=>"100001100",
  3278=>"001100101",
  3279=>"000000000",
  3280=>"010111011",
  3281=>"111001001",
  3282=>"111101111",
  3283=>"011011111",
  3284=>"111110001",
  3285=>"001000111",
  3286=>"101001010",
  3287=>"111110000",
  3288=>"000011101",
  3289=>"000100111",
  3290=>"011110111",
  3291=>"000011011",
  3292=>"011010000",
  3293=>"100001011",
  3294=>"000111110",
  3295=>"110001110",
  3296=>"001111000",
  3297=>"011101010",
  3298=>"110001000",
  3299=>"011001011",
  3300=>"001000000",
  3301=>"110101111",
  3302=>"010000111",
  3303=>"101101011",
  3304=>"000100011",
  3305=>"110100100",
  3306=>"110000110",
  3307=>"000010111",
  3308=>"100100000",
  3309=>"001101011",
  3310=>"011000000",
  3311=>"111110001",
  3312=>"111000101",
  3313=>"001011111",
  3314=>"001001110",
  3315=>"011100001",
  3316=>"000010100",
  3317=>"101110011",
  3318=>"100011110",
  3319=>"001000111",
  3320=>"011011011",
  3321=>"001110011",
  3322=>"110000011",
  3323=>"001110010",
  3324=>"010100001",
  3325=>"001001010",
  3326=>"011010011",
  3327=>"100010010",
  3328=>"011001001",
  3329=>"010000001",
  3330=>"001111001",
  3331=>"100010101",
  3332=>"000011110",
  3333=>"110100101",
  3334=>"111010010",
  3335=>"100011001",
  3336=>"000010111",
  3337=>"100110100",
  3338=>"010011111",
  3339=>"100000110",
  3340=>"111010110",
  3341=>"000001010",
  3342=>"100111100",
  3343=>"100111111",
  3344=>"110100011",
  3345=>"110011000",
  3346=>"011011001",
  3347=>"111110101",
  3348=>"010110001",
  3349=>"110010001",
  3350=>"010010101",
  3351=>"110010011",
  3352=>"110101100",
  3353=>"011111110",
  3354=>"010100000",
  3355=>"100011000",
  3356=>"000110100",
  3357=>"100000101",
  3358=>"000011000",
  3359=>"011010111",
  3360=>"000100101",
  3361=>"101010111",
  3362=>"100001001",
  3363=>"000000010",
  3364=>"110000110",
  3365=>"010000001",
  3366=>"000010011",
  3367=>"100010110",
  3368=>"010011100",
  3369=>"100011010",
  3370=>"010010011",
  3371=>"100010000",
  3372=>"000011110",
  3373=>"101111110",
  3374=>"000100101",
  3375=>"011011111",
  3376=>"100111000",
  3377=>"001100101",
  3378=>"101000100",
  3379=>"100001111",
  3380=>"001000011",
  3381=>"111111111",
  3382=>"010101011",
  3383=>"101000000",
  3384=>"010111111",
  3385=>"010001000",
  3386=>"001000011",
  3387=>"010111001",
  3388=>"110000001",
  3389=>"011000000",
  3390=>"110000000",
  3391=>"100100100",
  3392=>"111001001",
  3393=>"010100011",
  3394=>"011011000",
  3395=>"101000000",
  3396=>"101011010",
  3397=>"101111011",
  3398=>"010010101",
  3399=>"000011001",
  3400=>"101101110",
  3401=>"000000011",
  3402=>"011110111",
  3403=>"010011111",
  3404=>"111111010",
  3405=>"011010100",
  3406=>"100110000",
  3407=>"011000101",
  3408=>"001100001",
  3409=>"100100101",
  3410=>"110101010",
  3411=>"100000011",
  3412=>"010000011",
  3413=>"001001111",
  3414=>"001110000",
  3415=>"011001111",
  3416=>"000110101",
  3417=>"011001011",
  3418=>"110101011",
  3419=>"100000000",
  3420=>"000111000",
  3421=>"010000010",
  3422=>"010110001",
  3423=>"101000100",
  3424=>"110111100",
  3425=>"100000111",
  3426=>"111110011",
  3427=>"001111111",
  3428=>"100111000",
  3429=>"001100110",
  3430=>"100111001",
  3431=>"110100100",
  3432=>"100101101",
  3433=>"001010100",
  3434=>"000010000",
  3435=>"000011011",
  3436=>"001001100",
  3437=>"010011100",
  3438=>"111010000",
  3439=>"111111111",
  3440=>"010011111",
  3441=>"011011011",
  3442=>"101101010",
  3443=>"100111001",
  3444=>"101010000",
  3445=>"100011011",
  3446=>"001001001",
  3447=>"010110110",
  3448=>"011011000",
  3449=>"010111001",
  3450=>"110110011",
  3451=>"001010010",
  3452=>"001100100",
  3453=>"000111110",
  3454=>"001110010",
  3455=>"110010000",
  3456=>"111000011",
  3457=>"011110100",
  3458=>"011010000",
  3459=>"101001111",
  3460=>"101111010",
  3461=>"100001110",
  3462=>"010110111",
  3463=>"001000101",
  3464=>"011100000",
  3465=>"001011000",
  3466=>"111011101",
  3467=>"010001001",
  3468=>"010011011",
  3469=>"100110000",
  3470=>"101000111",
  3471=>"110000010",
  3472=>"000010001",
  3473=>"001001111",
  3474=>"111001011",
  3475=>"111010101",
  3476=>"000001001",
  3477=>"011001011",
  3478=>"100101111",
  3479=>"101100000",
  3480=>"110001000",
  3481=>"011010010",
  3482=>"001111111",
  3483=>"101011001",
  3484=>"000001111",
  3485=>"111111111",
  3486=>"111011000",
  3487=>"110010001",
  3488=>"010100010",
  3489=>"010001010",
  3490=>"011000000",
  3491=>"000010110",
  3492=>"101100011",
  3493=>"100110000",
  3494=>"100000000",
  3495=>"011110010",
  3496=>"010001010",
  3497=>"110010100",
  3498=>"100110111",
  3499=>"111010100",
  3500=>"111001110",
  3501=>"000001001",
  3502=>"010010010",
  3503=>"010010001",
  3504=>"100111011",
  3505=>"000010000",
  3506=>"101111000",
  3507=>"111100001",
  3508=>"010011100",
  3509=>"010101000",
  3510=>"100011111",
  3511=>"000011101",
  3512=>"000110000",
  3513=>"000011100",
  3514=>"000000010",
  3515=>"011010000",
  3516=>"010010010",
  3517=>"100001100",
  3518=>"010001101",
  3519=>"100101010",
  3520=>"001100111",
  3521=>"000001000",
  3522=>"000111011",
  3523=>"100101110",
  3524=>"010111111",
  3525=>"101100001",
  3526=>"111101010",
  3527=>"110001010",
  3528=>"011110110",
  3529=>"111111111",
  3530=>"010010000",
  3531=>"010110010",
  3532=>"111111111",
  3533=>"110101010",
  3534=>"100001101",
  3535=>"010110000",
  3536=>"011111101",
  3537=>"010110010",
  3538=>"010100001",
  3539=>"000100000",
  3540=>"001110000",
  3541=>"110111011",
  3542=>"011001100",
  3543=>"010010011",
  3544=>"100101011",
  3545=>"100100010",
  3546=>"101001011",
  3547=>"110001101",
  3548=>"110001110",
  3549=>"111010011",
  3550=>"100011000",
  3551=>"110110010",
  3552=>"110100001",
  3553=>"111010011",
  3554=>"001001110",
  3555=>"110001000",
  3556=>"011001011",
  3557=>"011100111",
  3558=>"000000101",
  3559=>"100111000",
  3560=>"001101101",
  3561=>"011100011",
  3562=>"011000010",
  3563=>"010100000",
  3564=>"111111011",
  3565=>"011110000",
  3566=>"100100100",
  3567=>"100000000",
  3568=>"001000100",
  3569=>"010101111",
  3570=>"100100010",
  3571=>"001001110",
  3572=>"011000000",
  3573=>"101110011",
  3574=>"011100000",
  3575=>"000101111",
  3576=>"100101111",
  3577=>"010100010",
  3578=>"101110101",
  3579=>"111111000",
  3580=>"110011111",
  3581=>"011100001",
  3582=>"001110000",
  3583=>"010011010",
  3584=>"001010100",
  3585=>"011101101",
  3586=>"001010110",
  3587=>"001000111",
  3588=>"110000100",
  3589=>"000011111",
  3590=>"110000111",
  3591=>"010001010",
  3592=>"001101101",
  3593=>"000100010",
  3594=>"110111111",
  3595=>"101000000",
  3596=>"110000001",
  3597=>"001110001",
  3598=>"001000111",
  3599=>"011001100",
  3600=>"010101101",
  3601=>"101110000",
  3602=>"110000100",
  3603=>"101101100",
  3604=>"010000010",
  3605=>"001101001",
  3606=>"000110001",
  3607=>"011000111",
  3608=>"101000100",
  3609=>"000011111",
  3610=>"010100110",
  3611=>"010110111",
  3612=>"111000111",
  3613=>"010011101",
  3614=>"100100100",
  3615=>"011011001",
  3616=>"011010000",
  3617=>"001001000",
  3618=>"110100101",
  3619=>"001000000",
  3620=>"111111101",
  3621=>"000000110",
  3622=>"100111001",
  3623=>"000110111",
  3624=>"101110010",
  3625=>"011001110",
  3626=>"001011111",
  3627=>"000110011",
  3628=>"011010010",
  3629=>"100001100",
  3630=>"001101010",
  3631=>"111110001",
  3632=>"101010101",
  3633=>"111101000",
  3634=>"001001010",
  3635=>"101111101",
  3636=>"110000001",
  3637=>"011010000",
  3638=>"011101101",
  3639=>"111111110",
  3640=>"100000011",
  3641=>"011001011",
  3642=>"110110001",
  3643=>"110000111",
  3644=>"010010000",
  3645=>"100110100",
  3646=>"111100011",
  3647=>"101110010",
  3648=>"111011111",
  3649=>"100001110",
  3650=>"010110001",
  3651=>"111001000",
  3652=>"011101101",
  3653=>"111111110",
  3654=>"001010101",
  3655=>"011110011",
  3656=>"011000100",
  3657=>"001001001",
  3658=>"010101101",
  3659=>"111011111",
  3660=>"000011001",
  3661=>"001011010",
  3662=>"010101111",
  3663=>"101000111",
  3664=>"010001101",
  3665=>"100011111",
  3666=>"000011000",
  3667=>"000001100",
  3668=>"010100000",
  3669=>"101011111",
  3670=>"101001010",
  3671=>"000010111",
  3672=>"100010110",
  3673=>"010011110",
  3674=>"110110101",
  3675=>"101100010",
  3676=>"000000100",
  3677=>"010100101",
  3678=>"010101100",
  3679=>"011011100",
  3680=>"010110100",
  3681=>"101100111",
  3682=>"110101000",
  3683=>"000000111",
  3684=>"111111010",
  3685=>"100001000",
  3686=>"011100011",
  3687=>"100101111",
  3688=>"110000000",
  3689=>"111011001",
  3690=>"100001011",
  3691=>"000101110",
  3692=>"111110111",
  3693=>"100111111",
  3694=>"100011101",
  3695=>"000110010",
  3696=>"010000010",
  3697=>"011100001",
  3698=>"000010110",
  3699=>"100011010",
  3700=>"100101111",
  3701=>"000000111",
  3702=>"101000000",
  3703=>"011111111",
  3704=>"011010010",
  3705=>"010001111",
  3706=>"111100100",
  3707=>"010001101",
  3708=>"110011100",
  3709=>"010010011",
  3710=>"101001010",
  3711=>"011111101",
  3712=>"011001110",
  3713=>"111110111",
  3714=>"001001001",
  3715=>"010010100",
  3716=>"010111100",
  3717=>"000110101",
  3718=>"001010000",
  3719=>"100010010",
  3720=>"001001100",
  3721=>"000100111",
  3722=>"110100000",
  3723=>"101001010",
  3724=>"111010110",
  3725=>"111100011",
  3726=>"001000011",
  3727=>"101010010",
  3728=>"010111110",
  3729=>"010101111",
  3730=>"011110101",
  3731=>"001011010",
  3732=>"111100100",
  3733=>"001001100",
  3734=>"010111101",
  3735=>"010000000",
  3736=>"111001010",
  3737=>"000110101",
  3738=>"000011000",
  3739=>"110100000",
  3740=>"000110110",
  3741=>"111100100",
  3742=>"110111000",
  3743=>"000101110",
  3744=>"110111111",
  3745=>"001011110",
  3746=>"100111100",
  3747=>"000111100",
  3748=>"001001001",
  3749=>"111110101",
  3750=>"111000111",
  3751=>"111010000",
  3752=>"110000010",
  3753=>"011111111",
  3754=>"010101011",
  3755=>"000011000",
  3756=>"000111010",
  3757=>"110011110",
  3758=>"010101111",
  3759=>"111010000",
  3760=>"010001001",
  3761=>"000000111",
  3762=>"001000111",
  3763=>"010011101",
  3764=>"111010111",
  3765=>"110001000",
  3766=>"001000010",
  3767=>"110111000",
  3768=>"110111101",
  3769=>"100110110",
  3770=>"000000111",
  3771=>"100000111",
  3772=>"000000111",
  3773=>"011111101",
  3774=>"111010010",
  3775=>"011000000",
  3776=>"010001110",
  3777=>"100110000",
  3778=>"000000000",
  3779=>"111100000",
  3780=>"100011000",
  3781=>"101011001",
  3782=>"000111010",
  3783=>"111011111",
  3784=>"001010100",
  3785=>"110011001",
  3786=>"001011100",
  3787=>"000010100",
  3788=>"010001111",
  3789=>"100000000",
  3790=>"101110000",
  3791=>"111101011",
  3792=>"001101000",
  3793=>"010101000",
  3794=>"100110001",
  3795=>"010011111",
  3796=>"110101000",
  3797=>"100000010",
  3798=>"001111001",
  3799=>"100111010",
  3800=>"011111111",
  3801=>"101101101",
  3802=>"011010001",
  3803=>"000001111",
  3804=>"000010010",
  3805=>"010101000",
  3806=>"100110111",
  3807=>"110110101",
  3808=>"000001100",
  3809=>"000101011",
  3810=>"111011011",
  3811=>"000110101",
  3812=>"110101101",
  3813=>"101011000",
  3814=>"000111110",
  3815=>"010000111",
  3816=>"010011001",
  3817=>"111011011",
  3818=>"010010101",
  3819=>"010010001",
  3820=>"000011010",
  3821=>"011010000",
  3822=>"100000000",
  3823=>"111111100",
  3824=>"100011010",
  3825=>"100111011",
  3826=>"101101110",
  3827=>"000101010",
  3828=>"100000001",
  3829=>"101010000",
  3830=>"101010010",
  3831=>"010111111",
  3832=>"101110000",
  3833=>"110100100",
  3834=>"010111000",
  3835=>"000000000",
  3836=>"111010100",
  3837=>"000111101",
  3838=>"101011000",
  3839=>"001001100",
  3840=>"101010010",
  3841=>"001000101",
  3842=>"011000110",
  3843=>"010101000",
  3844=>"000101111",
  3845=>"100001010",
  3846=>"100011001",
  3847=>"010101000",
  3848=>"111110111",
  3849=>"101101101",
  3850=>"110011110",
  3851=>"110101001",
  3852=>"010010100",
  3853=>"111100110",
  3854=>"111100100",
  3855=>"001001010",
  3856=>"100000111",
  3857=>"001011000",
  3858=>"010101100",
  3859=>"111000000",
  3860=>"110100011",
  3861=>"010001011",
  3862=>"000001001",
  3863=>"000100100",
  3864=>"111111111",
  3865=>"101101011",
  3866=>"011010011",
  3867=>"111000101",
  3868=>"011011110",
  3869=>"111110010",
  3870=>"001001111",
  3871=>"110101001",
  3872=>"100111011",
  3873=>"100100101",
  3874=>"101000000",
  3875=>"111001111",
  3876=>"100001100",
  3877=>"000011111",
  3878=>"100111100",
  3879=>"101000111",
  3880=>"010101100",
  3881=>"001100101",
  3882=>"101010000",
  3883=>"010010001",
  3884=>"111100111",
  3885=>"110100001",
  3886=>"101111011",
  3887=>"001111111",
  3888=>"110110010",
  3889=>"001010111",
  3890=>"000110000",
  3891=>"000111011",
  3892=>"000110010",
  3893=>"001001000",
  3894=>"100010000",
  3895=>"000000011",
  3896=>"101110010",
  3897=>"001101011",
  3898=>"111111101",
  3899=>"010001000",
  3900=>"011100010",
  3901=>"001110111",
  3902=>"000000001",
  3903=>"100111111",
  3904=>"011111011",
  3905=>"001001110",
  3906=>"010000001",
  3907=>"100101111",
  3908=>"101101111",
  3909=>"011011101",
  3910=>"000101111",
  3911=>"101001001",
  3912=>"110100011",
  3913=>"100100100",
  3914=>"000110011",
  3915=>"001011100",
  3916=>"100100100",
  3917=>"110110100",
  3918=>"100000111",
  3919=>"101000011",
  3920=>"011011011",
  3921=>"100001111",
  3922=>"010010100",
  3923=>"000100110",
  3924=>"010000000",
  3925=>"010110110",
  3926=>"110001101",
  3927=>"000000111",
  3928=>"011010111",
  3929=>"101100101",
  3930=>"011000111",
  3931=>"101100000",
  3932=>"100101000",
  3933=>"011111111",
  3934=>"101001100",
  3935=>"000100010",
  3936=>"110111100",
  3937=>"010001111",
  3938=>"100100110",
  3939=>"111101100",
  3940=>"011000010",
  3941=>"101001100",
  3942=>"010001000",
  3943=>"001110000",
  3944=>"011000010",
  3945=>"001100001",
  3946=>"100110111",
  3947=>"110010101",
  3948=>"001101000",
  3949=>"101010111",
  3950=>"011011000",
  3951=>"101000100",
  3952=>"000000000",
  3953=>"011110000",
  3954=>"001011010",
  3955=>"111111101",
  3956=>"000101111",
  3957=>"010010100",
  3958=>"100001001",
  3959=>"010001001",
  3960=>"001000000",
  3961=>"111000111",
  3962=>"001101100",
  3963=>"111011100",
  3964=>"001010111",
  3965=>"111001110",
  3966=>"011001011",
  3967=>"100010001",
  3968=>"010010001",
  3969=>"001010110",
  3970=>"101000111",
  3971=>"000111101",
  3972=>"001101000",
  3973=>"111110110",
  3974=>"011110110",
  3975=>"100100111",
  3976=>"101111000",
  3977=>"100111000",
  3978=>"101101100",
  3979=>"010000011",
  3980=>"111001010",
  3981=>"001000010",
  3982=>"110000000",
  3983=>"111110101",
  3984=>"011110110",
  3985=>"110010100",
  3986=>"000011111",
  3987=>"001100001",
  3988=>"111100110",
  3989=>"100001110",
  3990=>"101000010",
  3991=>"100101010",
  3992=>"101000100",
  3993=>"001011111",
  3994=>"101110101",
  3995=>"010101011",
  3996=>"110010101",
  3997=>"001010111",
  3998=>"001010111",
  3999=>"100000110",
  4000=>"101010011",
  4001=>"011101000",
  4002=>"110000110",
  4003=>"101110011",
  4004=>"001101000",
  4005=>"110110111",
  4006=>"100110001",
  4007=>"101001000",
  4008=>"000110111",
  4009=>"000110110",
  4010=>"000011110",
  4011=>"011111111",
  4012=>"010101011",
  4013=>"000010000",
  4014=>"011000000",
  4015=>"101001101",
  4016=>"111010010",
  4017=>"000000011",
  4018=>"011011000",
  4019=>"001110010",
  4020=>"100101010",
  4021=>"110101111",
  4022=>"100100100",
  4023=>"010000101",
  4024=>"000110111",
  4025=>"111100000",
  4026=>"010010000",
  4027=>"111010110",
  4028=>"001101110",
  4029=>"001101011",
  4030=>"001111001",
  4031=>"000011000",
  4032=>"101111100",
  4033=>"110000010",
  4034=>"101101011",
  4035=>"100101101",
  4036=>"111001011",
  4037=>"001111010",
  4038=>"010001001",
  4039=>"111001010",
  4040=>"000010001",
  4041=>"010000101",
  4042=>"000010000",
  4043=>"100011001",
  4044=>"001111101",
  4045=>"110010000",
  4046=>"000000000",
  4047=>"001100101",
  4048=>"011010111",
  4049=>"110011101",
  4050=>"011001110",
  4051=>"000100100",
  4052=>"111110000",
  4053=>"111110111",
  4054=>"000101101",
  4055=>"110000111",
  4056=>"001111011",
  4057=>"000000111",
  4058=>"110010000",
  4059=>"110100110",
  4060=>"011001010",
  4061=>"000000011",
  4062=>"110011011",
  4063=>"011001111",
  4064=>"110100100",
  4065=>"110101110",
  4066=>"110010111",
  4067=>"010001111",
  4068=>"000000000",
  4069=>"001011111",
  4070=>"010101011",
  4071=>"011000000",
  4072=>"001001011",
  4073=>"111010000",
  4074=>"011000110",
  4075=>"011110111",
  4076=>"010010010",
  4077=>"101011001",
  4078=>"010000111",
  4079=>"001111000",
  4080=>"000111111",
  4081=>"010010110",
  4082=>"011100111",
  4083=>"011101000",
  4084=>"011001101",
  4085=>"101101111",
  4086=>"111110101",
  4087=>"111010111",
  4088=>"110110000",
  4089=>"100001111",
  4090=>"010100010",
  4091=>"100000011",
  4092=>"111001111",
  4093=>"001101010",
  4094=>"000010101",
  4095=>"111011111",
  4096=>"101101110",
  4097=>"110100000",
  4098=>"110010111",
  4099=>"011111001",
  4100=>"001110111",
  4101=>"111001010",
  4102=>"110011011",
  4103=>"100000001",
  4104=>"110010011",
  4105=>"001010100",
  4106=>"100000001",
  4107=>"111001100",
  4108=>"101110001",
  4109=>"000101101",
  4110=>"000000100",
  4111=>"001100110",
  4112=>"100101011",
  4113=>"010000100",
  4114=>"101011110",
  4115=>"001000100",
  4116=>"000100010",
  4117=>"100101011",
  4118=>"010011000",
  4119=>"010011111",
  4120=>"100101100",
  4121=>"010111101",
  4122=>"111110000",
  4123=>"000111010",
  4124=>"000000000",
  4125=>"001111001",
  4126=>"100010101",
  4127=>"011011000",
  4128=>"000010100",
  4129=>"100111100",
  4130=>"100110000",
  4131=>"100101011",
  4132=>"010100100",
  4133=>"101101111",
  4134=>"111011010",
  4135=>"010101000",
  4136=>"001111011",
  4137=>"001100000",
  4138=>"011111110",
  4139=>"100110001",
  4140=>"001110111",
  4141=>"111111100",
  4142=>"000011100",
  4143=>"110111010",
  4144=>"101001111",
  4145=>"001010000",
  4146=>"011011010",
  4147=>"000100000",
  4148=>"000111111",
  4149=>"101001111",
  4150=>"110101110",
  4151=>"001111001",
  4152=>"000111000",
  4153=>"001111101",
  4154=>"000001010",
  4155=>"001000101",
  4156=>"000100011",
  4157=>"100101101",
  4158=>"001111101",
  4159=>"101111101",
  4160=>"011010101",
  4161=>"001000011",
  4162=>"111100001",
  4163=>"101101100",
  4164=>"110100110",
  4165=>"000101110",
  4166=>"110010010",
  4167=>"011011100",
  4168=>"100000010",
  4169=>"110110101",
  4170=>"001110011",
  4171=>"000010110",
  4172=>"110111100",
  4173=>"101101101",
  4174=>"100101110",
  4175=>"110011010",
  4176=>"001100001",
  4177=>"010111010",
  4178=>"100000011",
  4179=>"000010001",
  4180=>"010000100",
  4181=>"101000001",
  4182=>"010111100",
  4183=>"001001001",
  4184=>"110100100",
  4185=>"000101000",
  4186=>"011000000",
  4187=>"100100101",
  4188=>"000000000",
  4189=>"000000010",
  4190=>"101010101",
  4191=>"000100101",
  4192=>"001110111",
  4193=>"101110110",
  4194=>"000011111",
  4195=>"110110000",
  4196=>"110000001",
  4197=>"011111010",
  4198=>"111110101",
  4199=>"001111101",
  4200=>"111111110",
  4201=>"001000011",
  4202=>"000000010",
  4203=>"101100100",
  4204=>"011010000",
  4205=>"000001110",
  4206=>"011110000",
  4207=>"111001100",
  4208=>"001111110",
  4209=>"101101010",
  4210=>"000000100",
  4211=>"100101011",
  4212=>"010110011",
  4213=>"111010010",
  4214=>"111100011",
  4215=>"000110001",
  4216=>"100100101",
  4217=>"110101001",
  4218=>"111010110",
  4219=>"110001000",
  4220=>"010000001",
  4221=>"001010011",
  4222=>"100110001",
  4223=>"110100000",
  4224=>"010101000",
  4225=>"000000110",
  4226=>"110110110",
  4227=>"111001111",
  4228=>"100110101",
  4229=>"001001111",
  4230=>"110010000",
  4231=>"110100100",
  4232=>"010010100",
  4233=>"010001111",
  4234=>"001010101",
  4235=>"010001001",
  4236=>"010101101",
  4237=>"111110000",
  4238=>"100100111",
  4239=>"100000000",
  4240=>"001100011",
  4241=>"110010001",
  4242=>"100011000",
  4243=>"110001101",
  4244=>"010010111",
  4245=>"101111100",
  4246=>"001101110",
  4247=>"000110101",
  4248=>"011011110",
  4249=>"000101011",
  4250=>"010011010",
  4251=>"011010110",
  4252=>"001100110",
  4253=>"100111011",
  4254=>"100001110",
  4255=>"010010001",
  4256=>"100101010",
  4257=>"110000111",
  4258=>"100001011",
  4259=>"001110000",
  4260=>"100101111",
  4261=>"000000111",
  4262=>"001101100",
  4263=>"101010000",
  4264=>"000111101",
  4265=>"010110111",
  4266=>"101100101",
  4267=>"110010000",
  4268=>"110000010",
  4269=>"001000001",
  4270=>"010010000",
  4271=>"110001101",
  4272=>"111100110",
  4273=>"000111010",
  4274=>"101101001",
  4275=>"000110010",
  4276=>"111110010",
  4277=>"110001111",
  4278=>"010000101",
  4279=>"111000111",
  4280=>"000000110",
  4281=>"110001101",
  4282=>"010000000",
  4283=>"000111100",
  4284=>"111010000",
  4285=>"011100010",
  4286=>"001100010",
  4287=>"010011101",
  4288=>"011011100",
  4289=>"000110110",
  4290=>"110101001",
  4291=>"001100011",
  4292=>"000001110",
  4293=>"100000000",
  4294=>"000111101",
  4295=>"110000101",
  4296=>"111011010",
  4297=>"110111110",
  4298=>"001110101",
  4299=>"101011110",
  4300=>"101101011",
  4301=>"010100000",
  4302=>"000111111",
  4303=>"000000010",
  4304=>"101001010",
  4305=>"000000101",
  4306=>"100001001",
  4307=>"101101110",
  4308=>"110010111",
  4309=>"101001111",
  4310=>"111110001",
  4311=>"011000010",
  4312=>"100000000",
  4313=>"000100001",
  4314=>"000110111",
  4315=>"110001100",
  4316=>"111111001",
  4317=>"001010011",
  4318=>"101000000",
  4319=>"101110111",
  4320=>"000000111",
  4321=>"001001100",
  4322=>"011000111",
  4323=>"100010010",
  4324=>"010011101",
  4325=>"000101001",
  4326=>"101010001",
  4327=>"001110110",
  4328=>"000000000",
  4329=>"111111011",
  4330=>"000001110",
  4331=>"101100011",
  4332=>"111010111",
  4333=>"111100111",
  4334=>"010110111",
  4335=>"000000101",
  4336=>"101100111",
  4337=>"111000110",
  4338=>"001101001",
  4339=>"000000111",
  4340=>"010100100",
  4341=>"110001001",
  4342=>"100000000",
  4343=>"100000100",
  4344=>"110010000",
  4345=>"011001011",
  4346=>"000000111",
  4347=>"000000001",
  4348=>"101100001",
  4349=>"011111000",
  4350=>"101100010",
  4351=>"001010010",
  4352=>"101000100",
  4353=>"011011000",
  4354=>"001111111",
  4355=>"011001110",
  4356=>"101000111",
  4357=>"000000000",
  4358=>"011111110",
  4359=>"001001000",
  4360=>"110110111",
  4361=>"111011110",
  4362=>"111011010",
  4363=>"111010111",
  4364=>"110110010",
  4365=>"001000011",
  4366=>"010001111",
  4367=>"001100010",
  4368=>"011110101",
  4369=>"101100111",
  4370=>"001010000",
  4371=>"101111101",
  4372=>"011010111",
  4373=>"011101100",
  4374=>"101101011",
  4375=>"010110101",
  4376=>"011010011",
  4377=>"001100100",
  4378=>"010001101",
  4379=>"101111010",
  4380=>"110001101",
  4381=>"011011101",
  4382=>"000100101",
  4383=>"010100101",
  4384=>"010110100",
  4385=>"010011111",
  4386=>"100011100",
  4387=>"110000010",
  4388=>"010011001",
  4389=>"111111000",
  4390=>"001011001",
  4391=>"101111011",
  4392=>"001101010",
  4393=>"011011001",
  4394=>"000000011",
  4395=>"101001101",
  4396=>"101011111",
  4397=>"101100000",
  4398=>"000000110",
  4399=>"000001001",
  4400=>"101011110",
  4401=>"000011010",
  4402=>"111110000",
  4403=>"100110001",
  4404=>"000101100",
  4405=>"111100011",
  4406=>"011110000",
  4407=>"000110011",
  4408=>"110101111",
  4409=>"001011010",
  4410=>"100100001",
  4411=>"101010010",
  4412=>"100111101",
  4413=>"010111101",
  4414=>"100110110",
  4415=>"101000101",
  4416=>"010110101",
  4417=>"101100100",
  4418=>"000110010",
  4419=>"011010000",
  4420=>"111000011",
  4421=>"010100110",
  4422=>"000000001",
  4423=>"010100111",
  4424=>"110101111",
  4425=>"011011000",
  4426=>"111001100",
  4427=>"011011000",
  4428=>"100111111",
  4429=>"111100001",
  4430=>"111001111",
  4431=>"110101100",
  4432=>"111001100",
  4433=>"010110111",
  4434=>"000000101",
  4435=>"011001111",
  4436=>"000001000",
  4437=>"001010011",
  4438=>"101000011",
  4439=>"011100001",
  4440=>"100011110",
  4441=>"010100010",
  4442=>"001000100",
  4443=>"001110011",
  4444=>"111110101",
  4445=>"000010000",
  4446=>"110100110",
  4447=>"100100011",
  4448=>"110001011",
  4449=>"011101001",
  4450=>"011110000",
  4451=>"000011110",
  4452=>"000111100",
  4453=>"001000111",
  4454=>"101100010",
  4455=>"101000000",
  4456=>"000000011",
  4457=>"111001000",
  4458=>"001100010",
  4459=>"011011010",
  4460=>"001010001",
  4461=>"011001010",
  4462=>"011111110",
  4463=>"000101110",
  4464=>"001000100",
  4465=>"111001010",
  4466=>"110001011",
  4467=>"111110000",
  4468=>"111010010",
  4469=>"010111111",
  4470=>"001001110",
  4471=>"101011100",
  4472=>"000100011",
  4473=>"000011010",
  4474=>"111111111",
  4475=>"011100100",
  4476=>"101000111",
  4477=>"111100000",
  4478=>"010001010",
  4479=>"010111011",
  4480=>"011000011",
  4481=>"100110010",
  4482=>"110111101",
  4483=>"011010100",
  4484=>"010000001",
  4485=>"000000010",
  4486=>"010101101",
  4487=>"100001000",
  4488=>"000101011",
  4489=>"111011101",
  4490=>"000010110",
  4491=>"010101100",
  4492=>"100111000",
  4493=>"101100111",
  4494=>"111000111",
  4495=>"111000010",
  4496=>"001100110",
  4497=>"000010001",
  4498=>"111001000",
  4499=>"001000000",
  4500=>"010010100",
  4501=>"000001110",
  4502=>"110100000",
  4503=>"111110011",
  4504=>"010000001",
  4505=>"000000000",
  4506=>"011101000",
  4507=>"100110100",
  4508=>"011001100",
  4509=>"001110001",
  4510=>"010100100",
  4511=>"111100000",
  4512=>"001100101",
  4513=>"010010001",
  4514=>"011111010",
  4515=>"101000001",
  4516=>"010010010",
  4517=>"000000100",
  4518=>"010010011",
  4519=>"011010000",
  4520=>"111000111",
  4521=>"110011000",
  4522=>"001011111",
  4523=>"110010011",
  4524=>"001100100",
  4525=>"110111110",
  4526=>"000000101",
  4527=>"001000010",
  4528=>"010000111",
  4529=>"100100111",
  4530=>"011100111",
  4531=>"011010100",
  4532=>"000101100",
  4533=>"101001101",
  4534=>"000101001",
  4535=>"000100101",
  4536=>"101110110",
  4537=>"011011001",
  4538=>"011010011",
  4539=>"001101110",
  4540=>"101000101",
  4541=>"010111111",
  4542=>"100000000",
  4543=>"111111110",
  4544=>"101100010",
  4545=>"110000100",
  4546=>"100010110",
  4547=>"100100001",
  4548=>"001010011",
  4549=>"111111111",
  4550=>"100011010",
  4551=>"000000100",
  4552=>"010101100",
  4553=>"011010110",
  4554=>"101111001",
  4555=>"000110001",
  4556=>"101011111",
  4557=>"100100110",
  4558=>"001011110",
  4559=>"011100101",
  4560=>"101001011",
  4561=>"011110001",
  4562=>"010111110",
  4563=>"101010110",
  4564=>"000011101",
  4565=>"011100010",
  4566=>"001000000",
  4567=>"000010010",
  4568=>"011110000",
  4569=>"110010000",
  4570=>"001110111",
  4571=>"001011000",
  4572=>"111011110",
  4573=>"111100111",
  4574=>"011111111",
  4575=>"010010011",
  4576=>"000000001",
  4577=>"101000111",
  4578=>"101111010",
  4579=>"001100110",
  4580=>"101111011",
  4581=>"111110111",
  4582=>"011001010",
  4583=>"101000001",
  4584=>"011000000",
  4585=>"111001111",
  4586=>"101101110",
  4587=>"100110010",
  4588=>"011101001",
  4589=>"101000000",
  4590=>"110010101",
  4591=>"111000000",
  4592=>"100100011",
  4593=>"011010100",
  4594=>"110100011",
  4595=>"011110100",
  4596=>"000010101",
  4597=>"011011000",
  4598=>"101011111",
  4599=>"011100000",
  4600=>"010111110",
  4601=>"011001011",
  4602=>"000100110",
  4603=>"000000000",
  4604=>"010101001",
  4605=>"000011110",
  4606=>"100100011",
  4607=>"000111100",
  4608=>"100001111",
  4609=>"000110111",
  4610=>"010101100",
  4611=>"111100011",
  4612=>"001111101",
  4613=>"000100001",
  4614=>"001000001",
  4615=>"000010100",
  4616=>"000101000",
  4617=>"010111001",
  4618=>"011110001",
  4619=>"111110011",
  4620=>"111101100",
  4621=>"110111111",
  4622=>"110100010",
  4623=>"001011011",
  4624=>"111111100",
  4625=>"010111111",
  4626=>"101001111",
  4627=>"101010011",
  4628=>"110001001",
  4629=>"101101100",
  4630=>"100010111",
  4631=>"101011001",
  4632=>"001000101",
  4633=>"000110010",
  4634=>"000010000",
  4635=>"111001000",
  4636=>"000000000",
  4637=>"110000010",
  4638=>"011100010",
  4639=>"111100001",
  4640=>"010011010",
  4641=>"111100000",
  4642=>"010101011",
  4643=>"100101110",
  4644=>"111100001",
  4645=>"110111001",
  4646=>"111101110",
  4647=>"100000111",
  4648=>"000010001",
  4649=>"000101101",
  4650=>"100110000",
  4651=>"100100011",
  4652=>"100001000",
  4653=>"110000000",
  4654=>"110010001",
  4655=>"001001101",
  4656=>"001001010",
  4657=>"101110000",
  4658=>"100010100",
  4659=>"010111100",
  4660=>"100000100",
  4661=>"001111011",
  4662=>"001011101",
  4663=>"101000001",
  4664=>"101011101",
  4665=>"110011000",
  4666=>"001010100",
  4667=>"001100001",
  4668=>"110011100",
  4669=>"101111000",
  4670=>"100000110",
  4671=>"000011101",
  4672=>"011100010",
  4673=>"100000101",
  4674=>"100000000",
  4675=>"010011101",
  4676=>"000001110",
  4677=>"100101001",
  4678=>"010001100",
  4679=>"001100101",
  4680=>"011011101",
  4681=>"010100010",
  4682=>"100000100",
  4683=>"011000000",
  4684=>"101100100",
  4685=>"111000000",
  4686=>"101100011",
  4687=>"100010101",
  4688=>"010101101",
  4689=>"110011110",
  4690=>"001001101",
  4691=>"000001011",
  4692=>"101100000",
  4693=>"100110010",
  4694=>"111011110",
  4695=>"010111111",
  4696=>"111000011",
  4697=>"000111101",
  4698=>"010110100",
  4699=>"000000000",
  4700=>"111111011",
  4701=>"100111001",
  4702=>"010101001",
  4703=>"011100001",
  4704=>"010010010",
  4705=>"001101010",
  4706=>"111000001",
  4707=>"111110110",
  4708=>"001101010",
  4709=>"010010101",
  4710=>"100000111",
  4711=>"011001010",
  4712=>"111001000",
  4713=>"111011101",
  4714=>"000000010",
  4715=>"001001000",
  4716=>"101011110",
  4717=>"101111001",
  4718=>"000000001",
  4719=>"100000011",
  4720=>"100001001",
  4721=>"001111110",
  4722=>"001011100",
  4723=>"111110111",
  4724=>"001011100",
  4725=>"100000010",
  4726=>"111100001",
  4727=>"110001100",
  4728=>"011111110",
  4729=>"100010111",
  4730=>"011100010",
  4731=>"000110010",
  4732=>"101010001",
  4733=>"110000011",
  4734=>"100100100",
  4735=>"011010000",
  4736=>"100000110",
  4737=>"111000100",
  4738=>"011011000",
  4739=>"000111101",
  4740=>"111000010",
  4741=>"000010000",
  4742=>"110001011",
  4743=>"011010010",
  4744=>"111011111",
  4745=>"011000001",
  4746=>"011010111",
  4747=>"011100010",
  4748=>"100000010",
  4749=>"011111000",
  4750=>"110000111",
  4751=>"010011100",
  4752=>"010011011",
  4753=>"111011001",
  4754=>"111100000",
  4755=>"011110101",
  4756=>"000000010",
  4757=>"010110110",
  4758=>"011010101",
  4759=>"101110001",
  4760=>"110110111",
  4761=>"111101111",
  4762=>"011010001",
  4763=>"110000100",
  4764=>"111101000",
  4765=>"000110110",
  4766=>"111100100",
  4767=>"000010110",
  4768=>"111100011",
  4769=>"100111100",
  4770=>"111111111",
  4771=>"010000100",
  4772=>"001101011",
  4773=>"011000111",
  4774=>"011000101",
  4775=>"101101101",
  4776=>"111011011",
  4777=>"001010001",
  4778=>"010110111",
  4779=>"110101110",
  4780=>"110101100",
  4781=>"011011010",
  4782=>"111000011",
  4783=>"100000001",
  4784=>"111000100",
  4785=>"000011110",
  4786=>"001111011",
  4787=>"000111100",
  4788=>"010111011",
  4789=>"111001101",
  4790=>"101011010",
  4791=>"111111000",
  4792=>"100000001",
  4793=>"101010000",
  4794=>"111000110",
  4795=>"011111000",
  4796=>"100000100",
  4797=>"010000010",
  4798=>"110100000",
  4799=>"000111010",
  4800=>"111110011",
  4801=>"001110110",
  4802=>"000010100",
  4803=>"100101101",
  4804=>"001111011",
  4805=>"001111111",
  4806=>"011000111",
  4807=>"101000000",
  4808=>"000011000",
  4809=>"100001011",
  4810=>"101010001",
  4811=>"000011111",
  4812=>"000100000",
  4813=>"111110001",
  4814=>"100001011",
  4815=>"110001001",
  4816=>"001010000",
  4817=>"010011111",
  4818=>"111011011",
  4819=>"001110100",
  4820=>"001011100",
  4821=>"010001000",
  4822=>"110100011",
  4823=>"110101111",
  4824=>"000010011",
  4825=>"011011111",
  4826=>"000010000",
  4827=>"101000011",
  4828=>"101001010",
  4829=>"101110010",
  4830=>"101010000",
  4831=>"010000100",
  4832=>"010010000",
  4833=>"010100010",
  4834=>"010101010",
  4835=>"001111110",
  4836=>"101010111",
  4837=>"000111111",
  4838=>"110101100",
  4839=>"010100010",
  4840=>"011011100",
  4841=>"011001101",
  4842=>"011001010",
  4843=>"111111010",
  4844=>"110000110",
  4845=>"101111111",
  4846=>"000010001",
  4847=>"101000001",
  4848=>"100010110",
  4849=>"101000111",
  4850=>"100111000",
  4851=>"111101101",
  4852=>"100110101",
  4853=>"111111000",
  4854=>"010000110",
  4855=>"110001100",
  4856=>"010100011",
  4857=>"100001100",
  4858=>"101011100",
  4859=>"011101000",
  4860=>"010000010",
  4861=>"100101100",
  4862=>"101001001",
  4863=>"001010000",
  4864=>"100101001",
  4865=>"010010011",
  4866=>"101010000",
  4867=>"100111111",
  4868=>"001001010",
  4869=>"110001010",
  4870=>"111101110",
  4871=>"010100101",
  4872=>"000001110",
  4873=>"001001101",
  4874=>"001101101",
  4875=>"001110001",
  4876=>"111001110",
  4877=>"111111011",
  4878=>"010111110",
  4879=>"111111111",
  4880=>"111010100",
  4881=>"001011011",
  4882=>"010110100",
  4883=>"000111111",
  4884=>"001011000",
  4885=>"101000110",
  4886=>"011001001",
  4887=>"010101001",
  4888=>"011010000",
  4889=>"000100000",
  4890=>"000100101",
  4891=>"110011111",
  4892=>"101011011",
  4893=>"110010101",
  4894=>"011100110",
  4895=>"100110000",
  4896=>"011000011",
  4897=>"101111010",
  4898=>"111011001",
  4899=>"100011000",
  4900=>"110111000",
  4901=>"110011110",
  4902=>"110001011",
  4903=>"000001000",
  4904=>"100100101",
  4905=>"101010111",
  4906=>"101010010",
  4907=>"001001110",
  4908=>"011100011",
  4909=>"100011100",
  4910=>"110010000",
  4911=>"100101110",
  4912=>"101110010",
  4913=>"100010011",
  4914=>"100010010",
  4915=>"110110001",
  4916=>"000010111",
  4917=>"101110100",
  4918=>"101011010",
  4919=>"000101001",
  4920=>"011011011",
  4921=>"001000010",
  4922=>"101001110",
  4923=>"000010111",
  4924=>"100101011",
  4925=>"110010000",
  4926=>"000010011",
  4927=>"111101110",
  4928=>"000010000",
  4929=>"000000110",
  4930=>"000001111",
  4931=>"110101010",
  4932=>"111100011",
  4933=>"001110110",
  4934=>"000011101",
  4935=>"011011011",
  4936=>"011001111",
  4937=>"010001000",
  4938=>"000001110",
  4939=>"111001101",
  4940=>"100001010",
  4941=>"110110101",
  4942=>"001110111",
  4943=>"011100010",
  4944=>"110111000",
  4945=>"110000000",
  4946=>"000001000",
  4947=>"001011110",
  4948=>"101111000",
  4949=>"110000001",
  4950=>"010011110",
  4951=>"100110110",
  4952=>"011010110",
  4953=>"101000110",
  4954=>"000100011",
  4955=>"110110001",
  4956=>"011101111",
  4957=>"011111111",
  4958=>"111100101",
  4959=>"000101000",
  4960=>"011000010",
  4961=>"100011010",
  4962=>"000011000",
  4963=>"111001111",
  4964=>"010110110",
  4965=>"100101000",
  4966=>"111011111",
  4967=>"110000011",
  4968=>"010101101",
  4969=>"100100001",
  4970=>"001010100",
  4971=>"111111111",
  4972=>"100010111",
  4973=>"001000110",
  4974=>"000101011",
  4975=>"011011001",
  4976=>"111001000",
  4977=>"010000001",
  4978=>"101110011",
  4979=>"110101000",
  4980=>"010010011",
  4981=>"111111100",
  4982=>"101100110",
  4983=>"101101101",
  4984=>"101011100",
  4985=>"111011111",
  4986=>"000100101",
  4987=>"011011000",
  4988=>"000110010",
  4989=>"110101000",
  4990=>"110110111",
  4991=>"110110011",
  4992=>"011110101",
  4993=>"100100101",
  4994=>"001000100",
  4995=>"011100101",
  4996=>"000000010",
  4997=>"111010110",
  4998=>"001000111",
  4999=>"001000010",
  5000=>"110110111",
  5001=>"110001011",
  5002=>"100001011",
  5003=>"011101000",
  5004=>"001111001",
  5005=>"000110010",
  5006=>"011001001",
  5007=>"010000000",
  5008=>"010000011",
  5009=>"101011110",
  5010=>"000000110",
  5011=>"100000010",
  5012=>"100100000",
  5013=>"001010010",
  5014=>"001001101",
  5015=>"011010001",
  5016=>"110010011",
  5017=>"011110001",
  5018=>"110110001",
  5019=>"001010010",
  5020=>"110101111",
  5021=>"111111101",
  5022=>"101010001",
  5023=>"011011101",
  5024=>"011110100",
  5025=>"011101001",
  5026=>"110111111",
  5027=>"100110010",
  5028=>"000111000",
  5029=>"110001100",
  5030=>"010101001",
  5031=>"001111011",
  5032=>"000000101",
  5033=>"011000111",
  5034=>"111000110",
  5035=>"101000110",
  5036=>"001001001",
  5037=>"110111010",
  5038=>"100110100",
  5039=>"010001001",
  5040=>"110000111",
  5041=>"100101110",
  5042=>"101000010",
  5043=>"011110011",
  5044=>"001110000",
  5045=>"100001110",
  5046=>"100001111",
  5047=>"001001001",
  5048=>"111111100",
  5049=>"111111111",
  5050=>"111011100",
  5051=>"100011100",
  5052=>"101101010",
  5053=>"111000000",
  5054=>"000011000",
  5055=>"000101111",
  5056=>"000000010",
  5057=>"100001101",
  5058=>"110101111",
  5059=>"101000000",
  5060=>"000100001",
  5061=>"000111001",
  5062=>"101100111",
  5063=>"100000001",
  5064=>"110110100",
  5065=>"111011111",
  5066=>"001101101",
  5067=>"111010001",
  5068=>"010001010",
  5069=>"101110100",
  5070=>"001000100",
  5071=>"110001110",
  5072=>"011110111",
  5073=>"000111011",
  5074=>"100100110",
  5075=>"111101110",
  5076=>"111010000",
  5077=>"011101000",
  5078=>"101010011",
  5079=>"111000111",
  5080=>"110111000",
  5081=>"010010000",
  5082=>"101000001",
  5083=>"100001010",
  5084=>"011001100",
  5085=>"101000100",
  5086=>"011101011",
  5087=>"001001011",
  5088=>"001110000",
  5089=>"100100000",
  5090=>"010011101",
  5091=>"111011010",
  5092=>"001110111",
  5093=>"100001010",
  5094=>"011100000",
  5095=>"000110101",
  5096=>"100000101",
  5097=>"111110111",
  5098=>"000011101",
  5099=>"110110101",
  5100=>"100110010",
  5101=>"101001010",
  5102=>"100100111",
  5103=>"000000111",
  5104=>"100111110",
  5105=>"001100011",
  5106=>"010000010",
  5107=>"000010110",
  5108=>"110110111",
  5109=>"111000010",
  5110=>"111101011",
  5111=>"100011001",
  5112=>"110100000",
  5113=>"111001000",
  5114=>"101101101",
  5115=>"101000101",
  5116=>"110000001",
  5117=>"111000110",
  5118=>"111010011",
  5119=>"001100001",
  5120=>"010111110",
  5121=>"010110011",
  5122=>"001100001",
  5123=>"101011010",
  5124=>"101111010",
  5125=>"000110011",
  5126=>"101110111",
  5127=>"100111110",
  5128=>"011100110",
  5129=>"001100001",
  5130=>"101111011",
  5131=>"101011101",
  5132=>"000000010",
  5133=>"101001111",
  5134=>"110011010",
  5135=>"111101111",
  5136=>"001010100",
  5137=>"100110100",
  5138=>"000111100",
  5139=>"011000110",
  5140=>"100000100",
  5141=>"110101111",
  5142=>"101011111",
  5143=>"001010011",
  5144=>"110110000",
  5145=>"101000111",
  5146=>"001000101",
  5147=>"011000111",
  5148=>"110110111",
  5149=>"100000101",
  5150=>"001111101",
  5151=>"111101110",
  5152=>"011100011",
  5153=>"000110111",
  5154=>"001100001",
  5155=>"001000000",
  5156=>"000111101",
  5157=>"100001000",
  5158=>"111011100",
  5159=>"100001000",
  5160=>"011111000",
  5161=>"001010000",
  5162=>"010010011",
  5163=>"001101010",
  5164=>"011101011",
  5165=>"111000000",
  5166=>"010110111",
  5167=>"110100100",
  5168=>"010100000",
  5169=>"010111111",
  5170=>"011101001",
  5171=>"001100101",
  5172=>"100111001",
  5173=>"001000000",
  5174=>"001100100",
  5175=>"010111000",
  5176=>"000100011",
  5177=>"100000001",
  5178=>"100100001",
  5179=>"100001001",
  5180=>"010010001",
  5181=>"100100101",
  5182=>"101100001",
  5183=>"000101111",
  5184=>"101000001",
  5185=>"011010100",
  5186=>"000001001",
  5187=>"001111110",
  5188=>"000110111",
  5189=>"110101000",
  5190=>"001000111",
  5191=>"111111101",
  5192=>"111110000",
  5193=>"110011001",
  5194=>"011100001",
  5195=>"000000101",
  5196=>"100001001",
  5197=>"011011100",
  5198=>"000111011",
  5199=>"011100110",
  5200=>"101000010",
  5201=>"100011010",
  5202=>"010000010",
  5203=>"010111000",
  5204=>"011110010",
  5205=>"101000111",
  5206=>"110010101",
  5207=>"010100010",
  5208=>"110110101",
  5209=>"010111001",
  5210=>"010001010",
  5211=>"010111111",
  5212=>"110100101",
  5213=>"101001101",
  5214=>"010100111",
  5215=>"101101110",
  5216=>"010100111",
  5217=>"110000000",
  5218=>"000000001",
  5219=>"111000011",
  5220=>"111000111",
  5221=>"100010001",
  5222=>"101011101",
  5223=>"000000101",
  5224=>"010110111",
  5225=>"011111011",
  5226=>"011100000",
  5227=>"001001010",
  5228=>"000010001",
  5229=>"011010101",
  5230=>"001101001",
  5231=>"000110001",
  5232=>"000101000",
  5233=>"100010100",
  5234=>"110001001",
  5235=>"000010011",
  5236=>"111110011",
  5237=>"100100000",
  5238=>"010011011",
  5239=>"010110111",
  5240=>"111100100",
  5241=>"111010011",
  5242=>"000000101",
  5243=>"010010101",
  5244=>"000001001",
  5245=>"000000000",
  5246=>"000000111",
  5247=>"011011000",
  5248=>"000111001",
  5249=>"100111010",
  5250=>"101100100",
  5251=>"011111111",
  5252=>"111000000",
  5253=>"110011101",
  5254=>"010100000",
  5255=>"111100001",
  5256=>"110010111",
  5257=>"010000011",
  5258=>"011010101",
  5259=>"010010101",
  5260=>"110111011",
  5261=>"001101010",
  5262=>"110101100",
  5263=>"111010110",
  5264=>"011010011",
  5265=>"100000010",
  5266=>"010110000",
  5267=>"011011101",
  5268=>"000011101",
  5269=>"110110001",
  5270=>"011111100",
  5271=>"111101111",
  5272=>"001110011",
  5273=>"010000001",
  5274=>"101000011",
  5275=>"110100110",
  5276=>"001111010",
  5277=>"000101000",
  5278=>"111111100",
  5279=>"001001001",
  5280=>"001011101",
  5281=>"000000011",
  5282=>"110010001",
  5283=>"101110011",
  5284=>"010010100",
  5285=>"100101110",
  5286=>"111010101",
  5287=>"010101101",
  5288=>"001010100",
  5289=>"011100000",
  5290=>"011010101",
  5291=>"000000010",
  5292=>"011110111",
  5293=>"001110011",
  5294=>"000010101",
  5295=>"001000101",
  5296=>"011001011",
  5297=>"010001000",
  5298=>"000101000",
  5299=>"000000010",
  5300=>"001100010",
  5301=>"001001010",
  5302=>"000011100",
  5303=>"100100011",
  5304=>"010010011",
  5305=>"001011011",
  5306=>"001100010",
  5307=>"000010001",
  5308=>"101001111",
  5309=>"100001001",
  5310=>"001001101",
  5311=>"111000110",
  5312=>"110000111",
  5313=>"011011100",
  5314=>"111010000",
  5315=>"011110100",
  5316=>"011101000",
  5317=>"101110000",
  5318=>"100110011",
  5319=>"101101111",
  5320=>"000100110",
  5321=>"000001111",
  5322=>"010110111",
  5323=>"001111011",
  5324=>"001100100",
  5325=>"001101111",
  5326=>"000001101",
  5327=>"100110110",
  5328=>"100101111",
  5329=>"001011011",
  5330=>"011101010",
  5331=>"001011110",
  5332=>"101100011",
  5333=>"101000001",
  5334=>"110011000",
  5335=>"100001000",
  5336=>"011001010",
  5337=>"011111110",
  5338=>"010110001",
  5339=>"110111101",
  5340=>"101011000",
  5341=>"100100100",
  5342=>"011000001",
  5343=>"110110111",
  5344=>"010101001",
  5345=>"001010001",
  5346=>"011011010",
  5347=>"000010100",
  5348=>"010100110",
  5349=>"011100100",
  5350=>"000111001",
  5351=>"000101001",
  5352=>"101000101",
  5353=>"011001111",
  5354=>"100000000",
  5355=>"000010101",
  5356=>"110111010",
  5357=>"011000010",
  5358=>"001100110",
  5359=>"010011011",
  5360=>"011000011",
  5361=>"110110000",
  5362=>"010000100",
  5363=>"111011000",
  5364=>"000011010",
  5365=>"000000000",
  5366=>"111010110",
  5367=>"110001011",
  5368=>"110110001",
  5369=>"110000111",
  5370=>"011001111",
  5371=>"010010011",
  5372=>"111110111",
  5373=>"110100000",
  5374=>"111000100",
  5375=>"111111100",
  5376=>"000000100",
  5377=>"100110101",
  5378=>"110110011",
  5379=>"110011010",
  5380=>"010100100",
  5381=>"100100101",
  5382=>"111111111",
  5383=>"001010100",
  5384=>"110111000",
  5385=>"010111001",
  5386=>"010101000",
  5387=>"110111001",
  5388=>"011011110",
  5389=>"110000000",
  5390=>"111101000",
  5391=>"101111100",
  5392=>"011100000",
  5393=>"010010110",
  5394=>"011110100",
  5395=>"110010100",
  5396=>"000111011",
  5397=>"111000110",
  5398=>"000010111",
  5399=>"000000010",
  5400=>"001111111",
  5401=>"000001110",
  5402=>"110111111",
  5403=>"011011000",
  5404=>"111100111",
  5405=>"100000111",
  5406=>"010011111",
  5407=>"011001011",
  5408=>"010011111",
  5409=>"011111010",
  5410=>"001101110",
  5411=>"100111001",
  5412=>"100001101",
  5413=>"010111100",
  5414=>"001110110",
  5415=>"111001111",
  5416=>"001000001",
  5417=>"010101100",
  5418=>"110101100",
  5419=>"111011101",
  5420=>"011001000",
  5421=>"110011010",
  5422=>"010000111",
  5423=>"110010010",
  5424=>"101011010",
  5425=>"000000100",
  5426=>"100101110",
  5427=>"110000011",
  5428=>"011010101",
  5429=>"111010000",
  5430=>"011010000",
  5431=>"001001010",
  5432=>"011100011",
  5433=>"010110000",
  5434=>"010101100",
  5435=>"001100010",
  5436=>"100111011",
  5437=>"000001101",
  5438=>"010000011",
  5439=>"001100111",
  5440=>"111101000",
  5441=>"000101010",
  5442=>"111100000",
  5443=>"100100010",
  5444=>"111101000",
  5445=>"001001111",
  5446=>"001010000",
  5447=>"110010000",
  5448=>"110110110",
  5449=>"011100000",
  5450=>"011010001",
  5451=>"001000000",
  5452=>"111101101",
  5453=>"010010101",
  5454=>"101110010",
  5455=>"101111111",
  5456=>"110111111",
  5457=>"000100100",
  5458=>"111100001",
  5459=>"010000001",
  5460=>"010001011",
  5461=>"110100101",
  5462=>"001011010",
  5463=>"101000000",
  5464=>"110011010",
  5465=>"100100111",
  5466=>"001111100",
  5467=>"101001100",
  5468=>"110011110",
  5469=>"001011011",
  5470=>"000100011",
  5471=>"000100000",
  5472=>"011000110",
  5473=>"110110001",
  5474=>"011011101",
  5475=>"011010011",
  5476=>"010100100",
  5477=>"100100011",
  5478=>"001111100",
  5479=>"100011100",
  5480=>"111111011",
  5481=>"010011011",
  5482=>"001101001",
  5483=>"110011101",
  5484=>"010110000",
  5485=>"001111111",
  5486=>"010001011",
  5487=>"001010110",
  5488=>"101001001",
  5489=>"110000001",
  5490=>"011110111",
  5491=>"111001110",
  5492=>"111100010",
  5493=>"001010110",
  5494=>"011101001",
  5495=>"000110000",
  5496=>"001110000",
  5497=>"100001011",
  5498=>"111111011",
  5499=>"011010010",
  5500=>"010000000",
  5501=>"100001011",
  5502=>"000111101",
  5503=>"000011010",
  5504=>"011110001",
  5505=>"111110111",
  5506=>"001010111",
  5507=>"101011110",
  5508=>"011010001",
  5509=>"000001010",
  5510=>"000001100",
  5511=>"001101010",
  5512=>"100110011",
  5513=>"001000010",
  5514=>"110000101",
  5515=>"111001101",
  5516=>"000010001",
  5517=>"010011000",
  5518=>"110001100",
  5519=>"110101010",
  5520=>"100000101",
  5521=>"100111101",
  5522=>"100110110",
  5523=>"010110001",
  5524=>"010010010",
  5525=>"011101010",
  5526=>"010110011",
  5527=>"111001000",
  5528=>"010111111",
  5529=>"110000011",
  5530=>"101011011",
  5531=>"110001010",
  5532=>"111001111",
  5533=>"011001111",
  5534=>"110010000",
  5535=>"001111110",
  5536=>"011011000",
  5537=>"111000110",
  5538=>"101001000",
  5539=>"111100100",
  5540=>"000100110",
  5541=>"001000010",
  5542=>"001000100",
  5543=>"000110101",
  5544=>"010010011",
  5545=>"010100011",
  5546=>"000101110",
  5547=>"010010111",
  5548=>"100100110",
  5549=>"000000110",
  5550=>"001010110",
  5551=>"100000100",
  5552=>"011001100",
  5553=>"101101110",
  5554=>"011000011",
  5555=>"111011101",
  5556=>"010010111",
  5557=>"101101110",
  5558=>"100111011",
  5559=>"101010111",
  5560=>"010101100",
  5561=>"001100111",
  5562=>"001100011",
  5563=>"111111010",
  5564=>"101100111",
  5565=>"100111111",
  5566=>"011110000",
  5567=>"001101100",
  5568=>"111010000",
  5569=>"000001101",
  5570=>"010111010",
  5571=>"010000111",
  5572=>"000010001",
  5573=>"101100000",
  5574=>"110000001",
  5575=>"010001001",
  5576=>"010110011",
  5577=>"110010000",
  5578=>"101001111",
  5579=>"100100001",
  5580=>"111011101",
  5581=>"001000110",
  5582=>"010011010",
  5583=>"010000011",
  5584=>"101000110",
  5585=>"001001000",
  5586=>"000010101",
  5587=>"100110001",
  5588=>"000101101",
  5589=>"000000010",
  5590=>"111111101",
  5591=>"010100001",
  5592=>"001110101",
  5593=>"001110001",
  5594=>"000101100",
  5595=>"001001000",
  5596=>"101011011",
  5597=>"011001010",
  5598=>"110101000",
  5599=>"010111100",
  5600=>"101000101",
  5601=>"111110011",
  5602=>"110100011",
  5603=>"111001100",
  5604=>"101010111",
  5605=>"010100010",
  5606=>"010111111",
  5607=>"110000110",
  5608=>"101110001",
  5609=>"110011111",
  5610=>"001010001",
  5611=>"010111001",
  5612=>"010010100",
  5613=>"110010110",
  5614=>"000111000",
  5615=>"000010101",
  5616=>"010101111",
  5617=>"001101111",
  5618=>"100001000",
  5619=>"110100100",
  5620=>"101001111",
  5621=>"111101010",
  5622=>"001110011",
  5623=>"001111000",
  5624=>"110111000",
  5625=>"011110000",
  5626=>"001001001",
  5627=>"101101111",
  5628=>"100111101",
  5629=>"101010110",
  5630=>"111101101",
  5631=>"111011000",
  5632=>"100011010",
  5633=>"010100011",
  5634=>"001010110",
  5635=>"000110100",
  5636=>"100101000",
  5637=>"111010111",
  5638=>"010010110",
  5639=>"000011110",
  5640=>"000101110",
  5641=>"000001011",
  5642=>"000111101",
  5643=>"010101010",
  5644=>"111010010",
  5645=>"001110101",
  5646=>"111000111",
  5647=>"111111010",
  5648=>"000111100",
  5649=>"100101101",
  5650=>"000111100",
  5651=>"010101001",
  5652=>"011110000",
  5653=>"101101000",
  5654=>"011100001",
  5655=>"000111111",
  5656=>"110010100",
  5657=>"101001111",
  5658=>"111111100",
  5659=>"010011000",
  5660=>"101111110",
  5661=>"110101111",
  5662=>"000000010",
  5663=>"010100001",
  5664=>"001001001",
  5665=>"011001000",
  5666=>"001011000",
  5667=>"110110001",
  5668=>"010011100",
  5669=>"101010100",
  5670=>"110111110",
  5671=>"001000000",
  5672=>"000101101",
  5673=>"101111010",
  5674=>"011111001",
  5675=>"010001011",
  5676=>"011101001",
  5677=>"010011001",
  5678=>"101101011",
  5679=>"011110111",
  5680=>"100001010",
  5681=>"001111110",
  5682=>"010010011",
  5683=>"011001010",
  5684=>"100000000",
  5685=>"101011101",
  5686=>"101110000",
  5687=>"000000111",
  5688=>"010011001",
  5689=>"011110000",
  5690=>"010111101",
  5691=>"001100000",
  5692=>"100000001",
  5693=>"001111010",
  5694=>"110110011",
  5695=>"100110001",
  5696=>"011100100",
  5697=>"001100110",
  5698=>"000000000",
  5699=>"101010010",
  5700=>"011010011",
  5701=>"011101100",
  5702=>"110000000",
  5703=>"110010000",
  5704=>"100011011",
  5705=>"010001000",
  5706=>"110010100",
  5707=>"010011011",
  5708=>"000001000",
  5709=>"011011001",
  5710=>"111100111",
  5711=>"011111110",
  5712=>"100100101",
  5713=>"011111010",
  5714=>"000000010",
  5715=>"000000010",
  5716=>"101000000",
  5717=>"100110100",
  5718=>"001000001",
  5719=>"110011100",
  5720=>"010101110",
  5721=>"010010001",
  5722=>"110101101",
  5723=>"011001110",
  5724=>"011110110",
  5725=>"101001000",
  5726=>"010110000",
  5727=>"000011011",
  5728=>"101111010",
  5729=>"001000110",
  5730=>"101110001",
  5731=>"000111000",
  5732=>"111111001",
  5733=>"111100101",
  5734=>"111011100",
  5735=>"010101011",
  5736=>"110011100",
  5737=>"001110100",
  5738=>"111001111",
  5739=>"010000010",
  5740=>"000011111",
  5741=>"110000010",
  5742=>"110001000",
  5743=>"100001001",
  5744=>"111101110",
  5745=>"000110100",
  5746=>"101011001",
  5747=>"001001110",
  5748=>"000000011",
  5749=>"011101011",
  5750=>"000001111",
  5751=>"101111110",
  5752=>"011001001",
  5753=>"010110011",
  5754=>"100000011",
  5755=>"011001000",
  5756=>"110010001",
  5757=>"011100010",
  5758=>"010000000",
  5759=>"100101011",
  5760=>"000000101",
  5761=>"001111101",
  5762=>"001111010",
  5763=>"010101001",
  5764=>"110110110",
  5765=>"010100010",
  5766=>"001001100",
  5767=>"100111110",
  5768=>"100100010",
  5769=>"000000001",
  5770=>"101110000",
  5771=>"001000000",
  5772=>"110010100",
  5773=>"001101111",
  5774=>"101100111",
  5775=>"101110100",
  5776=>"000100010",
  5777=>"010101001",
  5778=>"110000001",
  5779=>"100100111",
  5780=>"111000000",
  5781=>"100010100",
  5782=>"011001010",
  5783=>"111001101",
  5784=>"111011011",
  5785=>"011110110",
  5786=>"000101011",
  5787=>"000100001",
  5788=>"011000000",
  5789=>"010100000",
  5790=>"111110010",
  5791=>"101110011",
  5792=>"111100000",
  5793=>"100001111",
  5794=>"010001110",
  5795=>"001011010",
  5796=>"110001000",
  5797=>"001100011",
  5798=>"101001010",
  5799=>"100011001",
  5800=>"100100100",
  5801=>"011000111",
  5802=>"110011010",
  5803=>"100111110",
  5804=>"000011011",
  5805=>"111000110",
  5806=>"111111111",
  5807=>"010010000",
  5808=>"010101100",
  5809=>"101111101",
  5810=>"100001111",
  5811=>"001001001",
  5812=>"000000001",
  5813=>"000111000",
  5814=>"010110100",
  5815=>"010001010",
  5816=>"111111010",
  5817=>"100000000",
  5818=>"011100100",
  5819=>"111111001",
  5820=>"010000111",
  5821=>"011011101",
  5822=>"000101001",
  5823=>"110011101",
  5824=>"000101011",
  5825=>"010010001",
  5826=>"000100110",
  5827=>"111010101",
  5828=>"110011111",
  5829=>"100101000",
  5830=>"001110101",
  5831=>"110011111",
  5832=>"000000001",
  5833=>"000011000",
  5834=>"100110101",
  5835=>"110000110",
  5836=>"000010011",
  5837=>"000010100",
  5838=>"001110101",
  5839=>"110111110",
  5840=>"000100011",
  5841=>"110111010",
  5842=>"101110000",
  5843=>"100010111",
  5844=>"011000010",
  5845=>"000101111",
  5846=>"100000001",
  5847=>"110111001",
  5848=>"011100010",
  5849=>"100100100",
  5850=>"001010001",
  5851=>"000011001",
  5852=>"001111100",
  5853=>"110000000",
  5854=>"111111101",
  5855=>"101111001",
  5856=>"010010110",
  5857=>"100011101",
  5858=>"111000000",
  5859=>"000011001",
  5860=>"010110111",
  5861=>"110000001",
  5862=>"100101111",
  5863=>"010000101",
  5864=>"110101011",
  5865=>"010001011",
  5866=>"010100011",
  5867=>"001100011",
  5868=>"010100001",
  5869=>"101110001",
  5870=>"000101101",
  5871=>"001001101",
  5872=>"011111110",
  5873=>"100010110",
  5874=>"101110011",
  5875=>"000011001",
  5876=>"110111000",
  5877=>"100011110",
  5878=>"111110100",
  5879=>"111001100",
  5880=>"001111111",
  5881=>"010010000",
  5882=>"100010001",
  5883=>"010010000",
  5884=>"000011010",
  5885=>"101101010",
  5886=>"011010000",
  5887=>"111001000",
  5888=>"110000101",
  5889=>"000011000",
  5890=>"011001101",
  5891=>"111000011",
  5892=>"101001010",
  5893=>"101000001",
  5894=>"101000001",
  5895=>"010010011",
  5896=>"101001101",
  5897=>"111000010",
  5898=>"011000111",
  5899=>"111001011",
  5900=>"000101010",
  5901=>"111111110",
  5902=>"101100011",
  5903=>"110111110",
  5904=>"110110011",
  5905=>"001101011",
  5906=>"100000110",
  5907=>"111000010",
  5908=>"001001101",
  5909=>"001101000",
  5910=>"001000000",
  5911=>"100100001",
  5912=>"011000100",
  5913=>"101110010",
  5914=>"100011001",
  5915=>"111100000",
  5916=>"110001100",
  5917=>"110010000",
  5918=>"011001001",
  5919=>"111111010",
  5920=>"110011111",
  5921=>"111000011",
  5922=>"010101101",
  5923=>"010111000",
  5924=>"110110110",
  5925=>"100100000",
  5926=>"101011110",
  5927=>"001010011",
  5928=>"001001010",
  5929=>"110001001",
  5930=>"100010110",
  5931=>"011100100",
  5932=>"110001110",
  5933=>"111000111",
  5934=>"011010010",
  5935=>"001110111",
  5936=>"101000111",
  5937=>"000111011",
  5938=>"110001111",
  5939=>"000011101",
  5940=>"110010010",
  5941=>"000110000",
  5942=>"101110110",
  5943=>"000100000",
  5944=>"111110101",
  5945=>"001000000",
  5946=>"010000100",
  5947=>"101110100",
  5948=>"111101111",
  5949=>"101010001",
  5950=>"101011110",
  5951=>"011010101",
  5952=>"100011000",
  5953=>"100000100",
  5954=>"110011101",
  5955=>"011011111",
  5956=>"000110001",
  5957=>"001111001",
  5958=>"101001111",
  5959=>"110110110",
  5960=>"011001101",
  5961=>"101011001",
  5962=>"010110101",
  5963=>"000100000",
  5964=>"000110000",
  5965=>"001100100",
  5966=>"000000001",
  5967=>"010111001",
  5968=>"010010011",
  5969=>"110010001",
  5970=>"010010011",
  5971=>"010000011",
  5972=>"000001000",
  5973=>"110111011",
  5974=>"000000111",
  5975=>"111001011",
  5976=>"000001110",
  5977=>"010010011",
  5978=>"110101011",
  5979=>"100101111",
  5980=>"100010011",
  5981=>"001010001",
  5982=>"100100001",
  5983=>"100001100",
  5984=>"100110011",
  5985=>"100101010",
  5986=>"110011100",
  5987=>"110111101",
  5988=>"001001011",
  5989=>"001011000",
  5990=>"000000001",
  5991=>"100000100",
  5992=>"110010000",
  5993=>"100100000",
  5994=>"111011101",
  5995=>"100011001",
  5996=>"000011110",
  5997=>"001010100",
  5998=>"100100110",
  5999=>"111000101",
  6000=>"001000011",
  6001=>"011110101",
  6002=>"010100000",
  6003=>"010001010",
  6004=>"010100111",
  6005=>"011100011",
  6006=>"000001111",
  6007=>"001000000",
  6008=>"100000110",
  6009=>"011010001",
  6010=>"011001110",
  6011=>"110011110",
  6012=>"000100110",
  6013=>"100100000",
  6014=>"100100000",
  6015=>"101010011",
  6016=>"111111100",
  6017=>"011101001",
  6018=>"000010010",
  6019=>"001001000",
  6020=>"111010100",
  6021=>"000010000",
  6022=>"111110000",
  6023=>"000000110",
  6024=>"101010010",
  6025=>"100000000",
  6026=>"011110000",
  6027=>"001110101",
  6028=>"001001000",
  6029=>"111011000",
  6030=>"011101010",
  6031=>"111111010",
  6032=>"001100011",
  6033=>"110011100",
  6034=>"101001111",
  6035=>"000001000",
  6036=>"011010110",
  6037=>"111110111",
  6038=>"001111000",
  6039=>"100100111",
  6040=>"001010011",
  6041=>"000000100",
  6042=>"101001000",
  6043=>"001011001",
  6044=>"000010010",
  6045=>"010110111",
  6046=>"001010100",
  6047=>"100110111",
  6048=>"111001111",
  6049=>"000101000",
  6050=>"100110100",
  6051=>"000111100",
  6052=>"001000110",
  6053=>"001101011",
  6054=>"100110100",
  6055=>"101011101",
  6056=>"001110010",
  6057=>"011011010",
  6058=>"110111111",
  6059=>"010110101",
  6060=>"110010111",
  6061=>"001111010",
  6062=>"000101100",
  6063=>"000111011",
  6064=>"010011101",
  6065=>"000101100",
  6066=>"000001010",
  6067=>"100000000",
  6068=>"110011110",
  6069=>"000110110",
  6070=>"000100000",
  6071=>"010001111",
  6072=>"100010100",
  6073=>"100010010",
  6074=>"011100101",
  6075=>"001111001",
  6076=>"011001110",
  6077=>"010000011",
  6078=>"110100101",
  6079=>"100001001",
  6080=>"110100100",
  6081=>"110101110",
  6082=>"110100011",
  6083=>"011111011",
  6084=>"000001001",
  6085=>"101100101",
  6086=>"100000010",
  6087=>"111101110",
  6088=>"000110000",
  6089=>"010000111",
  6090=>"001101110",
  6091=>"010001000",
  6092=>"000100010",
  6093=>"101000000",
  6094=>"000010101",
  6095=>"011100010",
  6096=>"111110101",
  6097=>"011011001",
  6098=>"010010100",
  6099=>"010010111",
  6100=>"100110100",
  6101=>"010000001",
  6102=>"000101101",
  6103=>"101000000",
  6104=>"010000000",
  6105=>"111001011",
  6106=>"010111011",
  6107=>"001001110",
  6108=>"100110110",
  6109=>"010000101",
  6110=>"111111110",
  6111=>"111001001",
  6112=>"010100001",
  6113=>"111000100",
  6114=>"110101101",
  6115=>"100001110",
  6116=>"010000000",
  6117=>"010101100",
  6118=>"000110000",
  6119=>"111000001",
  6120=>"010011000",
  6121=>"010010110",
  6122=>"110010010",
  6123=>"001101011",
  6124=>"111101000",
  6125=>"110011110",
  6126=>"100000001",
  6127=>"101000110",
  6128=>"000100000",
  6129=>"011110011",
  6130=>"101111110",
  6131=>"010000110",
  6132=>"011000001",
  6133=>"001101111",
  6134=>"011110111",
  6135=>"011000001",
  6136=>"011010010",
  6137=>"100101010",
  6138=>"110000110",
  6139=>"001100010",
  6140=>"011110000",
  6141=>"110101010",
  6142=>"010110101",
  6143=>"110100100",
  6144=>"000110010",
  6145=>"100101010",
  6146=>"001100000",
  6147=>"000001101",
  6148=>"000010110",
  6149=>"010100011",
  6150=>"110000100",
  6151=>"001001111",
  6152=>"011100001",
  6153=>"110000110",
  6154=>"101011101",
  6155=>"110000010",
  6156=>"110011110",
  6157=>"101110110",
  6158=>"011100010",
  6159=>"110100111",
  6160=>"111010000",
  6161=>"011100010",
  6162=>"001111100",
  6163=>"000110001",
  6164=>"000110000",
  6165=>"000111100",
  6166=>"100100100",
  6167=>"110010011",
  6168=>"100010000",
  6169=>"101011000",
  6170=>"100101111",
  6171=>"001011010",
  6172=>"101101001",
  6173=>"011010110",
  6174=>"000010101",
  6175=>"111111000",
  6176=>"010001101",
  6177=>"000111111",
  6178=>"011000010",
  6179=>"101111011",
  6180=>"110010100",
  6181=>"010111110",
  6182=>"111010110",
  6183=>"011101010",
  6184=>"101111100",
  6185=>"010101111",
  6186=>"100000101",
  6187=>"111000001",
  6188=>"110001000",
  6189=>"111010111",
  6190=>"110101000",
  6191=>"100101110",
  6192=>"001110110",
  6193=>"001110111",
  6194=>"110111110",
  6195=>"001010100",
  6196=>"101101001",
  6197=>"010110101",
  6198=>"110111110",
  6199=>"101000011",
  6200=>"001110001",
  6201=>"001001000",
  6202=>"101011011",
  6203=>"101000000",
  6204=>"000000000",
  6205=>"111011100",
  6206=>"100111110",
  6207=>"010101010",
  6208=>"111011100",
  6209=>"101010111",
  6210=>"011000111",
  6211=>"001010100",
  6212=>"001011011",
  6213=>"111100110",
  6214=>"000100010",
  6215=>"110010101",
  6216=>"011111010",
  6217=>"011100100",
  6218=>"110101001",
  6219=>"011011010",
  6220=>"100101101",
  6221=>"111010000",
  6222=>"101010010",
  6223=>"111110011",
  6224=>"101100100",
  6225=>"011110001",
  6226=>"111001100",
  6227=>"101100010",
  6228=>"111011111",
  6229=>"011010101",
  6230=>"111010000",
  6231=>"000101011",
  6232=>"111011111",
  6233=>"011110111",
  6234=>"010011100",
  6235=>"001100101",
  6236=>"100000111",
  6237=>"000010001",
  6238=>"110000001",
  6239=>"000011100",
  6240=>"010100100",
  6241=>"101100111",
  6242=>"111111001",
  6243=>"101101101",
  6244=>"100100000",
  6245=>"110101101",
  6246=>"111001111",
  6247=>"000000111",
  6248=>"011111001",
  6249=>"100011001",
  6250=>"110001001",
  6251=>"101000001",
  6252=>"001000001",
  6253=>"101101001",
  6254=>"000100000",
  6255=>"000011101",
  6256=>"010001010",
  6257=>"010111111",
  6258=>"110111000",
  6259=>"011100000",
  6260=>"001001111",
  6261=>"011011001",
  6262=>"111011001",
  6263=>"011110100",
  6264=>"110010001",
  6265=>"101100111",
  6266=>"010000010",
  6267=>"010101101",
  6268=>"101100001",
  6269=>"111111000",
  6270=>"001000010",
  6271=>"001000001",
  6272=>"101000100",
  6273=>"110100111",
  6274=>"001110100",
  6275=>"010111100",
  6276=>"101010010",
  6277=>"111010110",
  6278=>"010000011",
  6279=>"010111111",
  6280=>"110001011",
  6281=>"000010111",
  6282=>"011010001",
  6283=>"110010111",
  6284=>"010010101",
  6285=>"001000001",
  6286=>"100110101",
  6287=>"010100100",
  6288=>"110111010",
  6289=>"011001111",
  6290=>"110111010",
  6291=>"001001111",
  6292=>"001111010",
  6293=>"001001001",
  6294=>"010001111",
  6295=>"101101000",
  6296=>"000001010",
  6297=>"110110101",
  6298=>"010111100",
  6299=>"110110011",
  6300=>"011010110",
  6301=>"100111111",
  6302=>"000001000",
  6303=>"011111111",
  6304=>"100101010",
  6305=>"000001000",
  6306=>"000001001",
  6307=>"010011110",
  6308=>"010101011",
  6309=>"100011001",
  6310=>"010101010",
  6311=>"000111100",
  6312=>"011000001",
  6313=>"010000000",
  6314=>"101110000",
  6315=>"010000001",
  6316=>"100010111",
  6317=>"101111111",
  6318=>"000000101",
  6319=>"100110101",
  6320=>"011111000",
  6321=>"000000110",
  6322=>"010010000",
  6323=>"000000111",
  6324=>"100101110",
  6325=>"010001001",
  6326=>"110000111",
  6327=>"000010010",
  6328=>"101100100",
  6329=>"111111111",
  6330=>"100011000",
  6331=>"110000101",
  6332=>"010010000",
  6333=>"011100101",
  6334=>"111000011",
  6335=>"111011100",
  6336=>"100111101",
  6337=>"101011011",
  6338=>"111011110",
  6339=>"000111110",
  6340=>"101010000",
  6341=>"110110111",
  6342=>"100111001",
  6343=>"100000110",
  6344=>"111101010",
  6345=>"001011111",
  6346=>"011111110",
  6347=>"010111000",
  6348=>"100000010",
  6349=>"001110111",
  6350=>"011110110",
  6351=>"101010000",
  6352=>"010001010",
  6353=>"010011110",
  6354=>"100010000",
  6355=>"101101001",
  6356=>"100111011",
  6357=>"100000110",
  6358=>"000011010",
  6359=>"011111010",
  6360=>"111001010",
  6361=>"101100010",
  6362=>"001001101",
  6363=>"010011010",
  6364=>"101010010",
  6365=>"011000111",
  6366=>"000110011",
  6367=>"011010111",
  6368=>"000100011",
  6369=>"100010111",
  6370=>"111111101",
  6371=>"111101100",
  6372=>"111010011",
  6373=>"010000000",
  6374=>"001101110",
  6375=>"000010011",
  6376=>"001000011",
  6377=>"000111011",
  6378=>"101101001",
  6379=>"001011101",
  6380=>"001010001",
  6381=>"010111011",
  6382=>"000111111",
  6383=>"111111010",
  6384=>"001001000",
  6385=>"011110010",
  6386=>"100011111",
  6387=>"001011010",
  6388=>"100001001",
  6389=>"000001111",
  6390=>"110011100",
  6391=>"101100010",
  6392=>"010001011",
  6393=>"111100110",
  6394=>"110101101",
  6395=>"100000100",
  6396=>"011000100",
  6397=>"001010001",
  6398=>"001010000",
  6399=>"100111010",
  6400=>"110101110",
  6401=>"101101101",
  6402=>"011000111",
  6403=>"011011111",
  6404=>"010010100",
  6405=>"011111101",
  6406=>"100110101",
  6407=>"011110110",
  6408=>"011110010",
  6409=>"110011101",
  6410=>"000001101",
  6411=>"001101011",
  6412=>"011111011",
  6413=>"011011000",
  6414=>"000110101",
  6415=>"000110011",
  6416=>"011101000",
  6417=>"000100000",
  6418=>"000011001",
  6419=>"000000110",
  6420=>"100111100",
  6421=>"011001100",
  6422=>"000111001",
  6423=>"011100000",
  6424=>"000010100",
  6425=>"100111000",
  6426=>"111100111",
  6427=>"100001000",
  6428=>"111101110",
  6429=>"101011110",
  6430=>"100100100",
  6431=>"111110100",
  6432=>"000010111",
  6433=>"111000101",
  6434=>"110011000",
  6435=>"011101110",
  6436=>"111100111",
  6437=>"101101100",
  6438=>"001101011",
  6439=>"110100101",
  6440=>"010011101",
  6441=>"101110001",
  6442=>"011110011",
  6443=>"000110011",
  6444=>"110000001",
  6445=>"110000011",
  6446=>"010001110",
  6447=>"010001010",
  6448=>"101010101",
  6449=>"000100000",
  6450=>"000100111",
  6451=>"000101010",
  6452=>"011100001",
  6453=>"101001011",
  6454=>"010101010",
  6455=>"000110110",
  6456=>"111111110",
  6457=>"110101010",
  6458=>"000101100",
  6459=>"011111101",
  6460=>"110010110",
  6461=>"010111111",
  6462=>"011011101",
  6463=>"011010011",
  6464=>"100111100",
  6465=>"100101111",
  6466=>"111011011",
  6467=>"000001100",
  6468=>"000000101",
  6469=>"000011101",
  6470=>"000111110",
  6471=>"000010101",
  6472=>"010101000",
  6473=>"000111001",
  6474=>"101010000",
  6475=>"110100100",
  6476=>"001111100",
  6477=>"000001000",
  6478=>"010001110",
  6479=>"010000111",
  6480=>"011010000",
  6481=>"000101110",
  6482=>"000101001",
  6483=>"011100110",
  6484=>"010001100",
  6485=>"111100011",
  6486=>"110110000",
  6487=>"111110001",
  6488=>"111111101",
  6489=>"101000101",
  6490=>"011000000",
  6491=>"000000010",
  6492=>"100001001",
  6493=>"000101010",
  6494=>"010100100",
  6495=>"111000111",
  6496=>"010000011",
  6497=>"111101010",
  6498=>"000000111",
  6499=>"000001100",
  6500=>"101100001",
  6501=>"100110000",
  6502=>"101110110",
  6503=>"100101100",
  6504=>"100001000",
  6505=>"111001100",
  6506=>"110001100",
  6507=>"010001111",
  6508=>"000011110",
  6509=>"110010000",
  6510=>"101000001",
  6511=>"101101100",
  6512=>"000101000",
  6513=>"010101101",
  6514=>"111111111",
  6515=>"001110010",
  6516=>"010100001",
  6517=>"111111010",
  6518=>"111000011",
  6519=>"101110011",
  6520=>"001001100",
  6521=>"001101001",
  6522=>"111001101",
  6523=>"011000001",
  6524=>"100011011",
  6525=>"101111101",
  6526=>"101011111",
  6527=>"010110010",
  6528=>"111111001",
  6529=>"000110110",
  6530=>"111011010",
  6531=>"110100101",
  6532=>"110000001",
  6533=>"011001010",
  6534=>"111011110",
  6535=>"000000111",
  6536=>"110001001",
  6537=>"010100010",
  6538=>"001001011",
  6539=>"001000101",
  6540=>"011001111",
  6541=>"100011011",
  6542=>"000000000",
  6543=>"011111001",
  6544=>"010111111",
  6545=>"101000010",
  6546=>"000110010",
  6547=>"100011010",
  6548=>"101000100",
  6549=>"100001001",
  6550=>"011101111",
  6551=>"111011011",
  6552=>"110011101",
  6553=>"000010110",
  6554=>"110000001",
  6555=>"011000111",
  6556=>"001110110",
  6557=>"010110000",
  6558=>"110011000",
  6559=>"111010001",
  6560=>"011011011",
  6561=>"110000010",
  6562=>"010101011",
  6563=>"101011111",
  6564=>"001010111",
  6565=>"100001111",
  6566=>"010100100",
  6567=>"100110000",
  6568=>"111110100",
  6569=>"011011010",
  6570=>"111001001",
  6571=>"010011000",
  6572=>"001100101",
  6573=>"110101011",
  6574=>"001111111",
  6575=>"001111110",
  6576=>"111101111",
  6577=>"100101011",
  6578=>"001101101",
  6579=>"110111000",
  6580=>"001001001",
  6581=>"110010011",
  6582=>"101111110",
  6583=>"110000000",
  6584=>"001010100",
  6585=>"001100111",
  6586=>"000000011",
  6587=>"110111101",
  6588=>"000000001",
  6589=>"111110000",
  6590=>"000010110",
  6591=>"011110101",
  6592=>"011100010",
  6593=>"000010010",
  6594=>"100111100",
  6595=>"111010100",
  6596=>"000010000",
  6597=>"111010111",
  6598=>"101110001",
  6599=>"011011001",
  6600=>"010011000",
  6601=>"011100001",
  6602=>"000111101",
  6603=>"010111010",
  6604=>"110000011",
  6605=>"001010010",
  6606=>"010011010",
  6607=>"010110101",
  6608=>"011111010",
  6609=>"011000000",
  6610=>"000000011",
  6611=>"011100010",
  6612=>"110000000",
  6613=>"010100010",
  6614=>"011001101",
  6615=>"000010100",
  6616=>"101101101",
  6617=>"111111111",
  6618=>"011111111",
  6619=>"100010000",
  6620=>"100111101",
  6621=>"111011110",
  6622=>"100110101",
  6623=>"100100100",
  6624=>"100000000",
  6625=>"110010000",
  6626=>"100001111",
  6627=>"111110000",
  6628=>"110100111",
  6629=>"100101011",
  6630=>"101011000",
  6631=>"111100011",
  6632=>"010001110",
  6633=>"011111110",
  6634=>"000010100",
  6635=>"000010110",
  6636=>"110110111",
  6637=>"110110101",
  6638=>"001001100",
  6639=>"010111100",
  6640=>"001111111",
  6641=>"101101011",
  6642=>"000011000",
  6643=>"101000001",
  6644=>"010110000",
  6645=>"110011101",
  6646=>"100000001",
  6647=>"010111011",
  6648=>"100101011",
  6649=>"101001100",
  6650=>"000001001",
  6651=>"101010000",
  6652=>"111100110",
  6653=>"000000101",
  6654=>"111111101",
  6655=>"110101100",
  6656=>"011010101",
  6657=>"000101100",
  6658=>"111000001",
  6659=>"101000110",
  6660=>"011110111",
  6661=>"000100100",
  6662=>"011111010",
  6663=>"110011111",
  6664=>"101000000",
  6665=>"010000101",
  6666=>"110010011",
  6667=>"000111010",
  6668=>"000100000",
  6669=>"101010111",
  6670=>"100000000",
  6671=>"110111000",
  6672=>"111101001",
  6673=>"101101010",
  6674=>"111011100",
  6675=>"000010010",
  6676=>"011100000",
  6677=>"001110000",
  6678=>"010001110",
  6679=>"100001000",
  6680=>"011000000",
  6681=>"000011100",
  6682=>"010110000",
  6683=>"001110001",
  6684=>"101111110",
  6685=>"100011011",
  6686=>"101001000",
  6687=>"111111000",
  6688=>"101100000",
  6689=>"111100011",
  6690=>"010100010",
  6691=>"101110110",
  6692=>"110111101",
  6693=>"100001100",
  6694=>"011111111",
  6695=>"000011100",
  6696=>"111101100",
  6697=>"101100111",
  6698=>"000011111",
  6699=>"000100010",
  6700=>"001101111",
  6701=>"111111101",
  6702=>"100011110",
  6703=>"111010100",
  6704=>"110101011",
  6705=>"111110111",
  6706=>"100111000",
  6707=>"100010000",
  6708=>"001000011",
  6709=>"010000010",
  6710=>"000010010",
  6711=>"011110000",
  6712=>"000001110",
  6713=>"000000110",
  6714=>"010100010",
  6715=>"010000100",
  6716=>"101000011",
  6717=>"000110000",
  6718=>"110010111",
  6719=>"100100110",
  6720=>"111111111",
  6721=>"011110000",
  6722=>"001010101",
  6723=>"101111000",
  6724=>"011111100",
  6725=>"010010001",
  6726=>"010100000",
  6727=>"100101110",
  6728=>"001011111",
  6729=>"010001110",
  6730=>"111100010",
  6731=>"011101011",
  6732=>"100100111",
  6733=>"101100110",
  6734=>"100111111",
  6735=>"110011101",
  6736=>"000111111",
  6737=>"101001011",
  6738=>"101010100",
  6739=>"111011010",
  6740=>"001110000",
  6741=>"000000110",
  6742=>"111010110",
  6743=>"001100100",
  6744=>"010110101",
  6745=>"010011100",
  6746=>"101111011",
  6747=>"000000111",
  6748=>"000000010",
  6749=>"100100110",
  6750=>"000001100",
  6751=>"011100001",
  6752=>"110011001",
  6753=>"101110011",
  6754=>"011000011",
  6755=>"001001100",
  6756=>"111011011",
  6757=>"001101001",
  6758=>"110101101",
  6759=>"010001110",
  6760=>"000010010",
  6761=>"110011000",
  6762=>"010010000",
  6763=>"011110100",
  6764=>"101001000",
  6765=>"011000101",
  6766=>"111011100",
  6767=>"011000110",
  6768=>"011010000",
  6769=>"000000000",
  6770=>"001111011",
  6771=>"011110010",
  6772=>"110111100",
  6773=>"101101111",
  6774=>"110001111",
  6775=>"010000111",
  6776=>"111100000",
  6777=>"100110101",
  6778=>"110100010",
  6779=>"000011001",
  6780=>"011000111",
  6781=>"111011001",
  6782=>"100111110",
  6783=>"110001011",
  6784=>"001100000",
  6785=>"110101010",
  6786=>"110000010",
  6787=>"111100010",
  6788=>"000101110",
  6789=>"100010000",
  6790=>"110101111",
  6791=>"101001000",
  6792=>"010110110",
  6793=>"010011110",
  6794=>"111110010",
  6795=>"000110111",
  6796=>"110111000",
  6797=>"010001110",
  6798=>"101010000",
  6799=>"111010111",
  6800=>"010100011",
  6801=>"101001100",
  6802=>"000010110",
  6803=>"011011111",
  6804=>"010110110",
  6805=>"011111000",
  6806=>"100111111",
  6807=>"100010011",
  6808=>"001101001",
  6809=>"101001110",
  6810=>"010100000",
  6811=>"111100011",
  6812=>"111010111",
  6813=>"100010000",
  6814=>"000000010",
  6815=>"100110101",
  6816=>"001010110",
  6817=>"111101010",
  6818=>"110100110",
  6819=>"010110111",
  6820=>"101100101",
  6821=>"111100010",
  6822=>"010010011",
  6823=>"000001101",
  6824=>"100111000",
  6825=>"111011101",
  6826=>"000101010",
  6827=>"101101110",
  6828=>"001010110",
  6829=>"010111110",
  6830=>"111010110",
  6831=>"111110101",
  6832=>"010100110",
  6833=>"111101000",
  6834=>"101111111",
  6835=>"111011001",
  6836=>"111100111",
  6837=>"000011110",
  6838=>"101100101",
  6839=>"010011010",
  6840=>"100001111",
  6841=>"010111001",
  6842=>"010011011",
  6843=>"010000110",
  6844=>"011010000",
  6845=>"001010011",
  6846=>"001101110",
  6847=>"001101111",
  6848=>"111000101",
  6849=>"000010101",
  6850=>"001010000",
  6851=>"111111011",
  6852=>"010101100",
  6853=>"111100001",
  6854=>"110110101",
  6855=>"000100000",
  6856=>"111111111",
  6857=>"111110010",
  6858=>"001101000",
  6859=>"000010110",
  6860=>"000011110",
  6861=>"111110000",
  6862=>"011111010",
  6863=>"001110101",
  6864=>"110000011",
  6865=>"001001010",
  6866=>"111000011",
  6867=>"010110000",
  6868=>"110010100",
  6869=>"010000000",
  6870=>"000000000",
  6871=>"010001111",
  6872=>"010101110",
  6873=>"010001000",
  6874=>"100110001",
  6875=>"001000011",
  6876=>"000010100",
  6877=>"010000111",
  6878=>"011101001",
  6879=>"011011001",
  6880=>"011011101",
  6881=>"100100000",
  6882=>"100111111",
  6883=>"101101010",
  6884=>"011100001",
  6885=>"011000000",
  6886=>"100000000",
  6887=>"001010001",
  6888=>"010010000",
  6889=>"011010110",
  6890=>"100010010",
  6891=>"101011110",
  6892=>"010100011",
  6893=>"001100001",
  6894=>"101100011",
  6895=>"111001111",
  6896=>"110101111",
  6897=>"111100010",
  6898=>"001011011",
  6899=>"100000101",
  6900=>"011011000",
  6901=>"111110110",
  6902=>"101110001",
  6903=>"111100001",
  6904=>"000011010",
  6905=>"100110001",
  6906=>"000010110",
  6907=>"011001001",
  6908=>"010101100",
  6909=>"011001011",
  6910=>"010000000",
  6911=>"011100010",
  6912=>"101010010",
  6913=>"111011101",
  6914=>"010011000",
  6915=>"011111110",
  6916=>"011010000",
  6917=>"100111111",
  6918=>"110101110",
  6919=>"010010111",
  6920=>"010011010",
  6921=>"100111100",
  6922=>"010011000",
  6923=>"101111111",
  6924=>"110110100",
  6925=>"111100010",
  6926=>"111101110",
  6927=>"010000011",
  6928=>"111101111",
  6929=>"001110011",
  6930=>"000110100",
  6931=>"101010110",
  6932=>"000000100",
  6933=>"100110100",
  6934=>"110011101",
  6935=>"000111010",
  6936=>"110000010",
  6937=>"110110010",
  6938=>"000000010",
  6939=>"001000001",
  6940=>"111100100",
  6941=>"001010000",
  6942=>"000011011",
  6943=>"000111100",
  6944=>"100111101",
  6945=>"011110001",
  6946=>"101011100",
  6947=>"101110011",
  6948=>"111111000",
  6949=>"000001010",
  6950=>"001111001",
  6951=>"101100010",
  6952=>"011100000",
  6953=>"000110010",
  6954=>"000001111",
  6955=>"001111001",
  6956=>"110001011",
  6957=>"100100000",
  6958=>"110101111",
  6959=>"000111000",
  6960=>"101000111",
  6961=>"010111001",
  6962=>"011111111",
  6963=>"101110110",
  6964=>"011111111",
  6965=>"111001111",
  6966=>"101001111",
  6967=>"110110100",
  6968=>"101111101",
  6969=>"111001101",
  6970=>"011110110",
  6971=>"001111111",
  6972=>"001000101",
  6973=>"110100000",
  6974=>"110111111",
  6975=>"100011111",
  6976=>"000001000",
  6977=>"010101001",
  6978=>"010000011",
  6979=>"111100101",
  6980=>"001111010",
  6981=>"010010110",
  6982=>"011110011",
  6983=>"111000100",
  6984=>"111111110",
  6985=>"110010010",
  6986=>"010001011",
  6987=>"000011000",
  6988=>"100001101",
  6989=>"111001000",
  6990=>"111111001",
  6991=>"001010010",
  6992=>"100000101",
  6993=>"100101001",
  6994=>"000111000",
  6995=>"111000100",
  6996=>"100011110",
  6997=>"100000100",
  6998=>"010110111",
  6999=>"101110000",
  7000=>"011001000",
  7001=>"000110001",
  7002=>"111001101",
  7003=>"101100100",
  7004=>"101110001",
  7005=>"011010101",
  7006=>"110010011",
  7007=>"000000001",
  7008=>"101010000",
  7009=>"010000011",
  7010=>"111100000",
  7011=>"111010001",
  7012=>"001000011",
  7013=>"100100001",
  7014=>"010100101",
  7015=>"111110101",
  7016=>"100000000",
  7017=>"011101101",
  7018=>"010111101",
  7019=>"111110110",
  7020=>"111100000",
  7021=>"011010110",
  7022=>"000100101",
  7023=>"110001011",
  7024=>"100011100",
  7025=>"010101100",
  7026=>"010110010",
  7027=>"000110001",
  7028=>"001100101",
  7029=>"000000101",
  7030=>"001001001",
  7031=>"001001000",
  7032=>"100110010",
  7033=>"100101000",
  7034=>"011101000",
  7035=>"011011100",
  7036=>"011001000",
  7037=>"110011110",
  7038=>"001100111",
  7039=>"110010001",
  7040=>"011100100",
  7041=>"111101000",
  7042=>"110110101",
  7043=>"101011010",
  7044=>"111101001",
  7045=>"110100010",
  7046=>"010110000",
  7047=>"001111011",
  7048=>"100111111",
  7049=>"011111010",
  7050=>"110101101",
  7051=>"000001001",
  7052=>"000001110",
  7053=>"011011110",
  7054=>"110001101",
  7055=>"110000000",
  7056=>"110010111",
  7057=>"100111101",
  7058=>"000000010",
  7059=>"101000000",
  7060=>"101111111",
  7061=>"111111001",
  7062=>"011101001",
  7063=>"100000010",
  7064=>"001110010",
  7065=>"000011010",
  7066=>"100101111",
  7067=>"010010100",
  7068=>"011010100",
  7069=>"101110110",
  7070=>"010011010",
  7071=>"110110000",
  7072=>"000001001",
  7073=>"111111111",
  7074=>"100011011",
  7075=>"011110000",
  7076=>"100011110",
  7077=>"110010001",
  7078=>"000000001",
  7079=>"100100010",
  7080=>"010010111",
  7081=>"011000000",
  7082=>"110010010",
  7083=>"100101111",
  7084=>"110100011",
  7085=>"100110101",
  7086=>"011111001",
  7087=>"011010101",
  7088=>"101010111",
  7089=>"110011000",
  7090=>"101101000",
  7091=>"101001011",
  7092=>"000010000",
  7093=>"101011010",
  7094=>"011101000",
  7095=>"010111100",
  7096=>"100101110",
  7097=>"110111001",
  7098=>"010010011",
  7099=>"000110100",
  7100=>"011000111",
  7101=>"000111001",
  7102=>"000010000",
  7103=>"111111001",
  7104=>"011010000",
  7105=>"010110100",
  7106=>"001010101",
  7107=>"111111000",
  7108=>"010000010",
  7109=>"111111011",
  7110=>"010001010",
  7111=>"011111011",
  7112=>"001001111",
  7113=>"100000000",
  7114=>"111000110",
  7115=>"110000101",
  7116=>"101000110",
  7117=>"100000100",
  7118=>"111111010",
  7119=>"001001010",
  7120=>"000110010",
  7121=>"110100111",
  7122=>"001110011",
  7123=>"001010000",
  7124=>"010000100",
  7125=>"110111000",
  7126=>"001010101",
  7127=>"110110011",
  7128=>"011101100",
  7129=>"000011001",
  7130=>"111110101",
  7131=>"001010100",
  7132=>"101100010",
  7133=>"000110101",
  7134=>"100100001",
  7135=>"100100001",
  7136=>"111111100",
  7137=>"110011110",
  7138=>"110110100",
  7139=>"100010101",
  7140=>"000110001",
  7141=>"010001101",
  7142=>"101000010",
  7143=>"101111001",
  7144=>"011111100",
  7145=>"111110110",
  7146=>"101100010",
  7147=>"011110111",
  7148=>"000101111",
  7149=>"111100100",
  7150=>"010010111",
  7151=>"101100111",
  7152=>"101111110",
  7153=>"110011001",
  7154=>"001001100",
  7155=>"001110010",
  7156=>"011001110",
  7157=>"111001110",
  7158=>"000010000",
  7159=>"000111100",
  7160=>"111001011",
  7161=>"010001000",
  7162=>"101010001",
  7163=>"000111000",
  7164=>"100101001",
  7165=>"111011110",
  7166=>"111100110",
  7167=>"100101110",
  7168=>"101001010",
  7169=>"111001101",
  7170=>"001010000",
  7171=>"010101100",
  7172=>"000101000",
  7173=>"001101100",
  7174=>"110001000",
  7175=>"000101101",
  7176=>"110010010",
  7177=>"000010110",
  7178=>"101101010",
  7179=>"110110011",
  7180=>"001000010",
  7181=>"111001100",
  7182=>"100001000",
  7183=>"001000010",
  7184=>"100111110",
  7185=>"010101111",
  7186=>"101010000",
  7187=>"010000100",
  7188=>"111111111",
  7189=>"100100100",
  7190=>"110010101",
  7191=>"011001001",
  7192=>"001000101",
  7193=>"010001100",
  7194=>"011100000",
  7195=>"010101110",
  7196=>"000100100",
  7197=>"110010100",
  7198=>"111110010",
  7199=>"001000111",
  7200=>"011001001",
  7201=>"111000000",
  7202=>"111111111",
  7203=>"101101010",
  7204=>"001110010",
  7205=>"011000001",
  7206=>"101100111",
  7207=>"101101101",
  7208=>"111010111",
  7209=>"110100000",
  7210=>"000010010",
  7211=>"000101000",
  7212=>"101001111",
  7213=>"000101111",
  7214=>"000101100",
  7215=>"101010001",
  7216=>"110100000",
  7217=>"101111111",
  7218=>"110110100",
  7219=>"100011100",
  7220=>"001101111",
  7221=>"101100100",
  7222=>"010011000",
  7223=>"010100011",
  7224=>"010000101",
  7225=>"001101010",
  7226=>"110000000",
  7227=>"010010001",
  7228=>"001001100",
  7229=>"001101000",
  7230=>"010101001",
  7231=>"010010110",
  7232=>"110101101",
  7233=>"000000010",
  7234=>"010000011",
  7235=>"101011000",
  7236=>"100100110",
  7237=>"100100011",
  7238=>"000001000",
  7239=>"010010101",
  7240=>"110010111",
  7241=>"110100101",
  7242=>"001100010",
  7243=>"000100001",
  7244=>"010110010",
  7245=>"000010110",
  7246=>"010000100",
  7247=>"101000100",
  7248=>"100011001",
  7249=>"111101111",
  7250=>"001000001",
  7251=>"101100110",
  7252=>"010100001",
  7253=>"000010001",
  7254=>"010101111",
  7255=>"000111100",
  7256=>"010110010",
  7257=>"101000100",
  7258=>"010111000",
  7259=>"101001000",
  7260=>"001011100",
  7261=>"100000100",
  7262=>"000111100",
  7263=>"010000011",
  7264=>"110100111",
  7265=>"001010101",
  7266=>"100101111",
  7267=>"100101011",
  7268=>"010010011",
  7269=>"010011000",
  7270=>"110110011",
  7271=>"111100101",
  7272=>"001011110",
  7273=>"000000011",
  7274=>"000010110",
  7275=>"101110111",
  7276=>"101101001",
  7277=>"011100001",
  7278=>"111011111",
  7279=>"000011000",
  7280=>"011111110",
  7281=>"001011100",
  7282=>"111100101",
  7283=>"011000111",
  7284=>"001111011",
  7285=>"111010100",
  7286=>"010100111",
  7287=>"111111110",
  7288=>"010110111",
  7289=>"011011110",
  7290=>"101100110",
  7291=>"101101001",
  7292=>"011101110",
  7293=>"100100011",
  7294=>"011111101",
  7295=>"001100000",
  7296=>"100010111",
  7297=>"000101110",
  7298=>"000110001",
  7299=>"011110001",
  7300=>"111011110",
  7301=>"111110101",
  7302=>"111001001",
  7303=>"101011101",
  7304=>"111101111",
  7305=>"001100111",
  7306=>"001110110",
  7307=>"000001101",
  7308=>"000001100",
  7309=>"001111110",
  7310=>"110001000",
  7311=>"011000110",
  7312=>"111011001",
  7313=>"001110100",
  7314=>"100110111",
  7315=>"111000110",
  7316=>"000000010",
  7317=>"011101001",
  7318=>"111110010",
  7319=>"100100010",
  7320=>"110100010",
  7321=>"000110001",
  7322=>"110010101",
  7323=>"101111001",
  7324=>"000111011",
  7325=>"101010000",
  7326=>"101011011",
  7327=>"101111000",
  7328=>"110100011",
  7329=>"100011001",
  7330=>"010100111",
  7331=>"010111010",
  7332=>"111001111",
  7333=>"001000000",
  7334=>"010001111",
  7335=>"000110110",
  7336=>"000000001",
  7337=>"111101000",
  7338=>"101010101",
  7339=>"001010010",
  7340=>"100011001",
  7341=>"000000010",
  7342=>"011111101",
  7343=>"100110000",
  7344=>"011000101",
  7345=>"010011111",
  7346=>"001110010",
  7347=>"111101001",
  7348=>"011010110",
  7349=>"111111111",
  7350=>"110000110",
  7351=>"000100111",
  7352=>"001000010",
  7353=>"010111010",
  7354=>"010110010",
  7355=>"101100011",
  7356=>"111010000",
  7357=>"010100111",
  7358=>"001010000",
  7359=>"110111111",
  7360=>"000110001",
  7361=>"000010111",
  7362=>"010101100",
  7363=>"110010011",
  7364=>"100001000",
  7365=>"011011000",
  7366=>"101110100",
  7367=>"011010100",
  7368=>"001010001",
  7369=>"110010111",
  7370=>"001010000",
  7371=>"010101000",
  7372=>"001000010",
  7373=>"001001000",
  7374=>"011111111",
  7375=>"100001101",
  7376=>"000011011",
  7377=>"110001111",
  7378=>"010100000",
  7379=>"101101110",
  7380=>"011100001",
  7381=>"001110011",
  7382=>"011110100",
  7383=>"011110011",
  7384=>"010101001",
  7385=>"000111111",
  7386=>"010010000",
  7387=>"111101001",
  7388=>"111110111",
  7389=>"010111011",
  7390=>"011110000",
  7391=>"001011101",
  7392=>"011100111",
  7393=>"101110111",
  7394=>"111001101",
  7395=>"000000010",
  7396=>"110111010",
  7397=>"101111100",
  7398=>"100010101",
  7399=>"011111100",
  7400=>"100110100",
  7401=>"100110000",
  7402=>"111000110",
  7403=>"000101011",
  7404=>"010111100",
  7405=>"000011111",
  7406=>"110100100",
  7407=>"000111000",
  7408=>"010011010",
  7409=>"100110111",
  7410=>"010001011",
  7411=>"010110001",
  7412=>"111011011",
  7413=>"010100001",
  7414=>"010110000",
  7415=>"000001010",
  7416=>"110100001",
  7417=>"111110010",
  7418=>"001111011",
  7419=>"000000011",
  7420=>"010101111",
  7421=>"100000100",
  7422=>"010010100",
  7423=>"000011010",
  7424=>"000100000",
  7425=>"001010010",
  7426=>"111110011",
  7427=>"111011010",
  7428=>"000000101",
  7429=>"011001110",
  7430=>"111111010",
  7431=>"000001111",
  7432=>"010011101",
  7433=>"000011011",
  7434=>"000111001",
  7435=>"111010110",
  7436=>"010010100",
  7437=>"010110010",
  7438=>"110111111",
  7439=>"000111001",
  7440=>"100111011",
  7441=>"010011111",
  7442=>"000000001",
  7443=>"101111110",
  7444=>"111001011",
  7445=>"001110101",
  7446=>"010110100",
  7447=>"001111100",
  7448=>"000001011",
  7449=>"000010000",
  7450=>"111001101",
  7451=>"111101110",
  7452=>"101100011",
  7453=>"100001001",
  7454=>"101001111",
  7455=>"010010001",
  7456=>"010101010",
  7457=>"000101111",
  7458=>"111101100",
  7459=>"001001110",
  7460=>"011001100",
  7461=>"110000010",
  7462=>"111000001",
  7463=>"010000010",
  7464=>"110010010",
  7465=>"100010111",
  7466=>"011111110",
  7467=>"111011000",
  7468=>"000100001",
  7469=>"100001100",
  7470=>"100101001",
  7471=>"011100101",
  7472=>"011000101",
  7473=>"011110110",
  7474=>"000000000",
  7475=>"001100110",
  7476=>"110000011",
  7477=>"001001110",
  7478=>"111011111",
  7479=>"000010001",
  7480=>"000011100",
  7481=>"110010100",
  7482=>"101101100",
  7483=>"011101011",
  7484=>"101000110",
  7485=>"101111001",
  7486=>"000101000",
  7487=>"100001101",
  7488=>"110101010",
  7489=>"101101011",
  7490=>"010010101",
  7491=>"101111000",
  7492=>"101101111",
  7493=>"001110000",
  7494=>"111011001",
  7495=>"111100011",
  7496=>"001010110",
  7497=>"010001011",
  7498=>"010011011",
  7499=>"000000001",
  7500=>"001011001",
  7501=>"001011010",
  7502=>"000110001",
  7503=>"100101010",
  7504=>"100100011",
  7505=>"111010110",
  7506=>"000000111",
  7507=>"010011000",
  7508=>"101001010",
  7509=>"000001001",
  7510=>"110000101",
  7511=>"011100000",
  7512=>"100010111",
  7513=>"000100000",
  7514=>"011110110",
  7515=>"001110101",
  7516=>"011010010",
  7517=>"111011111",
  7518=>"110010111",
  7519=>"000111111",
  7520=>"000011011",
  7521=>"111000010",
  7522=>"010010011",
  7523=>"100010100",
  7524=>"110111011",
  7525=>"100000000",
  7526=>"110111101",
  7527=>"111111110",
  7528=>"100110001",
  7529=>"010111001",
  7530=>"101111000",
  7531=>"011111001",
  7532=>"100010011",
  7533=>"110100001",
  7534=>"011110000",
  7535=>"011010111",
  7536=>"001111110",
  7537=>"001111111",
  7538=>"011001110",
  7539=>"000101110",
  7540=>"011110000",
  7541=>"101101010",
  7542=>"000101001",
  7543=>"101111100",
  7544=>"010010000",
  7545=>"101110111",
  7546=>"010101000",
  7547=>"111001010",
  7548=>"001110111",
  7549=>"111110001",
  7550=>"100101100",
  7551=>"001110001",
  7552=>"000001100",
  7553=>"101010010",
  7554=>"000000111",
  7555=>"100101011",
  7556=>"011100110",
  7557=>"011010111",
  7558=>"011011010",
  7559=>"111010000",
  7560=>"110101100",
  7561=>"110100011",
  7562=>"010000001",
  7563=>"111111101",
  7564=>"001001110",
  7565=>"101000110",
  7566=>"110100001",
  7567=>"110110100",
  7568=>"100110110",
  7569=>"000000100",
  7570=>"110101100",
  7571=>"011111001",
  7572=>"000111111",
  7573=>"011010001",
  7574=>"001000000",
  7575=>"101011000",
  7576=>"100011001",
  7577=>"001010001",
  7578=>"111100011",
  7579=>"110010100",
  7580=>"111000010",
  7581=>"010100100",
  7582=>"101001001",
  7583=>"110011110",
  7584=>"011000111",
  7585=>"110000011",
  7586=>"001101100",
  7587=>"100100000",
  7588=>"110011100",
  7589=>"100000001",
  7590=>"100010010",
  7591=>"100110110",
  7592=>"110100011",
  7593=>"001110000",
  7594=>"011111111",
  7595=>"000111110",
  7596=>"010110111",
  7597=>"110100000",
  7598=>"001111101",
  7599=>"110000010",
  7600=>"111111011",
  7601=>"100100000",
  7602=>"000000000",
  7603=>"000111001",
  7604=>"000100001",
  7605=>"111100010",
  7606=>"000011001",
  7607=>"011110010",
  7608=>"100010110",
  7609=>"010100001",
  7610=>"001111110",
  7611=>"100100010",
  7612=>"001110111",
  7613=>"100101000",
  7614=>"111001111",
  7615=>"010001001",
  7616=>"000011001",
  7617=>"110001101",
  7618=>"100110011",
  7619=>"000110010",
  7620=>"110111111",
  7621=>"110010100",
  7622=>"111100111",
  7623=>"010010000",
  7624=>"101011001",
  7625=>"110100010",
  7626=>"111011110",
  7627=>"011001001",
  7628=>"010100111",
  7629=>"100101010",
  7630=>"000001110",
  7631=>"101100011",
  7632=>"100010011",
  7633=>"001000101",
  7634=>"111001100",
  7635=>"000100000",
  7636=>"110110011",
  7637=>"001110111",
  7638=>"011110110",
  7639=>"010100111",
  7640=>"110010101",
  7641=>"001100000",
  7642=>"001010100",
  7643=>"000110000",
  7644=>"000000001",
  7645=>"010101010",
  7646=>"001100100",
  7647=>"110100111",
  7648=>"000110100",
  7649=>"111001111",
  7650=>"111000000",
  7651=>"000111101",
  7652=>"110001101",
  7653=>"000000100",
  7654=>"110011110",
  7655=>"000100101",
  7656=>"101000101",
  7657=>"001101010",
  7658=>"100111001",
  7659=>"000110101",
  7660=>"100010001",
  7661=>"100011010",
  7662=>"011001011",
  7663=>"111110001",
  7664=>"010001010",
  7665=>"100100001",
  7666=>"000110111",
  7667=>"011000101",
  7668=>"010111011",
  7669=>"011110000",
  7670=>"001111010",
  7671=>"100110111",
  7672=>"110101011",
  7673=>"101100000",
  7674=>"001000111",
  7675=>"100000111",
  7676=>"000110101",
  7677=>"111110101",
  7678=>"110111001",
  7679=>"111001010",
  7680=>"111110001",
  7681=>"011111000",
  7682=>"100110010",
  7683=>"110001110",
  7684=>"111101100",
  7685=>"111001111",
  7686=>"111011001",
  7687=>"011111001",
  7688=>"101100010",
  7689=>"111011111",
  7690=>"101101110",
  7691=>"011001000",
  7692=>"011001011",
  7693=>"100111011",
  7694=>"010100100",
  7695=>"001010101",
  7696=>"000101010",
  7697=>"010111011",
  7698=>"000111001",
  7699=>"101011101",
  7700=>"011111111",
  7701=>"110100110",
  7702=>"111011100",
  7703=>"001000001",
  7704=>"100010011",
  7705=>"111001001",
  7706=>"111101111",
  7707=>"111110101",
  7708=>"011100010",
  7709=>"011111111",
  7710=>"101010010",
  7711=>"010000111",
  7712=>"101000100",
  7713=>"011010111",
  7714=>"010110010",
  7715=>"000001110",
  7716=>"001100011",
  7717=>"111000100",
  7718=>"100011111",
  7719=>"110111000",
  7720=>"001101001",
  7721=>"110011000",
  7722=>"100111001",
  7723=>"101111111",
  7724=>"001011001",
  7725=>"101011111",
  7726=>"010000000",
  7727=>"111111001",
  7728=>"001100100",
  7729=>"101011110",
  7730=>"000001111",
  7731=>"100111111",
  7732=>"100110010",
  7733=>"010011000",
  7734=>"000000010",
  7735=>"111100111",
  7736=>"001010110",
  7737=>"001011001",
  7738=>"011010000",
  7739=>"000111100",
  7740=>"010000001",
  7741=>"110100101",
  7742=>"001000001",
  7743=>"001101010",
  7744=>"111010100",
  7745=>"101010011",
  7746=>"000100110",
  7747=>"000111001",
  7748=>"110000001",
  7749=>"011010010",
  7750=>"000111100",
  7751=>"001010001",
  7752=>"100001001",
  7753=>"010111011",
  7754=>"101000110",
  7755=>"110001010",
  7756=>"011100101",
  7757=>"000100101",
  7758=>"011011111",
  7759=>"011001001",
  7760=>"101010010",
  7761=>"111110000",
  7762=>"111101001",
  7763=>"011101111",
  7764=>"110000100",
  7765=>"000100000",
  7766=>"010010011",
  7767=>"000000011",
  7768=>"111110000",
  7769=>"111101011",
  7770=>"100100011",
  7771=>"110100101",
  7772=>"000011001",
  7773=>"000000010",
  7774=>"000101000",
  7775=>"010000010",
  7776=>"001000110",
  7777=>"110010011",
  7778=>"011001110",
  7779=>"001011011",
  7780=>"111111100",
  7781=>"111011001",
  7782=>"011011000",
  7783=>"010101000",
  7784=>"100010110",
  7785=>"101100010",
  7786=>"011011100",
  7787=>"000110010",
  7788=>"111101010",
  7789=>"111011000",
  7790=>"101110011",
  7791=>"100101111",
  7792=>"000110100",
  7793=>"000010110",
  7794=>"000110111",
  7795=>"100000100",
  7796=>"000111101",
  7797=>"111001011",
  7798=>"110010011",
  7799=>"110000011",
  7800=>"011101101",
  7801=>"001111001",
  7802=>"001101101",
  7803=>"000001001",
  7804=>"110101000",
  7805=>"001001100",
  7806=>"100001001",
  7807=>"010101100",
  7808=>"110110001",
  7809=>"011101011",
  7810=>"110111011",
  7811=>"011001001",
  7812=>"101010111",
  7813=>"000000100",
  7814=>"110001110",
  7815=>"010010011",
  7816=>"010001110",
  7817=>"111010000",
  7818=>"010000001",
  7819=>"111101001",
  7820=>"101000011",
  7821=>"001110000",
  7822=>"111011001",
  7823=>"111110110",
  7824=>"011101100",
  7825=>"101011101",
  7826=>"111000101",
  7827=>"001001001",
  7828=>"010001100",
  7829=>"100111110",
  7830=>"001011100",
  7831=>"000001000",
  7832=>"101010010",
  7833=>"111110000",
  7834=>"000011101",
  7835=>"010110110",
  7836=>"000001100",
  7837=>"001100010",
  7838=>"100000001",
  7839=>"010011100",
  7840=>"111010011",
  7841=>"111111010",
  7842=>"001001111",
  7843=>"011100000",
  7844=>"110101110",
  7845=>"110010100",
  7846=>"010101010",
  7847=>"101000000",
  7848=>"011100100",
  7849=>"100110000",
  7850=>"110111011",
  7851=>"001100011",
  7852=>"100000101",
  7853=>"001011010",
  7854=>"110100011",
  7855=>"011110110",
  7856=>"011110001",
  7857=>"111111001",
  7858=>"100100000",
  7859=>"100001001",
  7860=>"001010100",
  7861=>"111010101",
  7862=>"010000101",
  7863=>"100011000",
  7864=>"101111010",
  7865=>"101010000",
  7866=>"100011110",
  7867=>"101111100",
  7868=>"011000100",
  7869=>"010101110",
  7870=>"010100011",
  7871=>"100000110",
  7872=>"010111000",
  7873=>"110111011",
  7874=>"010011010",
  7875=>"011110100",
  7876=>"110000000",
  7877=>"101111010",
  7878=>"000001001",
  7879=>"100001100",
  7880=>"000000110",
  7881=>"000110101",
  7882=>"100010100",
  7883=>"110010000",
  7884=>"000110111",
  7885=>"011100110",
  7886=>"010111111",
  7887=>"000000011",
  7888=>"010101110",
  7889=>"110101100",
  7890=>"111101100",
  7891=>"101101001",
  7892=>"101011011",
  7893=>"110010101",
  7894=>"111110101",
  7895=>"000000100",
  7896=>"001100011",
  7897=>"110111111",
  7898=>"111000111",
  7899=>"110111110",
  7900=>"011001000",
  7901=>"000100101",
  7902=>"000111011",
  7903=>"111111100",
  7904=>"000001100",
  7905=>"110101101",
  7906=>"000011101",
  7907=>"101101000",
  7908=>"001010101",
  7909=>"011101110",
  7910=>"001010000",
  7911=>"011111111",
  7912=>"111000110",
  7913=>"011011001",
  7914=>"000001001",
  7915=>"011110110",
  7916=>"010000101",
  7917=>"101101010",
  7918=>"001111111",
  7919=>"101000111",
  7920=>"110111110",
  7921=>"110111010",
  7922=>"000101100",
  7923=>"000000100",
  7924=>"011000010",
  7925=>"111011101",
  7926=>"010101101",
  7927=>"111110101",
  7928=>"111000111",
  7929=>"101000111",
  7930=>"000001111",
  7931=>"001100001",
  7932=>"100010101",
  7933=>"101010010",
  7934=>"110000011",
  7935=>"000011101",
  7936=>"000011110",
  7937=>"000101011",
  7938=>"001001011",
  7939=>"110111110",
  7940=>"010101111",
  7941=>"001011000",
  7942=>"001000010",
  7943=>"110111100",
  7944=>"101010001",
  7945=>"001000000",
  7946=>"111001011",
  7947=>"011100001",
  7948=>"011011000",
  7949=>"010001001",
  7950=>"111100111",
  7951=>"100101001",
  7952=>"010010111",
  7953=>"100111010",
  7954=>"111111100",
  7955=>"101010101",
  7956=>"011111100",
  7957=>"100111100",
  7958=>"110111101",
  7959=>"010010011",
  7960=>"010110110",
  7961=>"001101001",
  7962=>"111101111",
  7963=>"010000010",
  7964=>"011000101",
  7965=>"011111111",
  7966=>"111000101",
  7967=>"000111010",
  7968=>"000010001",
  7969=>"110000000",
  7970=>"001110001",
  7971=>"000000010",
  7972=>"011010100",
  7973=>"001010011",
  7974=>"011011100",
  7975=>"000010011",
  7976=>"000110000",
  7977=>"100011111",
  7978=>"110101000",
  7979=>"110011001",
  7980=>"101010011",
  7981=>"011001101",
  7982=>"010000111",
  7983=>"111111110",
  7984=>"011000001",
  7985=>"110111000",
  7986=>"010011100",
  7987=>"101101101",
  7988=>"000100101",
  7989=>"100000111",
  7990=>"000000000",
  7991=>"010011011",
  7992=>"111011100",
  7993=>"110100010",
  7994=>"010000000",
  7995=>"010100011",
  7996=>"010101101",
  7997=>"000010101",
  7998=>"010010000",
  7999=>"110101010",
  8000=>"111111000",
  8001=>"101101000",
  8002=>"100000011",
  8003=>"001100001",
  8004=>"100001000",
  8005=>"111001101",
  8006=>"111001111",
  8007=>"111110001",
  8008=>"101011100",
  8009=>"001011101",
  8010=>"100101100",
  8011=>"101101101",
  8012=>"010000010",
  8013=>"111101111",
  8014=>"001000100",
  8015=>"111001010",
  8016=>"011110010",
  8017=>"100000010",
  8018=>"011101111",
  8019=>"111001011",
  8020=>"111111000",
  8021=>"010111110",
  8022=>"111001100",
  8023=>"010000011",
  8024=>"001011011",
  8025=>"001010000",
  8026=>"011111111",
  8027=>"000010101",
  8028=>"101101010",
  8029=>"010000011",
  8030=>"010100110",
  8031=>"000111101",
  8032=>"000110001",
  8033=>"101000100",
  8034=>"101010001",
  8035=>"111110000",
  8036=>"111011111",
  8037=>"110100110",
  8038=>"010100011",
  8039=>"111001011",
  8040=>"001100111",
  8041=>"010011011",
  8042=>"011011010",
  8043=>"101110000",
  8044=>"100100011",
  8045=>"011110000",
  8046=>"010000010",
  8047=>"101101010",
  8048=>"001001000",
  8049=>"111000010",
  8050=>"110111001",
  8051=>"100011110",
  8052=>"000010010",
  8053=>"000110011",
  8054=>"000000000",
  8055=>"111101011",
  8056=>"001011101",
  8057=>"110111100",
  8058=>"100010110",
  8059=>"110010001",
  8060=>"100000110",
  8061=>"100000000",
  8062=>"001111001",
  8063=>"001011101",
  8064=>"011000100",
  8065=>"001011011",
  8066=>"111001101",
  8067=>"000011001",
  8068=>"001100101",
  8069=>"110010001",
  8070=>"100111001",
  8071=>"110110110",
  8072=>"101010100",
  8073=>"000100110",
  8074=>"100001010",
  8075=>"111000110",
  8076=>"111111011",
  8077=>"101111101",
  8078=>"111110110",
  8079=>"100001111",
  8080=>"011010000",
  8081=>"001111110",
  8082=>"101010111",
  8083=>"010110101",
  8084=>"111001100",
  8085=>"001001000",
  8086=>"111100110",
  8087=>"111100000",
  8088=>"110110110",
  8089=>"011001001",
  8090=>"111110001",
  8091=>"111010001",
  8092=>"001001010",
  8093=>"100110000",
  8094=>"111001000",
  8095=>"011001010",
  8096=>"010011010",
  8097=>"001000101",
  8098=>"110000111",
  8099=>"000001101",
  8100=>"000011001",
  8101=>"101110111",
  8102=>"100110110",
  8103=>"110011111",
  8104=>"110010100",
  8105=>"001000110",
  8106=>"110101011",
  8107=>"011000000",
  8108=>"111111100",
  8109=>"110111000",
  8110=>"010010111",
  8111=>"011011101",
  8112=>"110001101",
  8113=>"000111110",
  8114=>"010110110",
  8115=>"010110110",
  8116=>"101010001",
  8117=>"101100000",
  8118=>"010110011",
  8119=>"011110011",
  8120=>"001010010",
  8121=>"110010000",
  8122=>"010011011",
  8123=>"100101110",
  8124=>"100101101",
  8125=>"110000111",
  8126=>"011101000",
  8127=>"010000000",
  8128=>"011010000",
  8129=>"001001010",
  8130=>"111000000",
  8131=>"111110111",
  8132=>"101111110",
  8133=>"101110000",
  8134=>"001110010",
  8135=>"001111010",
  8136=>"000000000",
  8137=>"010011000",
  8138=>"000010000",
  8139=>"101000011",
  8140=>"100011000",
  8141=>"011000100",
  8142=>"011010011",
  8143=>"101011110",
  8144=>"111111101",
  8145=>"110010111",
  8146=>"100111000",
  8147=>"000101111",
  8148=>"111100001",
  8149=>"001100011",
  8150=>"000100111",
  8151=>"110010111",
  8152=>"110111111",
  8153=>"001000010",
  8154=>"010010010",
  8155=>"001000100",
  8156=>"011000010",
  8157=>"100111010",
  8158=>"001011001",
  8159=>"011101110",
  8160=>"110001001",
  8161=>"101011101",
  8162=>"101011010",
  8163=>"001101101",
  8164=>"101010101",
  8165=>"110010000",
  8166=>"101000100",
  8167=>"010110110",
  8168=>"110110100",
  8169=>"000000000",
  8170=>"010000011",
  8171=>"010010110",
  8172=>"000010011",
  8173=>"111111001",
  8174=>"011111001",
  8175=>"111101100",
  8176=>"011100101",
  8177=>"001000000",
  8178=>"000000011",
  8179=>"111010111",
  8180=>"100110001",
  8181=>"001000110",
  8182=>"000010011",
  8183=>"100000000",
  8184=>"100101100",
  8185=>"010110001",
  8186=>"001011100",
  8187=>"111110010",
  8188=>"001110101",
  8189=>"101100011",
  8190=>"000011101",
  8191=>"110100001",
  8192=>"101011000",
  8193=>"101100100",
  8194=>"111011001",
  8195=>"011110101",
  8196=>"111001000",
  8197=>"010000001",
  8198=>"001011010",
  8199=>"000100100",
  8200=>"010100011",
  8201=>"011000100",
  8202=>"110101100",
  8203=>"101010100",
  8204=>"010101100",
  8205=>"010101100",
  8206=>"011111001",
  8207=>"101011001",
  8208=>"001001000",
  8209=>"010111101",
  8210=>"010100111",
  8211=>"000010101",
  8212=>"111001000",
  8213=>"110001000",
  8214=>"100111110",
  8215=>"111100010",
  8216=>"100110011",
  8217=>"000000110",
  8218=>"100101110",
  8219=>"001010111",
  8220=>"001100010",
  8221=>"111101100",
  8222=>"110010110",
  8223=>"010110110",
  8224=>"110101011",
  8225=>"010110111",
  8226=>"101111110",
  8227=>"000000010",
  8228=>"101100011",
  8229=>"001000101",
  8230=>"000101101",
  8231=>"010011010",
  8232=>"000011111",
  8233=>"010100111",
  8234=>"111010010",
  8235=>"111100110",
  8236=>"011011111",
  8237=>"010101101",
  8238=>"000010011",
  8239=>"111101101",
  8240=>"010101000",
  8241=>"010101011",
  8242=>"001010100",
  8243=>"011100110",
  8244=>"100000110",
  8245=>"100000010",
  8246=>"000110010",
  8247=>"110101101",
  8248=>"111001110",
  8249=>"111000110",
  8250=>"000011101",
  8251=>"111001110",
  8252=>"001001001",
  8253=>"101000011",
  8254=>"111001000",
  8255=>"011100001",
  8256=>"010000100",
  8257=>"011010010",
  8258=>"101101110",
  8259=>"111000001",
  8260=>"001100101",
  8261=>"010111010",
  8262=>"101011001",
  8263=>"111100010",
  8264=>"000010100",
  8265=>"111111101",
  8266=>"111100100",
  8267=>"100111010",
  8268=>"000001101",
  8269=>"001000111",
  8270=>"001100111",
  8271=>"101101111",
  8272=>"010100100",
  8273=>"000000010",
  8274=>"010000001",
  8275=>"111000011",
  8276=>"111011100",
  8277=>"000110110",
  8278=>"011011011",
  8279=>"100000010",
  8280=>"000111110",
  8281=>"111001110",
  8282=>"010101011",
  8283=>"111110100",
  8284=>"010000000",
  8285=>"011101111",
  8286=>"111100011",
  8287=>"001110001",
  8288=>"011001001",
  8289=>"101111001",
  8290=>"111000101",
  8291=>"001000010",
  8292=>"101111111",
  8293=>"011011111",
  8294=>"011000101",
  8295=>"000100110",
  8296=>"011100100",
  8297=>"000010011",
  8298=>"111010101",
  8299=>"000010010",
  8300=>"111110001",
  8301=>"111000101",
  8302=>"001101010",
  8303=>"110001001",
  8304=>"111100001",
  8305=>"010100111",
  8306=>"000100010",
  8307=>"111110000",
  8308=>"111110110",
  8309=>"011101001",
  8310=>"001101010",
  8311=>"111010111",
  8312=>"101100100",
  8313=>"101001000",
  8314=>"101001100",
  8315=>"111010000",
  8316=>"101011110",
  8317=>"010111011",
  8318=>"111001000",
  8319=>"001101101",
  8320=>"011100110",
  8321=>"000001000",
  8322=>"110001000",
  8323=>"100000011",
  8324=>"110101101",
  8325=>"010111110",
  8326=>"010111011",
  8327=>"111000110",
  8328=>"001010101",
  8329=>"111111101",
  8330=>"111100110",
  8331=>"110001010",
  8332=>"100111100",
  8333=>"001110011",
  8334=>"101001000",
  8335=>"111111011",
  8336=>"111001111",
  8337=>"000000001",
  8338=>"111110111",
  8339=>"111001101",
  8340=>"000001001",
  8341=>"000000101",
  8342=>"000110001",
  8343=>"010011111",
  8344=>"101001111",
  8345=>"111011101",
  8346=>"011101110",
  8347=>"111000111",
  8348=>"000101011",
  8349=>"001011000",
  8350=>"101011011",
  8351=>"001110100",
  8352=>"101000001",
  8353=>"011001010",
  8354=>"110101110",
  8355=>"111001010",
  8356=>"001101110",
  8357=>"111011001",
  8358=>"101011100",
  8359=>"101010000",
  8360=>"111101100",
  8361=>"011011110",
  8362=>"001001010",
  8363=>"001111110",
  8364=>"001001000",
  8365=>"001010101",
  8366=>"111011101",
  8367=>"010110001",
  8368=>"000001000",
  8369=>"101011010",
  8370=>"010100100",
  8371=>"110011011",
  8372=>"001110101",
  8373=>"111111011",
  8374=>"001010100",
  8375=>"111000111",
  8376=>"110101100",
  8377=>"001010000",
  8378=>"000100110",
  8379=>"101111101",
  8380=>"001100110",
  8381=>"110100001",
  8382=>"010011000",
  8383=>"111101110",
  8384=>"111001010",
  8385=>"111101101",
  8386=>"101000110",
  8387=>"100001011",
  8388=>"111011001",
  8389=>"100000101",
  8390=>"000111110",
  8391=>"111111100",
  8392=>"000101001",
  8393=>"011101111",
  8394=>"011000110",
  8395=>"011011110",
  8396=>"010000000",
  8397=>"111110010",
  8398=>"111011111",
  8399=>"111100101",
  8400=>"001101100",
  8401=>"101001110",
  8402=>"001111011",
  8403=>"111010101",
  8404=>"111110010",
  8405=>"110100100",
  8406=>"001000000",
  8407=>"101011101",
  8408=>"110001000",
  8409=>"100011001",
  8410=>"001011111",
  8411=>"111000111",
  8412=>"100111110",
  8413=>"110001010",
  8414=>"010101010",
  8415=>"101111111",
  8416=>"111100011",
  8417=>"010111110",
  8418=>"001110001",
  8419=>"001110011",
  8420=>"111111101",
  8421=>"010100010",
  8422=>"011011010",
  8423=>"011100110",
  8424=>"010100010",
  8425=>"000001111",
  8426=>"011000111",
  8427=>"001110011",
  8428=>"000111000",
  8429=>"110110000",
  8430=>"100011100",
  8431=>"011110011",
  8432=>"110011011",
  8433=>"100111100",
  8434=>"000101001",
  8435=>"111111111",
  8436=>"101011000",
  8437=>"100110011",
  8438=>"010011100",
  8439=>"111000000",
  8440=>"110000100",
  8441=>"001011010",
  8442=>"000001010",
  8443=>"010101110",
  8444=>"000011110",
  8445=>"001000000",
  8446=>"010001010",
  8447=>"010000000",
  8448=>"000010101",
  8449=>"100011101",
  8450=>"001111011",
  8451=>"000101101",
  8452=>"001101100",
  8453=>"111000011",
  8454=>"110110010",
  8455=>"101011010",
  8456=>"110000011",
  8457=>"000001011",
  8458=>"110011111",
  8459=>"100100001",
  8460=>"110010010",
  8461=>"010100010",
  8462=>"000100100",
  8463=>"100000110",
  8464=>"001110101",
  8465=>"010011110",
  8466=>"110111001",
  8467=>"111101110",
  8468=>"010110001",
  8469=>"111000011",
  8470=>"101001101",
  8471=>"010000111",
  8472=>"100101000",
  8473=>"001011011",
  8474=>"111001101",
  8475=>"101111001",
  8476=>"110000000",
  8477=>"110000000",
  8478=>"001111111",
  8479=>"111110110",
  8480=>"111011001",
  8481=>"011111011",
  8482=>"101110100",
  8483=>"010111101",
  8484=>"010011011",
  8485=>"110101001",
  8486=>"110100111",
  8487=>"111110100",
  8488=>"001001011",
  8489=>"000010010",
  8490=>"010001010",
  8491=>"110010111",
  8492=>"111111111",
  8493=>"000111000",
  8494=>"101000001",
  8495=>"101110101",
  8496=>"111001001",
  8497=>"001010000",
  8498=>"000000000",
  8499=>"000111110",
  8500=>"000001111",
  8501=>"010000101",
  8502=>"001011000",
  8503=>"011001000",
  8504=>"001000110",
  8505=>"011100001",
  8506=>"110001001",
  8507=>"000001111",
  8508=>"011011001",
  8509=>"110110110",
  8510=>"111010100",
  8511=>"001000010",
  8512=>"101101111",
  8513=>"101001011",
  8514=>"001011011",
  8515=>"011110010",
  8516=>"101001011",
  8517=>"100001010",
  8518=>"110000001",
  8519=>"001000000",
  8520=>"011010101",
  8521=>"101010101",
  8522=>"111110010",
  8523=>"000010101",
  8524=>"100110000",
  8525=>"110000010",
  8526=>"001100011",
  8527=>"100000110",
  8528=>"101110001",
  8529=>"011101000",
  8530=>"110001111",
  8531=>"001011101",
  8532=>"010100111",
  8533=>"110101111",
  8534=>"111000000",
  8535=>"001100001",
  8536=>"010001001",
  8537=>"010001011",
  8538=>"010000111",
  8539=>"101111110",
  8540=>"100100101",
  8541=>"111010010",
  8542=>"110000001",
  8543=>"100010001",
  8544=>"010001000",
  8545=>"111000101",
  8546=>"001001101",
  8547=>"010001000",
  8548=>"110011100",
  8549=>"111011111",
  8550=>"110011011",
  8551=>"100001100",
  8552=>"000110000",
  8553=>"110111001",
  8554=>"100110101",
  8555=>"010100000",
  8556=>"101101010",
  8557=>"010111001",
  8558=>"100010010",
  8559=>"101010110",
  8560=>"001101111",
  8561=>"010001111",
  8562=>"100011001",
  8563=>"010000000",
  8564=>"010100010",
  8565=>"110100110",
  8566=>"010000110",
  8567=>"100101011",
  8568=>"010000101",
  8569=>"011011111",
  8570=>"111000111",
  8571=>"101101110",
  8572=>"110110001",
  8573=>"111111111",
  8574=>"101101011",
  8575=>"111000100",
  8576=>"100100101",
  8577=>"001000100",
  8578=>"100111010",
  8579=>"101101010",
  8580=>"110001000",
  8581=>"100111111",
  8582=>"110000110",
  8583=>"100000000",
  8584=>"000011010",
  8585=>"111000101",
  8586=>"000100000",
  8587=>"010001111",
  8588=>"010111100",
  8589=>"010100010",
  8590=>"110000000",
  8591=>"111001000",
  8592=>"111000101",
  8593=>"100000101",
  8594=>"011101001",
  8595=>"011111011",
  8596=>"100001100",
  8597=>"000110101",
  8598=>"100000011",
  8599=>"111111110",
  8600=>"001010111",
  8601=>"100000111",
  8602=>"111110001",
  8603=>"011000001",
  8604=>"011110111",
  8605=>"101100000",
  8606=>"101000010",
  8607=>"000000110",
  8608=>"001100001",
  8609=>"111101000",
  8610=>"110100011",
  8611=>"111010111",
  8612=>"101111101",
  8613=>"101100001",
  8614=>"010011101",
  8615=>"100000011",
  8616=>"010000101",
  8617=>"000011000",
  8618=>"011010101",
  8619=>"010001010",
  8620=>"000011000",
  8621=>"110000100",
  8622=>"001101100",
  8623=>"111110010",
  8624=>"111111010",
  8625=>"111100011",
  8626=>"111001000",
  8627=>"100011001",
  8628=>"111001001",
  8629=>"000101110",
  8630=>"000110111",
  8631=>"110010011",
  8632=>"100000101",
  8633=>"010100110",
  8634=>"001110000",
  8635=>"101011110",
  8636=>"100010101",
  8637=>"010000000",
  8638=>"010000011",
  8639=>"001010110",
  8640=>"000110000",
  8641=>"001110111",
  8642=>"000000110",
  8643=>"111110111",
  8644=>"111000111",
  8645=>"010110111",
  8646=>"011010111",
  8647=>"100100110",
  8648=>"110001101",
  8649=>"101100011",
  8650=>"000000100",
  8651=>"110010000",
  8652=>"000111001",
  8653=>"100011100",
  8654=>"111110010",
  8655=>"000000100",
  8656=>"010001011",
  8657=>"011001100",
  8658=>"000000011",
  8659=>"111101001",
  8660=>"100110111",
  8661=>"100011011",
  8662=>"111111011",
  8663=>"001001000",
  8664=>"110001000",
  8665=>"011001111",
  8666=>"000100010",
  8667=>"000111001",
  8668=>"110010001",
  8669=>"000110100",
  8670=>"011101101",
  8671=>"000011111",
  8672=>"101111100",
  8673=>"001011001",
  8674=>"011011001",
  8675=>"000111000",
  8676=>"000011001",
  8677=>"110111001",
  8678=>"001101001",
  8679=>"110101011",
  8680=>"100011111",
  8681=>"001100110",
  8682=>"101110000",
  8683=>"001001001",
  8684=>"011101110",
  8685=>"110010111",
  8686=>"000000011",
  8687=>"011000101",
  8688=>"110110111",
  8689=>"111111001",
  8690=>"000011110",
  8691=>"010101111",
  8692=>"100000101",
  8693=>"101110011",
  8694=>"010011001",
  8695=>"001101000",
  8696=>"000101110",
  8697=>"100011111",
  8698=>"001010000",
  8699=>"111111010",
  8700=>"101000001",
  8701=>"001100111",
  8702=>"110001110",
  8703=>"101111101",
  8704=>"010111010",
  8705=>"011010010",
  8706=>"110100000",
  8707=>"010011001",
  8708=>"000000101",
  8709=>"011000000",
  8710=>"110110010",
  8711=>"111111010",
  8712=>"011010000",
  8713=>"011000101",
  8714=>"101100111",
  8715=>"101110100",
  8716=>"101000100",
  8717=>"101101110",
  8718=>"101010111",
  8719=>"001011000",
  8720=>"100011111",
  8721=>"100110101",
  8722=>"101101000",
  8723=>"111101111",
  8724=>"000000000",
  8725=>"100000110",
  8726=>"001010101",
  8727=>"100011111",
  8728=>"100110011",
  8729=>"010101000",
  8730=>"101010111",
  8731=>"001001100",
  8732=>"110011000",
  8733=>"010101000",
  8734=>"101110011",
  8735=>"000001101",
  8736=>"100100010",
  8737=>"110101100",
  8738=>"001100000",
  8739=>"111101000",
  8740=>"010101000",
  8741=>"100101100",
  8742=>"100000000",
  8743=>"101000001",
  8744=>"100110111",
  8745=>"001100111",
  8746=>"010010011",
  8747=>"100100010",
  8748=>"011100101",
  8749=>"101000010",
  8750=>"000000010",
  8751=>"100000101",
  8752=>"011011101",
  8753=>"100110110",
  8754=>"000010101",
  8755=>"111001101",
  8756=>"011111001",
  8757=>"000110001",
  8758=>"010100010",
  8759=>"011011010",
  8760=>"110001100",
  8761=>"001100101",
  8762=>"001110110",
  8763=>"100010000",
  8764=>"010001110",
  8765=>"111011010",
  8766=>"111110110",
  8767=>"100000010",
  8768=>"110011001",
  8769=>"100000011",
  8770=>"111101000",
  8771=>"101000000",
  8772=>"011100010",
  8773=>"100011111",
  8774=>"111101001",
  8775=>"101101110",
  8776=>"110100001",
  8777=>"001110001",
  8778=>"011011100",
  8779=>"100110110",
  8780=>"011110000",
  8781=>"101111110",
  8782=>"111101111",
  8783=>"110111011",
  8784=>"100011100",
  8785=>"010101001",
  8786=>"111011000",
  8787=>"010010110",
  8788=>"000110101",
  8789=>"101100110",
  8790=>"011100101",
  8791=>"011011111",
  8792=>"111000011",
  8793=>"010111001",
  8794=>"100111001",
  8795=>"011101011",
  8796=>"111000010",
  8797=>"001000011",
  8798=>"001101011",
  8799=>"001011101",
  8800=>"011011011",
  8801=>"000001001",
  8802=>"111111011",
  8803=>"110011000",
  8804=>"110100101",
  8805=>"011100011",
  8806=>"000011101",
  8807=>"010101101",
  8808=>"010101010",
  8809=>"000000010",
  8810=>"001011000",
  8811=>"100000110",
  8812=>"100100100",
  8813=>"001100101",
  8814=>"010000110",
  8815=>"010100000",
  8816=>"000010101",
  8817=>"110101110",
  8818=>"100011110",
  8819=>"111001010",
  8820=>"010000111",
  8821=>"010000010",
  8822=>"001011101",
  8823=>"101101111",
  8824=>"100101111",
  8825=>"000001011",
  8826=>"111000000",
  8827=>"011011100",
  8828=>"111001110",
  8829=>"111001011",
  8830=>"011011000",
  8831=>"010000110",
  8832=>"101100101",
  8833=>"010011111",
  8834=>"111010111",
  8835=>"011010000",
  8836=>"001010000",
  8837=>"111000111",
  8838=>"001000011",
  8839=>"111101010",
  8840=>"100111001",
  8841=>"011000101",
  8842=>"011101000",
  8843=>"011000100",
  8844=>"111010001",
  8845=>"010010111",
  8846=>"101001010",
  8847=>"110101011",
  8848=>"010000110",
  8849=>"110101111",
  8850=>"001010011",
  8851=>"010000001",
  8852=>"101100010",
  8853=>"100001000",
  8854=>"101101110",
  8855=>"011001101",
  8856=>"011101111",
  8857=>"010110101",
  8858=>"100110011",
  8859=>"011010111",
  8860=>"100000011",
  8861=>"010101010",
  8862=>"000001011",
  8863=>"111001001",
  8864=>"111100100",
  8865=>"000000110",
  8866=>"001000101",
  8867=>"110000010",
  8868=>"010011100",
  8869=>"011010110",
  8870=>"001010001",
  8871=>"001010100",
  8872=>"111110111",
  8873=>"110001101",
  8874=>"000110000",
  8875=>"100110010",
  8876=>"000101000",
  8877=>"000100000",
  8878=>"000011110",
  8879=>"001110100",
  8880=>"111110101",
  8881=>"000000011",
  8882=>"111001110",
  8883=>"111001010",
  8884=>"011101100",
  8885=>"110111111",
  8886=>"111111110",
  8887=>"010001000",
  8888=>"100000011",
  8889=>"110101000",
  8890=>"011011100",
  8891=>"101100100",
  8892=>"011110010",
  8893=>"110100110",
  8894=>"100101000",
  8895=>"111000111",
  8896=>"111011111",
  8897=>"100000111",
  8898=>"001011001",
  8899=>"111111010",
  8900=>"011100010",
  8901=>"000110100",
  8902=>"111111001",
  8903=>"100000101",
  8904=>"000001100",
  8905=>"001011000",
  8906=>"001001001",
  8907=>"001100010",
  8908=>"111011011",
  8909=>"111000111",
  8910=>"011100101",
  8911=>"111000000",
  8912=>"011111101",
  8913=>"111000000",
  8914=>"111011100",
  8915=>"010111111",
  8916=>"000000110",
  8917=>"010000010",
  8918=>"011010011",
  8919=>"001001110",
  8920=>"001001110",
  8921=>"101100010",
  8922=>"001001111",
  8923=>"110100101",
  8924=>"101101100",
  8925=>"101011010",
  8926=>"010101000",
  8927=>"100101100",
  8928=>"000000001",
  8929=>"101000011",
  8930=>"001010111",
  8931=>"100100010",
  8932=>"000001010",
  8933=>"101000010",
  8934=>"101111100",
  8935=>"001101010",
  8936=>"011111000",
  8937=>"101101010",
  8938=>"111000110",
  8939=>"100101010",
  8940=>"010001010",
  8941=>"001001001",
  8942=>"101011010",
  8943=>"001111000",
  8944=>"110010110",
  8945=>"101111101",
  8946=>"000101000",
  8947=>"000001000",
  8948=>"100010010",
  8949=>"101111001",
  8950=>"111110000",
  8951=>"111011001",
  8952=>"100000111",
  8953=>"100011111",
  8954=>"110010001",
  8955=>"001100000",
  8956=>"000010101",
  8957=>"111011100",
  8958=>"110101111",
  8959=>"110101010",
  8960=>"000110110",
  8961=>"100001011",
  8962=>"001001111",
  8963=>"100000000",
  8964=>"011110100",
  8965=>"110111000",
  8966=>"010001110",
  8967=>"010000010",
  8968=>"011110110",
  8969=>"000111110",
  8970=>"000110001",
  8971=>"101011100",
  8972=>"101100001",
  8973=>"110111101",
  8974=>"001101100",
  8975=>"011011110",
  8976=>"010110111",
  8977=>"100001101",
  8978=>"100010011",
  8979=>"110010001",
  8980=>"100110101",
  8981=>"011011010",
  8982=>"010111010",
  8983=>"001010000",
  8984=>"010101100",
  8985=>"100110010",
  8986=>"011100101",
  8987=>"110101100",
  8988=>"110001100",
  8989=>"001001001",
  8990=>"110011011",
  8991=>"011010010",
  8992=>"011010001",
  8993=>"101011110",
  8994=>"010010101",
  8995=>"001100010",
  8996=>"110001110",
  8997=>"101011111",
  8998=>"100111000",
  8999=>"100011110",
  9000=>"010000000",
  9001=>"111010101",
  9002=>"110000010",
  9003=>"011000011",
  9004=>"100101100",
  9005=>"101100011",
  9006=>"011010000",
  9007=>"110111111",
  9008=>"100101101",
  9009=>"111110000",
  9010=>"111011100",
  9011=>"010100101",
  9012=>"110110101",
  9013=>"001101010",
  9014=>"101000011",
  9015=>"110101111",
  9016=>"111000111",
  9017=>"101111001",
  9018=>"111000011",
  9019=>"001100101",
  9020=>"111011001",
  9021=>"011100100",
  9022=>"010111111",
  9023=>"000001111",
  9024=>"111011010",
  9025=>"110111011",
  9026=>"100001101",
  9027=>"111110001",
  9028=>"100110111",
  9029=>"110000111",
  9030=>"111001111",
  9031=>"110001101",
  9032=>"000110000",
  9033=>"110101010",
  9034=>"001001010",
  9035=>"011101101",
  9036=>"010011100",
  9037=>"111100101",
  9038=>"010111000",
  9039=>"101000010",
  9040=>"111100011",
  9041=>"111010111",
  9042=>"100011010",
  9043=>"100001011",
  9044=>"001110000",
  9045=>"010010100",
  9046=>"000011001",
  9047=>"001111100",
  9048=>"000010100",
  9049=>"010101100",
  9050=>"011010011",
  9051=>"100000100",
  9052=>"101000000",
  9053=>"011101110",
  9054=>"111000011",
  9055=>"000000000",
  9056=>"010100111",
  9057=>"011000011",
  9058=>"000000010",
  9059=>"111001111",
  9060=>"111110000",
  9061=>"011110000",
  9062=>"111000000",
  9063=>"110110110",
  9064=>"010101001",
  9065=>"100111100",
  9066=>"001100010",
  9067=>"001011101",
  9068=>"010010000",
  9069=>"010001111",
  9070=>"011001000",
  9071=>"011001000",
  9072=>"010100100",
  9073=>"000011001",
  9074=>"010100000",
  9075=>"110001110",
  9076=>"110001000",
  9077=>"010000110",
  9078=>"101001000",
  9079=>"011011111",
  9080=>"001101111",
  9081=>"101101000",
  9082=>"010010001",
  9083=>"110010001",
  9084=>"101000100",
  9085=>"111110101",
  9086=>"000001101",
  9087=>"010001100",
  9088=>"001000100",
  9089=>"100111101",
  9090=>"010001001",
  9091=>"000000100",
  9092=>"011001101",
  9093=>"100111110",
  9094=>"100101110",
  9095=>"011111000",
  9096=>"110100101",
  9097=>"101011100",
  9098=>"001000111",
  9099=>"111111010",
  9100=>"010010110",
  9101=>"101101101",
  9102=>"111110000",
  9103=>"011101010",
  9104=>"001101010",
  9105=>"101101001",
  9106=>"101100101",
  9107=>"001011011",
  9108=>"011010000",
  9109=>"011101100",
  9110=>"001001111",
  9111=>"010010001",
  9112=>"000000001",
  9113=>"111001000",
  9114=>"000101011",
  9115=>"011101010",
  9116=>"010100110",
  9117=>"110110111",
  9118=>"010110010",
  9119=>"000001100",
  9120=>"100011011",
  9121=>"001000000",
  9122=>"111011101",
  9123=>"000000000",
  9124=>"111111011",
  9125=>"101000111",
  9126=>"010100010",
  9127=>"001010110",
  9128=>"101010110",
  9129=>"010000010",
  9130=>"101011110",
  9131=>"110110000",
  9132=>"100101100",
  9133=>"111100101",
  9134=>"001111000",
  9135=>"000110100",
  9136=>"101110010",
  9137=>"001010101",
  9138=>"000110100",
  9139=>"011101010",
  9140=>"010100101",
  9141=>"100100110",
  9142=>"010100011",
  9143=>"000110110",
  9144=>"011101100",
  9145=>"000010110",
  9146=>"000111101",
  9147=>"000111100",
  9148=>"100111001",
  9149=>"010010101",
  9150=>"000101000",
  9151=>"011001101",
  9152=>"000100010",
  9153=>"111011110",
  9154=>"001001111",
  9155=>"100010111",
  9156=>"011011111",
  9157=>"100010111",
  9158=>"010011011",
  9159=>"110110111",
  9160=>"010111010",
  9161=>"000010100",
  9162=>"010011010",
  9163=>"000110000",
  9164=>"100010001",
  9165=>"110001111",
  9166=>"010001100",
  9167=>"100001111",
  9168=>"111111110",
  9169=>"101001101",
  9170=>"010111000",
  9171=>"111111000",
  9172=>"101101110",
  9173=>"010000001",
  9174=>"111000111",
  9175=>"100011111",
  9176=>"111111010",
  9177=>"001110011",
  9178=>"111110100",
  9179=>"111010100",
  9180=>"001001001",
  9181=>"001001110",
  9182=>"010000111",
  9183=>"100100111",
  9184=>"111000101",
  9185=>"000110110",
  9186=>"001110110",
  9187=>"000001010",
  9188=>"111111001",
  9189=>"011111011",
  9190=>"000010011",
  9191=>"000001100",
  9192=>"110110110",
  9193=>"111010110",
  9194=>"010010001",
  9195=>"100001011",
  9196=>"110101111",
  9197=>"000000000",
  9198=>"110011111",
  9199=>"111001001",
  9200=>"100100111",
  9201=>"000011001",
  9202=>"110001000",
  9203=>"110010001",
  9204=>"100000000",
  9205=>"000100001",
  9206=>"010000101",
  9207=>"101000100",
  9208=>"011010011",
  9209=>"110001101",
  9210=>"110011011",
  9211=>"100011101",
  9212=>"000000010",
  9213=>"000010000",
  9214=>"010110010",
  9215=>"110101001",
  9216=>"010111001",
  9217=>"101011000",
  9218=>"110010000",
  9219=>"101010100",
  9220=>"110111111",
  9221=>"100001100",
  9222=>"111111001",
  9223=>"100101000",
  9224=>"010110111",
  9225=>"000110011",
  9226=>"001110010",
  9227=>"100100101",
  9228=>"010001000",
  9229=>"100010010",
  9230=>"011100000",
  9231=>"000000100",
  9232=>"110101011",
  9233=>"000010011",
  9234=>"110010110",
  9235=>"000001100",
  9236=>"000011101",
  9237=>"110000001",
  9238=>"101110001",
  9239=>"101010011",
  9240=>"000010100",
  9241=>"110000100",
  9242=>"011110011",
  9243=>"101001111",
  9244=>"110001010",
  9245=>"101011100",
  9246=>"000110001",
  9247=>"010010011",
  9248=>"100011001",
  9249=>"110110110",
  9250=>"000000100",
  9251=>"000100010",
  9252=>"100110010",
  9253=>"001010111",
  9254=>"001000000",
  9255=>"100100111",
  9256=>"110000111",
  9257=>"111011000",
  9258=>"100011011",
  9259=>"001000000",
  9260=>"011001011",
  9261=>"001110000",
  9262=>"101110011",
  9263=>"000100001",
  9264=>"010101101",
  9265=>"101111000",
  9266=>"010110111",
  9267=>"100000000",
  9268=>"011101111",
  9269=>"000111101",
  9270=>"011011100",
  9271=>"110001101",
  9272=>"011000010",
  9273=>"010001111",
  9274=>"101101100",
  9275=>"100110110",
  9276=>"000010010",
  9277=>"010100100",
  9278=>"100111000",
  9279=>"010100100",
  9280=>"101010011",
  9281=>"001101001",
  9282=>"011001011",
  9283=>"110111100",
  9284=>"010101110",
  9285=>"100000010",
  9286=>"100101111",
  9287=>"111010010",
  9288=>"110001110",
  9289=>"100100111",
  9290=>"110000011",
  9291=>"111111010",
  9292=>"101001011",
  9293=>"011111000",
  9294=>"001111111",
  9295=>"011010000",
  9296=>"000011110",
  9297=>"000101111",
  9298=>"100000010",
  9299=>"011101101",
  9300=>"100111000",
  9301=>"001111000",
  9302=>"100111101",
  9303=>"110000001",
  9304=>"010010111",
  9305=>"001111100",
  9306=>"101101110",
  9307=>"011110101",
  9308=>"111101001",
  9309=>"000101111",
  9310=>"110110010",
  9311=>"001000111",
  9312=>"100010111",
  9313=>"001011100",
  9314=>"001010111",
  9315=>"000000000",
  9316=>"101011101",
  9317=>"011100111",
  9318=>"101010110",
  9319=>"000001011",
  9320=>"100010010",
  9321=>"101110000",
  9322=>"000110010",
  9323=>"000111010",
  9324=>"111001001",
  9325=>"101110001",
  9326=>"111000001",
  9327=>"101001100",
  9328=>"110101111",
  9329=>"101011100",
  9330=>"000111000",
  9331=>"111110100",
  9332=>"011000110",
  9333=>"110001011",
  9334=>"010011100",
  9335=>"101011011",
  9336=>"011010111",
  9337=>"000101010",
  9338=>"000101011",
  9339=>"000010000",
  9340=>"111001100",
  9341=>"001001111",
  9342=>"100111001",
  9343=>"001111001",
  9344=>"011010101",
  9345=>"111101101",
  9346=>"000001101",
  9347=>"011001001",
  9348=>"101001010",
  9349=>"010101001",
  9350=>"010010010",
  9351=>"111100001",
  9352=>"011110100",
  9353=>"010000001",
  9354=>"010010101",
  9355=>"010000110",
  9356=>"111010101",
  9357=>"110101000",
  9358=>"001111111",
  9359=>"010011110",
  9360=>"100101110",
  9361=>"111001111",
  9362=>"000110010",
  9363=>"101001011",
  9364=>"000000101",
  9365=>"100010111",
  9366=>"000001001",
  9367=>"011101011",
  9368=>"000000010",
  9369=>"111110001",
  9370=>"110110000",
  9371=>"001010111",
  9372=>"111110001",
  9373=>"001101010",
  9374=>"001110001",
  9375=>"110111010",
  9376=>"000001001",
  9377=>"101100111",
  9378=>"001001110",
  9379=>"011101111",
  9380=>"000000101",
  9381=>"111111101",
  9382=>"111110001",
  9383=>"111100100",
  9384=>"011110110",
  9385=>"110111101",
  9386=>"001101001",
  9387=>"001101001",
  9388=>"111100010",
  9389=>"110011100",
  9390=>"110101101",
  9391=>"011100000",
  9392=>"000000110",
  9393=>"110000110",
  9394=>"100111000",
  9395=>"000000010",
  9396=>"111110010",
  9397=>"000010101",
  9398=>"101110010",
  9399=>"110110001",
  9400=>"000010000",
  9401=>"001101101",
  9402=>"001011010",
  9403=>"100110011",
  9404=>"100110101",
  9405=>"001010011",
  9406=>"101001110",
  9407=>"110000100",
  9408=>"011101001",
  9409=>"011000110",
  9410=>"011000011",
  9411=>"100101100",
  9412=>"011100011",
  9413=>"100110100",
  9414=>"010011010",
  9415=>"100000101",
  9416=>"001110111",
  9417=>"110010111",
  9418=>"111111110",
  9419=>"101101001",
  9420=>"001010000",
  9421=>"101011011",
  9422=>"101000111",
  9423=>"100000000",
  9424=>"011011000",
  9425=>"000010110",
  9426=>"011000011",
  9427=>"101000110",
  9428=>"110100100",
  9429=>"000100110",
  9430=>"101111001",
  9431=>"000000100",
  9432=>"010011000",
  9433=>"111001111",
  9434=>"001101010",
  9435=>"010010100",
  9436=>"111100000",
  9437=>"011110111",
  9438=>"101110110",
  9439=>"110111001",
  9440=>"000011111",
  9441=>"111100111",
  9442=>"011000000",
  9443=>"001100011",
  9444=>"101100111",
  9445=>"001100011",
  9446=>"100001001",
  9447=>"100100010",
  9448=>"000001100",
  9449=>"110010011",
  9450=>"101111001",
  9451=>"011110001",
  9452=>"111000111",
  9453=>"111110000",
  9454=>"100111001",
  9455=>"101000001",
  9456=>"110111100",
  9457=>"101100011",
  9458=>"000110111",
  9459=>"000000000",
  9460=>"001101010",
  9461=>"000000001",
  9462=>"110011100",
  9463=>"100101111",
  9464=>"001111110",
  9465=>"010100110",
  9466=>"000101101",
  9467=>"011000111",
  9468=>"010001100",
  9469=>"111010000",
  9470=>"101110010",
  9471=>"000101011",
  9472=>"001000010",
  9473=>"010111010",
  9474=>"001101100",
  9475=>"111011010",
  9476=>"101111001",
  9477=>"101101010",
  9478=>"001011011",
  9479=>"101110110",
  9480=>"011011100",
  9481=>"110110110",
  9482=>"100110110",
  9483=>"111111010",
  9484=>"001011010",
  9485=>"000110100",
  9486=>"001010001",
  9487=>"000110111",
  9488=>"000110100",
  9489=>"001001111",
  9490=>"010110100",
  9491=>"011101011",
  9492=>"000100111",
  9493=>"111011000",
  9494=>"001001011",
  9495=>"010100101",
  9496=>"010000010",
  9497=>"011100110",
  9498=>"100100000",
  9499=>"000110011",
  9500=>"010000001",
  9501=>"101111101",
  9502=>"000000101",
  9503=>"000110001",
  9504=>"001010001",
  9505=>"100111110",
  9506=>"010111010",
  9507=>"111001001",
  9508=>"010011011",
  9509=>"010010001",
  9510=>"111000101",
  9511=>"111011100",
  9512=>"110011110",
  9513=>"101101000",
  9514=>"101010000",
  9515=>"001000101",
  9516=>"011011010",
  9517=>"111111010",
  9518=>"100011110",
  9519=>"111110000",
  9520=>"001010110",
  9521=>"100001111",
  9522=>"101001110",
  9523=>"000110100",
  9524=>"001110100",
  9525=>"011001001",
  9526=>"001110101",
  9527=>"111001111",
  9528=>"000000110",
  9529=>"111101010",
  9530=>"011011011",
  9531=>"110011100",
  9532=>"100010111",
  9533=>"101110110",
  9534=>"011111000",
  9535=>"000100000",
  9536=>"101010011",
  9537=>"101101000",
  9538=>"111011101",
  9539=>"111000011",
  9540=>"010111100",
  9541=>"010111010",
  9542=>"101000001",
  9543=>"110010011",
  9544=>"000000100",
  9545=>"010001001",
  9546=>"110000110",
  9547=>"100110000",
  9548=>"011101010",
  9549=>"100110101",
  9550=>"011111011",
  9551=>"111011100",
  9552=>"011110000",
  9553=>"100111000",
  9554=>"111110111",
  9555=>"000010001",
  9556=>"001010001",
  9557=>"010010111",
  9558=>"100010101",
  9559=>"100001110",
  9560=>"001000110",
  9561=>"101000010",
  9562=>"110111110",
  9563=>"101010001",
  9564=>"110111100",
  9565=>"000001100",
  9566=>"100110110",
  9567=>"110000001",
  9568=>"011010001",
  9569=>"011001001",
  9570=>"111100011",
  9571=>"010000011",
  9572=>"001001001",
  9573=>"011101111",
  9574=>"010100100",
  9575=>"011100110",
  9576=>"111110110",
  9577=>"001111000",
  9578=>"000100100",
  9579=>"100100010",
  9580=>"001000001",
  9581=>"010001111",
  9582=>"111010110",
  9583=>"111101010",
  9584=>"101000110",
  9585=>"000001000",
  9586=>"011001100",
  9587=>"110000101",
  9588=>"010000100",
  9589=>"101001010",
  9590=>"010000010",
  9591=>"101111100",
  9592=>"011110100",
  9593=>"101100011",
  9594=>"111101011",
  9595=>"111001000",
  9596=>"101111011",
  9597=>"100111110",
  9598=>"010110011",
  9599=>"001110011",
  9600=>"001000011",
  9601=>"000010001",
  9602=>"111001011",
  9603=>"010011011",
  9604=>"001110011",
  9605=>"110100000",
  9606=>"001011111",
  9607=>"011011110",
  9608=>"000010000",
  9609=>"000101000",
  9610=>"100100111",
  9611=>"011111110",
  9612=>"010001000",
  9613=>"001001100",
  9614=>"101110011",
  9615=>"010110001",
  9616=>"100100011",
  9617=>"000000111",
  9618=>"101100111",
  9619=>"011001001",
  9620=>"110101101",
  9621=>"001001110",
  9622=>"111111010",
  9623=>"000000111",
  9624=>"000000010",
  9625=>"001000000",
  9626=>"101010010",
  9627=>"100011011",
  9628=>"101100100",
  9629=>"011001110",
  9630=>"011100101",
  9631=>"001011110",
  9632=>"100001001",
  9633=>"011010000",
  9634=>"001101011",
  9635=>"000001110",
  9636=>"111100011",
  9637=>"010110010",
  9638=>"001010101",
  9639=>"011000101",
  9640=>"001110011",
  9641=>"000011110",
  9642=>"111000011",
  9643=>"111100010",
  9644=>"101010110",
  9645=>"001100011",
  9646=>"101111011",
  9647=>"101011000",
  9648=>"010000111",
  9649=>"101111101",
  9650=>"110000100",
  9651=>"111011011",
  9652=>"111011100",
  9653=>"001100011",
  9654=>"111000110",
  9655=>"010100000",
  9656=>"101001110",
  9657=>"110101000",
  9658=>"001010010",
  9659=>"001000001",
  9660=>"110011011",
  9661=>"101110000",
  9662=>"001101101",
  9663=>"000111001",
  9664=>"001011010",
  9665=>"100000100",
  9666=>"100110110",
  9667=>"110111011",
  9668=>"010010111",
  9669=>"000001000",
  9670=>"111001010",
  9671=>"011111110",
  9672=>"000111000",
  9673=>"100001011",
  9674=>"110010101",
  9675=>"001100101",
  9676=>"000101001",
  9677=>"010010110",
  9678=>"011010000",
  9679=>"001011010",
  9680=>"111111000",
  9681=>"010101011",
  9682=>"110101101",
  9683=>"100101111",
  9684=>"010100010",
  9685=>"100111110",
  9686=>"100001011",
  9687=>"011010011",
  9688=>"010101101",
  9689=>"101110010",
  9690=>"101010110",
  9691=>"000101010",
  9692=>"011111001",
  9693=>"101101101",
  9694=>"000000101",
  9695=>"011110010",
  9696=>"001111111",
  9697=>"000101010",
  9698=>"111111011",
  9699=>"100011010",
  9700=>"000000101",
  9701=>"111101011",
  9702=>"101001101",
  9703=>"010110100",
  9704=>"011100010",
  9705=>"000101111",
  9706=>"011110110",
  9707=>"110010011",
  9708=>"000100010",
  9709=>"100001000",
  9710=>"000110000",
  9711=>"101011101",
  9712=>"101010101",
  9713=>"100010100",
  9714=>"110101010",
  9715=>"011001011",
  9716=>"001011000",
  9717=>"011000111",
  9718=>"010001101",
  9719=>"001110110",
  9720=>"110000000",
  9721=>"010110000",
  9722=>"110101001",
  9723=>"010000010",
  9724=>"111001100",
  9725=>"101111001",
  9726=>"011111100",
  9727=>"111011111",
  9728=>"010100000",
  9729=>"011110001",
  9730=>"110111000",
  9731=>"010001000",
  9732=>"110011100",
  9733=>"111100110",
  9734=>"000100110",
  9735=>"110110111",
  9736=>"010101001",
  9737=>"101001010",
  9738=>"000100010",
  9739=>"000001100",
  9740=>"101001101",
  9741=>"101110111",
  9742=>"011000000",
  9743=>"100101011",
  9744=>"011010110",
  9745=>"001100011",
  9746=>"011111010",
  9747=>"100101100",
  9748=>"101101010",
  9749=>"111001000",
  9750=>"101000010",
  9751=>"001001000",
  9752=>"111111010",
  9753=>"110010001",
  9754=>"011111111",
  9755=>"101101110",
  9756=>"001111011",
  9757=>"110000111",
  9758=>"100010001",
  9759=>"011001010",
  9760=>"010010011",
  9761=>"010000000",
  9762=>"010100001",
  9763=>"000011110",
  9764=>"010100111",
  9765=>"000001100",
  9766=>"010010111",
  9767=>"101101101",
  9768=>"010101111",
  9769=>"100111011",
  9770=>"001000101",
  9771=>"111011111",
  9772=>"100000110",
  9773=>"010100111",
  9774=>"000110101",
  9775=>"001011101",
  9776=>"011101100",
  9777=>"011110011",
  9778=>"000110000",
  9779=>"000100110",
  9780=>"000010010",
  9781=>"011000000",
  9782=>"111111000",
  9783=>"001010100",
  9784=>"001000001",
  9785=>"111000001",
  9786=>"100100101",
  9787=>"001110011",
  9788=>"101001001",
  9789=>"001000101",
  9790=>"101100110",
  9791=>"010011101",
  9792=>"000001001",
  9793=>"110000000",
  9794=>"010110101",
  9795=>"000010001",
  9796=>"011101010",
  9797=>"010010100",
  9798=>"100011101",
  9799=>"111011010",
  9800=>"011010100",
  9801=>"110111111",
  9802=>"001101010",
  9803=>"000001111",
  9804=>"001001111",
  9805=>"000011101",
  9806=>"111011001",
  9807=>"010111111",
  9808=>"111000001",
  9809=>"101101010",
  9810=>"101011110",
  9811=>"110001010",
  9812=>"000010100",
  9813=>"010001101",
  9814=>"000110000",
  9815=>"100110010",
  9816=>"011101000",
  9817=>"100010111",
  9818=>"100000100",
  9819=>"001010001",
  9820=>"111111010",
  9821=>"011010000",
  9822=>"001100111",
  9823=>"010011000",
  9824=>"110110001",
  9825=>"100101111",
  9826=>"100110100",
  9827=>"111010010",
  9828=>"000011101",
  9829=>"011010110",
  9830=>"000001101",
  9831=>"111111000",
  9832=>"011001100",
  9833=>"011001101",
  9834=>"000000101",
  9835=>"000001101",
  9836=>"000100010",
  9837=>"010101001",
  9838=>"011010001",
  9839=>"111100111",
  9840=>"110000000",
  9841=>"000010011",
  9842=>"000101110",
  9843=>"011111110",
  9844=>"100011000",
  9845=>"111101111",
  9846=>"111010000",
  9847=>"101101001",
  9848=>"100011101",
  9849=>"011001111",
  9850=>"011010101",
  9851=>"110010011",
  9852=>"011100101",
  9853=>"010111001",
  9854=>"110110101",
  9855=>"001110110",
  9856=>"000100100",
  9857=>"110011000",
  9858=>"100101000",
  9859=>"111011110",
  9860=>"010100001",
  9861=>"110110000",
  9862=>"101101111",
  9863=>"010011011",
  9864=>"110111111",
  9865=>"110101000",
  9866=>"110111101",
  9867=>"101111110",
  9868=>"111000101",
  9869=>"001001010",
  9870=>"011101011",
  9871=>"110100100",
  9872=>"100010010",
  9873=>"000001001",
  9874=>"011000101",
  9875=>"000100000",
  9876=>"000101111",
  9877=>"111110000",
  9878=>"110000011",
  9879=>"111000110",
  9880=>"000101111",
  9881=>"111000110",
  9882=>"100100010",
  9883=>"001000100",
  9884=>"101010000",
  9885=>"110011000",
  9886=>"001110001",
  9887=>"110100110",
  9888=>"001110101",
  9889=>"110101011",
  9890=>"010101100",
  9891=>"111010001",
  9892=>"100101110",
  9893=>"111111100",
  9894=>"000100000",
  9895=>"000000111",
  9896=>"100100001",
  9897=>"000010011",
  9898=>"000001111",
  9899=>"011011111",
  9900=>"101110101",
  9901=>"001011010",
  9902=>"111101000",
  9903=>"010100100",
  9904=>"100101110",
  9905=>"110101100",
  9906=>"001110101",
  9907=>"001001100",
  9908=>"001100111",
  9909=>"101101110",
  9910=>"110111000",
  9911=>"011010010",
  9912=>"101000101",
  9913=>"110110001",
  9914=>"011100010",
  9915=>"110110100",
  9916=>"111001100",
  9917=>"110100011",
  9918=>"100010001",
  9919=>"101100011",
  9920=>"101011111",
  9921=>"111011000",
  9922=>"010011101",
  9923=>"110000000",
  9924=>"001101101",
  9925=>"011011100",
  9926=>"111110001",
  9927=>"111011011",
  9928=>"111000000",
  9929=>"100000010",
  9930=>"110111110",
  9931=>"111011001",
  9932=>"110011011",
  9933=>"111100101",
  9934=>"000000000",
  9935=>"111010110",
  9936=>"011101011",
  9937=>"010011101",
  9938=>"101001101",
  9939=>"111111110",
  9940=>"010001100",
  9941=>"011110110",
  9942=>"001000110",
  9943=>"111111101",
  9944=>"010010111",
  9945=>"001010110",
  9946=>"010010000",
  9947=>"110100101",
  9948=>"101101001",
  9949=>"101100111",
  9950=>"000000111",
  9951=>"101101101",
  9952=>"010000011",
  9953=>"001010000",
  9954=>"101000111",
  9955=>"111000100",
  9956=>"010001101",
  9957=>"011011010",
  9958=>"010101111",
  9959=>"101000010",
  9960=>"011111010",
  9961=>"010001100",
  9962=>"110111000",
  9963=>"000011100",
  9964=>"111100011",
  9965=>"111011101",
  9966=>"000001000",
  9967=>"001110010",
  9968=>"111011010",
  9969=>"000011011",
  9970=>"101111101",
  9971=>"100011000",
  9972=>"100111110",
  9973=>"010111000",
  9974=>"000101001",
  9975=>"101101010",
  9976=>"000000101",
  9977=>"011011111",
  9978=>"010110111",
  9979=>"010111110",
  9980=>"110111111",
  9981=>"001110110",
  9982=>"000011100",
  9983=>"010011111",
  9984=>"100001101",
  9985=>"000111110",
  9986=>"110010000",
  9987=>"001001010",
  9988=>"010110100",
  9989=>"010011111",
  9990=>"101000001",
  9991=>"000011111",
  9992=>"101001000",
  9993=>"010010000",
  9994=>"100001100",
  9995=>"111010001",
  9996=>"110011001",
  9997=>"101011110",
  9998=>"000100100",
  9999=>"100101111",
  10000=>"101010001",
  10001=>"001010110",
  10002=>"101100111",
  10003=>"010100110",
  10004=>"111111010",
  10005=>"101101001",
  10006=>"101010011",
  10007=>"001000110",
  10008=>"010001100",
  10009=>"100101111",
  10010=>"010110001",
  10011=>"100010101",
  10012=>"111011110",
  10013=>"100011001",
  10014=>"111010100",
  10015=>"000110111",
  10016=>"001000101",
  10017=>"110111001",
  10018=>"001101101",
  10019=>"100110000",
  10020=>"000101100",
  10021=>"111011000",
  10022=>"001111001",
  10023=>"011100100",
  10024=>"111011100",
  10025=>"000100110",
  10026=>"001110100",
  10027=>"111011010",
  10028=>"010000110",
  10029=>"001001001",
  10030=>"010010110",
  10031=>"001111010",
  10032=>"011001000",
  10033=>"000100101",
  10034=>"010001010",
  10035=>"001010000",
  10036=>"111100011",
  10037=>"011001100",
  10038=>"111111010",
  10039=>"100111110",
  10040=>"000011010",
  10041=>"000010010",
  10042=>"101111111",
  10043=>"011111100",
  10044=>"100111011",
  10045=>"011011101",
  10046=>"010000111",
  10047=>"111000101",
  10048=>"001001000",
  10049=>"101111000",
  10050=>"100011000",
  10051=>"010010001",
  10052=>"100001011",
  10053=>"011001111",
  10054=>"111110100",
  10055=>"011001111",
  10056=>"111011101",
  10057=>"010000010",
  10058=>"110101000",
  10059=>"000011111",
  10060=>"011001110",
  10061=>"111101001",
  10062=>"010011110",
  10063=>"010000100",
  10064=>"010110111",
  10065=>"011010100",
  10066=>"010101001",
  10067=>"100011010",
  10068=>"101001010",
  10069=>"110100010",
  10070=>"101111110",
  10071=>"111001000",
  10072=>"110011111",
  10073=>"100001101",
  10074=>"000001001",
  10075=>"111110111",
  10076=>"000001000",
  10077=>"000010100",
  10078=>"100011011",
  10079=>"000001110",
  10080=>"100011001",
  10081=>"101110000",
  10082=>"111101011",
  10083=>"010011010",
  10084=>"000111111",
  10085=>"111110001",
  10086=>"000011110",
  10087=>"010000110",
  10088=>"101001001",
  10089=>"001000001",
  10090=>"011011001",
  10091=>"111001100",
  10092=>"100001001",
  10093=>"011001101",
  10094=>"111000111",
  10095=>"110101111",
  10096=>"110001000",
  10097=>"011000001",
  10098=>"000010010",
  10099=>"110101111",
  10100=>"000100010",
  10101=>"100001101",
  10102=>"100100010",
  10103=>"000010110",
  10104=>"101010100",
  10105=>"111111111",
  10106=>"101011011",
  10107=>"000001010",
  10108=>"100000110",
  10109=>"110100011",
  10110=>"011100011",
  10111=>"110011111",
  10112=>"011010001",
  10113=>"110010110",
  10114=>"011000111",
  10115=>"001001100",
  10116=>"111101110",
  10117=>"111011110",
  10118=>"000010101",
  10119=>"010110000",
  10120=>"101000001",
  10121=>"110010000",
  10122=>"110111001",
  10123=>"010011011",
  10124=>"011101011",
  10125=>"110110010",
  10126=>"000111000",
  10127=>"000000100",
  10128=>"010010100",
  10129=>"111110110",
  10130=>"111001100",
  10131=>"111011010",
  10132=>"111000111",
  10133=>"010111001",
  10134=>"110010101",
  10135=>"010010110",
  10136=>"000010101",
  10137=>"001001101",
  10138=>"011101000",
  10139=>"001100100",
  10140=>"010101111",
  10141=>"100011101",
  10142=>"010000011",
  10143=>"010110000",
  10144=>"100010000",
  10145=>"111011001",
  10146=>"111101110",
  10147=>"011000000",
  10148=>"000010000",
  10149=>"011100000",
  10150=>"110001110",
  10151=>"001110111",
  10152=>"000101010",
  10153=>"001110111",
  10154=>"110101010",
  10155=>"101101000",
  10156=>"000110000",
  10157=>"011111010",
  10158=>"100010101",
  10159=>"111111011",
  10160=>"011000111",
  10161=>"000001000",
  10162=>"000001101",
  10163=>"100000110",
  10164=>"010011001",
  10165=>"101111001",
  10166=>"010000010",
  10167=>"110011101",
  10168=>"101001100",
  10169=>"101100101",
  10170=>"001100100",
  10171=>"010011001",
  10172=>"100011111",
  10173=>"110111011",
  10174=>"000111111",
  10175=>"111101101",
  10176=>"001001111",
  10177=>"000110101",
  10178=>"101111111",
  10179=>"000001011",
  10180=>"000000000",
  10181=>"100001011",
  10182=>"100111100",
  10183=>"001011000",
  10184=>"101100011",
  10185=>"011100000",
  10186=>"111111111",
  10187=>"001110110",
  10188=>"000011111",
  10189=>"100000001",
  10190=>"001111011",
  10191=>"000001100",
  10192=>"111010100",
  10193=>"001001101",
  10194=>"001110010",
  10195=>"101000101",
  10196=>"010000101",
  10197=>"101110011",
  10198=>"111111011",
  10199=>"110110110",
  10200=>"100101011",
  10201=>"000111101",
  10202=>"111100111",
  10203=>"010001010",
  10204=>"001111100",
  10205=>"101111011",
  10206=>"000001010",
  10207=>"010010010",
  10208=>"100000000",
  10209=>"101010111",
  10210=>"100000000",
  10211=>"111111111",
  10212=>"010100011",
  10213=>"000000011",
  10214=>"110101100",
  10215=>"000100111",
  10216=>"100110001",
  10217=>"111000101",
  10218=>"111000010",
  10219=>"111011101",
  10220=>"011001111",
  10221=>"001011011",
  10222=>"001111010",
  10223=>"111100000",
  10224=>"101100111",
  10225=>"111101110",
  10226=>"010100100",
  10227=>"100001001",
  10228=>"001010000",
  10229=>"010101110",
  10230=>"100101011",
  10231=>"000101000",
  10232=>"111000000",
  10233=>"101011111",
  10234=>"110000101",
  10235=>"101101101",
  10236=>"000101001",
  10237=>"000110111",
  10238=>"011110100",
  10239=>"010011111",
  10240=>"111001011",
  10241=>"010010101",
  10242=>"001001111",
  10243=>"110110000",
  10244=>"001110110",
  10245=>"111011000",
  10246=>"111000000",
  10247=>"110011011",
  10248=>"100100100",
  10249=>"000001101",
  10250=>"010000110",
  10251=>"001110000",
  10252=>"011111110",
  10253=>"010110100",
  10254=>"110110011",
  10255=>"110101011",
  10256=>"000010110",
  10257=>"000000100",
  10258=>"111101100",
  10259=>"001000110",
  10260=>"000001100",
  10261=>"100010111",
  10262=>"101110101",
  10263=>"010011101",
  10264=>"111111011",
  10265=>"010011100",
  10266=>"001100011",
  10267=>"111001001",
  10268=>"011001110",
  10269=>"001001000",
  10270=>"101000101",
  10271=>"011100001",
  10272=>"111010101",
  10273=>"001000000",
  10274=>"100111011",
  10275=>"100101100",
  10276=>"111000010",
  10277=>"001000011",
  10278=>"000111111",
  10279=>"110010010",
  10280=>"100011011",
  10281=>"011011111",
  10282=>"010001010",
  10283=>"010100001",
  10284=>"101111010",
  10285=>"000100000",
  10286=>"000110110",
  10287=>"011011100",
  10288=>"010110011",
  10289=>"011111110",
  10290=>"101001110",
  10291=>"000110011",
  10292=>"101000010",
  10293=>"111011011",
  10294=>"000111011",
  10295=>"100010001",
  10296=>"001000011",
  10297=>"010100100",
  10298=>"011100010",
  10299=>"110000100",
  10300=>"010010100",
  10301=>"001000100",
  10302=>"110111001",
  10303=>"101100011",
  10304=>"011110010",
  10305=>"000000001",
  10306=>"010010110",
  10307=>"101100001",
  10308=>"111110001",
  10309=>"101011001",
  10310=>"010110110",
  10311=>"110110110",
  10312=>"100111100",
  10313=>"010110001",
  10314=>"111111110",
  10315=>"000000100",
  10316=>"011110101",
  10317=>"000010100",
  10318=>"000111101",
  10319=>"010001110",
  10320=>"011011111",
  10321=>"110011010",
  10322=>"100110111",
  10323=>"000011011",
  10324=>"101100100",
  10325=>"011100011",
  10326=>"000011000",
  10327=>"011100100",
  10328=>"111000111",
  10329=>"010001101",
  10330=>"010110011",
  10331=>"011101110",
  10332=>"111011100",
  10333=>"111000100",
  10334=>"100111110",
  10335=>"100111101",
  10336=>"010110101",
  10337=>"111010000",
  10338=>"001101111",
  10339=>"111011100",
  10340=>"101010101",
  10341=>"000110001",
  10342=>"010110100",
  10343=>"111011111",
  10344=>"011100101",
  10345=>"010100001",
  10346=>"010010001",
  10347=>"011111111",
  10348=>"010010011",
  10349=>"011100010",
  10350=>"000100000",
  10351=>"001100010",
  10352=>"000011110",
  10353=>"110011111",
  10354=>"100101101",
  10355=>"100011011",
  10356=>"000110110",
  10357=>"100110100",
  10358=>"010011001",
  10359=>"001110011",
  10360=>"100010001",
  10361=>"000110010",
  10362=>"110101011",
  10363=>"000110100",
  10364=>"101100001",
  10365=>"100110001",
  10366=>"010111000",
  10367=>"000101111",
  10368=>"001000101",
  10369=>"000111011",
  10370=>"110000100",
  10371=>"010000000",
  10372=>"011000001",
  10373=>"111010010",
  10374=>"000110100",
  10375=>"001111111",
  10376=>"110101000",
  10377=>"110101011",
  10378=>"101011110",
  10379=>"111001100",
  10380=>"001110110",
  10381=>"001111000",
  10382=>"011000111",
  10383=>"101110001",
  10384=>"011001001",
  10385=>"101111110",
  10386=>"011110101",
  10387=>"101110011",
  10388=>"001110111",
  10389=>"101011110",
  10390=>"001011000",
  10391=>"110110110",
  10392=>"110101100",
  10393=>"100100000",
  10394=>"001101111",
  10395=>"010001000",
  10396=>"011010111",
  10397=>"011000100",
  10398=>"100001001",
  10399=>"100100100",
  10400=>"010110100",
  10401=>"111001001",
  10402=>"110100100",
  10403=>"111010010",
  10404=>"110111110",
  10405=>"100110111",
  10406=>"001111001",
  10407=>"110000001",
  10408=>"010000110",
  10409=>"111010011",
  10410=>"100001000",
  10411=>"010111010",
  10412=>"111111111",
  10413=>"100101111",
  10414=>"110111100",
  10415=>"110101110",
  10416=>"000111001",
  10417=>"100010001",
  10418=>"111000100",
  10419=>"110001111",
  10420=>"010000111",
  10421=>"101111001",
  10422=>"000111100",
  10423=>"011001001",
  10424=>"000011111",
  10425=>"101110111",
  10426=>"010001010",
  10427=>"110100010",
  10428=>"111101111",
  10429=>"100011101",
  10430=>"001000101",
  10431=>"001000010",
  10432=>"101011011",
  10433=>"001001010",
  10434=>"000001111",
  10435=>"100001000",
  10436=>"010100001",
  10437=>"010001001",
  10438=>"011111100",
  10439=>"001000001",
  10440=>"101111111",
  10441=>"001011010",
  10442=>"001001000",
  10443=>"110101011",
  10444=>"101100001",
  10445=>"111011111",
  10446=>"100101111",
  10447=>"011010000",
  10448=>"111110001",
  10449=>"111100100",
  10450=>"101111001",
  10451=>"010101011",
  10452=>"101111010",
  10453=>"001101001",
  10454=>"010001011",
  10455=>"001101111",
  10456=>"101101111",
  10457=>"111010000",
  10458=>"000101101",
  10459=>"101010111",
  10460=>"101110000",
  10461=>"110011110",
  10462=>"001011100",
  10463=>"001011011",
  10464=>"011111010",
  10465=>"001010110",
  10466=>"110000100",
  10467=>"111000000",
  10468=>"111010111",
  10469=>"101100001",
  10470=>"110111011",
  10471=>"100001000",
  10472=>"000010011",
  10473=>"101011000",
  10474=>"100111111",
  10475=>"011101111",
  10476=>"001101001",
  10477=>"001000100",
  10478=>"100011011",
  10479=>"000101101",
  10480=>"110011111",
  10481=>"001010111",
  10482=>"001001000",
  10483=>"010101011",
  10484=>"110010000",
  10485=>"100000010",
  10486=>"100000101",
  10487=>"111000011",
  10488=>"100110101",
  10489=>"101001000",
  10490=>"000011010",
  10491=>"000000111",
  10492=>"010000010",
  10493=>"001011110",
  10494=>"110101011",
  10495=>"001010111",
  10496=>"100011110",
  10497=>"100011110",
  10498=>"011010100",
  10499=>"111100011",
  10500=>"111000101",
  10501=>"100100000",
  10502=>"000000011",
  10503=>"110111110",
  10504=>"111101011",
  10505=>"000010101",
  10506=>"110010111",
  10507=>"001011011",
  10508=>"111110001",
  10509=>"110010100",
  10510=>"101110100",
  10511=>"011000001",
  10512=>"110101101",
  10513=>"001011111",
  10514=>"111001110",
  10515=>"100111101",
  10516=>"100000000",
  10517=>"000101100",
  10518=>"011010111",
  10519=>"000010101",
  10520=>"001010100",
  10521=>"111100101",
  10522=>"010000110",
  10523=>"111010001",
  10524=>"011101110",
  10525=>"000100011",
  10526=>"101000110",
  10527=>"111001011",
  10528=>"000001100",
  10529=>"010001101",
  10530=>"000110101",
  10531=>"011110001",
  10532=>"010000100",
  10533=>"000010110",
  10534=>"000001001",
  10535=>"011111000",
  10536=>"010100110",
  10537=>"001011100",
  10538=>"110011010",
  10539=>"000010010",
  10540=>"101101011",
  10541=>"000010000",
  10542=>"001001110",
  10543=>"111110111",
  10544=>"000101010",
  10545=>"101101010",
  10546=>"001001001",
  10547=>"011101011",
  10548=>"101010110",
  10549=>"000101110",
  10550=>"101000000",
  10551=>"100101100",
  10552=>"111000101",
  10553=>"101000100",
  10554=>"101000100",
  10555=>"010010001",
  10556=>"110101111",
  10557=>"101001011",
  10558=>"000010111",
  10559=>"000011011",
  10560=>"100000001",
  10561=>"100110110",
  10562=>"011001001",
  10563=>"001110100",
  10564=>"000101100",
  10565=>"000100000",
  10566=>"000001100",
  10567=>"110111010",
  10568=>"010010100",
  10569=>"111010010",
  10570=>"011101100",
  10571=>"100100000",
  10572=>"011111000",
  10573=>"110101111",
  10574=>"000001100",
  10575=>"000111100",
  10576=>"011101001",
  10577=>"111110101",
  10578=>"000101000",
  10579=>"001010000",
  10580=>"000000100",
  10581=>"001011001",
  10582=>"100001110",
  10583=>"001100001",
  10584=>"011001100",
  10585=>"011010110",
  10586=>"010010001",
  10587=>"110010100",
  10588=>"100000011",
  10589=>"111001111",
  10590=>"011111110",
  10591=>"111011110",
  10592=>"100111001",
  10593=>"110010111",
  10594=>"010110011",
  10595=>"010001011",
  10596=>"101111100",
  10597=>"000100000",
  10598=>"111011111",
  10599=>"001100010",
  10600=>"010110111",
  10601=>"001010000",
  10602=>"110110110",
  10603=>"100101111",
  10604=>"011111101",
  10605=>"001101110",
  10606=>"101010000",
  10607=>"011111101",
  10608=>"011100110",
  10609=>"101000000",
  10610=>"011010011",
  10611=>"111001011",
  10612=>"001101110",
  10613=>"111100001",
  10614=>"010010101",
  10615=>"111101111",
  10616=>"000100010",
  10617=>"001011110",
  10618=>"101000110",
  10619=>"100010010",
  10620=>"010010001",
  10621=>"110100010",
  10622=>"111101101",
  10623=>"010101101",
  10624=>"111000001",
  10625=>"100000000",
  10626=>"001110000",
  10627=>"111011001",
  10628=>"011010101",
  10629=>"101101010",
  10630=>"010100110",
  10631=>"010101100",
  10632=>"010101100",
  10633=>"011011000",
  10634=>"111111010",
  10635=>"110101100",
  10636=>"010111110",
  10637=>"101010010",
  10638=>"000011100",
  10639=>"010011000",
  10640=>"000110000",
  10641=>"111111101",
  10642=>"111110100",
  10643=>"111011000",
  10644=>"000011001",
  10645=>"001000010",
  10646=>"011111000",
  10647=>"011100111",
  10648=>"110001001",
  10649=>"000100111",
  10650=>"111010000",
  10651=>"001011100",
  10652=>"001110000",
  10653=>"011011101",
  10654=>"000100110",
  10655=>"010010110",
  10656=>"001011000",
  10657=>"010101111",
  10658=>"000101111",
  10659=>"110100000",
  10660=>"110111010",
  10661=>"101010000",
  10662=>"110000110",
  10663=>"101110110",
  10664=>"100011111",
  10665=>"000101001",
  10666=>"001001001",
  10667=>"111011011",
  10668=>"010111111",
  10669=>"000011101",
  10670=>"001011011",
  10671=>"100100100",
  10672=>"111011111",
  10673=>"111111101",
  10674=>"000000101",
  10675=>"111100010",
  10676=>"010101111",
  10677=>"101011011",
  10678=>"101000000",
  10679=>"001010011",
  10680=>"000011110",
  10681=>"100101011",
  10682=>"111100111",
  10683=>"001111001",
  10684=>"011110111",
  10685=>"110000001",
  10686=>"011010011",
  10687=>"100000011",
  10688=>"010100010",
  10689=>"111000100",
  10690=>"110101111",
  10691=>"101111011",
  10692=>"111010110",
  10693=>"010000100",
  10694=>"000100100",
  10695=>"000010111",
  10696=>"011011100",
  10697=>"001101100",
  10698=>"110001000",
  10699=>"100000011",
  10700=>"100110111",
  10701=>"001111011",
  10702=>"100010001",
  10703=>"010001101",
  10704=>"010001111",
  10705=>"110011010",
  10706=>"111001011",
  10707=>"110011111",
  10708=>"011000110",
  10709=>"000110100",
  10710=>"010000011",
  10711=>"001011100",
  10712=>"111101001",
  10713=>"011000101",
  10714=>"110110000",
  10715=>"011001111",
  10716=>"111101100",
  10717=>"100110100",
  10718=>"110010110",
  10719=>"010111100",
  10720=>"010010100",
  10721=>"001011010",
  10722=>"000010011",
  10723=>"001011110",
  10724=>"011101111",
  10725=>"101111011",
  10726=>"111000001",
  10727=>"100111111",
  10728=>"101010111",
  10729=>"100010001",
  10730=>"001101010",
  10731=>"111001011",
  10732=>"000010100",
  10733=>"011111000",
  10734=>"010001010",
  10735=>"101011011",
  10736=>"101000101",
  10737=>"111110011",
  10738=>"001000001",
  10739=>"011010010",
  10740=>"000010111",
  10741=>"001101101",
  10742=>"010000101",
  10743=>"101010100",
  10744=>"110110010",
  10745=>"111110011",
  10746=>"011101110",
  10747=>"100010001",
  10748=>"111111000",
  10749=>"110000010",
  10750=>"101111011",
  10751=>"000011000",
  10752=>"111010101",
  10753=>"100001101",
  10754=>"100000011",
  10755=>"000000011",
  10756=>"101110010",
  10757=>"110001100",
  10758=>"111111001",
  10759=>"000100000",
  10760=>"100101011",
  10761=>"100111111",
  10762=>"110011110",
  10763=>"001000100",
  10764=>"001000100",
  10765=>"001011001",
  10766=>"010111100",
  10767=>"101000011",
  10768=>"001011110",
  10769=>"100000011",
  10770=>"010100111",
  10771=>"010110111",
  10772=>"111010111",
  10773=>"001110010",
  10774=>"011000110",
  10775=>"010100001",
  10776=>"111010111",
  10777=>"011011001",
  10778=>"101100000",
  10779=>"011100111",
  10780=>"111110101",
  10781=>"010001000",
  10782=>"101100001",
  10783=>"011010110",
  10784=>"000010000",
  10785=>"001101111",
  10786=>"000100111",
  10787=>"101001101",
  10788=>"011010000",
  10789=>"101101101",
  10790=>"110110011",
  10791=>"000010101",
  10792=>"100010010",
  10793=>"101000011",
  10794=>"101110111",
  10795=>"100100100",
  10796=>"101111000",
  10797=>"111000011",
  10798=>"000011011",
  10799=>"100110110",
  10800=>"101101110",
  10801=>"011000111",
  10802=>"011001001",
  10803=>"111001101",
  10804=>"001110001",
  10805=>"010011100",
  10806=>"101000101",
  10807=>"111100110",
  10808=>"000101111",
  10809=>"111100110",
  10810=>"100111000",
  10811=>"101101100",
  10812=>"100111110",
  10813=>"101011101",
  10814=>"011001011",
  10815=>"000100101",
  10816=>"110011101",
  10817=>"111011101",
  10818=>"000010001",
  10819=>"100001101",
  10820=>"101011011",
  10821=>"111110000",
  10822=>"001111101",
  10823=>"100110011",
  10824=>"001100010",
  10825=>"100111011",
  10826=>"011001001",
  10827=>"010111001",
  10828=>"110001100",
  10829=>"110101101",
  10830=>"110101011",
  10831=>"000100101",
  10832=>"000010010",
  10833=>"111110111",
  10834=>"101100101",
  10835=>"110011011",
  10836=>"000001011",
  10837=>"111010000",
  10838=>"101011100",
  10839=>"001010100",
  10840=>"110000011",
  10841=>"000010011",
  10842=>"011100101",
  10843=>"010101110",
  10844=>"111111100",
  10845=>"110101010",
  10846=>"000110101",
  10847=>"100110001",
  10848=>"001110100",
  10849=>"111010100",
  10850=>"010101000",
  10851=>"011011101",
  10852=>"100100101",
  10853=>"011011110",
  10854=>"010101000",
  10855=>"001110010",
  10856=>"000000110",
  10857=>"100100010",
  10858=>"001111110",
  10859=>"001000101",
  10860=>"001011000",
  10861=>"010111010",
  10862=>"000010000",
  10863=>"110110000",
  10864=>"011101001",
  10865=>"110110000",
  10866=>"110100011",
  10867=>"001011000",
  10868=>"110001001",
  10869=>"011100011",
  10870=>"010100101",
  10871=>"010011000",
  10872=>"111000110",
  10873=>"101110011",
  10874=>"000010000",
  10875=>"001111011",
  10876=>"010011111",
  10877=>"010110010",
  10878=>"001101001",
  10879=>"100010011",
  10880=>"000101101",
  10881=>"001111000",
  10882=>"001101001",
  10883=>"011011010",
  10884=>"000100111",
  10885=>"011110010",
  10886=>"011001101",
  10887=>"010110010",
  10888=>"101011000",
  10889=>"110111011",
  10890=>"010101101",
  10891=>"100001000",
  10892=>"101000010",
  10893=>"011010001",
  10894=>"011111010",
  10895=>"011110110",
  10896=>"110100101",
  10897=>"001100100",
  10898=>"011110000",
  10899=>"011111111",
  10900=>"111110111",
  10901=>"001000010",
  10902=>"111101010",
  10903=>"000101101",
  10904=>"111000010",
  10905=>"111101111",
  10906=>"011100110",
  10907=>"111111001",
  10908=>"000000000",
  10909=>"110111010",
  10910=>"111011100",
  10911=>"010001101",
  10912=>"101001001",
  10913=>"010001000",
  10914=>"111000001",
  10915=>"010001010",
  10916=>"110111100",
  10917=>"000010100",
  10918=>"010101010",
  10919=>"111011000",
  10920=>"001011111",
  10921=>"011011111",
  10922=>"110010110",
  10923=>"001011101",
  10924=>"011000110",
  10925=>"111000100",
  10926=>"000011110",
  10927=>"110010010",
  10928=>"011000011",
  10929=>"101110110",
  10930=>"011011111",
  10931=>"111100111",
  10932=>"011100111",
  10933=>"111101111",
  10934=>"011011101",
  10935=>"001100000",
  10936=>"000011111",
  10937=>"010010111",
  10938=>"100100001",
  10939=>"010110110",
  10940=>"110001110",
  10941=>"101100111",
  10942=>"001000000",
  10943=>"111100101",
  10944=>"100001011",
  10945=>"010101100",
  10946=>"110100100",
  10947=>"010111010",
  10948=>"110101000",
  10949=>"100110110",
  10950=>"111010100",
  10951=>"001101100",
  10952=>"100100000",
  10953=>"000011100",
  10954=>"001000101",
  10955=>"111110110",
  10956=>"001011111",
  10957=>"110110111",
  10958=>"111111111",
  10959=>"000100000",
  10960=>"010101110",
  10961=>"011111101",
  10962=>"010111010",
  10963=>"000101101",
  10964=>"101110011",
  10965=>"001010000",
  10966=>"101010011",
  10967=>"010101101",
  10968=>"100000111",
  10969=>"110110100",
  10970=>"000100000",
  10971=>"100011100",
  10972=>"111001100",
  10973=>"010011100",
  10974=>"111000101",
  10975=>"011111001",
  10976=>"100001111",
  10977=>"110111110",
  10978=>"110101100",
  10979=>"011001010",
  10980=>"000111011",
  10981=>"111010010",
  10982=>"111101101",
  10983=>"111110110",
  10984=>"111011111",
  10985=>"000001001",
  10986=>"110101001",
  10987=>"111111111",
  10988=>"000001011",
  10989=>"010011010",
  10990=>"000011100",
  10991=>"010110010",
  10992=>"000000011",
  10993=>"111001000",
  10994=>"010101011",
  10995=>"101001100",
  10996=>"101101001",
  10997=>"101011100",
  10998=>"001010110",
  10999=>"111101110",
  11000=>"001101100",
  11001=>"100111110",
  11002=>"110101010",
  11003=>"001100000",
  11004=>"100011101",
  11005=>"010101011",
  11006=>"101111100",
  11007=>"001000110",
  11008=>"001110111",
  11009=>"110000001",
  11010=>"110110011",
  11011=>"100011010",
  11012=>"110101111",
  11013=>"000001001",
  11014=>"000001001",
  11015=>"010111000",
  11016=>"101100101",
  11017=>"101010111",
  11018=>"110110011",
  11019=>"110010001",
  11020=>"100001011",
  11021=>"100001111",
  11022=>"110110101",
  11023=>"000010100",
  11024=>"100000011",
  11025=>"001001111",
  11026=>"111110100",
  11027=>"000110101",
  11028=>"011000000",
  11029=>"111111000",
  11030=>"101001001",
  11031=>"101110011",
  11032=>"101111100",
  11033=>"001101100",
  11034=>"000001010",
  11035=>"000010000",
  11036=>"001100001",
  11037=>"011000101",
  11038=>"000101010",
  11039=>"101001010",
  11040=>"000101110",
  11041=>"100111110",
  11042=>"001111001",
  11043=>"101110011",
  11044=>"010011101",
  11045=>"001001001",
  11046=>"100100001",
  11047=>"100010111",
  11048=>"000010101",
  11049=>"101110100",
  11050=>"110111110",
  11051=>"000010111",
  11052=>"110110000",
  11053=>"000100011",
  11054=>"011111111",
  11055=>"100110111",
  11056=>"000010010",
  11057=>"110100111",
  11058=>"001001011",
  11059=>"110110110",
  11060=>"011001101",
  11061=>"111101001",
  11062=>"011111010",
  11063=>"100111110",
  11064=>"000001100",
  11065=>"100110010",
  11066=>"111111111",
  11067=>"101100001",
  11068=>"011000011",
  11069=>"100000000",
  11070=>"111001000",
  11071=>"001000110",
  11072=>"000000010",
  11073=>"111000101",
  11074=>"001110011",
  11075=>"110011000",
  11076=>"001101000",
  11077=>"000001110",
  11078=>"101011101",
  11079=>"001000000",
  11080=>"001000000",
  11081=>"110111111",
  11082=>"111001010",
  11083=>"010011111",
  11084=>"101001100",
  11085=>"100111001",
  11086=>"010100001",
  11087=>"111010000",
  11088=>"001111101",
  11089=>"011011010",
  11090=>"010010000",
  11091=>"010111000",
  11092=>"101111011",
  11093=>"110001010",
  11094=>"111010010",
  11095=>"011011000",
  11096=>"100000001",
  11097=>"010110011",
  11098=>"001100110",
  11099=>"001011000",
  11100=>"110010101",
  11101=>"100100000",
  11102=>"010100010",
  11103=>"011011111",
  11104=>"111001110",
  11105=>"101010001",
  11106=>"000110010",
  11107=>"000101011",
  11108=>"001101001",
  11109=>"110111100",
  11110=>"111010010",
  11111=>"001011101",
  11112=>"110010001",
  11113=>"110011110",
  11114=>"101101100",
  11115=>"001000111",
  11116=>"010111111",
  11117=>"010111111",
  11118=>"010101011",
  11119=>"111111111",
  11120=>"110010111",
  11121=>"001111010",
  11122=>"001010010",
  11123=>"101000110",
  11124=>"001100000",
  11125=>"111000000",
  11126=>"101100100",
  11127=>"001010000",
  11128=>"011110000",
  11129=>"000010010",
  11130=>"110111100",
  11131=>"100010100",
  11132=>"010001110",
  11133=>"000111011",
  11134=>"111101010",
  11135=>"111100110",
  11136=>"010111110",
  11137=>"110011100",
  11138=>"011100001",
  11139=>"111000011",
  11140=>"110000001",
  11141=>"111101010",
  11142=>"110100110",
  11143=>"110011001",
  11144=>"000001000",
  11145=>"111110010",
  11146=>"011011011",
  11147=>"111101100",
  11148=>"101101110",
  11149=>"010100001",
  11150=>"011111001",
  11151=>"000010010",
  11152=>"110010000",
  11153=>"011010111",
  11154=>"010110000",
  11155=>"001110000",
  11156=>"101110100",
  11157=>"111101110",
  11158=>"100101101",
  11159=>"001011111",
  11160=>"001101111",
  11161=>"011011100",
  11162=>"100001101",
  11163=>"100101111",
  11164=>"011011111",
  11165=>"111111111",
  11166=>"010000001",
  11167=>"111100101",
  11168=>"011001000",
  11169=>"101111110",
  11170=>"100100010",
  11171=>"011110011",
  11172=>"001001000",
  11173=>"100100010",
  11174=>"010100011",
  11175=>"001001101",
  11176=>"111011110",
  11177=>"111001111",
  11178=>"101000011",
  11179=>"110101010",
  11180=>"001001011",
  11181=>"101011000",
  11182=>"100000001",
  11183=>"001110110",
  11184=>"101011001",
  11185=>"010111011",
  11186=>"100001000",
  11187=>"000010001",
  11188=>"000110100",
  11189=>"111001010",
  11190=>"101000010",
  11191=>"100100100",
  11192=>"011000010",
  11193=>"000100101",
  11194=>"111101000",
  11195=>"100100111",
  11196=>"110100100",
  11197=>"011000001",
  11198=>"011011001",
  11199=>"010100001",
  11200=>"101010100",
  11201=>"000000100",
  11202=>"110100001",
  11203=>"110010011",
  11204=>"000110010",
  11205=>"011110100",
  11206=>"111011011",
  11207=>"100000000",
  11208=>"001101010",
  11209=>"110001011",
  11210=>"011110001",
  11211=>"001011000",
  11212=>"111011011",
  11213=>"110010001",
  11214=>"110110000",
  11215=>"011011010",
  11216=>"100100110",
  11217=>"011000000",
  11218=>"001110111",
  11219=>"000000100",
  11220=>"000101111",
  11221=>"011100001",
  11222=>"010000100",
  11223=>"001100101",
  11224=>"111010001",
  11225=>"100010010",
  11226=>"011011000",
  11227=>"100101010",
  11228=>"111001100",
  11229=>"100001111",
  11230=>"000101111",
  11231=>"010110001",
  11232=>"010111011",
  11233=>"111101011",
  11234=>"111001100",
  11235=>"100110001",
  11236=>"100100001",
  11237=>"000011100",
  11238=>"000011110",
  11239=>"100001110",
  11240=>"000100101",
  11241=>"100000010",
  11242=>"111100011",
  11243=>"110011000",
  11244=>"011001111",
  11245=>"110001100",
  11246=>"001100100",
  11247=>"001110101",
  11248=>"011100011",
  11249=>"011000010",
  11250=>"001110111",
  11251=>"100011110",
  11252=>"000000110",
  11253=>"101010010",
  11254=>"000010010",
  11255=>"011111101",
  11256=>"100110100",
  11257=>"001000111",
  11258=>"011101110",
  11259=>"000100000",
  11260=>"111001010",
  11261=>"001000101",
  11262=>"100101001",
  11263=>"010111011",
  11264=>"101111100",
  11265=>"100110111",
  11266=>"110101111",
  11267=>"010000101",
  11268=>"111110000",
  11269=>"001011001",
  11270=>"010100001",
  11271=>"100011010",
  11272=>"110101000",
  11273=>"110111000",
  11274=>"010011100",
  11275=>"001110010",
  11276=>"011000100",
  11277=>"001111000",
  11278=>"010001011",
  11279=>"010000110",
  11280=>"011001010",
  11281=>"100101110",
  11282=>"101011110",
  11283=>"101011101",
  11284=>"001111100",
  11285=>"100110100",
  11286=>"011011010",
  11287=>"111100010",
  11288=>"010111111",
  11289=>"001011000",
  11290=>"100001010",
  11291=>"001011001",
  11292=>"000001001",
  11293=>"001010100",
  11294=>"000100110",
  11295=>"001001011",
  11296=>"000100000",
  11297=>"100111011",
  11298=>"000110011",
  11299=>"110100110",
  11300=>"001011101",
  11301=>"111001010",
  11302=>"011111011",
  11303=>"011111000",
  11304=>"011100010",
  11305=>"001101101",
  11306=>"000011101",
  11307=>"011010001",
  11308=>"110101111",
  11309=>"011110001",
  11310=>"010101111",
  11311=>"111000010",
  11312=>"000001001",
  11313=>"001011011",
  11314=>"000000000",
  11315=>"110100100",
  11316=>"100100110",
  11317=>"001100010",
  11318=>"101110101",
  11319=>"100001000",
  11320=>"000110111",
  11321=>"110000100",
  11322=>"000100101",
  11323=>"100110001",
  11324=>"010100000",
  11325=>"111111110",
  11326=>"101011110",
  11327=>"010000010",
  11328=>"111001110",
  11329=>"111100010",
  11330=>"111011101",
  11331=>"011000001",
  11332=>"111111100",
  11333=>"011010010",
  11334=>"000011100",
  11335=>"000110111",
  11336=>"010000011",
  11337=>"011001100",
  11338=>"110111011",
  11339=>"100010100",
  11340=>"001100110",
  11341=>"011110100",
  11342=>"010101010",
  11343=>"100100000",
  11344=>"101000111",
  11345=>"010011011",
  11346=>"100011000",
  11347=>"111001110",
  11348=>"000001111",
  11349=>"000010111",
  11350=>"100011110",
  11351=>"111001010",
  11352=>"111001011",
  11353=>"000001001",
  11354=>"100000111",
  11355=>"011001000",
  11356=>"111101001",
  11357=>"010110011",
  11358=>"110011000",
  11359=>"001001011",
  11360=>"001101010",
  11361=>"100011011",
  11362=>"101000111",
  11363=>"000000101",
  11364=>"011101101",
  11365=>"111011000",
  11366=>"110111101",
  11367=>"000101100",
  11368=>"101011101",
  11369=>"101000000",
  11370=>"111101110",
  11371=>"111101110",
  11372=>"000101100",
  11373=>"101001101",
  11374=>"001110011",
  11375=>"000111110",
  11376=>"010011011",
  11377=>"100110000",
  11378=>"111100101",
  11379=>"000010101",
  11380=>"000001011",
  11381=>"111110101",
  11382=>"111100100",
  11383=>"100110011",
  11384=>"100010001",
  11385=>"101001011",
  11386=>"110111100",
  11387=>"001100011",
  11388=>"000010000",
  11389=>"100100111",
  11390=>"111100111",
  11391=>"100010000",
  11392=>"001100110",
  11393=>"100110010",
  11394=>"101010000",
  11395=>"100100011",
  11396=>"110111100",
  11397=>"110010111",
  11398=>"001101100",
  11399=>"011000010",
  11400=>"100000101",
  11401=>"001110001",
  11402=>"001000011",
  11403=>"110011100",
  11404=>"000011101",
  11405=>"011101110",
  11406=>"001101101",
  11407=>"100100001",
  11408=>"001100001",
  11409=>"011010000",
  11410=>"111001100",
  11411=>"000111100",
  11412=>"010001111",
  11413=>"010011001",
  11414=>"011010110",
  11415=>"100010101",
  11416=>"101001000",
  11417=>"111111100",
  11418=>"000011110",
  11419=>"100000011",
  11420=>"001101010",
  11421=>"110110010",
  11422=>"111010101",
  11423=>"000100011",
  11424=>"010011101",
  11425=>"111011011",
  11426=>"001000101",
  11427=>"111011100",
  11428=>"111111010",
  11429=>"011000001",
  11430=>"101101111",
  11431=>"011101110",
  11432=>"111101111",
  11433=>"101001010",
  11434=>"000111110",
  11435=>"001101110",
  11436=>"010000010",
  11437=>"100111111",
  11438=>"100110111",
  11439=>"101111110",
  11440=>"101010011",
  11441=>"010101000",
  11442=>"011100001",
  11443=>"010010010",
  11444=>"000111000",
  11445=>"000000111",
  11446=>"001111010",
  11447=>"010101000",
  11448=>"101010100",
  11449=>"010011010",
  11450=>"010000100",
  11451=>"000101001",
  11452=>"101010010",
  11453=>"100001010",
  11454=>"011001111",
  11455=>"010100000",
  11456=>"010110011",
  11457=>"010001101",
  11458=>"101010001",
  11459=>"110011001",
  11460=>"000000111",
  11461=>"010000110",
  11462=>"001101000",
  11463=>"101010110",
  11464=>"000111010",
  11465=>"011111011",
  11466=>"011110001",
  11467=>"001110011",
  11468=>"010011111",
  11469=>"111110000",
  11470=>"110110001",
  11471=>"000101011",
  11472=>"000000100",
  11473=>"001010100",
  11474=>"011110011",
  11475=>"000011111",
  11476=>"101000110",
  11477=>"100001101",
  11478=>"111001001",
  11479=>"010011110",
  11480=>"000000101",
  11481=>"100111001",
  11482=>"100110011",
  11483=>"010010001",
  11484=>"110100010",
  11485=>"000011000",
  11486=>"010011101",
  11487=>"010111010",
  11488=>"010110100",
  11489=>"000110100",
  11490=>"100101000",
  11491=>"110111101",
  11492=>"101100001",
  11493=>"101110010",
  11494=>"000101101",
  11495=>"100010101",
  11496=>"011101101",
  11497=>"101001101",
  11498=>"010011010",
  11499=>"000100011",
  11500=>"001010100",
  11501=>"011000101",
  11502=>"001100001",
  11503=>"000010000",
  11504=>"011100110",
  11505=>"100110010",
  11506=>"010000011",
  11507=>"001011110",
  11508=>"101110000",
  11509=>"011111110",
  11510=>"001000011",
  11511=>"010000110",
  11512=>"011001010",
  11513=>"101111101",
  11514=>"111000011",
  11515=>"001000010",
  11516=>"111111100",
  11517=>"001111000",
  11518=>"111101010",
  11519=>"110010111",
  11520=>"000111011",
  11521=>"101011111",
  11522=>"110001001",
  11523=>"000010100",
  11524=>"001111101",
  11525=>"111000000",
  11526=>"010001001",
  11527=>"010100010",
  11528=>"100100011",
  11529=>"000100000",
  11530=>"111101011",
  11531=>"110011101",
  11532=>"001001100",
  11533=>"111110001",
  11534=>"110010100",
  11535=>"001010110",
  11536=>"110101001",
  11537=>"110110010",
  11538=>"111111000",
  11539=>"110111001",
  11540=>"010111000",
  11541=>"000011101",
  11542=>"001011010",
  11543=>"010000011",
  11544=>"111100101",
  11545=>"111001010",
  11546=>"011101001",
  11547=>"000110110",
  11548=>"110101011",
  11549=>"100010100",
  11550=>"100010110",
  11551=>"111001001",
  11552=>"000101000",
  11553=>"000011110",
  11554=>"100000101",
  11555=>"001000101",
  11556=>"101100011",
  11557=>"100011011",
  11558=>"110101111",
  11559=>"011101100",
  11560=>"001111101",
  11561=>"001001000",
  11562=>"001111010",
  11563=>"000010100",
  11564=>"010010010",
  11565=>"101000001",
  11566=>"000001100",
  11567=>"000011101",
  11568=>"000001010",
  11569=>"110100101",
  11570=>"101100000",
  11571=>"100101010",
  11572=>"001010010",
  11573=>"010000001",
  11574=>"000010110",
  11575=>"011111001",
  11576=>"000011010",
  11577=>"110101100",
  11578=>"111101101",
  11579=>"011110111",
  11580=>"011001101",
  11581=>"111111101",
  11582=>"111000001",
  11583=>"000000010",
  11584=>"100110010",
  11585=>"001000110",
  11586=>"000101010",
  11587=>"110111010",
  11588=>"011100001",
  11589=>"101110001",
  11590=>"110000010",
  11591=>"111101111",
  11592=>"000000100",
  11593=>"010110010",
  11594=>"011001001",
  11595=>"001000000",
  11596=>"011000100",
  11597=>"101011001",
  11598=>"111111011",
  11599=>"000101000",
  11600=>"000001100",
  11601=>"110001110",
  11602=>"111010111",
  11603=>"110101001",
  11604=>"100110001",
  11605=>"101000110",
  11606=>"001111101",
  11607=>"011000000",
  11608=>"100100111",
  11609=>"000011100",
  11610=>"001011011",
  11611=>"001000111",
  11612=>"010010101",
  11613=>"110001000",
  11614=>"110010000",
  11615=>"100111011",
  11616=>"011000011",
  11617=>"000000011",
  11618=>"101101110",
  11619=>"101000110",
  11620=>"000000110",
  11621=>"100100000",
  11622=>"010100011",
  11623=>"100001010",
  11624=>"111101101",
  11625=>"000100100",
  11626=>"011000111",
  11627=>"000000001",
  11628=>"100101010",
  11629=>"010101101",
  11630=>"100111001",
  11631=>"000100010",
  11632=>"100001101",
  11633=>"000100111",
  11634=>"111111110",
  11635=>"110010111",
  11636=>"001110100",
  11637=>"100001001",
  11638=>"000000111",
  11639=>"000100011",
  11640=>"010100110",
  11641=>"100111011",
  11642=>"000011011",
  11643=>"101100101",
  11644=>"000101110",
  11645=>"001000111",
  11646=>"000011000",
  11647=>"101000010",
  11648=>"110101110",
  11649=>"101110000",
  11650=>"011101011",
  11651=>"111111010",
  11652=>"111100100",
  11653=>"110101010",
  11654=>"000010111",
  11655=>"111100101",
  11656=>"010001000",
  11657=>"110110010",
  11658=>"010010110",
  11659=>"101010011",
  11660=>"111101101",
  11661=>"001000011",
  11662=>"001101000",
  11663=>"010001010",
  11664=>"110000101",
  11665=>"010000111",
  11666=>"100001100",
  11667=>"100100100",
  11668=>"011110000",
  11669=>"010111101",
  11670=>"100011001",
  11671=>"000100001",
  11672=>"110110111",
  11673=>"010100001",
  11674=>"111101110",
  11675=>"000000000",
  11676=>"001111111",
  11677=>"111110000",
  11678=>"110100010",
  11679=>"000100111",
  11680=>"000000100",
  11681=>"110001100",
  11682=>"000111111",
  11683=>"001101001",
  11684=>"010110101",
  11685=>"110000000",
  11686=>"001000100",
  11687=>"100010100",
  11688=>"000100110",
  11689=>"001110100",
  11690=>"101011101",
  11691=>"000001000",
  11692=>"011100010",
  11693=>"010100000",
  11694=>"000110001",
  11695=>"101111101",
  11696=>"011000001",
  11697=>"111001000",
  11698=>"101010011",
  11699=>"010111001",
  11700=>"101101000",
  11701=>"110110000",
  11702=>"010010010",
  11703=>"010111101",
  11704=>"100111000",
  11705=>"101110011",
  11706=>"101111101",
  11707=>"001110011",
  11708=>"010110001",
  11709=>"011001010",
  11710=>"100101000",
  11711=>"010010111",
  11712=>"011000101",
  11713=>"010001100",
  11714=>"001110101",
  11715=>"100000000",
  11716=>"110000110",
  11717=>"110000110",
  11718=>"010000100",
  11719=>"000110101",
  11720=>"101000000",
  11721=>"000000101",
  11722=>"001101011",
  11723=>"011110100",
  11724=>"000110110",
  11725=>"000111100",
  11726=>"000010011",
  11727=>"011010001",
  11728=>"100010101",
  11729=>"110001011",
  11730=>"010001111",
  11731=>"011110010",
  11732=>"000010001",
  11733=>"000110011",
  11734=>"110010001",
  11735=>"001110111",
  11736=>"010010110",
  11737=>"011010000",
  11738=>"101100000",
  11739=>"111111111",
  11740=>"110000101",
  11741=>"010111111",
  11742=>"101010000",
  11743=>"111111011",
  11744=>"110100101",
  11745=>"010110010",
  11746=>"011111110",
  11747=>"000110000",
  11748=>"011110010",
  11749=>"110010101",
  11750=>"011111110",
  11751=>"110010111",
  11752=>"010110111",
  11753=>"001010010",
  11754=>"110101001",
  11755=>"001001000",
  11756=>"010011000",
  11757=>"101011111",
  11758=>"010011110",
  11759=>"000010101",
  11760=>"011000001",
  11761=>"100111011",
  11762=>"100110000",
  11763=>"000100000",
  11764=>"011000100",
  11765=>"001100101",
  11766=>"000000101",
  11767=>"010101100",
  11768=>"001100000",
  11769=>"100001110",
  11770=>"100000000",
  11771=>"011101010",
  11772=>"110001111",
  11773=>"010010100",
  11774=>"111011111",
  11775=>"000000111",
  11776=>"001010000",
  11777=>"100001011",
  11778=>"000010000",
  11779=>"001100111",
  11780=>"000010001",
  11781=>"010111010",
  11782=>"000000001",
  11783=>"000100111",
  11784=>"011011010",
  11785=>"111100011",
  11786=>"110001101",
  11787=>"000100010",
  11788=>"111011110",
  11789=>"011011111",
  11790=>"111011110",
  11791=>"111111110",
  11792=>"010001011",
  11793=>"101110111",
  11794=>"000100111",
  11795=>"000100110",
  11796=>"101011101",
  11797=>"001000000",
  11798=>"111000111",
  11799=>"111011111",
  11800=>"100010001",
  11801=>"000000010",
  11802=>"010010011",
  11803=>"010100010",
  11804=>"100001111",
  11805=>"110001110",
  11806=>"111000101",
  11807=>"100101111",
  11808=>"111001111",
  11809=>"001101111",
  11810=>"101010010",
  11811=>"101110011",
  11812=>"101111000",
  11813=>"110010000",
  11814=>"011000001",
  11815=>"111001101",
  11816=>"101100000",
  11817=>"111110111",
  11818=>"101100111",
  11819=>"000000011",
  11820=>"110011001",
  11821=>"001011110",
  11822=>"001011000",
  11823=>"101101110",
  11824=>"111001001",
  11825=>"100111011",
  11826=>"000001000",
  11827=>"101011111",
  11828=>"001000101",
  11829=>"101010000",
  11830=>"010001000",
  11831=>"100101000",
  11832=>"100011101",
  11833=>"110011100",
  11834=>"111011100",
  11835=>"010110110",
  11836=>"111110100",
  11837=>"000011100",
  11838=>"111100011",
  11839=>"110000101",
  11840=>"011001001",
  11841=>"001000101",
  11842=>"110001010",
  11843=>"010010000",
  11844=>"001110111",
  11845=>"010100011",
  11846=>"101000100",
  11847=>"010011010",
  11848=>"100101000",
  11849=>"001100000",
  11850=>"101000010",
  11851=>"000100111",
  11852=>"110010010",
  11853=>"000010111",
  11854=>"001111100",
  11855=>"001001001",
  11856=>"100011010",
  11857=>"010001100",
  11858=>"100101111",
  11859=>"000000110",
  11860=>"100000111",
  11861=>"000101000",
  11862=>"111000011",
  11863=>"110101100",
  11864=>"111000011",
  11865=>"110110101",
  11866=>"011100001",
  11867=>"100001110",
  11868=>"010100001",
  11869=>"111000010",
  11870=>"100011000",
  11871=>"001000111",
  11872=>"100010100",
  11873=>"000010110",
  11874=>"110110101",
  11875=>"000110100",
  11876=>"010010000",
  11877=>"010101100",
  11878=>"111111110",
  11879=>"011010110",
  11880=>"000010001",
  11881=>"111110010",
  11882=>"111011110",
  11883=>"101000000",
  11884=>"011100011",
  11885=>"101101101",
  11886=>"010010011",
  11887=>"101101011",
  11888=>"000111111",
  11889=>"000011001",
  11890=>"001111110",
  11891=>"000000100",
  11892=>"010001110",
  11893=>"010001000",
  11894=>"101011011",
  11895=>"001101000",
  11896=>"010001100",
  11897=>"100100000",
  11898=>"000011001",
  11899=>"010101110",
  11900=>"011100111",
  11901=>"000111010",
  11902=>"011101001",
  11903=>"000011000",
  11904=>"000100000",
  11905=>"111111111",
  11906=>"001001110",
  11907=>"000010011",
  11908=>"111000100",
  11909=>"000000100",
  11910=>"011000110",
  11911=>"100100001",
  11912=>"101110000",
  11913=>"000010011",
  11914=>"101000010",
  11915=>"001110110",
  11916=>"110011001",
  11917=>"011101001",
  11918=>"000111110",
  11919=>"010101011",
  11920=>"110111010",
  11921=>"100111011",
  11922=>"110010001",
  11923=>"000111110",
  11924=>"101101010",
  11925=>"101110001",
  11926=>"010111110",
  11927=>"011000101",
  11928=>"101101111",
  11929=>"111100100",
  11930=>"001000000",
  11931=>"001001110",
  11932=>"111001011",
  11933=>"111111000",
  11934=>"101110001",
  11935=>"010001010",
  11936=>"011000101",
  11937=>"110100110",
  11938=>"100010101",
  11939=>"010110001",
  11940=>"111110111",
  11941=>"111011011",
  11942=>"001000000",
  11943=>"110000010",
  11944=>"110001111",
  11945=>"111000000",
  11946=>"001001110",
  11947=>"110001010",
  11948=>"000100001",
  11949=>"010110101",
  11950=>"111101100",
  11951=>"000110000",
  11952=>"111000100",
  11953=>"010001001",
  11954=>"000111010",
  11955=>"000101100",
  11956=>"001101111",
  11957=>"101111101",
  11958=>"000111111",
  11959=>"111011110",
  11960=>"001010011",
  11961=>"100111010",
  11962=>"010110011",
  11963=>"010101001",
  11964=>"100000001",
  11965=>"001000101",
  11966=>"110101011",
  11967=>"100110101",
  11968=>"011010101",
  11969=>"101011100",
  11970=>"110111111",
  11971=>"011011110",
  11972=>"011111000",
  11973=>"011001100",
  11974=>"101000111",
  11975=>"001101001",
  11976=>"101011100",
  11977=>"101011010",
  11978=>"011011000",
  11979=>"000111010",
  11980=>"011011111",
  11981=>"110000001",
  11982=>"110100110",
  11983=>"000100000",
  11984=>"011101111",
  11985=>"110000111",
  11986=>"010111111",
  11987=>"001001000",
  11988=>"111100011",
  11989=>"101010100",
  11990=>"001010011",
  11991=>"000101010",
  11992=>"000111101",
  11993=>"101001100",
  11994=>"010100110",
  11995=>"100000000",
  11996=>"000101010",
  11997=>"011110010",
  11998=>"010111010",
  11999=>"000110110",
  12000=>"001000100",
  12001=>"000111010",
  12002=>"010111000",
  12003=>"111101100",
  12004=>"000111111",
  12005=>"100100101",
  12006=>"001000011",
  12007=>"000011000",
  12008=>"010101110",
  12009=>"110010001",
  12010=>"110000111",
  12011=>"000000010",
  12012=>"100101011",
  12013=>"110010101",
  12014=>"011001011",
  12015=>"001110111",
  12016=>"110110111",
  12017=>"000111010",
  12018=>"000010100",
  12019=>"001101000",
  12020=>"111110011",
  12021=>"000101100",
  12022=>"100100100",
  12023=>"110001111",
  12024=>"010111111",
  12025=>"111110001",
  12026=>"100111110",
  12027=>"111011001",
  12028=>"011101110",
  12029=>"110111100",
  12030=>"000010010",
  12031=>"111110000",
  12032=>"010010101",
  12033=>"010100011",
  12034=>"011110001",
  12035=>"011101100",
  12036=>"100000010",
  12037=>"100001010",
  12038=>"001111110",
  12039=>"000100111",
  12040=>"001111100",
  12041=>"000000001",
  12042=>"001000100",
  12043=>"010100110",
  12044=>"101111101",
  12045=>"001100001",
  12046=>"110000011",
  12047=>"110101011",
  12048=>"011111110",
  12049=>"110010110",
  12050=>"000101010",
  12051=>"101111001",
  12052=>"011000111",
  12053=>"001111010",
  12054=>"100000111",
  12055=>"011000101",
  12056=>"111001111",
  12057=>"110010011",
  12058=>"010010110",
  12059=>"101001110",
  12060=>"110000100",
  12061=>"000111000",
  12062=>"011100000",
  12063=>"001110101",
  12064=>"110111010",
  12065=>"111001011",
  12066=>"000000010",
  12067=>"010100000",
  12068=>"101000101",
  12069=>"000010101",
  12070=>"000101011",
  12071=>"011000000",
  12072=>"111001100",
  12073=>"000111110",
  12074=>"111001011",
  12075=>"010110101",
  12076=>"010111110",
  12077=>"110000111",
  12078=>"010100101",
  12079=>"001111111",
  12080=>"111110110",
  12081=>"111011010",
  12082=>"110011010",
  12083=>"110000101",
  12084=>"100011101",
  12085=>"111100010",
  12086=>"100110100",
  12087=>"100110110",
  12088=>"111111010",
  12089=>"111111101",
  12090=>"110011101",
  12091=>"001110111",
  12092=>"001001110",
  12093=>"110110001",
  12094=>"010000010",
  12095=>"101100111",
  12096=>"111110010",
  12097=>"000000010",
  12098=>"000100001",
  12099=>"111010100",
  12100=>"111010111",
  12101=>"000110101",
  12102=>"011110101",
  12103=>"110100110",
  12104=>"110011001",
  12105=>"100000100",
  12106=>"000110111",
  12107=>"011100111",
  12108=>"011100110",
  12109=>"010101001",
  12110=>"000010101",
  12111=>"100001000",
  12112=>"001010101",
  12113=>"111000101",
  12114=>"100010001",
  12115=>"001000001",
  12116=>"000010101",
  12117=>"010110100",
  12118=>"010111110",
  12119=>"110101100",
  12120=>"001101100",
  12121=>"010011111",
  12122=>"000010100",
  12123=>"100000001",
  12124=>"011101011",
  12125=>"100101011",
  12126=>"011000100",
  12127=>"010000011",
  12128=>"100110111",
  12129=>"010100101",
  12130=>"100001111",
  12131=>"101001011",
  12132=>"100110000",
  12133=>"011011000",
  12134=>"011000110",
  12135=>"100101011",
  12136=>"101011101",
  12137=>"101101100",
  12138=>"001101101",
  12139=>"101000001",
  12140=>"101000001",
  12141=>"101000111",
  12142=>"111100000",
  12143=>"000001000",
  12144=>"000000100",
  12145=>"000111000",
  12146=>"011110001",
  12147=>"001000111",
  12148=>"011111101",
  12149=>"111100000",
  12150=>"000011100",
  12151=>"000001011",
  12152=>"110001001",
  12153=>"000111110",
  12154=>"111011000",
  12155=>"010101010",
  12156=>"110101110",
  12157=>"010101000",
  12158=>"000000111",
  12159=>"010010100",
  12160=>"011000011",
  12161=>"000111101",
  12162=>"110001110",
  12163=>"100100110",
  12164=>"000111000",
  12165=>"110010001",
  12166=>"101100001",
  12167=>"000000001",
  12168=>"110000101",
  12169=>"001000001",
  12170=>"010101001",
  12171=>"100001100",
  12172=>"100111010",
  12173=>"111110110",
  12174=>"010001000",
  12175=>"111110101",
  12176=>"111000100",
  12177=>"010001100",
  12178=>"101000000",
  12179=>"001100001",
  12180=>"101001011",
  12181=>"011111111",
  12182=>"111011111",
  12183=>"000101101",
  12184=>"001011111",
  12185=>"001110100",
  12186=>"000000001",
  12187=>"111110000",
  12188=>"110001001",
  12189=>"101100010",
  12190=>"010111101",
  12191=>"111001100",
  12192=>"001000001",
  12193=>"001011000",
  12194=>"001000100",
  12195=>"100001011",
  12196=>"011110101",
  12197=>"111001100",
  12198=>"100010100",
  12199=>"001011010",
  12200=>"100010010",
  12201=>"111001111",
  12202=>"001010101",
  12203=>"010000110",
  12204=>"001000100",
  12205=>"010001101",
  12206=>"001100010",
  12207=>"101110111",
  12208=>"110000100",
  12209=>"010101011",
  12210=>"000110100",
  12211=>"011111011",
  12212=>"111101101",
  12213=>"001111011",
  12214=>"101011110",
  12215=>"010001000",
  12216=>"000101101",
  12217=>"100001101",
  12218=>"000111000",
  12219=>"111010100",
  12220=>"001000000",
  12221=>"011110100",
  12222=>"110101111",
  12223=>"101010110",
  12224=>"101000010",
  12225=>"111000001",
  12226=>"010110011",
  12227=>"111000111",
  12228=>"010000010",
  12229=>"000000101",
  12230=>"111110111",
  12231=>"100000100",
  12232=>"011011100",
  12233=>"110100001",
  12234=>"110011001",
  12235=>"101100100",
  12236=>"110110011",
  12237=>"111000100",
  12238=>"010000100",
  12239=>"011000100",
  12240=>"111000000",
  12241=>"011000111",
  12242=>"011011000",
  12243=>"111110000",
  12244=>"101011100",
  12245=>"011110100",
  12246=>"000010011",
  12247=>"111001010",
  12248=>"100010111",
  12249=>"001100100",
  12250=>"011001100",
  12251=>"100000101",
  12252=>"000101100",
  12253=>"111111110",
  12254=>"011000010",
  12255=>"001000111",
  12256=>"100001000",
  12257=>"001110010",
  12258=>"010101001",
  12259=>"101100101",
  12260=>"000000011",
  12261=>"000100101",
  12262=>"000000011",
  12263=>"011000000",
  12264=>"100000000",
  12265=>"101000101",
  12266=>"001010111",
  12267=>"000110000",
  12268=>"001110100",
  12269=>"111101001",
  12270=>"101100100",
  12271=>"000110010",
  12272=>"000000110",
  12273=>"000010000",
  12274=>"101110001",
  12275=>"101100010",
  12276=>"000011000",
  12277=>"000000000",
  12278=>"000001111",
  12279=>"110001111",
  12280=>"000111110",
  12281=>"010011111",
  12282=>"000000111",
  12283=>"110111111",
  12284=>"111111101",
  12285=>"000101010",
  12286=>"101010100",
  12287=>"100011101",
  12288=>"110000100",
  12289=>"001010000",
  12290=>"100110100",
  12291=>"100010101",
  12292=>"111000100",
  12293=>"011011111",
  12294=>"111111111",
  12295=>"000111011",
  12296=>"110101111",
  12297=>"000000011",
  12298=>"010010000",
  12299=>"010110110",
  12300=>"110000011",
  12301=>"100001010",
  12302=>"111011111",
  12303=>"110100000",
  12304=>"111000100",
  12305=>"110110101",
  12306=>"010100100",
  12307=>"011010011",
  12308=>"010011100",
  12309=>"100110001",
  12310=>"001101110",
  12311=>"110110101",
  12312=>"101010111",
  12313=>"110001000",
  12314=>"011010000",
  12315=>"000010000",
  12316=>"011011101",
  12317=>"100101011",
  12318=>"100110010",
  12319=>"100110101",
  12320=>"011010111",
  12321=>"100011010",
  12322=>"010100001",
  12323=>"001011000",
  12324=>"010000101",
  12325=>"011111110",
  12326=>"011101101",
  12327=>"101011011",
  12328=>"010000111",
  12329=>"010010010",
  12330=>"000110010",
  12331=>"000001111",
  12332=>"111101010",
  12333=>"101111111",
  12334=>"001001011",
  12335=>"001000101",
  12336=>"000001000",
  12337=>"011101010",
  12338=>"110110000",
  12339=>"101000110",
  12340=>"100100110",
  12341=>"101001011",
  12342=>"001001100",
  12343=>"000111111",
  12344=>"011111011",
  12345=>"011000110",
  12346=>"100010101",
  12347=>"011111110",
  12348=>"001001100",
  12349=>"101001110",
  12350=>"101101100",
  12351=>"011101100",
  12352=>"011010010",
  12353=>"100000111",
  12354=>"000111110",
  12355=>"100000110",
  12356=>"011110011",
  12357=>"000011011",
  12358=>"010100100",
  12359=>"000010110",
  12360=>"011000110",
  12361=>"100011100",
  12362=>"100101101",
  12363=>"001000011",
  12364=>"010101110",
  12365=>"111001011",
  12366=>"010110001",
  12367=>"000100001",
  12368=>"100101000",
  12369=>"010100010",
  12370=>"110010111",
  12371=>"011101001",
  12372=>"000000100",
  12373=>"110101111",
  12374=>"011110000",
  12375=>"001001100",
  12376=>"000100110",
  12377=>"111110001",
  12378=>"111101010",
  12379=>"011000110",
  12380=>"110011110",
  12381=>"100111100",
  12382=>"001001011",
  12383=>"011011110",
  12384=>"000100000",
  12385=>"001010111",
  12386=>"000010111",
  12387=>"000011111",
  12388=>"000000111",
  12389=>"101101000",
  12390=>"001101011",
  12391=>"010000101",
  12392=>"001100111",
  12393=>"110111010",
  12394=>"000100111",
  12395=>"011010110",
  12396=>"011101011",
  12397=>"111001111",
  12398=>"111000000",
  12399=>"010111110",
  12400=>"011111000",
  12401=>"011101111",
  12402=>"000011001",
  12403=>"110111111",
  12404=>"101101100",
  12405=>"010000011",
  12406=>"000001111",
  12407=>"111101100",
  12408=>"011000111",
  12409=>"100111101",
  12410=>"101010011",
  12411=>"001011110",
  12412=>"010100000",
  12413=>"100111101",
  12414=>"001101110",
  12415=>"100111110",
  12416=>"101101110",
  12417=>"000011111",
  12418=>"110101011",
  12419=>"010101011",
  12420=>"111000101",
  12421=>"000011010",
  12422=>"011101010",
  12423=>"011011010",
  12424=>"001010111",
  12425=>"100000011",
  12426=>"000010010",
  12427=>"000111110",
  12428=>"000000111",
  12429=>"010100011",
  12430=>"001101110",
  12431=>"110001011",
  12432=>"000100100",
  12433=>"000110010",
  12434=>"000001101",
  12435=>"010101010",
  12436=>"010110100",
  12437=>"001100101",
  12438=>"110101101",
  12439=>"101110001",
  12440=>"101101111",
  12441=>"010100110",
  12442=>"110101001",
  12443=>"110100100",
  12444=>"111011111",
  12445=>"100010111",
  12446=>"001010011",
  12447=>"010100110",
  12448=>"001101100",
  12449=>"011001000",
  12450=>"001011100",
  12451=>"010110111",
  12452=>"111111011",
  12453=>"110111111",
  12454=>"101110100",
  12455=>"100111110",
  12456=>"100000101",
  12457=>"010101000",
  12458=>"101000001",
  12459=>"011101101",
  12460=>"001101110",
  12461=>"001001000",
  12462=>"110100101",
  12463=>"000000110",
  12464=>"101001011",
  12465=>"100000110",
  12466=>"001101101",
  12467=>"101101100",
  12468=>"000000100",
  12469=>"000000101",
  12470=>"000000100",
  12471=>"011011100",
  12472=>"011100000",
  12473=>"010001010",
  12474=>"110001111",
  12475=>"100101110",
  12476=>"110000111",
  12477=>"000010100",
  12478=>"111100100",
  12479=>"100110001",
  12480=>"111101011",
  12481=>"011000101",
  12482=>"110010100",
  12483=>"110111000",
  12484=>"000111000",
  12485=>"110100101",
  12486=>"001011010",
  12487=>"111110111",
  12488=>"100001011",
  12489=>"111011000",
  12490=>"010000010",
  12491=>"111001000",
  12492=>"011000010",
  12493=>"001000111",
  12494=>"110101110",
  12495=>"100100100",
  12496=>"010111110",
  12497=>"101011010",
  12498=>"010000000",
  12499=>"011111001",
  12500=>"101100101",
  12501=>"111010011",
  12502=>"101010111",
  12503=>"110011011",
  12504=>"001000111",
  12505=>"011101111",
  12506=>"100110101",
  12507=>"000101000",
  12508=>"101111000",
  12509=>"000010010",
  12510=>"110010011",
  12511=>"000000011",
  12512=>"000110110",
  12513=>"001000000",
  12514=>"110011101",
  12515=>"110001110",
  12516=>"010000011",
  12517=>"110010001",
  12518=>"110101001",
  12519=>"101001011",
  12520=>"100000101",
  12521=>"111111101",
  12522=>"101100100",
  12523=>"010000010",
  12524=>"111000011",
  12525=>"111100110",
  12526=>"000100011",
  12527=>"010001111",
  12528=>"110111101",
  12529=>"000001110",
  12530=>"110000111",
  12531=>"000000011",
  12532=>"001110000",
  12533=>"111110111",
  12534=>"101111011",
  12535=>"000101101",
  12536=>"110011111",
  12537=>"101110011",
  12538=>"111011110",
  12539=>"110011101",
  12540=>"010010111",
  12541=>"011100110",
  12542=>"111100110",
  12543=>"100000100",
  12544=>"101101001",
  12545=>"000110000",
  12546=>"111101010",
  12547=>"101011110",
  12548=>"011000110",
  12549=>"000010011",
  12550=>"000000000",
  12551=>"100011110",
  12552=>"111110100",
  12553=>"100011001",
  12554=>"100000001",
  12555=>"011101111",
  12556=>"001010110",
  12557=>"100111100",
  12558=>"000000010",
  12559=>"100010011",
  12560=>"111001101",
  12561=>"011001100",
  12562=>"011100111",
  12563=>"100110011",
  12564=>"111101011",
  12565=>"001101001",
  12566=>"110000110",
  12567=>"010110100",
  12568=>"011000011",
  12569=>"101100011",
  12570=>"001011010",
  12571=>"001000000",
  12572=>"011010110",
  12573=>"011010110",
  12574=>"111111100",
  12575=>"100110011",
  12576=>"010100010",
  12577=>"111110011",
  12578=>"101100011",
  12579=>"111100111",
  12580=>"000100000",
  12581=>"000000010",
  12582=>"000010111",
  12583=>"000110111",
  12584=>"011001101",
  12585=>"111110110",
  12586=>"101100100",
  12587=>"011110100",
  12588=>"111110001",
  12589=>"010101010",
  12590=>"010011110",
  12591=>"101101110",
  12592=>"111000110",
  12593=>"010111111",
  12594=>"010100101",
  12595=>"011000111",
  12596=>"100111000",
  12597=>"110101001",
  12598=>"110011100",
  12599=>"001110110",
  12600=>"010110000",
  12601=>"101100100",
  12602=>"101001101",
  12603=>"010000100",
  12604=>"101000110",
  12605=>"011011101",
  12606=>"010111000",
  12607=>"011001001",
  12608=>"001110001",
  12609=>"101110111",
  12610=>"101110001",
  12611=>"010111000",
  12612=>"010001101",
  12613=>"110101101",
  12614=>"010110000",
  12615=>"111001101",
  12616=>"001010101",
  12617=>"010101100",
  12618=>"000101110",
  12619=>"000100110",
  12620=>"001001001",
  12621=>"010100100",
  12622=>"101110011",
  12623=>"100100101",
  12624=>"011111011",
  12625=>"000111010",
  12626=>"111001100",
  12627=>"010110000",
  12628=>"010001111",
  12629=>"000010111",
  12630=>"101101100",
  12631=>"110101100",
  12632=>"011010000",
  12633=>"110001000",
  12634=>"110010111",
  12635=>"001010010",
  12636=>"010000100",
  12637=>"011011100",
  12638=>"010100010",
  12639=>"110011001",
  12640=>"010001110",
  12641=>"000010000",
  12642=>"011010010",
  12643=>"000100011",
  12644=>"110010111",
  12645=>"110011111",
  12646=>"000000101",
  12647=>"111000110",
  12648=>"101100101",
  12649=>"101000000",
  12650=>"101110010",
  12651=>"110011000",
  12652=>"000011101",
  12653=>"110010000",
  12654=>"001101100",
  12655=>"100100000",
  12656=>"101010000",
  12657=>"001001101",
  12658=>"010010101",
  12659=>"100110110",
  12660=>"100110111",
  12661=>"011001010",
  12662=>"100011010",
  12663=>"100101100",
  12664=>"010101101",
  12665=>"010001110",
  12666=>"000111001",
  12667=>"101010110",
  12668=>"101011101",
  12669=>"011101011",
  12670=>"101110110",
  12671=>"010110000",
  12672=>"010001100",
  12673=>"100000011",
  12674=>"001110100",
  12675=>"000000011",
  12676=>"001001001",
  12677=>"001011101",
  12678=>"001001100",
  12679=>"101000010",
  12680=>"110000000",
  12681=>"100000000",
  12682=>"101100011",
  12683=>"010100110",
  12684=>"000011101",
  12685=>"011101111",
  12686=>"110000110",
  12687=>"000010100",
  12688=>"001001111",
  12689=>"010001011",
  12690=>"011110000",
  12691=>"110000001",
  12692=>"101111111",
  12693=>"010000000",
  12694=>"010010111",
  12695=>"010010111",
  12696=>"000110001",
  12697=>"100000111",
  12698=>"011001000",
  12699=>"100101101",
  12700=>"011111011",
  12701=>"111011111",
  12702=>"001111010",
  12703=>"000110101",
  12704=>"000111110",
  12705=>"011111011",
  12706=>"010001010",
  12707=>"000101001",
  12708=>"110101011",
  12709=>"001011000",
  12710=>"101101000",
  12711=>"101001101",
  12712=>"111110010",
  12713=>"000101000",
  12714=>"001100001",
  12715=>"111110110",
  12716=>"110110010",
  12717=>"100000100",
  12718=>"000100001",
  12719=>"010001001",
  12720=>"100001110",
  12721=>"000001100",
  12722=>"011101011",
  12723=>"101011010",
  12724=>"101110010",
  12725=>"001010111",
  12726=>"110100100",
  12727=>"101110110",
  12728=>"011101010",
  12729=>"101000101",
  12730=>"000000111",
  12731=>"001001111",
  12732=>"100010101",
  12733=>"000000101",
  12734=>"100000011",
  12735=>"101001000",
  12736=>"001011001",
  12737=>"011000111",
  12738=>"100111001",
  12739=>"111001100",
  12740=>"011000011",
  12741=>"100001010",
  12742=>"111000011",
  12743=>"010100000",
  12744=>"110000000",
  12745=>"111011100",
  12746=>"001110001",
  12747=>"010101100",
  12748=>"111011010",
  12749=>"110011110",
  12750=>"011110101",
  12751=>"110111100",
  12752=>"000001101",
  12753=>"001110100",
  12754=>"100100100",
  12755=>"010110001",
  12756=>"011100111",
  12757=>"000101001",
  12758=>"111100010",
  12759=>"100001010",
  12760=>"001110010",
  12761=>"111000100",
  12762=>"100110100",
  12763=>"101101000",
  12764=>"100000101",
  12765=>"010001110",
  12766=>"011011100",
  12767=>"101010100",
  12768=>"000001000",
  12769=>"100000111",
  12770=>"110100000",
  12771=>"111011101",
  12772=>"000100111",
  12773=>"110101111",
  12774=>"110100101",
  12775=>"011000010",
  12776=>"110011111",
  12777=>"011110001",
  12778=>"110010010",
  12779=>"000110000",
  12780=>"101111110",
  12781=>"111001111",
  12782=>"110000100",
  12783=>"100101100",
  12784=>"010000111",
  12785=>"000100000",
  12786=>"001100111",
  12787=>"111010001",
  12788=>"111110110",
  12789=>"010101001",
  12790=>"000110101",
  12791=>"000001111",
  12792=>"111111010",
  12793=>"100010110",
  12794=>"101111111",
  12795=>"111100111",
  12796=>"001000100",
  12797=>"000101001",
  12798=>"001010011",
  12799=>"001110101",
  12800=>"100110101",
  12801=>"111101011",
  12802=>"011110110",
  12803=>"010101011",
  12804=>"111011101",
  12805=>"001110110",
  12806=>"001101001",
  12807=>"110110011",
  12808=>"001010110",
  12809=>"001010011",
  12810=>"000100000",
  12811=>"000111111",
  12812=>"111010000",
  12813=>"011010001",
  12814=>"111000100",
  12815=>"100011111",
  12816=>"000001110",
  12817=>"111110111",
  12818=>"011110100",
  12819=>"101101111",
  12820=>"001101110",
  12821=>"111111001",
  12822=>"101110110",
  12823=>"001111111",
  12824=>"001000110",
  12825=>"000011001",
  12826=>"010011000",
  12827=>"001111101",
  12828=>"111110001",
  12829=>"100100101",
  12830=>"010010110",
  12831=>"100111111",
  12832=>"101100111",
  12833=>"100000001",
  12834=>"110100010",
  12835=>"000110101",
  12836=>"000011000",
  12837=>"111100100",
  12838=>"001100100",
  12839=>"000000000",
  12840=>"100010100",
  12841=>"101101000",
  12842=>"000001110",
  12843=>"010111111",
  12844=>"101001110",
  12845=>"100110001",
  12846=>"000010100",
  12847=>"000101111",
  12848=>"001110010",
  12849=>"001001101",
  12850=>"011100110",
  12851=>"011010001",
  12852=>"001011000",
  12853=>"101101101",
  12854=>"111101111",
  12855=>"100101011",
  12856=>"010010001",
  12857=>"011001101",
  12858=>"101011110",
  12859=>"100010100",
  12860=>"100110011",
  12861=>"000010000",
  12862=>"011100111",
  12863=>"101111010",
  12864=>"011010100",
  12865=>"110110111",
  12866=>"100000010",
  12867=>"101011000",
  12868=>"000000110",
  12869=>"111001001",
  12870=>"001000001",
  12871=>"001111011",
  12872=>"101100111",
  12873=>"101100110",
  12874=>"100001010",
  12875=>"100111101",
  12876=>"000111101",
  12877=>"111001110",
  12878=>"000100011",
  12879=>"000100010",
  12880=>"100100001",
  12881=>"011001101",
  12882=>"100111110",
  12883=>"010010111",
  12884=>"001001110",
  12885=>"000000110",
  12886=>"101001011",
  12887=>"101011111",
  12888=>"101110100",
  12889=>"000011010",
  12890=>"001110010",
  12891=>"111101011",
  12892=>"110110000",
  12893=>"001010101",
  12894=>"010010100",
  12895=>"110001111",
  12896=>"110100110",
  12897=>"101100011",
  12898=>"001010100",
  12899=>"100010010",
  12900=>"110111011",
  12901=>"110011111",
  12902=>"001110100",
  12903=>"111001001",
  12904=>"111100001",
  12905=>"111111110",
  12906=>"010011010",
  12907=>"011111001",
  12908=>"000100111",
  12909=>"110100011",
  12910=>"001101010",
  12911=>"100101000",
  12912=>"011011011",
  12913=>"011111000",
  12914=>"111000011",
  12915=>"001001101",
  12916=>"110111001",
  12917=>"010011011",
  12918=>"001111110",
  12919=>"011100001",
  12920=>"100110111",
  12921=>"011000011",
  12922=>"010000001",
  12923=>"101000111",
  12924=>"111100000",
  12925=>"110011100",
  12926=>"010000010",
  12927=>"100001011",
  12928=>"000101011",
  12929=>"000011101",
  12930=>"100011111",
  12931=>"101110111",
  12932=>"010000010",
  12933=>"000111001",
  12934=>"111011000",
  12935=>"010111010",
  12936=>"100000000",
  12937=>"011100011",
  12938=>"110110111",
  12939=>"010001000",
  12940=>"000001101",
  12941=>"000000111",
  12942=>"101010101",
  12943=>"100011111",
  12944=>"011001111",
  12945=>"101111101",
  12946=>"111110110",
  12947=>"000011011",
  12948=>"010010100",
  12949=>"111111100",
  12950=>"111001011",
  12951=>"111110010",
  12952=>"111011100",
  12953=>"010010011",
  12954=>"000110011",
  12955=>"111101000",
  12956=>"011001000",
  12957=>"110110110",
  12958=>"011110111",
  12959=>"101101101",
  12960=>"010110101",
  12961=>"010010111",
  12962=>"001111001",
  12963=>"000111000",
  12964=>"000000100",
  12965=>"101100011",
  12966=>"000101100",
  12967=>"100010001",
  12968=>"111101100",
  12969=>"111000100",
  12970=>"101100001",
  12971=>"111000101",
  12972=>"001100100",
  12973=>"101011001",
  12974=>"110101111",
  12975=>"110000011",
  12976=>"101001101",
  12977=>"100110111",
  12978=>"100010000",
  12979=>"000001001",
  12980=>"000110000",
  12981=>"000100010",
  12982=>"110001110",
  12983=>"111001110",
  12984=>"001110110",
  12985=>"011001100",
  12986=>"001011111",
  12987=>"001111101",
  12988=>"110001100",
  12989=>"010001010",
  12990=>"110111000",
  12991=>"100010010",
  12992=>"111111100",
  12993=>"011110100",
  12994=>"011001000",
  12995=>"110011111",
  12996=>"000001010",
  12997=>"101101010",
  12998=>"001101101",
  12999=>"111001010",
  13000=>"001010001",
  13001=>"000001101",
  13002=>"011001110",
  13003=>"010110001",
  13004=>"010011010",
  13005=>"010100001",
  13006=>"010000000",
  13007=>"111100000",
  13008=>"100001111",
  13009=>"100010111",
  13010=>"101000111",
  13011=>"110110111",
  13012=>"101001100",
  13013=>"100011011",
  13014=>"011110000",
  13015=>"001111011",
  13016=>"001101101",
  13017=>"101110011",
  13018=>"000001010",
  13019=>"100001111",
  13020=>"100011000",
  13021=>"000111001",
  13022=>"001001010",
  13023=>"100101010",
  13024=>"111010110",
  13025=>"000001001",
  13026=>"000011000",
  13027=>"001100000",
  13028=>"110100001",
  13029=>"100100011",
  13030=>"000000001",
  13031=>"000001000",
  13032=>"011100011",
  13033=>"110001001",
  13034=>"101110111",
  13035=>"110101111",
  13036=>"110000100",
  13037=>"010111001",
  13038=>"100100101",
  13039=>"010111010",
  13040=>"111110000",
  13041=>"001111000",
  13042=>"100001111",
  13043=>"100110001",
  13044=>"110100000",
  13045=>"011001011",
  13046=>"001001011",
  13047=>"101011110",
  13048=>"010001110",
  13049=>"101010010",
  13050=>"000010001",
  13051=>"010010100",
  13052=>"101111110",
  13053=>"100001111",
  13054=>"101101011",
  13055=>"010000111",
  13056=>"101101011",
  13057=>"000101000",
  13058=>"000011010",
  13059=>"001000100",
  13060=>"101110001",
  13061=>"111000011",
  13062=>"010000100",
  13063=>"100001010",
  13064=>"011000111",
  13065=>"110101000",
  13066=>"001100000",
  13067=>"101000000",
  13068=>"111111011",
  13069=>"110100011",
  13070=>"011110000",
  13071=>"100010100",
  13072=>"110101100",
  13073=>"001111001",
  13074=>"111010110",
  13075=>"111100101",
  13076=>"111100111",
  13077=>"000101101",
  13078=>"100110111",
  13079=>"111001001",
  13080=>"000101001",
  13081=>"101000010",
  13082=>"011111100",
  13083=>"101001100",
  13084=>"001101101",
  13085=>"001000001",
  13086=>"101110001",
  13087=>"010001100",
  13088=>"000000011",
  13089=>"000000011",
  13090=>"101001011",
  13091=>"100010101",
  13092=>"101010101",
  13093=>"111101100",
  13094=>"101001001",
  13095=>"100000010",
  13096=>"000001001",
  13097=>"010000011",
  13098=>"000111100",
  13099=>"000011101",
  13100=>"110111000",
  13101=>"101100100",
  13102=>"110101111",
  13103=>"001000010",
  13104=>"000000011",
  13105=>"111101100",
  13106=>"001111100",
  13107=>"010100010",
  13108=>"110001010",
  13109=>"010011111",
  13110=>"001010111",
  13111=>"100000110",
  13112=>"000100110",
  13113=>"011101111",
  13114=>"000011010",
  13115=>"101010100",
  13116=>"110100111",
  13117=>"101010001",
  13118=>"001000001",
  13119=>"010110000",
  13120=>"110111101",
  13121=>"111110110",
  13122=>"101101000",
  13123=>"111011001",
  13124=>"011010110",
  13125=>"000000001",
  13126=>"110011100",
  13127=>"110010010",
  13128=>"111111110",
  13129=>"001111101",
  13130=>"011010101",
  13131=>"000010101",
  13132=>"011111001",
  13133=>"001111100",
  13134=>"010111101",
  13135=>"110000001",
  13136=>"101000001",
  13137=>"101101001",
  13138=>"000100001",
  13139=>"111000011",
  13140=>"111001101",
  13141=>"011001101",
  13142=>"000011000",
  13143=>"001001100",
  13144=>"111100100",
  13145=>"000111101",
  13146=>"110100101",
  13147=>"000010110",
  13148=>"001001011",
  13149=>"010000001",
  13150=>"111010010",
  13151=>"010001111",
  13152=>"111001100",
  13153=>"000101111",
  13154=>"111110000",
  13155=>"000110110",
  13156=>"000011001",
  13157=>"011100001",
  13158=>"111111011",
  13159=>"000001100",
  13160=>"011011110",
  13161=>"111010010",
  13162=>"011010110",
  13163=>"001011011",
  13164=>"100010101",
  13165=>"010011011",
  13166=>"001011000",
  13167=>"100001101",
  13168=>"111010100",
  13169=>"100001110",
  13170=>"100001100",
  13171=>"100011001",
  13172=>"011001111",
  13173=>"010010101",
  13174=>"100110000",
  13175=>"000010001",
  13176=>"011011010",
  13177=>"111001011",
  13178=>"000001000",
  13179=>"100100101",
  13180=>"001110011",
  13181=>"010000001",
  13182=>"011000101",
  13183=>"110110011",
  13184=>"011100100",
  13185=>"011011000",
  13186=>"100001111",
  13187=>"100110100",
  13188=>"000010000",
  13189=>"100100000",
  13190=>"010110011",
  13191=>"000001110",
  13192=>"010011101",
  13193=>"010110110",
  13194=>"011100010",
  13195=>"111011100",
  13196=>"010001111",
  13197=>"001000011",
  13198=>"111110010",
  13199=>"010000011",
  13200=>"000100011",
  13201=>"100001110",
  13202=>"111000101",
  13203=>"001101100",
  13204=>"000010001",
  13205=>"011110010",
  13206=>"110100001",
  13207=>"111101011",
  13208=>"001001101",
  13209=>"101100001",
  13210=>"011001101",
  13211=>"110010001",
  13212=>"011011111",
  13213=>"010001100",
  13214=>"101000110",
  13215=>"000000011",
  13216=>"010011000",
  13217=>"000110000",
  13218=>"100111011",
  13219=>"010000000",
  13220=>"000110000",
  13221=>"110101110",
  13222=>"100101010",
  13223=>"000111100",
  13224=>"001011100",
  13225=>"001100000",
  13226=>"000010101",
  13227=>"111111110",
  13228=>"000001000",
  13229=>"001101010",
  13230=>"010110110",
  13231=>"000111111",
  13232=>"101000101",
  13233=>"101010100",
  13234=>"010000011",
  13235=>"110101111",
  13236=>"010110111",
  13237=>"110010010",
  13238=>"000101010",
  13239=>"110111011",
  13240=>"000001101",
  13241=>"101011010",
  13242=>"011011111",
  13243=>"110000001",
  13244=>"001010111",
  13245=>"000000000",
  13246=>"010101111",
  13247=>"010100100",
  13248=>"110100010",
  13249=>"101000011",
  13250=>"110110011",
  13251=>"001101101",
  13252=>"000100101",
  13253=>"000000010",
  13254=>"111000001",
  13255=>"110100001",
  13256=>"100101001",
  13257=>"011111101",
  13258=>"111101100",
  13259=>"001101010",
  13260=>"110000110",
  13261=>"000001010",
  13262=>"100100110",
  13263=>"110000110",
  13264=>"000000000",
  13265=>"010001000",
  13266=>"100011000",
  13267=>"101100100",
  13268=>"011110101",
  13269=>"000000011",
  13270=>"100010110",
  13271=>"011110100",
  13272=>"100111111",
  13273=>"000001000",
  13274=>"000001000",
  13275=>"011000111",
  13276=>"011111011",
  13277=>"100100111",
  13278=>"011110101",
  13279=>"110100110",
  13280=>"000100111",
  13281=>"100011101",
  13282=>"100001110",
  13283=>"001110101",
  13284=>"100000000",
  13285=>"011110110",
  13286=>"111100100",
  13287=>"100001000",
  13288=>"110010011",
  13289=>"001001011",
  13290=>"111101111",
  13291=>"100001001",
  13292=>"111010010",
  13293=>"100111000",
  13294=>"101010010",
  13295=>"111110111",
  13296=>"001101101",
  13297=>"100100110",
  13298=>"110010111",
  13299=>"101111000",
  13300=>"000110111",
  13301=>"001110110",
  13302=>"111101000",
  13303=>"001100111",
  13304=>"010100110",
  13305=>"111111101",
  13306=>"001110100",
  13307=>"100000000",
  13308=>"110111100",
  13309=>"011000000",
  13310=>"111111000",
  13311=>"011110001",
  13312=>"010011010",
  13313=>"000000101",
  13314=>"101111010",
  13315=>"111010101",
  13316=>"100111010",
  13317=>"010101110",
  13318=>"000101101",
  13319=>"110000100",
  13320=>"001010100",
  13321=>"100110111",
  13322=>"100110101",
  13323=>"000011010",
  13324=>"101010111",
  13325=>"110111001",
  13326=>"001001010",
  13327=>"000010000",
  13328=>"111010111",
  13329=>"010100000",
  13330=>"010000010",
  13331=>"001110000",
  13332=>"010001110",
  13333=>"100100110",
  13334=>"000101010",
  13335=>"010100011",
  13336=>"100011100",
  13337=>"001110100",
  13338=>"000010111",
  13339=>"110010101",
  13340=>"111111101",
  13341=>"001010111",
  13342=>"111011111",
  13343=>"111001001",
  13344=>"000100110",
  13345=>"001011010",
  13346=>"001101100",
  13347=>"111010101",
  13348=>"010011101",
  13349=>"100101000",
  13350=>"001100001",
  13351=>"100001101",
  13352=>"001111000",
  13353=>"011010110",
  13354=>"011011011",
  13355=>"100010001",
  13356=>"001000010",
  13357=>"110110111",
  13358=>"110111100",
  13359=>"100001110",
  13360=>"001111110",
  13361=>"110000101",
  13362=>"010110101",
  13363=>"110111101",
  13364=>"010001000",
  13365=>"100010101",
  13366=>"110011101",
  13367=>"111001000",
  13368=>"011000111",
  13369=>"001111100",
  13370=>"100010110",
  13371=>"001111100",
  13372=>"111001011",
  13373=>"110110000",
  13374=>"111000011",
  13375=>"001011001",
  13376=>"000100100",
  13377=>"111010101",
  13378=>"000110010",
  13379=>"001100110",
  13380=>"010010001",
  13381=>"001110010",
  13382=>"011100100",
  13383=>"111111000",
  13384=>"001010011",
  13385=>"110101100",
  13386=>"110101101",
  13387=>"001011100",
  13388=>"100111110",
  13389=>"100111100",
  13390=>"100001100",
  13391=>"110001010",
  13392=>"010000001",
  13393=>"010000111",
  13394=>"010100011",
  13395=>"101100111",
  13396=>"101001000",
  13397=>"111000010",
  13398=>"100101111",
  13399=>"001111100",
  13400=>"000110100",
  13401=>"010010011",
  13402=>"100101001",
  13403=>"110000000",
  13404=>"010110100",
  13405=>"011110011",
  13406=>"111011010",
  13407=>"100111001",
  13408=>"110100101",
  13409=>"100000010",
  13410=>"100111011",
  13411=>"011111010",
  13412=>"000001010",
  13413=>"110110010",
  13414=>"010011010",
  13415=>"010000101",
  13416=>"101001000",
  13417=>"100000011",
  13418=>"001101111",
  13419=>"011010000",
  13420=>"000000111",
  13421=>"101101000",
  13422=>"100011001",
  13423=>"011011100",
  13424=>"010010101",
  13425=>"110110100",
  13426=>"111010101",
  13427=>"110100001",
  13428=>"000010011",
  13429=>"111100010",
  13430=>"001011011",
  13431=>"110000110",
  13432=>"101111010",
  13433=>"010101110",
  13434=>"000100110",
  13435=>"000000000",
  13436=>"101111010",
  13437=>"100111111",
  13438=>"101000001",
  13439=>"101001111",
  13440=>"110111000",
  13441=>"110100011",
  13442=>"101000000",
  13443=>"100000100",
  13444=>"100000111",
  13445=>"100010010",
  13446=>"101001011",
  13447=>"001111101",
  13448=>"101001110",
  13449=>"011111011",
  13450=>"011101011",
  13451=>"101100010",
  13452=>"100000000",
  13453=>"000111100",
  13454=>"111000011",
  13455=>"011000011",
  13456=>"110111100",
  13457=>"101000100",
  13458=>"110001000",
  13459=>"000010000",
  13460=>"011101101",
  13461=>"100001010",
  13462=>"110001110",
  13463=>"101100000",
  13464=>"011001011",
  13465=>"010110111",
  13466=>"001000001",
  13467=>"010100000",
  13468=>"010101011",
  13469=>"100011101",
  13470=>"011011011",
  13471=>"111001010",
  13472=>"100010100",
  13473=>"110001001",
  13474=>"110100100",
  13475=>"010000101",
  13476=>"010011111",
  13477=>"000001110",
  13478=>"101010001",
  13479=>"110111101",
  13480=>"110001111",
  13481=>"101000101",
  13482=>"010001001",
  13483=>"011101011",
  13484=>"101101100",
  13485=>"100100111",
  13486=>"110010010",
  13487=>"010001101",
  13488=>"110100011",
  13489=>"011111001",
  13490=>"011111111",
  13491=>"101100111",
  13492=>"001100000",
  13493=>"001110110",
  13494=>"001010100",
  13495=>"000000010",
  13496=>"100001110",
  13497=>"111111110",
  13498=>"111011000",
  13499=>"001111010",
  13500=>"010011110",
  13501=>"001010000",
  13502=>"001011011",
  13503=>"101000011",
  13504=>"100100110",
  13505=>"100000100",
  13506=>"110011111",
  13507=>"010110110",
  13508=>"000010110",
  13509=>"001010101",
  13510=>"011101011",
  13511=>"010111100",
  13512=>"011010000",
  13513=>"100100000",
  13514=>"000000101",
  13515=>"000101001",
  13516=>"100110010",
  13517=>"000101110",
  13518=>"110100010",
  13519=>"001101101",
  13520=>"000111001",
  13521=>"101100100",
  13522=>"001000000",
  13523=>"100101010",
  13524=>"111101000",
  13525=>"110110101",
  13526=>"001001100",
  13527=>"001101010",
  13528=>"000010110",
  13529=>"010111100",
  13530=>"110100110",
  13531=>"100101010",
  13532=>"000001101",
  13533=>"111111110",
  13534=>"101011110",
  13535=>"111110101",
  13536=>"100011010",
  13537=>"001010100",
  13538=>"101001000",
  13539=>"111011001",
  13540=>"010110010",
  13541=>"110011011",
  13542=>"111001110",
  13543=>"101000110",
  13544=>"101011101",
  13545=>"011001011",
  13546=>"000101001",
  13547=>"101101101",
  13548=>"111000100",
  13549=>"011010101",
  13550=>"110010000",
  13551=>"001101111",
  13552=>"101000000",
  13553=>"101010111",
  13554=>"101001010",
  13555=>"110011001",
  13556=>"100100011",
  13557=>"001001101",
  13558=>"111110010",
  13559=>"100111101",
  13560=>"000011111",
  13561=>"110011010",
  13562=>"100110011",
  13563=>"110110001",
  13564=>"011001011",
  13565=>"101010110",
  13566=>"011010000",
  13567=>"100100111",
  13568=>"110010110",
  13569=>"111110110",
  13570=>"000110111",
  13571=>"000111110",
  13572=>"000011011",
  13573=>"001101101",
  13574=>"110011000",
  13575=>"100000000",
  13576=>"001100110",
  13577=>"010011010",
  13578=>"001001001",
  13579=>"110101101",
  13580=>"010001001",
  13581=>"111111100",
  13582=>"100010110",
  13583=>"011110000",
  13584=>"001101010",
  13585=>"010001111",
  13586=>"000101000",
  13587=>"101001101",
  13588=>"111100110",
  13589=>"001001000",
  13590=>"000001001",
  13591=>"100111001",
  13592=>"100110111",
  13593=>"111100000",
  13594=>"011111111",
  13595=>"101010011",
  13596=>"101010010",
  13597=>"001001100",
  13598=>"101111011",
  13599=>"000000100",
  13600=>"101000010",
  13601=>"110110101",
  13602=>"101001101",
  13603=>"011011000",
  13604=>"001001100",
  13605=>"110101011",
  13606=>"010110110",
  13607=>"000101101",
  13608=>"011101100",
  13609=>"100101100",
  13610=>"010000101",
  13611=>"011001000",
  13612=>"000010001",
  13613=>"001001010",
  13614=>"100100110",
  13615=>"001001010",
  13616=>"111011000",
  13617=>"011011100",
  13618=>"101010110",
  13619=>"001011100",
  13620=>"100000111",
  13621=>"100100111",
  13622=>"100000100",
  13623=>"000100011",
  13624=>"000001010",
  13625=>"011111011",
  13626=>"110010000",
  13627=>"010110011",
  13628=>"000100000",
  13629=>"000101101",
  13630=>"000111111",
  13631=>"111111111",
  13632=>"100101101",
  13633=>"101011110",
  13634=>"010001010",
  13635=>"000011110",
  13636=>"011000101",
  13637=>"111100010",
  13638=>"111110001",
  13639=>"011100000",
  13640=>"110100101",
  13641=>"010001011",
  13642=>"001000100",
  13643=>"100000111",
  13644=>"111110110",
  13645=>"100000111",
  13646=>"001101101",
  13647=>"011110100",
  13648=>"000110111",
  13649=>"111110101",
  13650=>"001001100",
  13651=>"001001101",
  13652=>"000100110",
  13653=>"111011011",
  13654=>"011111010",
  13655=>"111011110",
  13656=>"100110000",
  13657=>"110010101",
  13658=>"010000011",
  13659=>"000001110",
  13660=>"001111100",
  13661=>"111101011",
  13662=>"100000111",
  13663=>"011101111",
  13664=>"010010110",
  13665=>"100010111",
  13666=>"111111001",
  13667=>"100000001",
  13668=>"000110010",
  13669=>"001100111",
  13670=>"111001011",
  13671=>"111001001",
  13672=>"101110010",
  13673=>"010010101",
  13674=>"011010110",
  13675=>"000010000",
  13676=>"011100101",
  13677=>"100000010",
  13678=>"010000001",
  13679=>"110111101",
  13680=>"000000001",
  13681=>"011111110",
  13682=>"101110111",
  13683=>"100000111",
  13684=>"110101111",
  13685=>"110101000",
  13686=>"100111000",
  13687=>"111010000",
  13688=>"010011010",
  13689=>"001101111",
  13690=>"101111011",
  13691=>"111001001",
  13692=>"010011101",
  13693=>"101011011",
  13694=>"000111000",
  13695=>"011110000",
  13696=>"111110101",
  13697=>"111011011",
  13698=>"001101000",
  13699=>"101001001",
  13700=>"011000101",
  13701=>"010110100",
  13702=>"010001110",
  13703=>"000011110",
  13704=>"110010010",
  13705=>"111110001",
  13706=>"000011111",
  13707=>"111100110",
  13708=>"100011110",
  13709=>"101110101",
  13710=>"001000101",
  13711=>"100000000",
  13712=>"111010001",
  13713=>"011100100",
  13714=>"101000100",
  13715=>"101001110",
  13716=>"011110011",
  13717=>"000001011",
  13718=>"000101000",
  13719=>"001100001",
  13720=>"111110110",
  13721=>"110101001",
  13722=>"110101110",
  13723=>"100111010",
  13724=>"010100110",
  13725=>"010011101",
  13726=>"101110000",
  13727=>"011110110",
  13728=>"110001111",
  13729=>"110100000",
  13730=>"101100111",
  13731=>"101111100",
  13732=>"110011000",
  13733=>"110101101",
  13734=>"001100010",
  13735=>"110100111",
  13736=>"100111010",
  13737=>"100100000",
  13738=>"110100001",
  13739=>"001001011",
  13740=>"111010001",
  13741=>"111010110",
  13742=>"010101001",
  13743=>"011101010",
  13744=>"011001010",
  13745=>"111110010",
  13746=>"101000001",
  13747=>"110000101",
  13748=>"011100100",
  13749=>"010100011",
  13750=>"100111111",
  13751=>"011100011",
  13752=>"000110101",
  13753=>"011001001",
  13754=>"101100000",
  13755=>"111101111",
  13756=>"011001100",
  13757=>"110100000",
  13758=>"111011101",
  13759=>"111010000",
  13760=>"111000001",
  13761=>"110100111",
  13762=>"011010100",
  13763=>"011110011",
  13764=>"101010011",
  13765=>"111111101",
  13766=>"111001110",
  13767=>"000100000",
  13768=>"101100110",
  13769=>"000100100",
  13770=>"001100100",
  13771=>"111111111",
  13772=>"001101001",
  13773=>"010000010",
  13774=>"000110011",
  13775=>"010010001",
  13776=>"111111001",
  13777=>"010110010",
  13778=>"011001000",
  13779=>"101101100",
  13780=>"100011101",
  13781=>"000010110",
  13782=>"001100000",
  13783=>"100011111",
  13784=>"111010110",
  13785=>"000111100",
  13786=>"010010100",
  13787=>"110111110",
  13788=>"000011111",
  13789=>"000001010",
  13790=>"101110111",
  13791=>"111010001",
  13792=>"001001000",
  13793=>"000010001",
  13794=>"001011001",
  13795=>"011011100",
  13796=>"100001000",
  13797=>"001001111",
  13798=>"111010000",
  13799=>"011011110",
  13800=>"010101010",
  13801=>"001011101",
  13802=>"001001010",
  13803=>"011111001",
  13804=>"110111111",
  13805=>"010000011",
  13806=>"100100110",
  13807=>"011000000",
  13808=>"110000000",
  13809=>"000100000",
  13810=>"110101000",
  13811=>"110011110",
  13812=>"110001010",
  13813=>"001111101",
  13814=>"110111010",
  13815=>"010010010",
  13816=>"110110010",
  13817=>"111001100",
  13818=>"000100101",
  13819=>"111111000",
  13820=>"111101110",
  13821=>"000110001",
  13822=>"001011110",
  13823=>"110001000",
  13824=>"111110110",
  13825=>"010110100",
  13826=>"101100011",
  13827=>"011010000",
  13828=>"101010111",
  13829=>"001000110",
  13830=>"101000101",
  13831=>"011000101",
  13832=>"001100000",
  13833=>"000010010",
  13834=>"111111111",
  13835=>"010100000",
  13836=>"111100111",
  13837=>"011001010",
  13838=>"000100100",
  13839=>"001110001",
  13840=>"000000110",
  13841=>"111011010",
  13842=>"101111001",
  13843=>"111010100",
  13844=>"100111110",
  13845=>"010000001",
  13846=>"010101111",
  13847=>"111001101",
  13848=>"010101110",
  13849=>"101010000",
  13850=>"110011110",
  13851=>"100110000",
  13852=>"010010001",
  13853=>"010100001",
  13854=>"010001100",
  13855=>"101000011",
  13856=>"110001100",
  13857=>"111111101",
  13858=>"111111101",
  13859=>"101110101",
  13860=>"001110000",
  13861=>"100010110",
  13862=>"110101000",
  13863=>"001110111",
  13864=>"110110001",
  13865=>"101110101",
  13866=>"001110111",
  13867=>"001000000",
  13868=>"000010001",
  13869=>"010011000",
  13870=>"010001110",
  13871=>"010001011",
  13872=>"110111111",
  13873=>"010100000",
  13874=>"100101000",
  13875=>"010100100",
  13876=>"100111101",
  13877=>"110100101",
  13878=>"000111000",
  13879=>"001101110",
  13880=>"111110100",
  13881=>"010100101",
  13882=>"100110000",
  13883=>"000111101",
  13884=>"101001100",
  13885=>"111000101",
  13886=>"101010001",
  13887=>"000110111",
  13888=>"011101010",
  13889=>"100001000",
  13890=>"011100011",
  13891=>"111010011",
  13892=>"100011111",
  13893=>"010100111",
  13894=>"100100111",
  13895=>"011011110",
  13896=>"000011111",
  13897=>"011111010",
  13898=>"010010111",
  13899=>"111100110",
  13900=>"110101101",
  13901=>"101011101",
  13902=>"100110010",
  13903=>"010000000",
  13904=>"000111001",
  13905=>"011111000",
  13906=>"101100001",
  13907=>"010100000",
  13908=>"011111010",
  13909=>"100100101",
  13910=>"011001011",
  13911=>"001100000",
  13912=>"111000011",
  13913=>"110110100",
  13914=>"010010100",
  13915=>"111010010",
  13916=>"100100101",
  13917=>"010001001",
  13918=>"010100111",
  13919=>"100010101",
  13920=>"101100110",
  13921=>"101111111",
  13922=>"101111101",
  13923=>"010101010",
  13924=>"011001000",
  13925=>"010010100",
  13926=>"100001100",
  13927=>"010011000",
  13928=>"100010100",
  13929=>"100101011",
  13930=>"100100011",
  13931=>"111011001",
  13932=>"110111001",
  13933=>"100100101",
  13934=>"100101000",
  13935=>"011100001",
  13936=>"100000010",
  13937=>"111010011",
  13938=>"101100001",
  13939=>"100110010",
  13940=>"011100010",
  13941=>"101101100",
  13942=>"110100101",
  13943=>"010110011",
  13944=>"110100101",
  13945=>"010111110",
  13946=>"111111011",
  13947=>"110100001",
  13948=>"110001011",
  13949=>"000001100",
  13950=>"111101111",
  13951=>"010101110",
  13952=>"100101010",
  13953=>"111011000",
  13954=>"101001110",
  13955=>"111100111",
  13956=>"010011100",
  13957=>"100101101",
  13958=>"111100101",
  13959=>"110110010",
  13960=>"100101010",
  13961=>"100100010",
  13962=>"001111011",
  13963=>"010101111",
  13964=>"111010000",
  13965=>"110010110",
  13966=>"011100001",
  13967=>"010000111",
  13968=>"000111110",
  13969=>"111111010",
  13970=>"000101000",
  13971=>"001000001",
  13972=>"111010110",
  13973=>"001001001",
  13974=>"010010011",
  13975=>"010010110",
  13976=>"011101000",
  13977=>"010011010",
  13978=>"101011111",
  13979=>"011000110",
  13980=>"110100000",
  13981=>"100001000",
  13982=>"100100000",
  13983=>"000111011",
  13984=>"010111011",
  13985=>"110010010",
  13986=>"111100111",
  13987=>"101101000",
  13988=>"100000010",
  13989=>"111111111",
  13990=>"111101001",
  13991=>"000111001",
  13992=>"011110001",
  13993=>"000101010",
  13994=>"000011011",
  13995=>"101101000",
  13996=>"101100000",
  13997=>"101100000",
  13998=>"111011010",
  13999=>"111010011",
  14000=>"001001001",
  14001=>"000011011",
  14002=>"010011000",
  14003=>"101100010",
  14004=>"010101110",
  14005=>"110111101",
  14006=>"111001110",
  14007=>"001101111",
  14008=>"010110100",
  14009=>"111000000",
  14010=>"100010100",
  14011=>"100010101",
  14012=>"101011101",
  14013=>"100000000",
  14014=>"110110001",
  14015=>"010110110",
  14016=>"000101001",
  14017=>"100111111",
  14018=>"101101100",
  14019=>"111100010",
  14020=>"110101001",
  14021=>"010111001",
  14022=>"000001000",
  14023=>"001001100",
  14024=>"000000101",
  14025=>"111001001",
  14026=>"011000011",
  14027=>"011100101",
  14028=>"001001111",
  14029=>"000111110",
  14030=>"001100000",
  14031=>"000001000",
  14032=>"111100111",
  14033=>"111111110",
  14034=>"111101011",
  14035=>"010011011",
  14036=>"001101001",
  14037=>"010100001",
  14038=>"111011010",
  14039=>"011000010",
  14040=>"001101000",
  14041=>"101110010",
  14042=>"100110010",
  14043=>"000100111",
  14044=>"000111011",
  14045=>"010101101",
  14046=>"010100111",
  14047=>"111011011",
  14048=>"010101000",
  14049=>"000100010",
  14050=>"100011101",
  14051=>"100000101",
  14052=>"001010101",
  14053=>"010100100",
  14054=>"101001110",
  14055=>"100011010",
  14056=>"011100011",
  14057=>"110101001",
  14058=>"000010101",
  14059=>"001111001",
  14060=>"100000110",
  14061=>"001000111",
  14062=>"000110110",
  14063=>"000010110",
  14064=>"001010000",
  14065=>"010011011",
  14066=>"101101001",
  14067=>"000001010",
  14068=>"010100001",
  14069=>"111110000",
  14070=>"010101011",
  14071=>"011101011",
  14072=>"000010010",
  14073=>"101101101",
  14074=>"100011111",
  14075=>"011001001",
  14076=>"011001110",
  14077=>"110000010",
  14078=>"111101001",
  14079=>"011011110",
  14080=>"000111011",
  14081=>"110110100",
  14082=>"100011010",
  14083=>"101110111",
  14084=>"111111101",
  14085=>"000110100",
  14086=>"101001001",
  14087=>"000010101",
  14088=>"101100001",
  14089=>"100100011",
  14090=>"011011011",
  14091=>"000110111",
  14092=>"000010000",
  14093=>"111001100",
  14094=>"011110110",
  14095=>"010010001",
  14096=>"101011011",
  14097=>"001010010",
  14098=>"100111011",
  14099=>"010010111",
  14100=>"011100111",
  14101=>"100111111",
  14102=>"110100101",
  14103=>"011000110",
  14104=>"100010110",
  14105=>"101001001",
  14106=>"001001111",
  14107=>"101101110",
  14108=>"010011010",
  14109=>"101110111",
  14110=>"001010010",
  14111=>"111010000",
  14112=>"001001010",
  14113=>"000110100",
  14114=>"101001001",
  14115=>"111101111",
  14116=>"111100110",
  14117=>"000000000",
  14118=>"001111001",
  14119=>"001011111",
  14120=>"111110001",
  14121=>"111110000",
  14122=>"111111011",
  14123=>"111010010",
  14124=>"111110011",
  14125=>"010011000",
  14126=>"010101011",
  14127=>"010100111",
  14128=>"111000110",
  14129=>"101100000",
  14130=>"011101110",
  14131=>"111111001",
  14132=>"101110010",
  14133=>"111111101",
  14134=>"001000110",
  14135=>"101111111",
  14136=>"101111100",
  14137=>"000011101",
  14138=>"001001000",
  14139=>"111000011",
  14140=>"111111011",
  14141=>"110101011",
  14142=>"111110110",
  14143=>"010101001",
  14144=>"111000110",
  14145=>"000111011",
  14146=>"010110101",
  14147=>"110011111",
  14148=>"101110001",
  14149=>"101000100",
  14150=>"011001010",
  14151=>"111111110",
  14152=>"010011000",
  14153=>"101100000",
  14154=>"101100111",
  14155=>"110000110",
  14156=>"010101110",
  14157=>"101010010",
  14158=>"100001101",
  14159=>"011000110",
  14160=>"010010100",
  14161=>"101000010",
  14162=>"000000100",
  14163=>"000000111",
  14164=>"111100110",
  14165=>"101000001",
  14166=>"101000011",
  14167=>"101000001",
  14168=>"011110111",
  14169=>"101011000",
  14170=>"011100100",
  14171=>"100010101",
  14172=>"001001011",
  14173=>"010001101",
  14174=>"110000110",
  14175=>"111100110",
  14176=>"111111111",
  14177=>"010111000",
  14178=>"110110011",
  14179=>"000101011",
  14180=>"001001100",
  14181=>"011110010",
  14182=>"011100000",
  14183=>"111110001",
  14184=>"101110110",
  14185=>"111101101",
  14186=>"101001110",
  14187=>"110011001",
  14188=>"011110000",
  14189=>"010110111",
  14190=>"010111010",
  14191=>"101111000",
  14192=>"011111010",
  14193=>"110001100",
  14194=>"100101110",
  14195=>"101110110",
  14196=>"001111101",
  14197=>"001101100",
  14198=>"011000101",
  14199=>"011011111",
  14200=>"111000000",
  14201=>"110000000",
  14202=>"000001101",
  14203=>"001110010",
  14204=>"010111010",
  14205=>"011011100",
  14206=>"010101110",
  14207=>"001111110",
  14208=>"110111001",
  14209=>"011001101",
  14210=>"011000010",
  14211=>"001101110",
  14212=>"101101111",
  14213=>"000011000",
  14214=>"010111111",
  14215=>"001100101",
  14216=>"110111111",
  14217=>"001100111",
  14218=>"000011111",
  14219=>"110000111",
  14220=>"100011001",
  14221=>"111100100",
  14222=>"010011000",
  14223=>"000111000",
  14224=>"010100000",
  14225=>"110010101",
  14226=>"000100100",
  14227=>"001000101",
  14228=>"110010010",
  14229=>"101011001",
  14230=>"110100011",
  14231=>"001111111",
  14232=>"000000111",
  14233=>"011001000",
  14234=>"101000101",
  14235=>"000000111",
  14236=>"111111001",
  14237=>"011000101",
  14238=>"000110011",
  14239=>"000001011",
  14240=>"101100111",
  14241=>"011010111",
  14242=>"101010100",
  14243=>"100111000",
  14244=>"111011010",
  14245=>"100000011",
  14246=>"010101010",
  14247=>"111011100",
  14248=>"010011000",
  14249=>"101110110",
  14250=>"101101101",
  14251=>"000111011",
  14252=>"100111111",
  14253=>"100011011",
  14254=>"101011011",
  14255=>"110110110",
  14256=>"001010110",
  14257=>"010011010",
  14258=>"011101000",
  14259=>"010000000",
  14260=>"100010001",
  14261=>"100000101",
  14262=>"001011000",
  14263=>"111011111",
  14264=>"101001100",
  14265=>"100011000",
  14266=>"101101100",
  14267=>"010100010",
  14268=>"011001100",
  14269=>"111111110",
  14270=>"010000010",
  14271=>"100000111",
  14272=>"001111111",
  14273=>"100100010",
  14274=>"100001101",
  14275=>"110001000",
  14276=>"011100000",
  14277=>"000100100",
  14278=>"011111001",
  14279=>"110011111",
  14280=>"111000000",
  14281=>"111000101",
  14282=>"100001000",
  14283=>"101001000",
  14284=>"100000000",
  14285=>"100011010",
  14286=>"011001011",
  14287=>"100111101",
  14288=>"000111110",
  14289=>"101001010",
  14290=>"110110000",
  14291=>"100000111",
  14292=>"011010000",
  14293=>"100001000",
  14294=>"001010001",
  14295=>"101100110",
  14296=>"110000001",
  14297=>"001011001",
  14298=>"011100010",
  14299=>"001010101",
  14300=>"010111010",
  14301=>"010101000",
  14302=>"001110000",
  14303=>"110101110",
  14304=>"000000110",
  14305=>"100111000",
  14306=>"111011111",
  14307=>"000100110",
  14308=>"100000111",
  14309=>"000000001",
  14310=>"010100101",
  14311=>"011010000",
  14312=>"111000111",
  14313=>"111101000",
  14314=>"110100010",
  14315=>"001010001",
  14316=>"001100111",
  14317=>"101111011",
  14318=>"111101101",
  14319=>"100100010",
  14320=>"110000000",
  14321=>"111101001",
  14322=>"110001101",
  14323=>"001111100",
  14324=>"011110101",
  14325=>"000001110",
  14326=>"011110110",
  14327=>"111011010",
  14328=>"110011111",
  14329=>"011010110",
  14330=>"111100001",
  14331=>"011110100",
  14332=>"000100001",
  14333=>"111111001",
  14334=>"010011100",
  14335=>"101100000",
  14336=>"010000001",
  14337=>"100010010",
  14338=>"110011110",
  14339=>"110000001",
  14340=>"111000101",
  14341=>"110100001",
  14342=>"110110010",
  14343=>"000111101",
  14344=>"101000111",
  14345=>"101011100",
  14346=>"010001001",
  14347=>"011110111",
  14348=>"011101011",
  14349=>"010111000",
  14350=>"010100111",
  14351=>"011100011",
  14352=>"100010111",
  14353=>"010000100",
  14354=>"110011011",
  14355=>"011110001",
  14356=>"011000011",
  14357=>"001000110",
  14358=>"011010110",
  14359=>"010000001",
  14360=>"110111000",
  14361=>"111110000",
  14362=>"000000100",
  14363=>"111011100",
  14364=>"010100001",
  14365=>"110000110",
  14366=>"101001010",
  14367=>"101110000",
  14368=>"011000010",
  14369=>"100000101",
  14370=>"000110100",
  14371=>"010011001",
  14372=>"110000000",
  14373=>"001010011",
  14374=>"000100010",
  14375=>"010001010",
  14376=>"110000010",
  14377=>"011001000",
  14378=>"101101100",
  14379=>"101111000",
  14380=>"101110111",
  14381=>"101111100",
  14382=>"001001001",
  14383=>"100001110",
  14384=>"011101101",
  14385=>"111100000",
  14386=>"010101101",
  14387=>"001100111",
  14388=>"101010010",
  14389=>"011000111",
  14390=>"110010000",
  14391=>"110101101",
  14392=>"100000000",
  14393=>"000000011",
  14394=>"010001000",
  14395=>"111011111",
  14396=>"111001110",
  14397=>"110100100",
  14398=>"010110001",
  14399=>"011111100",
  14400=>"011110111",
  14401=>"100010101",
  14402=>"110010011",
  14403=>"100110011",
  14404=>"100001010",
  14405=>"001011001",
  14406=>"000111011",
  14407=>"010111001",
  14408=>"101001001",
  14409=>"011110010",
  14410=>"111011010",
  14411=>"001011110",
  14412=>"011010100",
  14413=>"010001011",
  14414=>"100000100",
  14415=>"101111000",
  14416=>"111010011",
  14417=>"110011101",
  14418=>"010111001",
  14419=>"111010111",
  14420=>"001001011",
  14421=>"000110001",
  14422=>"101100000",
  14423=>"000000100",
  14424=>"110010110",
  14425=>"100011011",
  14426=>"101110110",
  14427=>"011101101",
  14428=>"011011101",
  14429=>"000000011",
  14430=>"011100011",
  14431=>"110001111",
  14432=>"011000100",
  14433=>"000010100",
  14434=>"011100100",
  14435=>"100011011",
  14436=>"110110010",
  14437=>"010000000",
  14438=>"111111100",
  14439=>"010000001",
  14440=>"101111001",
  14441=>"011101011",
  14442=>"111000101",
  14443=>"111110101",
  14444=>"110011001",
  14445=>"001000011",
  14446=>"110110101",
  14447=>"100111111",
  14448=>"000001110",
  14449=>"101001010",
  14450=>"011001110",
  14451=>"010000001",
  14452=>"100111110",
  14453=>"010001111",
  14454=>"011001011",
  14455=>"011110000",
  14456=>"100010011",
  14457=>"110110111",
  14458=>"011101100",
  14459=>"111110111",
  14460=>"111000101",
  14461=>"111111111",
  14462=>"110111101",
  14463=>"110110111",
  14464=>"101110010",
  14465=>"110111100",
  14466=>"000010101",
  14467=>"101110011",
  14468=>"101011010",
  14469=>"001100000",
  14470=>"000010100",
  14471=>"110110110",
  14472=>"011000110",
  14473=>"111101001",
  14474=>"100011000",
  14475=>"101111111",
  14476=>"010010010",
  14477=>"011011011",
  14478=>"100010111",
  14479=>"001000100",
  14480=>"011011010",
  14481=>"010111110",
  14482=>"111000101",
  14483=>"100101111",
  14484=>"111001010",
  14485=>"110101100",
  14486=>"110010111",
  14487=>"110100000",
  14488=>"110001101",
  14489=>"010011101",
  14490=>"000111010",
  14491=>"010111110",
  14492=>"000010000",
  14493=>"000100100",
  14494=>"101111000",
  14495=>"011000100",
  14496=>"110111010",
  14497=>"100001100",
  14498=>"111100111",
  14499=>"000001100",
  14500=>"111100000",
  14501=>"001111111",
  14502=>"000101110",
  14503=>"100100100",
  14504=>"111000001",
  14505=>"011100111",
  14506=>"110101100",
  14507=>"101001111",
  14508=>"011011101",
  14509=>"101111110",
  14510=>"000111001",
  14511=>"100101001",
  14512=>"011111001",
  14513=>"000011110",
  14514=>"000000011",
  14515=>"001001100",
  14516=>"111000001",
  14517=>"000000101",
  14518=>"110000101",
  14519=>"101001101",
  14520=>"000100110",
  14521=>"011101000",
  14522=>"101010010",
  14523=>"011111111",
  14524=>"101000001",
  14525=>"101110111",
  14526=>"101100001",
  14527=>"010010111",
  14528=>"101111111",
  14529=>"100101110",
  14530=>"000100001",
  14531=>"101100111",
  14532=>"001010101",
  14533=>"101101000",
  14534=>"001100010",
  14535=>"000010110",
  14536=>"000110010",
  14537=>"100011001",
  14538=>"000110111",
  14539=>"110100010",
  14540=>"011111011",
  14541=>"011100010",
  14542=>"001011111",
  14543=>"000110101",
  14544=>"010110010",
  14545=>"111101111",
  14546=>"111001010",
  14547=>"011011000",
  14548=>"100010111",
  14549=>"111100010",
  14550=>"011110010",
  14551=>"111101101",
  14552=>"100111111",
  14553=>"011000010",
  14554=>"110110001",
  14555=>"011111101",
  14556=>"100110010",
  14557=>"010101101",
  14558=>"110111001",
  14559=>"000000011",
  14560=>"010110011",
  14561=>"000101111",
  14562=>"101000000",
  14563=>"111101000",
  14564=>"000000001",
  14565=>"110011101",
  14566=>"011010000",
  14567=>"001011010",
  14568=>"100000101",
  14569=>"100001100",
  14570=>"110010110",
  14571=>"100000010",
  14572=>"100111100",
  14573=>"001010101",
  14574=>"101010010",
  14575=>"001110110",
  14576=>"000010111",
  14577=>"101101000",
  14578=>"010111011",
  14579=>"110111110",
  14580=>"110111100",
  14581=>"011100011",
  14582=>"100011100",
  14583=>"000110100",
  14584=>"111100110",
  14585=>"111101010",
  14586=>"111100011",
  14587=>"000110000",
  14588=>"001110111",
  14589=>"111010001",
  14590=>"011111101",
  14591=>"010000100",
  14592=>"011111101",
  14593=>"001100001",
  14594=>"001001011",
  14595=>"101101101",
  14596=>"111111110",
  14597=>"000110111",
  14598=>"011000010",
  14599=>"010000011",
  14600=>"110010011",
  14601=>"111000001",
  14602=>"001100001",
  14603=>"001000000",
  14604=>"100001011",
  14605=>"101110001",
  14606=>"001010110",
  14607=>"010000011",
  14608=>"001111110",
  14609=>"000001010",
  14610=>"010011100",
  14611=>"000000010",
  14612=>"011111100",
  14613=>"001100010",
  14614=>"001011000",
  14615=>"110101001",
  14616=>"111011000",
  14617=>"101100110",
  14618=>"101110010",
  14619=>"100110110",
  14620=>"011101101",
  14621=>"001101111",
  14622=>"100100111",
  14623=>"000110010",
  14624=>"100101111",
  14625=>"000110010",
  14626=>"010010100",
  14627=>"111010111",
  14628=>"101101101",
  14629=>"100010010",
  14630=>"010100111",
  14631=>"110001111",
  14632=>"100000000",
  14633=>"110100001",
  14634=>"010010110",
  14635=>"110011100",
  14636=>"011101110",
  14637=>"110000000",
  14638=>"101111010",
  14639=>"001111101",
  14640=>"011010110",
  14641=>"101110110",
  14642=>"001000111",
  14643=>"011011100",
  14644=>"100100110",
  14645=>"100100000",
  14646=>"100000001",
  14647=>"100010111",
  14648=>"100001000",
  14649=>"001101010",
  14650=>"011001010",
  14651=>"011110100",
  14652=>"011010010",
  14653=>"101000111",
  14654=>"010000011",
  14655=>"110111111",
  14656=>"011011010",
  14657=>"001001011",
  14658=>"011000000",
  14659=>"011011001",
  14660=>"010000001",
  14661=>"110100000",
  14662=>"110001011",
  14663=>"011110100",
  14664=>"001000010",
  14665=>"101101001",
  14666=>"011110000",
  14667=>"100000111",
  14668=>"000111101",
  14669=>"100000101",
  14670=>"010110111",
  14671=>"011111010",
  14672=>"101110001",
  14673=>"000011011",
  14674=>"110111010",
  14675=>"111010010",
  14676=>"010101010",
  14677=>"110011000",
  14678=>"100001011",
  14679=>"110010111",
  14680=>"010010001",
  14681=>"101011010",
  14682=>"011100010",
  14683=>"100000000",
  14684=>"010101110",
  14685=>"010000011",
  14686=>"110000010",
  14687=>"101100001",
  14688=>"001111101",
  14689=>"110010111",
  14690=>"000000111",
  14691=>"000000111",
  14692=>"010111010",
  14693=>"100010110",
  14694=>"000111001",
  14695=>"111101110",
  14696=>"000110100",
  14697=>"010011111",
  14698=>"011011011",
  14699=>"101111101",
  14700=>"001000010",
  14701=>"010101110",
  14702=>"010100000",
  14703=>"110001000",
  14704=>"111101111",
  14705=>"110001000",
  14706=>"100101011",
  14707=>"111110101",
  14708=>"001001000",
  14709=>"000011010",
  14710=>"001001100",
  14711=>"001100010",
  14712=>"011100000",
  14713=>"011000101",
  14714=>"101101000",
  14715=>"101111111",
  14716=>"000001011",
  14717=>"110000001",
  14718=>"011100101",
  14719=>"000010001",
  14720=>"011000000",
  14721=>"010000000",
  14722=>"000011111",
  14723=>"100111010",
  14724=>"001001101",
  14725=>"010111000",
  14726=>"101010011",
  14727=>"001000000",
  14728=>"010011001",
  14729=>"000000100",
  14730=>"010001111",
  14731=>"100110011",
  14732=>"000001001",
  14733=>"000001011",
  14734=>"101101010",
  14735=>"001001000",
  14736=>"111101110",
  14737=>"111010110",
  14738=>"001011010",
  14739=>"001000010",
  14740=>"101001110",
  14741=>"101010101",
  14742=>"111011000",
  14743=>"101001001",
  14744=>"101001001",
  14745=>"001010000",
  14746=>"010011010",
  14747=>"110001010",
  14748=>"011111001",
  14749=>"100000101",
  14750=>"111100001",
  14751=>"110111001",
  14752=>"110001010",
  14753=>"000010111",
  14754=>"101110100",
  14755=>"101110000",
  14756=>"100110010",
  14757=>"000000101",
  14758=>"110010110",
  14759=>"110001100",
  14760=>"000101100",
  14761=>"000011001",
  14762=>"000001100",
  14763=>"011000000",
  14764=>"000000010",
  14765=>"010101011",
  14766=>"000001010",
  14767=>"000001000",
  14768=>"111111111",
  14769=>"010110000",
  14770=>"100000111",
  14771=>"000100010",
  14772=>"000011111",
  14773=>"110111110",
  14774=>"001110000",
  14775=>"110110110",
  14776=>"101001110",
  14777=>"111110111",
  14778=>"101010010",
  14779=>"100001111",
  14780=>"111110100",
  14781=>"100010000",
  14782=>"101100000",
  14783=>"100010001",
  14784=>"110110000",
  14785=>"000001001",
  14786=>"101001111",
  14787=>"111111010",
  14788=>"010001010",
  14789=>"110011010",
  14790=>"000010111",
  14791=>"010001101",
  14792=>"001001110",
  14793=>"011111101",
  14794=>"011111001",
  14795=>"011000110",
  14796=>"001000001",
  14797=>"000001101",
  14798=>"001001001",
  14799=>"000101011",
  14800=>"000000000",
  14801=>"000111111",
  14802=>"110110101",
  14803=>"111011101",
  14804=>"000100001",
  14805=>"110110000",
  14806=>"001010100",
  14807=>"010100001",
  14808=>"111000001",
  14809=>"000000100",
  14810=>"100101001",
  14811=>"001000001",
  14812=>"011001010",
  14813=>"101101100",
  14814=>"000010111",
  14815=>"110000010",
  14816=>"101000011",
  14817=>"010001000",
  14818=>"110110001",
  14819=>"000110000",
  14820=>"100100110",
  14821=>"010010100",
  14822=>"010110100",
  14823=>"010110001",
  14824=>"010000011",
  14825=>"010111100",
  14826=>"011001011",
  14827=>"101101111",
  14828=>"111000110",
  14829=>"111111101",
  14830=>"111001100",
  14831=>"111111001",
  14832=>"011101001",
  14833=>"101111010",
  14834=>"110010101",
  14835=>"111010011",
  14836=>"000100111",
  14837=>"011010011",
  14838=>"010001001",
  14839=>"110111011",
  14840=>"000100000",
  14841=>"111101101",
  14842=>"010000101",
  14843=>"011011110",
  14844=>"100100111",
  14845=>"110001100",
  14846=>"111000100",
  14847=>"011001001",
  14848=>"001110110",
  14849=>"100000000",
  14850=>"111111000",
  14851=>"010010111",
  14852=>"111000010",
  14853=>"111100010",
  14854=>"100001001",
  14855=>"100111110",
  14856=>"100011110",
  14857=>"110110001",
  14858=>"010000010",
  14859=>"000110110",
  14860=>"110110010",
  14861=>"000011001",
  14862=>"010100110",
  14863=>"011010110",
  14864=>"110100001",
  14865=>"110100000",
  14866=>"110000001",
  14867=>"000111111",
  14868=>"110101010",
  14869=>"010111100",
  14870=>"001111000",
  14871=>"110111010",
  14872=>"111111000",
  14873=>"000000011",
  14874=>"000110111",
  14875=>"111110010",
  14876=>"011011110",
  14877=>"110110100",
  14878=>"101111001",
  14879=>"110010101",
  14880=>"011010001",
  14881=>"110110101",
  14882=>"000100011",
  14883=>"100110011",
  14884=>"001110001",
  14885=>"011001100",
  14886=>"101010101",
  14887=>"001100000",
  14888=>"100010010",
  14889=>"011001011",
  14890=>"101011101",
  14891=>"110100111",
  14892=>"111010100",
  14893=>"110000101",
  14894=>"010011110",
  14895=>"101100101",
  14896=>"001110111",
  14897=>"101111000",
  14898=>"110001111",
  14899=>"000110101",
  14900=>"010101101",
  14901=>"001101000",
  14902=>"010100101",
  14903=>"011101101",
  14904=>"010111111",
  14905=>"101101110",
  14906=>"010000100",
  14907=>"010010111",
  14908=>"000101100",
  14909=>"110100000",
  14910=>"000101011",
  14911=>"000010100",
  14912=>"111110000",
  14913=>"011011010",
  14914=>"011110010",
  14915=>"001100111",
  14916=>"000000010",
  14917=>"100101100",
  14918=>"111010101",
  14919=>"100101110",
  14920=>"011101100",
  14921=>"010011011",
  14922=>"101100100",
  14923=>"010100010",
  14924=>"010100110",
  14925=>"101000111",
  14926=>"011000010",
  14927=>"100110001",
  14928=>"101111011",
  14929=>"111111111",
  14930=>"001100111",
  14931=>"011100011",
  14932=>"000100110",
  14933=>"000011110",
  14934=>"001100101",
  14935=>"100101001",
  14936=>"101111110",
  14937=>"110011111",
  14938=>"011000101",
  14939=>"001110001",
  14940=>"000100101",
  14941=>"100001000",
  14942=>"000001011",
  14943=>"001100110",
  14944=>"001101100",
  14945=>"000100100",
  14946=>"001101101",
  14947=>"111011100",
  14948=>"000111001",
  14949=>"001110001",
  14950=>"011011111",
  14951=>"101010011",
  14952=>"010100101",
  14953=>"110010001",
  14954=>"110000110",
  14955=>"111111110",
  14956=>"001000110",
  14957=>"110011110",
  14958=>"011011001",
  14959=>"100011100",
  14960=>"110110101",
  14961=>"110010001",
  14962=>"100011111",
  14963=>"111100000",
  14964=>"010111011",
  14965=>"011011101",
  14966=>"001111110",
  14967=>"010110111",
  14968=>"101011001",
  14969=>"011101001",
  14970=>"010000110",
  14971=>"011000111",
  14972=>"100011000",
  14973=>"110000111",
  14974=>"100101100",
  14975=>"101110100",
  14976=>"101101001",
  14977=>"100101011",
  14978=>"010001000",
  14979=>"011111110",
  14980=>"011101001",
  14981=>"101110110",
  14982=>"010100100",
  14983=>"111100011",
  14984=>"101111000",
  14985=>"000110000",
  14986=>"011100010",
  14987=>"101001111",
  14988=>"101011010",
  14989=>"010100001",
  14990=>"101011101",
  14991=>"111110110",
  14992=>"001111100",
  14993=>"010111100",
  14994=>"000010001",
  14995=>"011101110",
  14996=>"000110110",
  14997=>"000110001",
  14998=>"110011110",
  14999=>"001010100",
  15000=>"111100011",
  15001=>"010001000",
  15002=>"001000011",
  15003=>"001001001",
  15004=>"001011010",
  15005=>"101101110",
  15006=>"111010001",
  15007=>"101111011",
  15008=>"111110001",
  15009=>"000001011",
  15010=>"010111000",
  15011=>"101011101",
  15012=>"010100100",
  15013=>"110111111",
  15014=>"001010011",
  15015=>"000101100",
  15016=>"000111101",
  15017=>"101001011",
  15018=>"000101100",
  15019=>"100110000",
  15020=>"001011100",
  15021=>"101000100",
  15022=>"101110011",
  15023=>"100110110",
  15024=>"011001011",
  15025=>"101001111",
  15026=>"001110011",
  15027=>"001110101",
  15028=>"110001001",
  15029=>"001001101",
  15030=>"000001100",
  15031=>"001111010",
  15032=>"001001110",
  15033=>"100110011",
  15034=>"000110111",
  15035=>"001001000",
  15036=>"101000011",
  15037=>"101110111",
  15038=>"110110000",
  15039=>"001100100",
  15040=>"111111000",
  15041=>"011110010",
  15042=>"101110101",
  15043=>"001110000",
  15044=>"110110100",
  15045=>"001111110",
  15046=>"000000101",
  15047=>"100001000",
  15048=>"101101001",
  15049=>"010100001",
  15050=>"011100111",
  15051=>"111111000",
  15052=>"111101101",
  15053=>"101100101",
  15054=>"101001100",
  15055=>"101001001",
  15056=>"110000001",
  15057=>"110100101",
  15058=>"001011111",
  15059=>"000010011",
  15060=>"101101101",
  15061=>"101101011",
  15062=>"011011000",
  15063=>"000000010",
  15064=>"000001100",
  15065=>"000001111",
  15066=>"011000010",
  15067=>"110011100",
  15068=>"111001101",
  15069=>"010100100",
  15070=>"110000001",
  15071=>"000111001",
  15072=>"001111110",
  15073=>"100000000",
  15074=>"101110100",
  15075=>"110101010",
  15076=>"011010110",
  15077=>"101011011",
  15078=>"000001000",
  15079=>"111010000",
  15080=>"011110010",
  15081=>"001100110",
  15082=>"101111100",
  15083=>"001000000",
  15084=>"000000111",
  15085=>"100000100",
  15086=>"000110011",
  15087=>"010100110",
  15088=>"100000011",
  15089=>"001101110",
  15090=>"010000000",
  15091=>"011100011",
  15092=>"000010001",
  15093=>"010100101",
  15094=>"100011001",
  15095=>"000011000",
  15096=>"110000110",
  15097=>"011111110",
  15098=>"101010111",
  15099=>"010101101",
  15100=>"001000101",
  15101=>"101111000",
  15102=>"100111100",
  15103=>"101100010",
  15104=>"101111111",
  15105=>"001110111",
  15106=>"101000110",
  15107=>"000011111",
  15108=>"000101011",
  15109=>"110001001",
  15110=>"000100110",
  15111=>"111010111",
  15112=>"000111000",
  15113=>"101010110",
  15114=>"010101100",
  15115=>"111100111",
  15116=>"111010101",
  15117=>"111000010",
  15118=>"111010000",
  15119=>"110010001",
  15120=>"111011001",
  15121=>"011000111",
  15122=>"001111111",
  15123=>"101011001",
  15124=>"101000011",
  15125=>"111011000",
  15126=>"010010001",
  15127=>"000110101",
  15128=>"111010101",
  15129=>"010000111",
  15130=>"111111111",
  15131=>"001000111",
  15132=>"000010000",
  15133=>"010110110",
  15134=>"111000001",
  15135=>"000101010",
  15136=>"010110010",
  15137=>"111110110",
  15138=>"111011110",
  15139=>"001111110",
  15140=>"010001010",
  15141=>"000000011",
  15142=>"011110011",
  15143=>"000010000",
  15144=>"000101110",
  15145=>"101101101",
  15146=>"111100101",
  15147=>"111010011",
  15148=>"111101001",
  15149=>"111010101",
  15150=>"011111110",
  15151=>"101000101",
  15152=>"001101100",
  15153=>"000100111",
  15154=>"000001100",
  15155=>"101000000",
  15156=>"011110010",
  15157=>"111110000",
  15158=>"011101010",
  15159=>"000010010",
  15160=>"100011010",
  15161=>"010001110",
  15162=>"000100000",
  15163=>"001110110",
  15164=>"001001001",
  15165=>"001110011",
  15166=>"011101111",
  15167=>"101111110",
  15168=>"101111101",
  15169=>"000011111",
  15170=>"101010111",
  15171=>"010001011",
  15172=>"001110010",
  15173=>"101100011",
  15174=>"001000001",
  15175=>"000101100",
  15176=>"000111111",
  15177=>"111101001",
  15178=>"111100101",
  15179=>"101101001",
  15180=>"110000111",
  15181=>"001001111",
  15182=>"010000101",
  15183=>"101011101",
  15184=>"111010010",
  15185=>"110111100",
  15186=>"000101101",
  15187=>"011111101",
  15188=>"101000010",
  15189=>"011000100",
  15190=>"111011010",
  15191=>"100000000",
  15192=>"000100111",
  15193=>"111011010",
  15194=>"100100011",
  15195=>"111000001",
  15196=>"110010011",
  15197=>"111001000",
  15198=>"000001110",
  15199=>"100011100",
  15200=>"100100011",
  15201=>"001001000",
  15202=>"000110101",
  15203=>"110011001",
  15204=>"000111111",
  15205=>"000010000",
  15206=>"000000101",
  15207=>"000110001",
  15208=>"101100010",
  15209=>"001110000",
  15210=>"000000010",
  15211=>"101111010",
  15212=>"111100100",
  15213=>"101111011",
  15214=>"001111011",
  15215=>"110010111",
  15216=>"001000101",
  15217=>"001110100",
  15218=>"011111010",
  15219=>"110011001",
  15220=>"111000001",
  15221=>"010001010",
  15222=>"101111000",
  15223=>"111100010",
  15224=>"011000010",
  15225=>"110010010",
  15226=>"111000010",
  15227=>"111000101",
  15228=>"011101100",
  15229=>"001010001",
  15230=>"010001100",
  15231=>"001001110",
  15232=>"010111101",
  15233=>"101000000",
  15234=>"001100011",
  15235=>"001010110",
  15236=>"000001110",
  15237=>"100011010",
  15238=>"000011111",
  15239=>"010001101",
  15240=>"000011101",
  15241=>"100010111",
  15242=>"110010100",
  15243=>"011000110",
  15244=>"101010101",
  15245=>"001001111",
  15246=>"101001111",
  15247=>"100011101",
  15248=>"011100100",
  15249=>"011011010",
  15250=>"010000010",
  15251=>"010110010",
  15252=>"000100001",
  15253=>"011001100",
  15254=>"001111100",
  15255=>"001010100",
  15256=>"111110010",
  15257=>"000111000",
  15258=>"000001001",
  15259=>"000101011",
  15260=>"111100000",
  15261=>"010110101",
  15262=>"100010000",
  15263=>"000101010",
  15264=>"101100011",
  15265=>"101000000",
  15266=>"100011011",
  15267=>"101101001",
  15268=>"100001000",
  15269=>"000110101",
  15270=>"000011000",
  15271=>"110100011",
  15272=>"010000001",
  15273=>"010111000",
  15274=>"001011110",
  15275=>"111011110",
  15276=>"100110101",
  15277=>"001100110",
  15278=>"111110101",
  15279=>"000011100",
  15280=>"001110110",
  15281=>"110110110",
  15282=>"100100010",
  15283=>"011110111",
  15284=>"101000000",
  15285=>"011011100",
  15286=>"010110001",
  15287=>"010011010",
  15288=>"110000111",
  15289=>"110011101",
  15290=>"111111000",
  15291=>"001010111",
  15292=>"010001010",
  15293=>"011011000",
  15294=>"011111011",
  15295=>"111001110",
  15296=>"010111111",
  15297=>"011100010",
  15298=>"010101111",
  15299=>"000000110",
  15300=>"001111111",
  15301=>"001000101",
  15302=>"010010100",
  15303=>"100111000",
  15304=>"000000010",
  15305=>"000010000",
  15306=>"111011010",
  15307=>"101101000",
  15308=>"010101011",
  15309=>"100100110",
  15310=>"001111010",
  15311=>"000101000",
  15312=>"000100001",
  15313=>"101011111",
  15314=>"101101000",
  15315=>"010011011",
  15316=>"111100000",
  15317=>"000000101",
  15318=>"101100001",
  15319=>"001000011",
  15320=>"100011011",
  15321=>"010101101",
  15322=>"001010101",
  15323=>"101000111",
  15324=>"000001000",
  15325=>"100100101",
  15326=>"000001111",
  15327=>"100000111",
  15328=>"111011110",
  15329=>"100110011",
  15330=>"000000111",
  15331=>"110100010",
  15332=>"001100111",
  15333=>"001001011",
  15334=>"000000110",
  15335=>"111000100",
  15336=>"000100100",
  15337=>"101110000",
  15338=>"010100010",
  15339=>"111110110",
  15340=>"100001011",
  15341=>"001111100",
  15342=>"111100101",
  15343=>"010110100",
  15344=>"100100011",
  15345=>"110001100",
  15346=>"000100010",
  15347=>"110110001",
  15348=>"011011011",
  15349=>"000001100",
  15350=>"011101100",
  15351=>"011010011",
  15352=>"101101111",
  15353=>"101111011",
  15354=>"011001101",
  15355=>"000110110",
  15356=>"001110101",
  15357=>"011111001",
  15358=>"000101001",
  15359=>"010100110",
  15360=>"000000100",
  15361=>"100110111",
  15362=>"111011011",
  15363=>"010111010",
  15364=>"010011100",
  15365=>"001111110",
  15366=>"000011101",
  15367=>"101111000",
  15368=>"001111101",
  15369=>"000011100",
  15370=>"100001000",
  15371=>"011111000",
  15372=>"011111111",
  15373=>"000100111",
  15374=>"110010000",
  15375=>"111111111",
  15376=>"111110101",
  15377=>"100011100",
  15378=>"111100010",
  15379=>"100101110",
  15380=>"000001111",
  15381=>"100000111",
  15382=>"010001101",
  15383=>"001111000",
  15384=>"001010010",
  15385=>"100111110",
  15386=>"110010110",
  15387=>"001000011",
  15388=>"011110001",
  15389=>"101010001",
  15390=>"111011000",
  15391=>"001011110",
  15392=>"110110111",
  15393=>"101101011",
  15394=>"011001001",
  15395=>"010110111",
  15396=>"000111101",
  15397=>"110000000",
  15398=>"000110100",
  15399=>"110111111",
  15400=>"110111101",
  15401=>"100101010",
  15402=>"010010000",
  15403=>"100111101",
  15404=>"110011111",
  15405=>"011100101",
  15406=>"100001011",
  15407=>"011101010",
  15408=>"101111001",
  15409=>"000000101",
  15410=>"000000111",
  15411=>"110010100",
  15412=>"000000000",
  15413=>"011001100",
  15414=>"001111110",
  15415=>"010001100",
  15416=>"101100010",
  15417=>"100110101",
  15418=>"000101111",
  15419=>"101110000",
  15420=>"000000100",
  15421=>"110100111",
  15422=>"110000000",
  15423=>"111110101",
  15424=>"011011001",
  15425=>"101000101",
  15426=>"010011001",
  15427=>"001111110",
  15428=>"000000110",
  15429=>"010010100",
  15430=>"100000100",
  15431=>"011100100",
  15432=>"100001110",
  15433=>"010001110",
  15434=>"010011000",
  15435=>"001111100",
  15436=>"011110001",
  15437=>"100001000",
  15438=>"011011101",
  15439=>"000010010",
  15440=>"100010111",
  15441=>"110111101",
  15442=>"010101010",
  15443=>"111101000",
  15444=>"110011111",
  15445=>"001101001",
  15446=>"110100000",
  15447=>"000001111",
  15448=>"100010001",
  15449=>"011101010",
  15450=>"100001000",
  15451=>"011001100",
  15452=>"011111101",
  15453=>"111011111",
  15454=>"111011110",
  15455=>"100000001",
  15456=>"001001110",
  15457=>"110111101",
  15458=>"111111110",
  15459=>"011101110",
  15460=>"000010110",
  15461=>"110100001",
  15462=>"001101101",
  15463=>"000111111",
  15464=>"001001100",
  15465=>"101111001",
  15466=>"110100011",
  15467=>"111101110",
  15468=>"100010101",
  15469=>"110110100",
  15470=>"000001110",
  15471=>"010111111",
  15472=>"001001010",
  15473=>"011100100",
  15474=>"111111111",
  15475=>"110010010",
  15476=>"010000000",
  15477=>"011111100",
  15478=>"010111001",
  15479=>"100100011",
  15480=>"111010100",
  15481=>"001110110",
  15482=>"110001011",
  15483=>"000110010",
  15484=>"111101110",
  15485=>"011000101",
  15486=>"010001110",
  15487=>"100001100",
  15488=>"011101111",
  15489=>"001110010",
  15490=>"100001101",
  15491=>"010001001",
  15492=>"110100001",
  15493=>"010110100",
  15494=>"010000011",
  15495=>"000100000",
  15496=>"110100010",
  15497=>"010110001",
  15498=>"101101000",
  15499=>"010111110",
  15500=>"101011011",
  15501=>"110011101",
  15502=>"000011100",
  15503=>"000001000",
  15504=>"010100000",
  15505=>"011000011",
  15506=>"110011111",
  15507=>"001000001",
  15508=>"111101110",
  15509=>"110111110",
  15510=>"010100101",
  15511=>"110111110",
  15512=>"001100100",
  15513=>"010111111",
  15514=>"000000011",
  15515=>"100110110",
  15516=>"000111011",
  15517=>"000001000",
  15518=>"000001100",
  15519=>"010001101",
  15520=>"101000100",
  15521=>"111000001",
  15522=>"111010001",
  15523=>"111010001",
  15524=>"101000100",
  15525=>"101011101",
  15526=>"001000010",
  15527=>"000101111",
  15528=>"011100000",
  15529=>"110001001",
  15530=>"000100000",
  15531=>"111111011",
  15532=>"111110011",
  15533=>"101111000",
  15534=>"100100110",
  15535=>"011101000",
  15536=>"001101010",
  15537=>"001110000",
  15538=>"100000000",
  15539=>"101110110",
  15540=>"000110100",
  15541=>"101000110",
  15542=>"111001101",
  15543=>"010110101",
  15544=>"000011000",
  15545=>"001111000",
  15546=>"101001111",
  15547=>"010010000",
  15548=>"001011000",
  15549=>"001101011",
  15550=>"101100001",
  15551=>"110111000",
  15552=>"010011001",
  15553=>"110101100",
  15554=>"100110011",
  15555=>"111111100",
  15556=>"000010000",
  15557=>"000001001",
  15558=>"100001010",
  15559=>"110001100",
  15560=>"111010110",
  15561=>"101011101",
  15562=>"001100001",
  15563=>"100010101",
  15564=>"101010111",
  15565=>"100000000",
  15566=>"001000100",
  15567=>"100110000",
  15568=>"011001011",
  15569=>"111100110",
  15570=>"000000110",
  15571=>"000010101",
  15572=>"100001110",
  15573=>"100111001",
  15574=>"111101101",
  15575=>"011100100",
  15576=>"100001000",
  15577=>"100100000",
  15578=>"011110000",
  15579=>"000101001",
  15580=>"111110001",
  15581=>"000110110",
  15582=>"101010110",
  15583=>"110110001",
  15584=>"001010101",
  15585=>"000110110",
  15586=>"111001010",
  15587=>"100001100",
  15588=>"001111101",
  15589=>"001000001",
  15590=>"110100001",
  15591=>"011111001",
  15592=>"000110011",
  15593=>"101011000",
  15594=>"111111000",
  15595=>"001110001",
  15596=>"111111111",
  15597=>"000001111",
  15598=>"101000001",
  15599=>"000001010",
  15600=>"001000011",
  15601=>"010100101",
  15602=>"001000010",
  15603=>"000010001",
  15604=>"010111011",
  15605=>"010010000",
  15606=>"000100011",
  15607=>"000010110",
  15608=>"110101100",
  15609=>"100011010",
  15610=>"110110001",
  15611=>"101010011",
  15612=>"101001010",
  15613=>"110010111",
  15614=>"010000000",
  15615=>"110010111",
  15616=>"001110100",
  15617=>"101111011",
  15618=>"010111110",
  15619=>"010010110",
  15620=>"001001000",
  15621=>"000010110",
  15622=>"111100000",
  15623=>"010101010",
  15624=>"000101001",
  15625=>"100010000",
  15626=>"100010000",
  15627=>"000001100",
  15628=>"110011111",
  15629=>"010000101",
  15630=>"110011111",
  15631=>"011000010",
  15632=>"011011000",
  15633=>"111110110",
  15634=>"111101110",
  15635=>"010011011",
  15636=>"001001100",
  15637=>"000010011",
  15638=>"000100111",
  15639=>"110011100",
  15640=>"010010110",
  15641=>"100010111",
  15642=>"010100010",
  15643=>"001100110",
  15644=>"000100110",
  15645=>"111010101",
  15646=>"011101010",
  15647=>"111110011",
  15648=>"000011001",
  15649=>"100010100",
  15650=>"111101110",
  15651=>"111010000",
  15652=>"010100011",
  15653=>"000101100",
  15654=>"000111111",
  15655=>"100000000",
  15656=>"111000101",
  15657=>"010100101",
  15658=>"111111010",
  15659=>"000010000",
  15660=>"110000011",
  15661=>"100000010",
  15662=>"001001011",
  15663=>"000110100",
  15664=>"010101011",
  15665=>"101101110",
  15666=>"011001110",
  15667=>"111010000",
  15668=>"100000010",
  15669=>"100100110",
  15670=>"001110011",
  15671=>"010101111",
  15672=>"100011110",
  15673=>"001011000",
  15674=>"111101110",
  15675=>"011101011",
  15676=>"001010101",
  15677=>"100000010",
  15678=>"100101100",
  15679=>"001000000",
  15680=>"000001101",
  15681=>"110001111",
  15682=>"101010101",
  15683=>"011010000",
  15684=>"010111011",
  15685=>"111000000",
  15686=>"101000001",
  15687=>"001100000",
  15688=>"100001010",
  15689=>"001000110",
  15690=>"010101111",
  15691=>"000011001",
  15692=>"110100111",
  15693=>"111011011",
  15694=>"100110100",
  15695=>"110001011",
  15696=>"000010011",
  15697=>"100100101",
  15698=>"100011011",
  15699=>"001111001",
  15700=>"001001000",
  15701=>"000101101",
  15702=>"000101100",
  15703=>"011101001",
  15704=>"001110000",
  15705=>"100011101",
  15706=>"010101100",
  15707=>"000011000",
  15708=>"011010101",
  15709=>"010000000",
  15710=>"001010011",
  15711=>"010101110",
  15712=>"110110010",
  15713=>"000000101",
  15714=>"111001101",
  15715=>"000011110",
  15716=>"010001001",
  15717=>"010110010",
  15718=>"100000011",
  15719=>"101010010",
  15720=>"011001011",
  15721=>"000111100",
  15722=>"111011000",
  15723=>"011111111",
  15724=>"001001001",
  15725=>"110111100",
  15726=>"000110001",
  15727=>"011100111",
  15728=>"001011111",
  15729=>"101001100",
  15730=>"011111110",
  15731=>"100010011",
  15732=>"110110000",
  15733=>"100001000",
  15734=>"101110001",
  15735=>"011010010",
  15736=>"011011010",
  15737=>"101011110",
  15738=>"011101001",
  15739=>"001100011",
  15740=>"011001101",
  15741=>"001111001",
  15742=>"001010110",
  15743=>"101101110",
  15744=>"011000111",
  15745=>"100010010",
  15746=>"111110000",
  15747=>"010001111",
  15748=>"011101110",
  15749=>"010001001",
  15750=>"101111110",
  15751=>"101000001",
  15752=>"000110001",
  15753=>"011111111",
  15754=>"010001100",
  15755=>"010110011",
  15756=>"010110011",
  15757=>"010111010",
  15758=>"100011111",
  15759=>"000010000",
  15760=>"101010000",
  15761=>"000001111",
  15762=>"101011111",
  15763=>"011010111",
  15764=>"010111101",
  15765=>"111110001",
  15766=>"100100111",
  15767=>"100010001",
  15768=>"100110001",
  15769=>"010100111",
  15770=>"100101101",
  15771=>"011010101",
  15772=>"010010010",
  15773=>"101110110",
  15774=>"101000010",
  15775=>"111011111",
  15776=>"100101101",
  15777=>"100011000",
  15778=>"100010000",
  15779=>"000001101",
  15780=>"010111100",
  15781=>"000111011",
  15782=>"111101011",
  15783=>"100001001",
  15784=>"111101001",
  15785=>"001000110",
  15786=>"001010101",
  15787=>"001101010",
  15788=>"111011111",
  15789=>"001001101",
  15790=>"011110010",
  15791=>"001010101",
  15792=>"001010011",
  15793=>"110110000",
  15794=>"010001001",
  15795=>"110100011",
  15796=>"011111101",
  15797=>"000010000",
  15798=>"000110101",
  15799=>"100100001",
  15800=>"110111100",
  15801=>"100001111",
  15802=>"001100000",
  15803=>"000000110",
  15804=>"000100011",
  15805=>"100001001",
  15806=>"111111001",
  15807=>"010011101",
  15808=>"001001010",
  15809=>"111100000",
  15810=>"110001111",
  15811=>"010011111",
  15812=>"000100101",
  15813=>"100001001",
  15814=>"011011011",
  15815=>"001000000",
  15816=>"111011111",
  15817=>"100100101",
  15818=>"101000010",
  15819=>"010110101",
  15820=>"110110101",
  15821=>"110111001",
  15822=>"000000010",
  15823=>"011100001",
  15824=>"111011011",
  15825=>"000011111",
  15826=>"101000001",
  15827=>"110101101",
  15828=>"011111000",
  15829=>"011011110",
  15830=>"011000010",
  15831=>"000100000",
  15832=>"111100001",
  15833=>"001101010",
  15834=>"011000000",
  15835=>"011101000",
  15836=>"101100011",
  15837=>"000000000",
  15838=>"101100010",
  15839=>"001111010",
  15840=>"110000110",
  15841=>"110010010",
  15842=>"000001110",
  15843=>"101111010",
  15844=>"000100110",
  15845=>"010111001",
  15846=>"111000001",
  15847=>"011000001",
  15848=>"101000010",
  15849=>"101110100",
  15850=>"100110100",
  15851=>"010111101",
  15852=>"000101001",
  15853=>"111010000",
  15854=>"000100000",
  15855=>"110111000",
  15856=>"000110001",
  15857=>"100011001",
  15858=>"110110111",
  15859=>"110101110",
  15860=>"001100101",
  15861=>"000000110",
  15862=>"111001101",
  15863=>"000101000",
  15864=>"000001011",
  15865=>"111101110",
  15866=>"001010101",
  15867=>"101111110",
  15868=>"100011111",
  15869=>"001111110",
  15870=>"111101011",
  15871=>"100011001",
  15872=>"110111010",
  15873=>"000101011",
  15874=>"010111011",
  15875=>"011010000",
  15876=>"010101111",
  15877=>"000011111",
  15878=>"100000110",
  15879=>"001100101",
  15880=>"010000010",
  15881=>"111000100",
  15882=>"001001110",
  15883=>"010111000",
  15884=>"001001010",
  15885=>"011011110",
  15886=>"101101101",
  15887=>"101000010",
  15888=>"100011001",
  15889=>"010010110",
  15890=>"010101010",
  15891=>"011100011",
  15892=>"101001000",
  15893=>"001110001",
  15894=>"111100011",
  15895=>"111011001",
  15896=>"101010001",
  15897=>"000101011",
  15898=>"001001110",
  15899=>"011101110",
  15900=>"011000100",
  15901=>"001000000",
  15902=>"111000111",
  15903=>"100000011",
  15904=>"001100111",
  15905=>"111011001",
  15906=>"001010111",
  15907=>"111100000",
  15908=>"110010010",
  15909=>"110100100",
  15910=>"001100011",
  15911=>"011000000",
  15912=>"110100100",
  15913=>"111100010",
  15914=>"100111011",
  15915=>"110101110",
  15916=>"101001001",
  15917=>"011011001",
  15918=>"101110000",
  15919=>"000110011",
  15920=>"100100001",
  15921=>"010110110",
  15922=>"100100000",
  15923=>"110100000",
  15924=>"001011010",
  15925=>"011000101",
  15926=>"001101100",
  15927=>"100001100",
  15928=>"010000001",
  15929=>"101010001",
  15930=>"111111010",
  15931=>"111111001",
  15932=>"010100100",
  15933=>"010110100",
  15934=>"111100111",
  15935=>"001100100",
  15936=>"100101001",
  15937=>"111100001",
  15938=>"011001110",
  15939=>"011001000",
  15940=>"000110000",
  15941=>"110100000",
  15942=>"000010011",
  15943=>"111001001",
  15944=>"000110100",
  15945=>"011111100",
  15946=>"000100000",
  15947=>"011000111",
  15948=>"010110000",
  15949=>"101000000",
  15950=>"101111110",
  15951=>"111101011",
  15952=>"000011000",
  15953=>"010111000",
  15954=>"101101110",
  15955=>"100100010",
  15956=>"110110001",
  15957=>"111010011",
  15958=>"100000001",
  15959=>"000100110",
  15960=>"101001000",
  15961=>"101000100",
  15962=>"000110101",
  15963=>"001001001",
  15964=>"100010101",
  15965=>"101010110",
  15966=>"001101010",
  15967=>"110110111",
  15968=>"011001100",
  15969=>"011011111",
  15970=>"111010101",
  15971=>"100110110",
  15972=>"011011001",
  15973=>"000000101",
  15974=>"110101011",
  15975=>"000110100",
  15976=>"000001101",
  15977=>"001001101",
  15978=>"100010111",
  15979=>"111100011",
  15980=>"110101001",
  15981=>"101110110",
  15982=>"011111100",
  15983=>"101101010",
  15984=>"100111000",
  15985=>"100101100",
  15986=>"011010000",
  15987=>"010001111",
  15988=>"001110101",
  15989=>"101001111",
  15990=>"011010101",
  15991=>"010000010",
  15992=>"011001110",
  15993=>"001010001",
  15994=>"000011001",
  15995=>"101010111",
  15996=>"011000101",
  15997=>"110000100",
  15998=>"010011110",
  15999=>"010110000",
  16000=>"000011011",
  16001=>"110110011",
  16002=>"111010101",
  16003=>"111000001",
  16004=>"100101111",
  16005=>"101100010",
  16006=>"101000001",
  16007=>"101001100",
  16008=>"011010110",
  16009=>"001000010",
  16010=>"111110100",
  16011=>"010000000",
  16012=>"000100111",
  16013=>"011000101",
  16014=>"000011101",
  16015=>"110101100",
  16016=>"011111001",
  16017=>"101100110",
  16018=>"110011110",
  16019=>"000000001",
  16020=>"110011001",
  16021=>"010000101",
  16022=>"100101010",
  16023=>"011100001",
  16024=>"110111001",
  16025=>"010000000",
  16026=>"001111111",
  16027=>"011000010",
  16028=>"010100001",
  16029=>"110101100",
  16030=>"010100100",
  16031=>"000110101",
  16032=>"011001111",
  16033=>"010000110",
  16034=>"100011000",
  16035=>"001110110",
  16036=>"000000000",
  16037=>"110111001",
  16038=>"110000110",
  16039=>"001110100",
  16040=>"110000000",
  16041=>"000001001",
  16042=>"101000011",
  16043=>"000000011",
  16044=>"010000001",
  16045=>"111010010",
  16046=>"000000010",
  16047=>"110100010",
  16048=>"111111000",
  16049=>"111001100",
  16050=>"100010010",
  16051=>"100000110",
  16052=>"011001001",
  16053=>"001110100",
  16054=>"110000000",
  16055=>"100111101",
  16056=>"000111000",
  16057=>"110001000",
  16058=>"011101010",
  16059=>"001101100",
  16060=>"100000111",
  16061=>"000011111",
  16062=>"101000111",
  16063=>"111101101",
  16064=>"010111101",
  16065=>"001111001",
  16066=>"100111000",
  16067=>"001000000",
  16068=>"110111110",
  16069=>"100100110",
  16070=>"101111010",
  16071=>"011110101",
  16072=>"010111001",
  16073=>"100011000",
  16074=>"011001010",
  16075=>"000010001",
  16076=>"011100011",
  16077=>"110000100",
  16078=>"000101111",
  16079=>"110010011",
  16080=>"110111011",
  16081=>"011001110",
  16082=>"101001011",
  16083=>"000101010",
  16084=>"010110000",
  16085=>"010001000",
  16086=>"111010100",
  16087=>"101010000",
  16088=>"110000111",
  16089=>"111101110",
  16090=>"101000101",
  16091=>"000000100",
  16092=>"001110111",
  16093=>"100101001",
  16094=>"111100110",
  16095=>"011000101",
  16096=>"001101111",
  16097=>"011001100",
  16098=>"100000111",
  16099=>"100101110",
  16100=>"011001000",
  16101=>"011011110",
  16102=>"110011100",
  16103=>"010101101",
  16104=>"011111000",
  16105=>"010010110",
  16106=>"011101111",
  16107=>"000001011",
  16108=>"000011111",
  16109=>"111000111",
  16110=>"111000000",
  16111=>"000101110",
  16112=>"100111000",
  16113=>"100111011",
  16114=>"010101111",
  16115=>"010011111",
  16116=>"010011000",
  16117=>"001101101",
  16118=>"000001010",
  16119=>"001101110",
  16120=>"011111000",
  16121=>"001101111",
  16122=>"000111000",
  16123=>"001000111",
  16124=>"101100001",
  16125=>"110101100",
  16126=>"011000011",
  16127=>"110101110",
  16128=>"100010101",
  16129=>"001111111",
  16130=>"101110010",
  16131=>"000010010",
  16132=>"100011001",
  16133=>"110000000",
  16134=>"011110000",
  16135=>"100111000",
  16136=>"001110101",
  16137=>"101100011",
  16138=>"110011010",
  16139=>"010110010",
  16140=>"000000101",
  16141=>"111110111",
  16142=>"010000100",
  16143=>"111000000",
  16144=>"010000111",
  16145=>"000001010",
  16146=>"000001000",
  16147=>"011101000",
  16148=>"001110011",
  16149=>"110001011",
  16150=>"010001101",
  16151=>"000011010",
  16152=>"011011111",
  16153=>"011001101",
  16154=>"100011001",
  16155=>"110001110",
  16156=>"011001011",
  16157=>"110000110",
  16158=>"000110111",
  16159=>"000011100",
  16160=>"100101100",
  16161=>"001011100",
  16162=>"100010110",
  16163=>"111010000",
  16164=>"001001110",
  16165=>"001101111",
  16166=>"011111010",
  16167=>"011110000",
  16168=>"000111001",
  16169=>"010001110",
  16170=>"101011110",
  16171=>"101110101",
  16172=>"010110110",
  16173=>"110100100",
  16174=>"001101010",
  16175=>"001010001",
  16176=>"001010110",
  16177=>"111011100",
  16178=>"101010101",
  16179=>"100100010",
  16180=>"000101000",
  16181=>"101100100",
  16182=>"000010111",
  16183=>"110011111",
  16184=>"000010100",
  16185=>"101101101",
  16186=>"010110010",
  16187=>"101100000",
  16188=>"110010100",
  16189=>"001010011",
  16190=>"000011011",
  16191=>"010101111",
  16192=>"100011001",
  16193=>"100011010",
  16194=>"010011000",
  16195=>"001000010",
  16196=>"100011010",
  16197=>"010100101",
  16198=>"111001110",
  16199=>"011001101",
  16200=>"000010100",
  16201=>"111111100",
  16202=>"111110111",
  16203=>"001100001",
  16204=>"011101010",
  16205=>"010001100",
  16206=>"010101101",
  16207=>"000010000",
  16208=>"110111010",
  16209=>"001010101",
  16210=>"001010010",
  16211=>"000110011",
  16212=>"011010000",
  16213=>"111000010",
  16214=>"000010111",
  16215=>"110110101",
  16216=>"000101010",
  16217=>"111111101",
  16218=>"100111110",
  16219=>"001111000",
  16220=>"000101011",
  16221=>"010110100",
  16222=>"101100000",
  16223=>"010001100",
  16224=>"111111110",
  16225=>"000000010",
  16226=>"111101011",
  16227=>"001011000",
  16228=>"110001101",
  16229=>"000010000",
  16230=>"111110111",
  16231=>"011111111",
  16232=>"011000001",
  16233=>"010110001",
  16234=>"001011100",
  16235=>"000001001",
  16236=>"000011001",
  16237=>"001010110",
  16238=>"001101100",
  16239=>"110010010",
  16240=>"100111101",
  16241=>"001100100",
  16242=>"111100100",
  16243=>"011100010",
  16244=>"100111011",
  16245=>"001110001",
  16246=>"100111101",
  16247=>"101000000",
  16248=>"011011100",
  16249=>"011110011",
  16250=>"101100100",
  16251=>"001011111",
  16252=>"000000001",
  16253=>"010100100",
  16254=>"010010011",
  16255=>"110111110",
  16256=>"101101101",
  16257=>"100111111",
  16258=>"000001010",
  16259=>"100100101",
  16260=>"111100101",
  16261=>"000100001",
  16262=>"110011000",
  16263=>"000010001",
  16264=>"011001001",
  16265=>"000110111",
  16266=>"111000001",
  16267=>"000111110",
  16268=>"010011000",
  16269=>"001110110",
  16270=>"001110000",
  16271=>"010000001",
  16272=>"101101111",
  16273=>"101000001",
  16274=>"000000010",
  16275=>"110110110",
  16276=>"001110001",
  16277=>"001010001",
  16278=>"000000101",
  16279=>"110000110",
  16280=>"110001011",
  16281=>"000010101",
  16282=>"011110011",
  16283=>"100000101",
  16284=>"100010100",
  16285=>"001100111",
  16286=>"001011000",
  16287=>"111101110",
  16288=>"011101011",
  16289=>"011001101",
  16290=>"111111000",
  16291=>"010100100",
  16292=>"000101011",
  16293=>"010011010",
  16294=>"110010000",
  16295=>"010001100",
  16296=>"010100101",
  16297=>"001000101",
  16298=>"111001011",
  16299=>"111001111",
  16300=>"000001100",
  16301=>"001110111",
  16302=>"000001011",
  16303=>"001111011",
  16304=>"111011101",
  16305=>"111000111",
  16306=>"101100001",
  16307=>"000000001",
  16308=>"000110111",
  16309=>"100101011",
  16310=>"001000101",
  16311=>"110110110",
  16312=>"001101110",
  16313=>"001011010",
  16314=>"110010010",
  16315=>"111111001",
  16316=>"000011010",
  16317=>"100001110",
  16318=>"101110100",
  16319=>"000010100",
  16320=>"110000001",
  16321=>"011110101",
  16322=>"011010010",
  16323=>"100101101",
  16324=>"001010001",
  16325=>"010000001",
  16326=>"111101101",
  16327=>"110101100",
  16328=>"001001011",
  16329=>"001000000",
  16330=>"100110100",
  16331=>"101101000",
  16332=>"111111001",
  16333=>"101101010",
  16334=>"101010110",
  16335=>"000100110",
  16336=>"110111110",
  16337=>"011010010",
  16338=>"010000100",
  16339=>"011001100",
  16340=>"101101111",
  16341=>"001100111",
  16342=>"101111100",
  16343=>"110101100",
  16344=>"100010111",
  16345=>"010101100",
  16346=>"100110001",
  16347=>"110001011",
  16348=>"111000100",
  16349=>"010001100",
  16350=>"000001000",
  16351=>"010111101",
  16352=>"111111101",
  16353=>"100110010",
  16354=>"001001001",
  16355=>"000111101",
  16356=>"000010000",
  16357=>"111010001",
  16358=>"000101000",
  16359=>"101001010",
  16360=>"100011101",
  16361=>"001010111",
  16362=>"001101110",
  16363=>"001100111",
  16364=>"100010011",
  16365=>"000111010",
  16366=>"000100101",
  16367=>"101100111",
  16368=>"011110011",
  16369=>"000011111",
  16370=>"000101101",
  16371=>"111110010",
  16372=>"001010101",
  16373=>"010011111",
  16374=>"011001101",
  16375=>"100111110",
  16376=>"111110110",
  16377=>"101110111",
  16378=>"001100101",
  16379=>"111010001",
  16380=>"001110111",
  16381=>"110001001",
  16382=>"010001001",
  16383=>"101100001",
  16384=>"010000000",
  16385=>"000001000",
  16386=>"010100101",
  16387=>"110100101",
  16388=>"011010010",
  16389=>"011110111",
  16390=>"001010000",
  16391=>"111010011",
  16392=>"001110000",
  16393=>"101011111",
  16394=>"000110101",
  16395=>"111110010",
  16396=>"100011111",
  16397=>"111100011",
  16398=>"000001101",
  16399=>"100101110",
  16400=>"001010111",
  16401=>"010000000",
  16402=>"011110110",
  16403=>"101111111",
  16404=>"010100000",
  16405=>"011111010",
  16406=>"000101011",
  16407=>"010110000",
  16408=>"111100111",
  16409=>"000000100",
  16410=>"111010110",
  16411=>"001111011",
  16412=>"100111110",
  16413=>"010100010",
  16414=>"011010101",
  16415=>"001111100",
  16416=>"011100111",
  16417=>"111111101",
  16418=>"011100110",
  16419=>"010100100",
  16420=>"011111000",
  16421=>"000000000",
  16422=>"010001000",
  16423=>"101101010",
  16424=>"101101010",
  16425=>"000100001",
  16426=>"111101110",
  16427=>"000010111",
  16428=>"010001101",
  16429=>"000110111",
  16430=>"110100100",
  16431=>"001101001",
  16432=>"111111111",
  16433=>"111011111",
  16434=>"110011111",
  16435=>"010111101",
  16436=>"101100110",
  16437=>"000001000",
  16438=>"111001001",
  16439=>"001110111",
  16440=>"000000010",
  16441=>"011111101",
  16442=>"110100101",
  16443=>"010101110",
  16444=>"000111010",
  16445=>"001001000",
  16446=>"000000100",
  16447=>"100001101",
  16448=>"001111110",
  16449=>"001110000",
  16450=>"001101000",
  16451=>"001010001",
  16452=>"010001011",
  16453=>"010000000",
  16454=>"111001000",
  16455=>"011100011",
  16456=>"010010001",
  16457=>"101000100",
  16458=>"011111001",
  16459=>"110001101",
  16460=>"010100101",
  16461=>"100010111",
  16462=>"110100110",
  16463=>"111100010",
  16464=>"010010110",
  16465=>"110111000",
  16466=>"001111011",
  16467=>"001100111",
  16468=>"001001010",
  16469=>"110110101",
  16470=>"100110011",
  16471=>"000011001",
  16472=>"100010111",
  16473=>"011110100",
  16474=>"001011101",
  16475=>"001001110",
  16476=>"000011111",
  16477=>"011010000",
  16478=>"110001010",
  16479=>"001000011",
  16480=>"111111011",
  16481=>"111110011",
  16482=>"110101110",
  16483=>"111100010",
  16484=>"101011111",
  16485=>"010110001",
  16486=>"101101111",
  16487=>"111101110",
  16488=>"110011010",
  16489=>"111011000",
  16490=>"101111010",
  16491=>"010101101",
  16492=>"000110111",
  16493=>"010010000",
  16494=>"010111111",
  16495=>"110001010",
  16496=>"000101011",
  16497=>"100011001",
  16498=>"100111101",
  16499=>"010110110",
  16500=>"100010101",
  16501=>"101011111",
  16502=>"001111011",
  16503=>"111101111",
  16504=>"101111111",
  16505=>"000001011",
  16506=>"000100001",
  16507=>"011111010",
  16508=>"011110000",
  16509=>"001001000",
  16510=>"101011011",
  16511=>"110000010",
  16512=>"000011010",
  16513=>"010111001",
  16514=>"110011010",
  16515=>"110100001",
  16516=>"110010000",
  16517=>"111010011",
  16518=>"001000011",
  16519=>"100001101",
  16520=>"011001100",
  16521=>"010111101",
  16522=>"101011111",
  16523=>"001100110",
  16524=>"111110010",
  16525=>"110011000",
  16526=>"110101010",
  16527=>"111100000",
  16528=>"111011000",
  16529=>"001100110",
  16530=>"100110111",
  16531=>"011011110",
  16532=>"100100010",
  16533=>"010100000",
  16534=>"011100100",
  16535=>"011000110",
  16536=>"010001110",
  16537=>"000010000",
  16538=>"100110101",
  16539=>"111000001",
  16540=>"101001110",
  16541=>"110011111",
  16542=>"001101011",
  16543=>"010111100",
  16544=>"001101000",
  16545=>"101000001",
  16546=>"000011111",
  16547=>"000011010",
  16548=>"101010111",
  16549=>"011100001",
  16550=>"100110000",
  16551=>"100000100",
  16552=>"001101101",
  16553=>"110101011",
  16554=>"000111010",
  16555=>"001011000",
  16556=>"001001011",
  16557=>"110001100",
  16558=>"110011100",
  16559=>"011111001",
  16560=>"111000011",
  16561=>"000101100",
  16562=>"010100001",
  16563=>"000001000",
  16564=>"001010001",
  16565=>"101000001",
  16566=>"111100101",
  16567=>"111101101",
  16568=>"011010001",
  16569=>"110100111",
  16570=>"010000001",
  16571=>"111011001",
  16572=>"011010111",
  16573=>"111111111",
  16574=>"011111101",
  16575=>"110011001",
  16576=>"010011100",
  16577=>"111001011",
  16578=>"010101111",
  16579=>"111101100",
  16580=>"101101111",
  16581=>"011001110",
  16582=>"111011000",
  16583=>"100000010",
  16584=>"010100100",
  16585=>"000110000",
  16586=>"001000110",
  16587=>"000001000",
  16588=>"011101010",
  16589=>"000001111",
  16590=>"101011011",
  16591=>"001111011",
  16592=>"110011000",
  16593=>"001001101",
  16594=>"001001000",
  16595=>"111100000",
  16596=>"001001101",
  16597=>"101010001",
  16598=>"110011000",
  16599=>"111010111",
  16600=>"000001011",
  16601=>"111111100",
  16602=>"001000000",
  16603=>"110000111",
  16604=>"111011001",
  16605=>"101110100",
  16606=>"100110110",
  16607=>"111111000",
  16608=>"100101000",
  16609=>"000000100",
  16610=>"001010001",
  16611=>"001000110",
  16612=>"000011100",
  16613=>"010011001",
  16614=>"011110101",
  16615=>"111001010",
  16616=>"111011010",
  16617=>"010110011",
  16618=>"001001000",
  16619=>"111011010",
  16620=>"001000110",
  16621=>"000100110",
  16622=>"010000011",
  16623=>"101111111",
  16624=>"011110111",
  16625=>"100000111",
  16626=>"000010101",
  16627=>"001001001",
  16628=>"100001011",
  16629=>"011110001",
  16630=>"110100001",
  16631=>"010101010",
  16632=>"101110000",
  16633=>"111010110",
  16634=>"000010010",
  16635=>"011000000",
  16636=>"011101111",
  16637=>"110010010",
  16638=>"001100000",
  16639=>"011100011",
  16640=>"000100101",
  16641=>"011001000",
  16642=>"101110010",
  16643=>"010001111",
  16644=>"100110001",
  16645=>"011100010",
  16646=>"010000000",
  16647=>"111000100",
  16648=>"010100110",
  16649=>"110001000",
  16650=>"010000010",
  16651=>"011010110",
  16652=>"101001001",
  16653=>"000001110",
  16654=>"110010101",
  16655=>"001001100",
  16656=>"010010001",
  16657=>"011010010",
  16658=>"110111101",
  16659=>"111111011",
  16660=>"111011000",
  16661=>"000101000",
  16662=>"101101100",
  16663=>"001110100",
  16664=>"000011101",
  16665=>"000101101",
  16666=>"110101010",
  16667=>"101001011",
  16668=>"011011001",
  16669=>"000110010",
  16670=>"110110011",
  16671=>"010101000",
  16672=>"010010111",
  16673=>"100000001",
  16674=>"100011111",
  16675=>"111000000",
  16676=>"111110100",
  16677=>"100100001",
  16678=>"100110010",
  16679=>"001010100",
  16680=>"000001110",
  16681=>"000100010",
  16682=>"000000100",
  16683=>"101101111",
  16684=>"101100000",
  16685=>"001110100",
  16686=>"011111011",
  16687=>"011010111",
  16688=>"010000000",
  16689=>"110010101",
  16690=>"111111010",
  16691=>"011110101",
  16692=>"001101101",
  16693=>"001010100",
  16694=>"000111111",
  16695=>"010011001",
  16696=>"100000011",
  16697=>"100101111",
  16698=>"110111100",
  16699=>"000000001",
  16700=>"111100000",
  16701=>"101110100",
  16702=>"000100100",
  16703=>"000011110",
  16704=>"110111101",
  16705=>"000010110",
  16706=>"000100111",
  16707=>"000110001",
  16708=>"101100100",
  16709=>"011000111",
  16710=>"101000011",
  16711=>"010110100",
  16712=>"001000011",
  16713=>"000000010",
  16714=>"111011111",
  16715=>"100010110",
  16716=>"111001011",
  16717=>"111100110",
  16718=>"110011010",
  16719=>"110000100",
  16720=>"010011001",
  16721=>"001110111",
  16722=>"000110100",
  16723=>"011000010",
  16724=>"011001110",
  16725=>"010000010",
  16726=>"110010101",
  16727=>"010011110",
  16728=>"000011110",
  16729=>"010011111",
  16730=>"111010011",
  16731=>"011010100",
  16732=>"010011010",
  16733=>"011111010",
  16734=>"101010110",
  16735=>"110111011",
  16736=>"101000001",
  16737=>"001010010",
  16738=>"000100101",
  16739=>"001010101",
  16740=>"100001010",
  16741=>"000110101",
  16742=>"101101101",
  16743=>"101101011",
  16744=>"110000110",
  16745=>"011100110",
  16746=>"101101110",
  16747=>"011101010",
  16748=>"100101010",
  16749=>"111101011",
  16750=>"000010111",
  16751=>"111101101",
  16752=>"000010100",
  16753=>"010011010",
  16754=>"110001100",
  16755=>"011001111",
  16756=>"010101101",
  16757=>"100010001",
  16758=>"001111111",
  16759=>"101010100",
  16760=>"000000010",
  16761=>"101101110",
  16762=>"001000101",
  16763=>"101110011",
  16764=>"000101011",
  16765=>"011110010",
  16766=>"110001000",
  16767=>"011000010",
  16768=>"010000111",
  16769=>"101101010",
  16770=>"101010101",
  16771=>"011010010",
  16772=>"101110110",
  16773=>"010110110",
  16774=>"110111001",
  16775=>"000000010",
  16776=>"001011000",
  16777=>"110111011",
  16778=>"011110001",
  16779=>"110100101",
  16780=>"000100011",
  16781=>"011100010",
  16782=>"011000101",
  16783=>"001010011",
  16784=>"110110010",
  16785=>"101001010",
  16786=>"111111111",
  16787=>"011111101",
  16788=>"110100111",
  16789=>"111100011",
  16790=>"000011100",
  16791=>"011110001",
  16792=>"001011100",
  16793=>"001110001",
  16794=>"011001100",
  16795=>"001101010",
  16796=>"011010010",
  16797=>"000000010",
  16798=>"111011100",
  16799=>"100011111",
  16800=>"001011110",
  16801=>"111011110",
  16802=>"000100111",
  16803=>"111011100",
  16804=>"100001001",
  16805=>"101100110",
  16806=>"101000000",
  16807=>"010011011",
  16808=>"011011010",
  16809=>"100111000",
  16810=>"011000100",
  16811=>"001010001",
  16812=>"000010110",
  16813=>"110101110",
  16814=>"011000100",
  16815=>"000110010",
  16816=>"001000111",
  16817=>"101010111",
  16818=>"000001000",
  16819=>"000110000",
  16820=>"010110110",
  16821=>"011011110",
  16822=>"000111110",
  16823=>"001100100",
  16824=>"010001001",
  16825=>"010000101",
  16826=>"000000001",
  16827=>"000001010",
  16828=>"000101100",
  16829=>"000111001",
  16830=>"111111101",
  16831=>"110110001",
  16832=>"011011000",
  16833=>"101001001",
  16834=>"011110111",
  16835=>"010111101",
  16836=>"001101101",
  16837=>"111011001",
  16838=>"100000000",
  16839=>"010111001",
  16840=>"000110010",
  16841=>"010000011",
  16842=>"100010101",
  16843=>"010010010",
  16844=>"110010010",
  16845=>"010010111",
  16846=>"111001000",
  16847=>"110011000",
  16848=>"000111000",
  16849=>"011100110",
  16850=>"101110110",
  16851=>"000111100",
  16852=>"111111010",
  16853=>"111001111",
  16854=>"111100011",
  16855=>"110000110",
  16856=>"100111000",
  16857=>"011011011",
  16858=>"110001010",
  16859=>"010000100",
  16860=>"100110100",
  16861=>"111011000",
  16862=>"000010001",
  16863=>"111110010",
  16864=>"110101001",
  16865=>"111110001",
  16866=>"000000110",
  16867=>"000010110",
  16868=>"001000100",
  16869=>"110011001",
  16870=>"101010111",
  16871=>"100010011",
  16872=>"100001001",
  16873=>"001110100",
  16874=>"110111011",
  16875=>"101000011",
  16876=>"010000000",
  16877=>"010110111",
  16878=>"001110101",
  16879=>"110111111",
  16880=>"101111100",
  16881=>"011110010",
  16882=>"100000001",
  16883=>"011001010",
  16884=>"111010010",
  16885=>"000110010",
  16886=>"100100001",
  16887=>"100000101",
  16888=>"010001110",
  16889=>"000000001",
  16890=>"000100011",
  16891=>"000011100",
  16892=>"001011101",
  16893=>"011111011",
  16894=>"000110000",
  16895=>"111111100",
  16896=>"111000100",
  16897=>"100100000",
  16898=>"100100100",
  16899=>"010011100",
  16900=>"100000011",
  16901=>"111010000",
  16902=>"111100100",
  16903=>"001001001",
  16904=>"111010010",
  16905=>"101111001",
  16906=>"110110100",
  16907=>"011000011",
  16908=>"110101110",
  16909=>"001110011",
  16910=>"000110001",
  16911=>"100000101",
  16912=>"010010000",
  16913=>"010001000",
  16914=>"001010100",
  16915=>"111000010",
  16916=>"111000101",
  16917=>"010100101",
  16918=>"110010000",
  16919=>"000110000",
  16920=>"111000010",
  16921=>"010010111",
  16922=>"010000010",
  16923=>"001110110",
  16924=>"010010101",
  16925=>"111101100",
  16926=>"011010001",
  16927=>"001100101",
  16928=>"011011100",
  16929=>"101010001",
  16930=>"000111010",
  16931=>"111010010",
  16932=>"111111100",
  16933=>"110100111",
  16934=>"101010111",
  16935=>"010001111",
  16936=>"000100111",
  16937=>"011111111",
  16938=>"100010110",
  16939=>"101100110",
  16940=>"000010011",
  16941=>"100001110",
  16942=>"010001001",
  16943=>"000100010",
  16944=>"011110000",
  16945=>"000111000",
  16946=>"010111011",
  16947=>"111110100",
  16948=>"111000010",
  16949=>"110111010",
  16950=>"001010100",
  16951=>"001110011",
  16952=>"100110010",
  16953=>"110000010",
  16954=>"101101011",
  16955=>"101111111",
  16956=>"010000001",
  16957=>"100010011",
  16958=>"010110010",
  16959=>"011110001",
  16960=>"000100110",
  16961=>"111101100",
  16962=>"010011000",
  16963=>"110110110",
  16964=>"001101011",
  16965=>"111011111",
  16966=>"010111111",
  16967=>"100111110",
  16968=>"000001111",
  16969=>"000100101",
  16970=>"110101110",
  16971=>"110110101",
  16972=>"111000101",
  16973=>"011010101",
  16974=>"001000110",
  16975=>"111001111",
  16976=>"111101010",
  16977=>"011011000",
  16978=>"110010101",
  16979=>"010010111",
  16980=>"101011110",
  16981=>"010110111",
  16982=>"000111001",
  16983=>"010110011",
  16984=>"111111000",
  16985=>"111100000",
  16986=>"000000000",
  16987=>"111010100",
  16988=>"010001011",
  16989=>"100010000",
  16990=>"100111110",
  16991=>"000111110",
  16992=>"001110000",
  16993=>"000000101",
  16994=>"001111101",
  16995=>"100111110",
  16996=>"100100010",
  16997=>"110010000",
  16998=>"000111100",
  16999=>"011110011",
  17000=>"010110010",
  17001=>"000110000",
  17002=>"101010011",
  17003=>"011100000",
  17004=>"000001101",
  17005=>"010011111",
  17006=>"111111111",
  17007=>"000000101",
  17008=>"110001100",
  17009=>"001110100",
  17010=>"100100101",
  17011=>"111111001",
  17012=>"100010100",
  17013=>"001110101",
  17014=>"111111100",
  17015=>"001001100",
  17016=>"001011000",
  17017=>"010110101",
  17018=>"010101001",
  17019=>"100100001",
  17020=>"111111010",
  17021=>"011000001",
  17022=>"110100100",
  17023=>"110101011",
  17024=>"001000011",
  17025=>"101111110",
  17026=>"000101110",
  17027=>"001001000",
  17028=>"011101011",
  17029=>"000000011",
  17030=>"011010001",
  17031=>"111010010",
  17032=>"011000101",
  17033=>"010010100",
  17034=>"110101111",
  17035=>"011111011",
  17036=>"000111011",
  17037=>"101000011",
  17038=>"000110010",
  17039=>"000010010",
  17040=>"011101110",
  17041=>"001100000",
  17042=>"011001100",
  17043=>"111111110",
  17044=>"110100101",
  17045=>"111000110",
  17046=>"111110110",
  17047=>"101110111",
  17048=>"000101111",
  17049=>"100010000",
  17050=>"110010111",
  17051=>"000111011",
  17052=>"110110010",
  17053=>"110111110",
  17054=>"000100101",
  17055=>"100000100",
  17056=>"001111010",
  17057=>"011100100",
  17058=>"101110000",
  17059=>"110101100",
  17060=>"010010100",
  17061=>"111001000",
  17062=>"000010100",
  17063=>"000100010",
  17064=>"001000011",
  17065=>"111110001",
  17066=>"110010011",
  17067=>"100011100",
  17068=>"101110110",
  17069=>"100001011",
  17070=>"000011110",
  17071=>"000000000",
  17072=>"000010000",
  17073=>"011101001",
  17074=>"111100001",
  17075=>"110100100",
  17076=>"011010010",
  17077=>"010000101",
  17078=>"110110100",
  17079=>"100001111",
  17080=>"100000111",
  17081=>"100110111",
  17082=>"000000001",
  17083=>"101011110",
  17084=>"000000010",
  17085=>"110110101",
  17086=>"000010000",
  17087=>"110101001",
  17088=>"111001010",
  17089=>"111010110",
  17090=>"111010000",
  17091=>"110001010",
  17092=>"101010101",
  17093=>"100000001",
  17094=>"101100010",
  17095=>"011111111",
  17096=>"110110010",
  17097=>"000011110",
  17098=>"011000011",
  17099=>"000100111",
  17100=>"101001011",
  17101=>"000000010",
  17102=>"111010100",
  17103=>"000100011",
  17104=>"000110110",
  17105=>"000100000",
  17106=>"101100000",
  17107=>"000100001",
  17108=>"111111011",
  17109=>"111111110",
  17110=>"110001010",
  17111=>"000011110",
  17112=>"011011010",
  17113=>"110101111",
  17114=>"111101001",
  17115=>"010001000",
  17116=>"100001010",
  17117=>"011011010",
  17118=>"101101011",
  17119=>"101011101",
  17120=>"010000001",
  17121=>"001000000",
  17122=>"100110011",
  17123=>"100001000",
  17124=>"011011110",
  17125=>"000000000",
  17126=>"001000110",
  17127=>"101101101",
  17128=>"001000110",
  17129=>"000011010",
  17130=>"000100010",
  17131=>"111001010",
  17132=>"000110111",
  17133=>"101100101",
  17134=>"100010100",
  17135=>"110000011",
  17136=>"111001111",
  17137=>"010100000",
  17138=>"000110000",
  17139=>"001000100",
  17140=>"001000001",
  17141=>"101010100",
  17142=>"110000001",
  17143=>"111000111",
  17144=>"101001011",
  17145=>"001100101",
  17146=>"101101001",
  17147=>"001011101",
  17148=>"000110000",
  17149=>"111110000",
  17150=>"110100000",
  17151=>"000011000",
  17152=>"111100000",
  17153=>"001101111",
  17154=>"010110110",
  17155=>"000100111",
  17156=>"001110010",
  17157=>"100001100",
  17158=>"010001101",
  17159=>"111100010",
  17160=>"101011011",
  17161=>"111111111",
  17162=>"001001100",
  17163=>"011000100",
  17164=>"010010011",
  17165=>"011101111",
  17166=>"101101000",
  17167=>"100110011",
  17168=>"001000001",
  17169=>"010000010",
  17170=>"100110011",
  17171=>"001000110",
  17172=>"101000011",
  17173=>"011100001",
  17174=>"000011110",
  17175=>"011100000",
  17176=>"111011111",
  17177=>"010101000",
  17178=>"101001010",
  17179=>"010111011",
  17180=>"010010010",
  17181=>"111111110",
  17182=>"001001110",
  17183=>"100001110",
  17184=>"110001001",
  17185=>"011000001",
  17186=>"001011000",
  17187=>"010111100",
  17188=>"000000110",
  17189=>"011100110",
  17190=>"011100110",
  17191=>"100110011",
  17192=>"010111111",
  17193=>"110010100",
  17194=>"010000000",
  17195=>"100101010",
  17196=>"101101000",
  17197=>"001001010",
  17198=>"010000100",
  17199=>"110001001",
  17200=>"110011010",
  17201=>"001001111",
  17202=>"110101111",
  17203=>"010001010",
  17204=>"010011100",
  17205=>"011010001",
  17206=>"000001010",
  17207=>"001101011",
  17208=>"111101111",
  17209=>"000000101",
  17210=>"011011001",
  17211=>"101101010",
  17212=>"011101100",
  17213=>"110011111",
  17214=>"111111100",
  17215=>"111111111",
  17216=>"110101001",
  17217=>"110000101",
  17218=>"100111111",
  17219=>"111000010",
  17220=>"010010011",
  17221=>"001001001",
  17222=>"011100010",
  17223=>"100010110",
  17224=>"001101111",
  17225=>"001001000",
  17226=>"010111010",
  17227=>"101110111",
  17228=>"000010001",
  17229=>"001001100",
  17230=>"001010011",
  17231=>"011111011",
  17232=>"011011000",
  17233=>"000000111",
  17234=>"100011000",
  17235=>"010110000",
  17236=>"000000001",
  17237=>"111010100",
  17238=>"111011010",
  17239=>"101101001",
  17240=>"111001110",
  17241=>"111100100",
  17242=>"001000010",
  17243=>"010000011",
  17244=>"111101001",
  17245=>"001100100",
  17246=>"100010111",
  17247=>"111111001",
  17248=>"100110111",
  17249=>"100000101",
  17250=>"100110010",
  17251=>"100010010",
  17252=>"110001110",
  17253=>"000001000",
  17254=>"000010000",
  17255=>"111001000",
  17256=>"001010101",
  17257=>"101010000",
  17258=>"010010011",
  17259=>"101001011",
  17260=>"000010110",
  17261=>"000001110",
  17262=>"010110110",
  17263=>"111000010",
  17264=>"100110001",
  17265=>"011110100",
  17266=>"000110000",
  17267=>"001100100",
  17268=>"000000101",
  17269=>"110010010",
  17270=>"010111000",
  17271=>"010011110",
  17272=>"100001101",
  17273=>"000100010",
  17274=>"101100010",
  17275=>"101110110",
  17276=>"110101011",
  17277=>"001110011",
  17278=>"010010001",
  17279=>"001111101",
  17280=>"001011101",
  17281=>"111001110",
  17282=>"110100110",
  17283=>"010000000",
  17284=>"101110001",
  17285=>"110110000",
  17286=>"110110111",
  17287=>"111111111",
  17288=>"111001100",
  17289=>"101000101",
  17290=>"011111001",
  17291=>"010111000",
  17292=>"001111100",
  17293=>"100101110",
  17294=>"011101010",
  17295=>"101001001",
  17296=>"010000010",
  17297=>"110110010",
  17298=>"010100111",
  17299=>"000001011",
  17300=>"001010000",
  17301=>"101000000",
  17302=>"011001100",
  17303=>"010101110",
  17304=>"101100101",
  17305=>"000010010",
  17306=>"111010001",
  17307=>"110011001",
  17308=>"000100111",
  17309=>"011110011",
  17310=>"001011100",
  17311=>"001000011",
  17312=>"011011100",
  17313=>"001000011",
  17314=>"101000000",
  17315=>"010011000",
  17316=>"001001010",
  17317=>"000000011",
  17318=>"011010100",
  17319=>"001101110",
  17320=>"000100001",
  17321=>"000101100",
  17322=>"011100011",
  17323=>"001000001",
  17324=>"110011110",
  17325=>"000110110",
  17326=>"111010101",
  17327=>"010001001",
  17328=>"100111000",
  17329=>"010100000",
  17330=>"001000001",
  17331=>"001100000",
  17332=>"101111010",
  17333=>"101111010",
  17334=>"100000000",
  17335=>"111101100",
  17336=>"110101100",
  17337=>"110101011",
  17338=>"110100101",
  17339=>"001110011",
  17340=>"111000110",
  17341=>"100110010",
  17342=>"111010100",
  17343=>"010100000",
  17344=>"111011111",
  17345=>"000101000",
  17346=>"001000010",
  17347=>"101000100",
  17348=>"010101001",
  17349=>"100110000",
  17350=>"111001111",
  17351=>"001001000",
  17352=>"000010111",
  17353=>"101010110",
  17354=>"101011010",
  17355=>"010010101",
  17356=>"100001001",
  17357=>"000100001",
  17358=>"011110111",
  17359=>"000100111",
  17360=>"011110010",
  17361=>"101000001",
  17362=>"011010010",
  17363=>"101110111",
  17364=>"111011101",
  17365=>"000010010",
  17366=>"010110000",
  17367=>"000111111",
  17368=>"101001111",
  17369=>"111110100",
  17370=>"011101110",
  17371=>"000001001",
  17372=>"110001001",
  17373=>"101110011",
  17374=>"101001101",
  17375=>"110111110",
  17376=>"111101011",
  17377=>"001000110",
  17378=>"101001111",
  17379=>"000101011",
  17380=>"111001001",
  17381=>"000111001",
  17382=>"010101100",
  17383=>"001011100",
  17384=>"011000110",
  17385=>"111110011",
  17386=>"000000100",
  17387=>"001100111",
  17388=>"110100011",
  17389=>"101100101",
  17390=>"011111001",
  17391=>"111001100",
  17392=>"100110000",
  17393=>"000100111",
  17394=>"110011000",
  17395=>"010101101",
  17396=>"000110110",
  17397=>"001001001",
  17398=>"010010101",
  17399=>"111000001",
  17400=>"111101111",
  17401=>"011110000",
  17402=>"101011011",
  17403=>"101011100",
  17404=>"000110111",
  17405=>"000110001",
  17406=>"100101101",
  17407=>"001111011",
  17408=>"100010100",
  17409=>"100000011",
  17410=>"010101111",
  17411=>"100011100",
  17412=>"010011100",
  17413=>"000000101",
  17414=>"001110001",
  17415=>"110101000",
  17416=>"001000001",
  17417=>"100111110",
  17418=>"110100100",
  17419=>"110010111",
  17420=>"010110010",
  17421=>"101110111",
  17422=>"100100010",
  17423=>"110110101",
  17424=>"000011101",
  17425=>"000111110",
  17426=>"001110100",
  17427=>"110101011",
  17428=>"111000001",
  17429=>"111101110",
  17430=>"011001101",
  17431=>"100000001",
  17432=>"000011111",
  17433=>"111010101",
  17434=>"000010111",
  17435=>"011001001",
  17436=>"100100001",
  17437=>"110100101",
  17438=>"001000001",
  17439=>"010101001",
  17440=>"011011000",
  17441=>"001000100",
  17442=>"011010111",
  17443=>"001010010",
  17444=>"110000011",
  17445=>"010011001",
  17446=>"010101100",
  17447=>"000000111",
  17448=>"010111000",
  17449=>"011111111",
  17450=>"111110101",
  17451=>"110010010",
  17452=>"010100110",
  17453=>"011001001",
  17454=>"001101010",
  17455=>"000000110",
  17456=>"100011010",
  17457=>"101011100",
  17458=>"001000110",
  17459=>"110000011",
  17460=>"011101000",
  17461=>"000101000",
  17462=>"100101100",
  17463=>"010101010",
  17464=>"011001111",
  17465=>"000011001",
  17466=>"000101101",
  17467=>"101001111",
  17468=>"000001110",
  17469=>"000000001",
  17470=>"000011100",
  17471=>"011000111",
  17472=>"000010011",
  17473=>"101000101",
  17474=>"000111000",
  17475=>"010111011",
  17476=>"010000010",
  17477=>"001011001",
  17478=>"011101100",
  17479=>"000111001",
  17480=>"101011111",
  17481=>"101000001",
  17482=>"011101101",
  17483=>"101000001",
  17484=>"100001000",
  17485=>"101111011",
  17486=>"011100111",
  17487=>"110010001",
  17488=>"100001000",
  17489=>"000011010",
  17490=>"001001010",
  17491=>"011110101",
  17492=>"101010111",
  17493=>"010001011",
  17494=>"111000111",
  17495=>"101000001",
  17496=>"011101011",
  17497=>"110111011",
  17498=>"001000001",
  17499=>"000010100",
  17500=>"011111100",
  17501=>"110000010",
  17502=>"101110111",
  17503=>"000001001",
  17504=>"000100111",
  17505=>"101010111",
  17506=>"011101010",
  17507=>"001000110",
  17508=>"001101101",
  17509=>"110001110",
  17510=>"110000111",
  17511=>"111110110",
  17512=>"000010100",
  17513=>"010110010",
  17514=>"111101010",
  17515=>"111110001",
  17516=>"000110111",
  17517=>"000011010",
  17518=>"100111100",
  17519=>"100110110",
  17520=>"001101011",
  17521=>"010010001",
  17522=>"100001111",
  17523=>"110111110",
  17524=>"010000101",
  17525=>"101110100",
  17526=>"110111111",
  17527=>"011101111",
  17528=>"101000011",
  17529=>"110100111",
  17530=>"101110001",
  17531=>"100111001",
  17532=>"010001101",
  17533=>"110011001",
  17534=>"011011001",
  17535=>"100010000",
  17536=>"001101010",
  17537=>"111000000",
  17538=>"000101000",
  17539=>"000111111",
  17540=>"110110000",
  17541=>"101110100",
  17542=>"000101001",
  17543=>"010010111",
  17544=>"111000111",
  17545=>"111110011",
  17546=>"010011001",
  17547=>"000100101",
  17548=>"110011011",
  17549=>"000000100",
  17550=>"110011001",
  17551=>"110001111",
  17552=>"010000111",
  17553=>"100111110",
  17554=>"001010011",
  17555=>"011011000",
  17556=>"000101100",
  17557=>"110000111",
  17558=>"011000000",
  17559=>"110110000",
  17560=>"001100101",
  17561=>"100110001",
  17562=>"100111000",
  17563=>"001100010",
  17564=>"111000011",
  17565=>"101111011",
  17566=>"110110101",
  17567=>"000001100",
  17568=>"110100000",
  17569=>"001100100",
  17570=>"001000110",
  17571=>"111111001",
  17572=>"111111111",
  17573=>"000111000",
  17574=>"101111111",
  17575=>"110000000",
  17576=>"001100110",
  17577=>"110100000",
  17578=>"100101111",
  17579=>"101101010",
  17580=>"011011100",
  17581=>"010111111",
  17582=>"101110110",
  17583=>"000001001",
  17584=>"010010101",
  17585=>"010000000",
  17586=>"011101111",
  17587=>"100001101",
  17588=>"100111100",
  17589=>"000010000",
  17590=>"100111101",
  17591=>"100111101",
  17592=>"101000111",
  17593=>"110110110",
  17594=>"011001001",
  17595=>"000110110",
  17596=>"111100111",
  17597=>"011101100",
  17598=>"110000110",
  17599=>"110001010",
  17600=>"110111011",
  17601=>"100001011",
  17602=>"101001001",
  17603=>"000010000",
  17604=>"001010010",
  17605=>"000010001",
  17606=>"100110010",
  17607=>"100101000",
  17608=>"011111101",
  17609=>"001110101",
  17610=>"011100111",
  17611=>"101111111",
  17612=>"100101011",
  17613=>"110100000",
  17614=>"010100100",
  17615=>"011100101",
  17616=>"011100001",
  17617=>"001011111",
  17618=>"011001010",
  17619=>"000111000",
  17620=>"110111100",
  17621=>"000000110",
  17622=>"100111000",
  17623=>"000001111",
  17624=>"010000101",
  17625=>"001010111",
  17626=>"010111111",
  17627=>"001011001",
  17628=>"101100011",
  17629=>"100000110",
  17630=>"010011001",
  17631=>"010100101",
  17632=>"101000110",
  17633=>"110101011",
  17634=>"000101010",
  17635=>"010000110",
  17636=>"001000110",
  17637=>"100100101",
  17638=>"000110100",
  17639=>"000100011",
  17640=>"010101000",
  17641=>"101000101",
  17642=>"000000000",
  17643=>"001110011",
  17644=>"010010001",
  17645=>"010000011",
  17646=>"001111001",
  17647=>"110110101",
  17648=>"001111100",
  17649=>"001110001",
  17650=>"000100111",
  17651=>"010011011",
  17652=>"001000101",
  17653=>"000000101",
  17654=>"111100110",
  17655=>"111010011",
  17656=>"011011110",
  17657=>"000110000",
  17658=>"001100011",
  17659=>"010111000",
  17660=>"110111111",
  17661=>"010000001",
  17662=>"000111001",
  17663=>"101001001",
  17664=>"001101101",
  17665=>"000110111",
  17666=>"110111011",
  17667=>"010110000",
  17668=>"110111111",
  17669=>"010000111",
  17670=>"101100111",
  17671=>"101010110",
  17672=>"101001001",
  17673=>"000111101",
  17674=>"101001001",
  17675=>"110101101",
  17676=>"010011110",
  17677=>"011101010",
  17678=>"010000100",
  17679=>"001000000",
  17680=>"100001100",
  17681=>"111111101",
  17682=>"001011000",
  17683=>"101001001",
  17684=>"111100100",
  17685=>"101000010",
  17686=>"111011111",
  17687=>"110110111",
  17688=>"001001011",
  17689=>"010110010",
  17690=>"111101100",
  17691=>"100101010",
  17692=>"011001100",
  17693=>"001010011",
  17694=>"100000000",
  17695=>"100010110",
  17696=>"000111001",
  17697=>"001111110",
  17698=>"000101101",
  17699=>"000110110",
  17700=>"010010110",
  17701=>"110010000",
  17702=>"101101111",
  17703=>"000011001",
  17704=>"000011011",
  17705=>"100100010",
  17706=>"011110111",
  17707=>"111101011",
  17708=>"001111110",
  17709=>"001010001",
  17710=>"001000001",
  17711=>"000111100",
  17712=>"000001000",
  17713=>"011001101",
  17714=>"101001101",
  17715=>"011110011",
  17716=>"010101100",
  17717=>"010111100",
  17718=>"010110111",
  17719=>"001011001",
  17720=>"110100101",
  17721=>"010011111",
  17722=>"000001100",
  17723=>"011101100",
  17724=>"110111111",
  17725=>"111001101",
  17726=>"000100111",
  17727=>"011111101",
  17728=>"101111000",
  17729=>"011001010",
  17730=>"010101010",
  17731=>"011011111",
  17732=>"111110000",
  17733=>"000010010",
  17734=>"001100000",
  17735=>"001100000",
  17736=>"110001110",
  17737=>"101110000",
  17738=>"001000100",
  17739=>"010011000",
  17740=>"101100101",
  17741=>"001011000",
  17742=>"101111011",
  17743=>"001000000",
  17744=>"011110000",
  17745=>"011100101",
  17746=>"000101111",
  17747=>"011111111",
  17748=>"101001111",
  17749=>"101100101",
  17750=>"010111101",
  17751=>"010111111",
  17752=>"111101010",
  17753=>"111010011",
  17754=>"110110110",
  17755=>"111001111",
  17756=>"111011111",
  17757=>"110100101",
  17758=>"001010011",
  17759=>"111011000",
  17760=>"110111101",
  17761=>"001101100",
  17762=>"100000110",
  17763=>"000101110",
  17764=>"001001100",
  17765=>"101000101",
  17766=>"100100000",
  17767=>"110001101",
  17768=>"110001111",
  17769=>"001110111",
  17770=>"011110011",
  17771=>"111111010",
  17772=>"000001110",
  17773=>"010100101",
  17774=>"001011100",
  17775=>"101110010",
  17776=>"111000101",
  17777=>"011001000",
  17778=>"111000110",
  17779=>"010101001",
  17780=>"111101000",
  17781=>"011111111",
  17782=>"110100111",
  17783=>"111101001",
  17784=>"000000000",
  17785=>"100000010",
  17786=>"011101110",
  17787=>"001011110",
  17788=>"110101101",
  17789=>"101000101",
  17790=>"000111111",
  17791=>"010000111",
  17792=>"001001100",
  17793=>"001011110",
  17794=>"110000100",
  17795=>"001100011",
  17796=>"010111000",
  17797=>"000110000",
  17798=>"001101110",
  17799=>"110111010",
  17800=>"101001101",
  17801=>"101110100",
  17802=>"110010000",
  17803=>"001000010",
  17804=>"110100000",
  17805=>"101111110",
  17806=>"011110011",
  17807=>"100001110",
  17808=>"101011010",
  17809=>"110110000",
  17810=>"101011011",
  17811=>"000001011",
  17812=>"110011011",
  17813=>"001111110",
  17814=>"000011001",
  17815=>"001110000",
  17816=>"101101001",
  17817=>"101001001",
  17818=>"111111111",
  17819=>"011011000",
  17820=>"011101000",
  17821=>"010000100",
  17822=>"100001110",
  17823=>"111011011",
  17824=>"000011010",
  17825=>"110110101",
  17826=>"100010000",
  17827=>"111010001",
  17828=>"011010110",
  17829=>"000000000",
  17830=>"110111011",
  17831=>"100101011",
  17832=>"000010111",
  17833=>"100011000",
  17834=>"010010011",
  17835=>"101010001",
  17836=>"111110110",
  17837=>"000000110",
  17838=>"001111101",
  17839=>"110111001",
  17840=>"001000110",
  17841=>"011010100",
  17842=>"111110100",
  17843=>"010001001",
  17844=>"001100000",
  17845=>"100000111",
  17846=>"000010110",
  17847=>"011111110",
  17848=>"010010111",
  17849=>"110001100",
  17850=>"001000100",
  17851=>"011011100",
  17852=>"011110000",
  17853=>"101001001",
  17854=>"000011011",
  17855=>"110010011",
  17856=>"111010000",
  17857=>"101111101",
  17858=>"101100000",
  17859=>"011111101",
  17860=>"101110111",
  17861=>"010000000",
  17862=>"111100100",
  17863=>"110000100",
  17864=>"011100000",
  17865=>"011001011",
  17866=>"000110111",
  17867=>"010011111",
  17868=>"010001110",
  17869=>"111010100",
  17870=>"000001000",
  17871=>"100111111",
  17872=>"111111111",
  17873=>"110000001",
  17874=>"111011001",
  17875=>"010100011",
  17876=>"101101100",
  17877=>"001101100",
  17878=>"111010101",
  17879=>"111110101",
  17880=>"001010001",
  17881=>"101111000",
  17882=>"111101000",
  17883=>"111001000",
  17884=>"110000000",
  17885=>"110100111",
  17886=>"001000001",
  17887=>"110101110",
  17888=>"110000110",
  17889=>"100011001",
  17890=>"000101000",
  17891=>"001001100",
  17892=>"011010101",
  17893=>"011111110",
  17894=>"101110010",
  17895=>"011100000",
  17896=>"111011111",
  17897=>"100011000",
  17898=>"000001000",
  17899=>"000101000",
  17900=>"100101100",
  17901=>"110110100",
  17902=>"101110000",
  17903=>"001001100",
  17904=>"111000001",
  17905=>"010110000",
  17906=>"111110001",
  17907=>"001011110",
  17908=>"110100110",
  17909=>"101011101",
  17910=>"111111010",
  17911=>"010011111",
  17912=>"001000001",
  17913=>"100000111",
  17914=>"001100101",
  17915=>"100100111",
  17916=>"111110011",
  17917=>"000010110",
  17918=>"001111011",
  17919=>"000110100",
  17920=>"000111110",
  17921=>"000000000",
  17922=>"011001101",
  17923=>"111000011",
  17924=>"010011000",
  17925=>"101000001",
  17926=>"010110110",
  17927=>"100101010",
  17928=>"001100000",
  17929=>"111011000",
  17930=>"100000011",
  17931=>"010111001",
  17932=>"010111111",
  17933=>"000110110",
  17934=>"100000100",
  17935=>"001111011",
  17936=>"000111100",
  17937=>"110011010",
  17938=>"100100100",
  17939=>"011110011",
  17940=>"101000011",
  17941=>"011000001",
  17942=>"000000000",
  17943=>"011110111",
  17944=>"100101110",
  17945=>"101100001",
  17946=>"001000101",
  17947=>"011101100",
  17948=>"011110110",
  17949=>"110111000",
  17950=>"101001011",
  17951=>"101011010",
  17952=>"000001110",
  17953=>"111101010",
  17954=>"011110100",
  17955=>"001110011",
  17956=>"111101001",
  17957=>"011010010",
  17958=>"100100100",
  17959=>"000101010",
  17960=>"101100011",
  17961=>"101001010",
  17962=>"110011001",
  17963=>"011011000",
  17964=>"010011111",
  17965=>"101110100",
  17966=>"000000011",
  17967=>"010100101",
  17968=>"001001111",
  17969=>"011000111",
  17970=>"110100011",
  17971=>"010010000",
  17972=>"110110110",
  17973=>"110111001",
  17974=>"000011001",
  17975=>"001100010",
  17976=>"010001011",
  17977=>"101000010",
  17978=>"101111011",
  17979=>"111100011",
  17980=>"011011010",
  17981=>"000100011",
  17982=>"110100001",
  17983=>"000100011",
  17984=>"010010000",
  17985=>"100101010",
  17986=>"010000101",
  17987=>"111111010",
  17988=>"100000010",
  17989=>"010001110",
  17990=>"000011000",
  17991=>"110101111",
  17992=>"010010000",
  17993=>"011101101",
  17994=>"100111000",
  17995=>"100000110",
  17996=>"101010000",
  17997=>"011001001",
  17998=>"010000010",
  17999=>"110110011",
  18000=>"101001100",
  18001=>"111100100",
  18002=>"000111110",
  18003=>"100010001",
  18004=>"000010010",
  18005=>"001000000",
  18006=>"000110100",
  18007=>"100110100",
  18008=>"101010111",
  18009=>"000100100",
  18010=>"011111111",
  18011=>"000001000",
  18012=>"000001100",
  18013=>"111000000",
  18014=>"000101011",
  18015=>"001111000",
  18016=>"010010111",
  18017=>"000010111",
  18018=>"001110101",
  18019=>"101010010",
  18020=>"111010011",
  18021=>"100110011",
  18022=>"110001100",
  18023=>"010000011",
  18024=>"001110000",
  18025=>"001000100",
  18026=>"011100001",
  18027=>"000010110",
  18028=>"011110111",
  18029=>"101011111",
  18030=>"010001101",
  18031=>"010100111",
  18032=>"110110010",
  18033=>"110101001",
  18034=>"111001011",
  18035=>"001000011",
  18036=>"000000010",
  18037=>"001010101",
  18038=>"110011101",
  18039=>"001100010",
  18040=>"100100000",
  18041=>"000101011",
  18042=>"111110100",
  18043=>"111001000",
  18044=>"111100000",
  18045=>"101101000",
  18046=>"011011010",
  18047=>"011000110",
  18048=>"010011011",
  18049=>"110001101",
  18050=>"110010100",
  18051=>"110010100",
  18052=>"000001000",
  18053=>"000110110",
  18054=>"100000010",
  18055=>"110101001",
  18056=>"011011011",
  18057=>"100000011",
  18058=>"101100011",
  18059=>"111100100",
  18060=>"101000101",
  18061=>"011001100",
  18062=>"001111101",
  18063=>"010001011",
  18064=>"100111010",
  18065=>"010000010",
  18066=>"001111001",
  18067=>"101101111",
  18068=>"000001011",
  18069=>"101100101",
  18070=>"001010100",
  18071=>"100000011",
  18072=>"000100101",
  18073=>"111101101",
  18074=>"111011010",
  18075=>"000001100",
  18076=>"110010100",
  18077=>"000001000",
  18078=>"011001100",
  18079=>"110110101",
  18080=>"011010111",
  18081=>"110000011",
  18082=>"000100110",
  18083=>"100100011",
  18084=>"110100100",
  18085=>"010101011",
  18086=>"110111000",
  18087=>"000101001",
  18088=>"110010101",
  18089=>"001100000",
  18090=>"000001101",
  18091=>"110001110",
  18092=>"001110000",
  18093=>"111100011",
  18094=>"010001011",
  18095=>"010111101",
  18096=>"110100000",
  18097=>"010011111",
  18098=>"001000001",
  18099=>"000100011",
  18100=>"011000010",
  18101=>"001011101",
  18102=>"010000101",
  18103=>"101001011",
  18104=>"010111011",
  18105=>"001100110",
  18106=>"011100011",
  18107=>"011101010",
  18108=>"100001100",
  18109=>"011111000",
  18110=>"010001100",
  18111=>"100010001",
  18112=>"101000001",
  18113=>"101001111",
  18114=>"001100001",
  18115=>"100000011",
  18116=>"111001010",
  18117=>"101110100",
  18118=>"111111110",
  18119=>"001110101",
  18120=>"011111100",
  18121=>"000110011",
  18122=>"011110011",
  18123=>"100011100",
  18124=>"101101011",
  18125=>"100010100",
  18126=>"011000011",
  18127=>"110000101",
  18128=>"011100000",
  18129=>"001000001",
  18130=>"010010011",
  18131=>"101110010",
  18132=>"000100010",
  18133=>"000100011",
  18134=>"001000010",
  18135=>"101111100",
  18136=>"000000001",
  18137=>"000011100",
  18138=>"001011100",
  18139=>"101001010",
  18140=>"110001101",
  18141=>"101101111",
  18142=>"000110110",
  18143=>"100000011",
  18144=>"001010000",
  18145=>"110101101",
  18146=>"100010111",
  18147=>"001111111",
  18148=>"110110001",
  18149=>"001111001",
  18150=>"110010000",
  18151=>"000111011",
  18152=>"000100100",
  18153=>"100111101",
  18154=>"100100000",
  18155=>"000111010",
  18156=>"000100111",
  18157=>"110101100",
  18158=>"000101101",
  18159=>"000010001",
  18160=>"100111100",
  18161=>"100100011",
  18162=>"001110101",
  18163=>"010000110",
  18164=>"011001100",
  18165=>"001110100",
  18166=>"100010010",
  18167=>"100101010",
  18168=>"110111100",
  18169=>"001101011",
  18170=>"010110101",
  18171=>"111100100",
  18172=>"101100110",
  18173=>"011101010",
  18174=>"101000100",
  18175=>"001010010",
  18176=>"110100100",
  18177=>"001011011",
  18178=>"011100110",
  18179=>"100010111",
  18180=>"001011001",
  18181=>"000100110",
  18182=>"100000010",
  18183=>"101100111",
  18184=>"010110011",
  18185=>"101100101",
  18186=>"010001000",
  18187=>"111001101",
  18188=>"110001111",
  18189=>"010101111",
  18190=>"011110001",
  18191=>"011111001",
  18192=>"001101001",
  18193=>"100010101",
  18194=>"010011111",
  18195=>"001001101",
  18196=>"011001111",
  18197=>"110101101",
  18198=>"100001010",
  18199=>"011110101",
  18200=>"010000110",
  18201=>"100000010",
  18202=>"101001101",
  18203=>"111010111",
  18204=>"110101111",
  18205=>"011011010",
  18206=>"110000000",
  18207=>"010011000",
  18208=>"100110000",
  18209=>"000000111",
  18210=>"110010001",
  18211=>"001100001",
  18212=>"111110110",
  18213=>"010011111",
  18214=>"101111010",
  18215=>"011000110",
  18216=>"110001100",
  18217=>"110111111",
  18218=>"101111111",
  18219=>"001000011",
  18220=>"001111100",
  18221=>"000100010",
  18222=>"000111100",
  18223=>"011111111",
  18224=>"111111010",
  18225=>"101111010",
  18226=>"011111010",
  18227=>"111100100",
  18228=>"101101111",
  18229=>"001100000",
  18230=>"111011011",
  18231=>"101110000",
  18232=>"010110011",
  18233=>"011010011",
  18234=>"101001000",
  18235=>"111110100",
  18236=>"010100110",
  18237=>"110000000",
  18238=>"111000000",
  18239=>"000000000",
  18240=>"011100100",
  18241=>"010010100",
  18242=>"001001110",
  18243=>"011001001",
  18244=>"100000111",
  18245=>"110010101",
  18246=>"101011011",
  18247=>"000100000",
  18248=>"100111101",
  18249=>"010110110",
  18250=>"000000001",
  18251=>"110100001",
  18252=>"011101000",
  18253=>"010110000",
  18254=>"101010011",
  18255=>"000000000",
  18256=>"000100101",
  18257=>"101000100",
  18258=>"110000110",
  18259=>"111011100",
  18260=>"111111101",
  18261=>"010011110",
  18262=>"011111000",
  18263=>"111011100",
  18264=>"000000000",
  18265=>"110101011",
  18266=>"101110001",
  18267=>"100010101",
  18268=>"110001011",
  18269=>"111011111",
  18270=>"011010010",
  18271=>"000000000",
  18272=>"111001010",
  18273=>"000100101",
  18274=>"110011110",
  18275=>"100011100",
  18276=>"111010101",
  18277=>"110010100",
  18278=>"101001101",
  18279=>"100111100",
  18280=>"111001000",
  18281=>"100100010",
  18282=>"000011001",
  18283=>"111111010",
  18284=>"111000101",
  18285=>"110110011",
  18286=>"100010001",
  18287=>"100101010",
  18288=>"100001000",
  18289=>"100000010",
  18290=>"010001001",
  18291=>"101001000",
  18292=>"110001001",
  18293=>"011010110",
  18294=>"001000100",
  18295=>"101100101",
  18296=>"001100000",
  18297=>"101100010",
  18298=>"100101011",
  18299=>"111010011",
  18300=>"100100111",
  18301=>"110100000",
  18302=>"100001011",
  18303=>"100011001",
  18304=>"010100110",
  18305=>"001110101",
  18306=>"111110011",
  18307=>"101010001",
  18308=>"001111000",
  18309=>"101001000",
  18310=>"100111110",
  18311=>"001110000",
  18312=>"011110111",
  18313=>"000101010",
  18314=>"000011000",
  18315=>"011110001",
  18316=>"111101110",
  18317=>"001100110",
  18318=>"010000110",
  18319=>"010010100",
  18320=>"100100111",
  18321=>"000011111",
  18322=>"011011111",
  18323=>"111111100",
  18324=>"001100011",
  18325=>"001010110",
  18326=>"000111000",
  18327=>"010010111",
  18328=>"010011011",
  18329=>"000110000",
  18330=>"110000101",
  18331=>"101100010",
  18332=>"110001001",
  18333=>"110100010",
  18334=>"001001110",
  18335=>"010011000",
  18336=>"111000101",
  18337=>"101001101",
  18338=>"101001010",
  18339=>"000000000",
  18340=>"100111000",
  18341=>"101111100",
  18342=>"001001110",
  18343=>"001010011",
  18344=>"010110010",
  18345=>"110000111",
  18346=>"010011001",
  18347=>"010010100",
  18348=>"110100011",
  18349=>"101000110",
  18350=>"011100010",
  18351=>"001000000",
  18352=>"100110010",
  18353=>"001111110",
  18354=>"111110000",
  18355=>"100111110",
  18356=>"010001000",
  18357=>"111000100",
  18358=>"011001101",
  18359=>"001100101",
  18360=>"001101100",
  18361=>"111000110",
  18362=>"100010100",
  18363=>"001110101",
  18364=>"010010111",
  18365=>"011001101",
  18366=>"000100111",
  18367=>"100001110",
  18368=>"100111001",
  18369=>"011101101",
  18370=>"011010001",
  18371=>"110011001",
  18372=>"001111001",
  18373=>"101111110",
  18374=>"110011110",
  18375=>"100001110",
  18376=>"110101100",
  18377=>"010001010",
  18378=>"000000100",
  18379=>"001111000",
  18380=>"011101101",
  18381=>"011110100",
  18382=>"010101011",
  18383=>"001001011",
  18384=>"100110011",
  18385=>"010010000",
  18386=>"110100010",
  18387=>"010101010",
  18388=>"010010000",
  18389=>"000000111",
  18390=>"100101100",
  18391=>"001111011",
  18392=>"001010111",
  18393=>"010100101",
  18394=>"111000001",
  18395=>"101001010",
  18396=>"010111101",
  18397=>"111101100",
  18398=>"110001100",
  18399=>"001011010",
  18400=>"011110111",
  18401=>"100101001",
  18402=>"100110100",
  18403=>"010010010",
  18404=>"111110100",
  18405=>"010001101",
  18406=>"101101000",
  18407=>"110101000",
  18408=>"101010011",
  18409=>"110100111",
  18410=>"010100001",
  18411=>"010010000",
  18412=>"101000010",
  18413=>"011111110",
  18414=>"010000101",
  18415=>"110110110",
  18416=>"000000000",
  18417=>"010010100",
  18418=>"111110110",
  18419=>"000010101",
  18420=>"001101010",
  18421=>"100001000",
  18422=>"010111100",
  18423=>"010101010",
  18424=>"000001001",
  18425=>"001011111",
  18426=>"001110100",
  18427=>"010111110",
  18428=>"000010101",
  18429=>"111000100",
  18430=>"001110000",
  18431=>"000000101",
  18432=>"101111001",
  18433=>"010101001",
  18434=>"101101011",
  18435=>"000011010",
  18436=>"110010001",
  18437=>"001110011",
  18438=>"010000010",
  18439=>"111111011",
  18440=>"100010000",
  18441=>"110100101",
  18442=>"010111100",
  18443=>"001010100",
  18444=>"101001111",
  18445=>"110001100",
  18446=>"000010010",
  18447=>"100001110",
  18448=>"101111101",
  18449=>"000110011",
  18450=>"001001000",
  18451=>"010000010",
  18452=>"111111110",
  18453=>"110100011",
  18454=>"001000010",
  18455=>"110111101",
  18456=>"000000010",
  18457=>"010001010",
  18458=>"101010001",
  18459=>"000011001",
  18460=>"001100000",
  18461=>"010010111",
  18462=>"001001010",
  18463=>"010111101",
  18464=>"011101101",
  18465=>"101101011",
  18466=>"111011010",
  18467=>"000000000",
  18468=>"101111010",
  18469=>"010010010",
  18470=>"000101000",
  18471=>"110010010",
  18472=>"000000011",
  18473=>"101101111",
  18474=>"000100100",
  18475=>"011101110",
  18476=>"110000111",
  18477=>"111101110",
  18478=>"111000101",
  18479=>"100000010",
  18480=>"100000111",
  18481=>"100100000",
  18482=>"011100000",
  18483=>"001110101",
  18484=>"010111111",
  18485=>"000001000",
  18486=>"001100101",
  18487=>"100000111",
  18488=>"000010111",
  18489=>"101111101",
  18490=>"110110111",
  18491=>"100001010",
  18492=>"101101000",
  18493=>"010110111",
  18494=>"010100000",
  18495=>"000011011",
  18496=>"110101001",
  18497=>"011001000",
  18498=>"100000000",
  18499=>"000001011",
  18500=>"101001010",
  18501=>"000011111",
  18502=>"010111110",
  18503=>"000000111",
  18504=>"110101100",
  18505=>"000001000",
  18506=>"110001011",
  18507=>"100100010",
  18508=>"101011000",
  18509=>"110000101",
  18510=>"010010000",
  18511=>"011110010",
  18512=>"001000100",
  18513=>"100011010",
  18514=>"010011111",
  18515=>"001111001",
  18516=>"010010100",
  18517=>"001110111",
  18518=>"111100001",
  18519=>"001011010",
  18520=>"011001000",
  18521=>"110010000",
  18522=>"011101001",
  18523=>"011111101",
  18524=>"001011101",
  18525=>"100000100",
  18526=>"100011001",
  18527=>"001100111",
  18528=>"110101111",
  18529=>"100101001",
  18530=>"100111110",
  18531=>"110111100",
  18532=>"011111010",
  18533=>"010111101",
  18534=>"010111110",
  18535=>"000010000",
  18536=>"111010010",
  18537=>"010110101",
  18538=>"011111100",
  18539=>"011010111",
  18540=>"010010100",
  18541=>"010100010",
  18542=>"000101000",
  18543=>"000000111",
  18544=>"001001101",
  18545=>"000011100",
  18546=>"001010000",
  18547=>"001000011",
  18548=>"111100001",
  18549=>"111001111",
  18550=>"110000001",
  18551=>"101000110",
  18552=>"011111101",
  18553=>"011010000",
  18554=>"010101111",
  18555=>"111011000",
  18556=>"110010110",
  18557=>"001000100",
  18558=>"010111011",
  18559=>"111010110",
  18560=>"010100110",
  18561=>"011101010",
  18562=>"010110000",
  18563=>"011101001",
  18564=>"010011001",
  18565=>"111110101",
  18566=>"111001100",
  18567=>"000000001",
  18568=>"010000111",
  18569=>"110100111",
  18570=>"011101100",
  18571=>"010100000",
  18572=>"011001010",
  18573=>"100111000",
  18574=>"001111101",
  18575=>"111100101",
  18576=>"000001111",
  18577=>"011100111",
  18578=>"000101101",
  18579=>"110001111",
  18580=>"100000000",
  18581=>"111010010",
  18582=>"000100111",
  18583=>"010010001",
  18584=>"000010000",
  18585=>"111010011",
  18586=>"101111110",
  18587=>"000111000",
  18588=>"001100100",
  18589=>"011010111",
  18590=>"001100100",
  18591=>"001000100",
  18592=>"011001001",
  18593=>"000001001",
  18594=>"011111111",
  18595=>"010110001",
  18596=>"001011010",
  18597=>"111110101",
  18598=>"010110010",
  18599=>"101011011",
  18600=>"000100011",
  18601=>"010011011",
  18602=>"010100001",
  18603=>"000011001",
  18604=>"011011011",
  18605=>"010010001",
  18606=>"111110011",
  18607=>"010100110",
  18608=>"000100101",
  18609=>"100110111",
  18610=>"000000001",
  18611=>"100010000",
  18612=>"101111111",
  18613=>"001010011",
  18614=>"100001100",
  18615=>"111111000",
  18616=>"000100110",
  18617=>"100010100",
  18618=>"011110100",
  18619=>"000011110",
  18620=>"011001011",
  18621=>"110011111",
  18622=>"000011101",
  18623=>"011000011",
  18624=>"001111111",
  18625=>"111101100",
  18626=>"100010011",
  18627=>"000000111",
  18628=>"111101001",
  18629=>"010000111",
  18630=>"011101110",
  18631=>"110011000",
  18632=>"010110100",
  18633=>"010111010",
  18634=>"000111101",
  18635=>"111001110",
  18636=>"110001011",
  18637=>"010111111",
  18638=>"111001001",
  18639=>"001101111",
  18640=>"101100001",
  18641=>"111010101",
  18642=>"101011000",
  18643=>"100110001",
  18644=>"010001101",
  18645=>"101010000",
  18646=>"101001111",
  18647=>"100001001",
  18648=>"000010101",
  18649=>"000001111",
  18650=>"101001100",
  18651=>"111001101",
  18652=>"101100100",
  18653=>"101010000",
  18654=>"001001100",
  18655=>"110011100",
  18656=>"101111111",
  18657=>"000100101",
  18658=>"101101010",
  18659=>"000011110",
  18660=>"101001100",
  18661=>"100111001",
  18662=>"110010100",
  18663=>"110011100",
  18664=>"100010101",
  18665=>"010010110",
  18666=>"000000001",
  18667=>"000000101",
  18668=>"111101001",
  18669=>"001100101",
  18670=>"101110101",
  18671=>"011111111",
  18672=>"110000110",
  18673=>"111000000",
  18674=>"000101000",
  18675=>"011100011",
  18676=>"011110001",
  18677=>"101111000",
  18678=>"010010011",
  18679=>"101000001",
  18680=>"011000100",
  18681=>"111000111",
  18682=>"000011100",
  18683=>"100001100",
  18684=>"111000101",
  18685=>"100100100",
  18686=>"110110001",
  18687=>"100011010",
  18688=>"001101010",
  18689=>"111001000",
  18690=>"101101111",
  18691=>"110110101",
  18692=>"100110000",
  18693=>"100001010",
  18694=>"011110110",
  18695=>"001011101",
  18696=>"110011111",
  18697=>"101101010",
  18698=>"111101111",
  18699=>"100100001",
  18700=>"011111101",
  18701=>"001011000",
  18702=>"001110000",
  18703=>"010110111",
  18704=>"011010000",
  18705=>"111110011",
  18706=>"111110010",
  18707=>"011001001",
  18708=>"101110110",
  18709=>"101110001",
  18710=>"010000010",
  18711=>"100011111",
  18712=>"010011100",
  18713=>"010110001",
  18714=>"011101111",
  18715=>"101010011",
  18716=>"010111011",
  18717=>"010001110",
  18718=>"010100000",
  18719=>"111101111",
  18720=>"000001010",
  18721=>"111011011",
  18722=>"011101010",
  18723=>"000100101",
  18724=>"110101101",
  18725=>"100011100",
  18726=>"001100111",
  18727=>"111011001",
  18728=>"010011010",
  18729=>"000010001",
  18730=>"111100101",
  18731=>"110101100",
  18732=>"110111110",
  18733=>"011000100",
  18734=>"001111101",
  18735=>"110000011",
  18736=>"011100001",
  18737=>"000100000",
  18738=>"001110011",
  18739=>"001100011",
  18740=>"101110110",
  18741=>"010000110",
  18742=>"000010001",
  18743=>"101111010",
  18744=>"100100100",
  18745=>"000110111",
  18746=>"101111001",
  18747=>"110001110",
  18748=>"011111110",
  18749=>"110011100",
  18750=>"101100010",
  18751=>"100011101",
  18752=>"100011001",
  18753=>"111011110",
  18754=>"111010010",
  18755=>"011101100",
  18756=>"110010000",
  18757=>"001000000",
  18758=>"010011100",
  18759=>"000000001",
  18760=>"111101011",
  18761=>"011000000",
  18762=>"111110000",
  18763=>"010001110",
  18764=>"011001011",
  18765=>"110111100",
  18766=>"111110001",
  18767=>"110010000",
  18768=>"101110110",
  18769=>"000101110",
  18770=>"100000101",
  18771=>"111110100",
  18772=>"010010010",
  18773=>"000000100",
  18774=>"001111111",
  18775=>"000000010",
  18776=>"100010101",
  18777=>"010110110",
  18778=>"010011000",
  18779=>"110001011",
  18780=>"101010100",
  18781=>"010101101",
  18782=>"001100101",
  18783=>"110000010",
  18784=>"100010000",
  18785=>"010101110",
  18786=>"000001010",
  18787=>"111100001",
  18788=>"011111001",
  18789=>"101110110",
  18790=>"100110101",
  18791=>"101010110",
  18792=>"000010100",
  18793=>"010010111",
  18794=>"001000011",
  18795=>"111001000",
  18796=>"000100010",
  18797=>"111111000",
  18798=>"000001011",
  18799=>"100001110",
  18800=>"100111100",
  18801=>"001110000",
  18802=>"001000101",
  18803=>"110011110",
  18804=>"101011101",
  18805=>"010101010",
  18806=>"111100010",
  18807=>"111000101",
  18808=>"001001101",
  18809=>"110111100",
  18810=>"100000101",
  18811=>"010101100",
  18812=>"100111011",
  18813=>"101100000",
  18814=>"110110010",
  18815=>"101011001",
  18816=>"100000000",
  18817=>"011000101",
  18818=>"010001011",
  18819=>"111110000",
  18820=>"001100111",
  18821=>"111100011",
  18822=>"110010001",
  18823=>"001110011",
  18824=>"000100110",
  18825=>"001011100",
  18826=>"010010011",
  18827=>"010110011",
  18828=>"100100100",
  18829=>"011000011",
  18830=>"001010110",
  18831=>"000000101",
  18832=>"010110000",
  18833=>"110010000",
  18834=>"111010101",
  18835=>"000101001",
  18836=>"000001101",
  18837=>"010101011",
  18838=>"000011000",
  18839=>"000001011",
  18840=>"010001001",
  18841=>"000011000",
  18842=>"111110010",
  18843=>"000101110",
  18844=>"110000100",
  18845=>"010101000",
  18846=>"000100011",
  18847=>"010000010",
  18848=>"101111101",
  18849=>"111101110",
  18850=>"010010100",
  18851=>"111000011",
  18852=>"011010000",
  18853=>"100101111",
  18854=>"100010011",
  18855=>"001011111",
  18856=>"100011000",
  18857=>"011111101",
  18858=>"111110011",
  18859=>"110000110",
  18860=>"111110111",
  18861=>"000010110",
  18862=>"110101110",
  18863=>"010101111",
  18864=>"110111111",
  18865=>"000101111",
  18866=>"111011010",
  18867=>"101000001",
  18868=>"110001110",
  18869=>"011000101",
  18870=>"001100111",
  18871=>"101010001",
  18872=>"011001100",
  18873=>"000010101",
  18874=>"000110110",
  18875=>"011001000",
  18876=>"100101011",
  18877=>"000010010",
  18878=>"101001010",
  18879=>"110111111",
  18880=>"000101000",
  18881=>"001000011",
  18882=>"000000111",
  18883=>"010110010",
  18884=>"100100011",
  18885=>"001101111",
  18886=>"001100000",
  18887=>"110110111",
  18888=>"011101011",
  18889=>"111101000",
  18890=>"000101110",
  18891=>"110010000",
  18892=>"110100010",
  18893=>"010001110",
  18894=>"101101101",
  18895=>"111000101",
  18896=>"101011011",
  18897=>"011010010",
  18898=>"110010011",
  18899=>"001000011",
  18900=>"111111111",
  18901=>"111111000",
  18902=>"001010101",
  18903=>"100110010",
  18904=>"001011111",
  18905=>"010001100",
  18906=>"010010010",
  18907=>"110110111",
  18908=>"110110010",
  18909=>"110000100",
  18910=>"010101101",
  18911=>"100110101",
  18912=>"011000100",
  18913=>"000101100",
  18914=>"000011111",
  18915=>"110111011",
  18916=>"011000110",
  18917=>"011101001",
  18918=>"000101010",
  18919=>"110001000",
  18920=>"001111001",
  18921=>"010110100",
  18922=>"110101011",
  18923=>"110000111",
  18924=>"111010001",
  18925=>"110111101",
  18926=>"101000101",
  18927=>"001111111",
  18928=>"011000111",
  18929=>"000010000",
  18930=>"010101010",
  18931=>"000101001",
  18932=>"111001101",
  18933=>"010010010",
  18934=>"101001001",
  18935=>"111011101",
  18936=>"100001000",
  18937=>"110100111",
  18938=>"101111111",
  18939=>"000000000",
  18940=>"110001000",
  18941=>"000100011",
  18942=>"000100100",
  18943=>"000000011",
  18944=>"010101110",
  18945=>"001101110",
  18946=>"111000101",
  18947=>"110110000",
  18948=>"000000101",
  18949=>"111111011",
  18950=>"000101110",
  18951=>"101101001",
  18952=>"101011000",
  18953=>"101111100",
  18954=>"010110010",
  18955=>"111110111",
  18956=>"010111000",
  18957=>"010000011",
  18958=>"011111101",
  18959=>"101101110",
  18960=>"100100000",
  18961=>"001000010",
  18962=>"111001000",
  18963=>"100000001",
  18964=>"011001011",
  18965=>"111110011",
  18966=>"001001001",
  18967=>"101010001",
  18968=>"000000111",
  18969=>"000101011",
  18970=>"001010101",
  18971=>"000010001",
  18972=>"111001111",
  18973=>"111101001",
  18974=>"011001001",
  18975=>"101011101",
  18976=>"111110110",
  18977=>"100100111",
  18978=>"110000001",
  18979=>"100110011",
  18980=>"111101101",
  18981=>"111000000",
  18982=>"100100101",
  18983=>"101010101",
  18984=>"100001010",
  18985=>"100111010",
  18986=>"100101010",
  18987=>"011001010",
  18988=>"100100000",
  18989=>"010101111",
  18990=>"001100010",
  18991=>"011010100",
  18992=>"010110100",
  18993=>"011001010",
  18994=>"111110011",
  18995=>"011111010",
  18996=>"011011011",
  18997=>"000011101",
  18998=>"011110010",
  18999=>"010111111",
  19000=>"111101101",
  19001=>"000101001",
  19002=>"111010011",
  19003=>"110000000",
  19004=>"111110011",
  19005=>"100010010",
  19006=>"101011110",
  19007=>"000001000",
  19008=>"000100010",
  19009=>"110010010",
  19010=>"010011100",
  19011=>"110000010",
  19012=>"110110111",
  19013=>"011000010",
  19014=>"011000111",
  19015=>"010000000",
  19016=>"100101001",
  19017=>"111001011",
  19018=>"000000011",
  19019=>"000110000",
  19020=>"111110110",
  19021=>"101101110",
  19022=>"111100101",
  19023=>"001000100",
  19024=>"011000000",
  19025=>"110100101",
  19026=>"101100011",
  19027=>"011110011",
  19028=>"111011011",
  19029=>"101000001",
  19030=>"101000000",
  19031=>"010111111",
  19032=>"100100001",
  19033=>"111101011",
  19034=>"111001011",
  19035=>"001100100",
  19036=>"101100001",
  19037=>"010111011",
  19038=>"111110111",
  19039=>"111000111",
  19040=>"011100010",
  19041=>"000101101",
  19042=>"001011000",
  19043=>"101001101",
  19044=>"101101100",
  19045=>"100000110",
  19046=>"101111010",
  19047=>"111101011",
  19048=>"110000111",
  19049=>"000000010",
  19050=>"000001110",
  19051=>"110111000",
  19052=>"011110000",
  19053=>"110011001",
  19054=>"001011001",
  19055=>"011000010",
  19056=>"101001101",
  19057=>"011011111",
  19058=>"100010000",
  19059=>"100010000",
  19060=>"111011000",
  19061=>"010110100",
  19062=>"010000100",
  19063=>"011111111",
  19064=>"111011001",
  19065=>"101000001",
  19066=>"110011000",
  19067=>"110011101",
  19068=>"110010110",
  19069=>"010100001",
  19070=>"010100100",
  19071=>"000011011",
  19072=>"010000101",
  19073=>"100110100",
  19074=>"011011010",
  19075=>"101000010",
  19076=>"011010001",
  19077=>"001101000",
  19078=>"011101001",
  19079=>"000000001",
  19080=>"000111110",
  19081=>"111011011",
  19082=>"110011110",
  19083=>"010000100",
  19084=>"000110000",
  19085=>"101110100",
  19086=>"111001000",
  19087=>"100110110",
  19088=>"010010000",
  19089=>"110110110",
  19090=>"001011100",
  19091=>"100000011",
  19092=>"100110011",
  19093=>"000111001",
  19094=>"000000001",
  19095=>"111001101",
  19096=>"110011101",
  19097=>"010110001",
  19098=>"011001100",
  19099=>"110111001",
  19100=>"010111010",
  19101=>"110001001",
  19102=>"000000110",
  19103=>"111010010",
  19104=>"001111100",
  19105=>"011111111",
  19106=>"101011000",
  19107=>"010110110",
  19108=>"011001010",
  19109=>"111100111",
  19110=>"100011100",
  19111=>"110000110",
  19112=>"111010111",
  19113=>"101111100",
  19114=>"111100100",
  19115=>"000000011",
  19116=>"000010100",
  19117=>"000111000",
  19118=>"001111000",
  19119=>"000111011",
  19120=>"001110100",
  19121=>"111000000",
  19122=>"111101101",
  19123=>"101110101",
  19124=>"100110100",
  19125=>"001000010",
  19126=>"010001100",
  19127=>"101101011",
  19128=>"000000101",
  19129=>"110000100",
  19130=>"101000010",
  19131=>"001100100",
  19132=>"000100000",
  19133=>"011010110",
  19134=>"110010011",
  19135=>"010011111",
  19136=>"100011110",
  19137=>"101001101",
  19138=>"111110000",
  19139=>"010110011",
  19140=>"011011010",
  19141=>"011110000",
  19142=>"110010001",
  19143=>"011010101",
  19144=>"111111000",
  19145=>"110110111",
  19146=>"010101111",
  19147=>"111110011",
  19148=>"001100001",
  19149=>"000000001",
  19150=>"011110110",
  19151=>"011101001",
  19152=>"111111000",
  19153=>"100101001",
  19154=>"100100111",
  19155=>"001000110",
  19156=>"100110001",
  19157=>"000110011",
  19158=>"000011001",
  19159=>"111011011",
  19160=>"101111011",
  19161=>"000101111",
  19162=>"111001000",
  19163=>"000111010",
  19164=>"011000111",
  19165=>"111000110",
  19166=>"101001001",
  19167=>"101011111",
  19168=>"001100011",
  19169=>"010001010",
  19170=>"010111010",
  19171=>"111010011",
  19172=>"101011000",
  19173=>"011011001",
  19174=>"010110100",
  19175=>"101111011",
  19176=>"101011100",
  19177=>"111001110",
  19178=>"100101111",
  19179=>"001000001",
  19180=>"100011010",
  19181=>"101000010",
  19182=>"010000000",
  19183=>"110111010",
  19184=>"100111111",
  19185=>"101110111",
  19186=>"001011100",
  19187=>"110010011",
  19188=>"001010111",
  19189=>"011111111",
  19190=>"010010110",
  19191=>"001001101",
  19192=>"010101010",
  19193=>"110110111",
  19194=>"001010010",
  19195=>"111011001",
  19196=>"011110101",
  19197=>"001011101",
  19198=>"011100100",
  19199=>"010011010",
  19200=>"000001100",
  19201=>"100100000",
  19202=>"111000010",
  19203=>"110000000",
  19204=>"000100110",
  19205=>"110000000",
  19206=>"100101000",
  19207=>"001011001",
  19208=>"011110010",
  19209=>"111110111",
  19210=>"100110011",
  19211=>"011101011",
  19212=>"000101001",
  19213=>"000111010",
  19214=>"110001010",
  19215=>"011110001",
  19216=>"101000100",
  19217=>"100111111",
  19218=>"100111100",
  19219=>"111001010",
  19220=>"110100001",
  19221=>"001100001",
  19222=>"110011000",
  19223=>"110100111",
  19224=>"101001111",
  19225=>"111010000",
  19226=>"111101110",
  19227=>"110111111",
  19228=>"010100000",
  19229=>"100001011",
  19230=>"111111011",
  19231=>"100011111",
  19232=>"111011100",
  19233=>"010101000",
  19234=>"100000100",
  19235=>"111111101",
  19236=>"000000100",
  19237=>"011110010",
  19238=>"111111011",
  19239=>"101000010",
  19240=>"100110110",
  19241=>"100000010",
  19242=>"011011001",
  19243=>"110111010",
  19244=>"110101101",
  19245=>"110110010",
  19246=>"010110000",
  19247=>"001111111",
  19248=>"001100010",
  19249=>"000100001",
  19250=>"001011001",
  19251=>"010001001",
  19252=>"000111000",
  19253=>"000111000",
  19254=>"000000100",
  19255=>"101011111",
  19256=>"110111011",
  19257=>"110011111",
  19258=>"101011100",
  19259=>"110011001",
  19260=>"000101111",
  19261=>"000111100",
  19262=>"111111110",
  19263=>"101000011",
  19264=>"010010111",
  19265=>"010111010",
  19266=>"010100001",
  19267=>"111101101",
  19268=>"101100101",
  19269=>"110000010",
  19270=>"111001001",
  19271=>"111011111",
  19272=>"110101001",
  19273=>"011101111",
  19274=>"101011111",
  19275=>"000101010",
  19276=>"100100001",
  19277=>"100101010",
  19278=>"101000000",
  19279=>"001000100",
  19280=>"101101001",
  19281=>"101101111",
  19282=>"100101100",
  19283=>"111010001",
  19284=>"000000000",
  19285=>"101111110",
  19286=>"110010110",
  19287=>"001001010",
  19288=>"010100010",
  19289=>"111111000",
  19290=>"011110110",
  19291=>"111001000",
  19292=>"010001011",
  19293=>"111001111",
  19294=>"110011001",
  19295=>"111100110",
  19296=>"101111010",
  19297=>"010111100",
  19298=>"000010111",
  19299=>"110110100",
  19300=>"110110101",
  19301=>"000110100",
  19302=>"111110101",
  19303=>"100000000",
  19304=>"000011011",
  19305=>"100101010",
  19306=>"101101101",
  19307=>"000111110",
  19308=>"100111101",
  19309=>"011111110",
  19310=>"000011000",
  19311=>"101010101",
  19312=>"010000110",
  19313=>"111110101",
  19314=>"000100111",
  19315=>"000001110",
  19316=>"110001001",
  19317=>"000011011",
  19318=>"011011000",
  19319=>"001001110",
  19320=>"010001001",
  19321=>"100110011",
  19322=>"100110101",
  19323=>"111111101",
  19324=>"111111111",
  19325=>"011100111",
  19326=>"001110110",
  19327=>"001101000",
  19328=>"001100010",
  19329=>"111010010",
  19330=>"101111100",
  19331=>"000100000",
  19332=>"110001011",
  19333=>"011000001",
  19334=>"100101010",
  19335=>"101111100",
  19336=>"101111111",
  19337=>"011011111",
  19338=>"111000110",
  19339=>"010110011",
  19340=>"001011010",
  19341=>"010101100",
  19342=>"110110011",
  19343=>"001111001",
  19344=>"111111111",
  19345=>"011111110",
  19346=>"110100010",
  19347=>"101000011",
  19348=>"111101111",
  19349=>"000010001",
  19350=>"011000100",
  19351=>"001011000",
  19352=>"011100111",
  19353=>"110100010",
  19354=>"101101101",
  19355=>"110110110",
  19356=>"001001110",
  19357=>"001110011",
  19358=>"111110110",
  19359=>"101001010",
  19360=>"110001110",
  19361=>"000110000",
  19362=>"100010001",
  19363=>"101011001",
  19364=>"100000100",
  19365=>"000001011",
  19366=>"111001101",
  19367=>"011101100",
  19368=>"110111110",
  19369=>"000100100",
  19370=>"001011001",
  19371=>"000000101",
  19372=>"010011111",
  19373=>"111100101",
  19374=>"011111101",
  19375=>"011010000",
  19376=>"101101001",
  19377=>"111110110",
  19378=>"000110010",
  19379=>"010110111",
  19380=>"000111111",
  19381=>"001111001",
  19382=>"000000111",
  19383=>"111011001",
  19384=>"010010101",
  19385=>"001111111",
  19386=>"011000101",
  19387=>"111001000",
  19388=>"101011001",
  19389=>"100000001",
  19390=>"000000010",
  19391=>"101111011",
  19392=>"011110001",
  19393=>"111010000",
  19394=>"101100110",
  19395=>"011110001",
  19396=>"100110010",
  19397=>"000011001",
  19398=>"010010010",
  19399=>"000011100",
  19400=>"001001010",
  19401=>"101101001",
  19402=>"100110000",
  19403=>"101101010",
  19404=>"001010011",
  19405=>"000111110",
  19406=>"001000101",
  19407=>"000110000",
  19408=>"000010000",
  19409=>"110110000",
  19410=>"010011100",
  19411=>"011001000",
  19412=>"101011011",
  19413=>"000010100",
  19414=>"100010011",
  19415=>"101011000",
  19416=>"101000101",
  19417=>"110111000",
  19418=>"000000000",
  19419=>"110000011",
  19420=>"001011011",
  19421=>"110101011",
  19422=>"010110001",
  19423=>"000000001",
  19424=>"010000001",
  19425=>"101111000",
  19426=>"000011100",
  19427=>"111000100",
  19428=>"111011111",
  19429=>"000001110",
  19430=>"001111001",
  19431=>"111010011",
  19432=>"110101000",
  19433=>"011100101",
  19434=>"111100001",
  19435=>"001011000",
  19436=>"000110000",
  19437=>"001010001",
  19438=>"101000001",
  19439=>"011101111",
  19440=>"000100110",
  19441=>"111010001",
  19442=>"110110101",
  19443=>"100100001",
  19444=>"110111000",
  19445=>"110001101",
  19446=>"011111001",
  19447=>"000011010",
  19448=>"001110001",
  19449=>"010101111",
  19450=>"110110011",
  19451=>"010001100",
  19452=>"000000000",
  19453=>"110101110",
  19454=>"000111110",
  19455=>"010101010",
  19456=>"010111010",
  19457=>"111010011",
  19458=>"011010100",
  19459=>"110110110",
  19460=>"111111101",
  19461=>"000111000",
  19462=>"111000001",
  19463=>"101111010",
  19464=>"110011000",
  19465=>"010100010",
  19466=>"101101001",
  19467=>"101100010",
  19468=>"101111010",
  19469=>"001100111",
  19470=>"001001000",
  19471=>"001011110",
  19472=>"101100000",
  19473=>"010101001",
  19474=>"011101011",
  19475=>"101011000",
  19476=>"110100000",
  19477=>"110101111",
  19478=>"010010101",
  19479=>"110100010",
  19480=>"100001001",
  19481=>"010000100",
  19482=>"101010110",
  19483=>"001011111",
  19484=>"010100000",
  19485=>"011101111",
  19486=>"010110010",
  19487=>"100000100",
  19488=>"010001010",
  19489=>"101011100",
  19490=>"000010101",
  19491=>"100101011",
  19492=>"101010100",
  19493=>"001101100",
  19494=>"011010001",
  19495=>"100101101",
  19496=>"001011110",
  19497=>"000110111",
  19498=>"110100001",
  19499=>"110000010",
  19500=>"101001101",
  19501=>"100001111",
  19502=>"111111100",
  19503=>"001001100",
  19504=>"100000001",
  19505=>"000100111",
  19506=>"010010010",
  19507=>"111110000",
  19508=>"111011001",
  19509=>"111001010",
  19510=>"110011001",
  19511=>"001011110",
  19512=>"011001100",
  19513=>"100011010",
  19514=>"011011100",
  19515=>"101010011",
  19516=>"111001010",
  19517=>"010111011",
  19518=>"000100001",
  19519=>"011110011",
  19520=>"100000001",
  19521=>"111110001",
  19522=>"111011110",
  19523=>"011011100",
  19524=>"110101000",
  19525=>"001000011",
  19526=>"110100100",
  19527=>"110111001",
  19528=>"110100101",
  19529=>"100001110",
  19530=>"000000110",
  19531=>"011011111",
  19532=>"101010100",
  19533=>"000001111",
  19534=>"011011100",
  19535=>"001001100",
  19536=>"011011101",
  19537=>"011001000",
  19538=>"101100000",
  19539=>"011000100",
  19540=>"110110010",
  19541=>"011101101",
  19542=>"000110100",
  19543=>"111001010",
  19544=>"111000111",
  19545=>"000111011",
  19546=>"101000101",
  19547=>"111111011",
  19548=>"100110110",
  19549=>"001110110",
  19550=>"101000111",
  19551=>"010111001",
  19552=>"110101110",
  19553=>"000100011",
  19554=>"101100110",
  19555=>"101111011",
  19556=>"111010000",
  19557=>"101001110",
  19558=>"011101101",
  19559=>"000101011",
  19560=>"001100010",
  19561=>"010011001",
  19562=>"000111001",
  19563=>"110000111",
  19564=>"100110100",
  19565=>"000011100",
  19566=>"011110011",
  19567=>"111011100",
  19568=>"110001100",
  19569=>"001100001",
  19570=>"001011100",
  19571=>"101110110",
  19572=>"101111101",
  19573=>"001110101",
  19574=>"010000011",
  19575=>"011000000",
  19576=>"000100100",
  19577=>"011100110",
  19578=>"110101111",
  19579=>"010011111",
  19580=>"011011110",
  19581=>"011011011",
  19582=>"011010100",
  19583=>"011011000",
  19584=>"000000111",
  19585=>"001000110",
  19586=>"001010100",
  19587=>"000101000",
  19588=>"011001101",
  19589=>"000001001",
  19590=>"100010110",
  19591=>"111100011",
  19592=>"001111110",
  19593=>"001011111",
  19594=>"110100011",
  19595=>"001101100",
  19596=>"010100001",
  19597=>"011101011",
  19598=>"111100010",
  19599=>"001110010",
  19600=>"101100001",
  19601=>"010100110",
  19602=>"111010110",
  19603=>"111111000",
  19604=>"010111010",
  19605=>"000101111",
  19606=>"100110100",
  19607=>"011000111",
  19608=>"011101111",
  19609=>"000010011",
  19610=>"100110010",
  19611=>"101111110",
  19612=>"001010010",
  19613=>"001000100",
  19614=>"100001011",
  19615=>"000010110",
  19616=>"010100111",
  19617=>"110000110",
  19618=>"110101110",
  19619=>"000110110",
  19620=>"100101110",
  19621=>"100000110",
  19622=>"011110000",
  19623=>"001110101",
  19624=>"100001101",
  19625=>"001010001",
  19626=>"111111111",
  19627=>"001101101",
  19628=>"100000111",
  19629=>"110101011",
  19630=>"100000111",
  19631=>"111001100",
  19632=>"001011000",
  19633=>"111011010",
  19634=>"001100111",
  19635=>"110110000",
  19636=>"011011010",
  19637=>"010001001",
  19638=>"101011000",
  19639=>"010011001",
  19640=>"101011011",
  19641=>"010000001",
  19642=>"110111001",
  19643=>"001100010",
  19644=>"101111011",
  19645=>"010001001",
  19646=>"001110101",
  19647=>"011011011",
  19648=>"110100001",
  19649=>"100101100",
  19650=>"110110000",
  19651=>"011101001",
  19652=>"101000010",
  19653=>"101000000",
  19654=>"001001001",
  19655=>"110100100",
  19656=>"110000110",
  19657=>"100100011",
  19658=>"011010000",
  19659=>"010100101",
  19660=>"110010011",
  19661=>"010011110",
  19662=>"101100010",
  19663=>"011101011",
  19664=>"101111011",
  19665=>"101101111",
  19666=>"101100100",
  19667=>"100010001",
  19668=>"100101000",
  19669=>"011011100",
  19670=>"000100101",
  19671=>"100101001",
  19672=>"000111011",
  19673=>"000000111",
  19674=>"011110011",
  19675=>"011001010",
  19676=>"111100111",
  19677=>"000100001",
  19678=>"100000110",
  19679=>"111111101",
  19680=>"010010111",
  19681=>"001100110",
  19682=>"101001000",
  19683=>"000100111",
  19684=>"011101110",
  19685=>"011011110",
  19686=>"001010100",
  19687=>"100101001",
  19688=>"111010101",
  19689=>"111101011",
  19690=>"110000101",
  19691=>"001011111",
  19692=>"101111011",
  19693=>"001110101",
  19694=>"000100001",
  19695=>"110010100",
  19696=>"010010000",
  19697=>"101100111",
  19698=>"100110101",
  19699=>"001110100",
  19700=>"001111010",
  19701=>"011110011",
  19702=>"110010011",
  19703=>"001000000",
  19704=>"100010110",
  19705=>"001110001",
  19706=>"000011000",
  19707=>"100100011",
  19708=>"000000000",
  19709=>"000011110",
  19710=>"010111100",
  19711=>"000101111",
  19712=>"010111001",
  19713=>"110001110",
  19714=>"001011101",
  19715=>"000010000",
  19716=>"000100100",
  19717=>"101010110",
  19718=>"111110000",
  19719=>"111111000",
  19720=>"000011010",
  19721=>"100001011",
  19722=>"001110001",
  19723=>"010000011",
  19724=>"100011001",
  19725=>"101011010",
  19726=>"001000000",
  19727=>"001000101",
  19728=>"101110000",
  19729=>"100010111",
  19730=>"011001001",
  19731=>"101010000",
  19732=>"000010010",
  19733=>"011000101",
  19734=>"111101111",
  19735=>"110101001",
  19736=>"001111000",
  19737=>"110011011",
  19738=>"110101101",
  19739=>"100110010",
  19740=>"101100100",
  19741=>"011010100",
  19742=>"001011111",
  19743=>"111011001",
  19744=>"010011000",
  19745=>"010100010",
  19746=>"011110011",
  19747=>"100110111",
  19748=>"111100101",
  19749=>"100000101",
  19750=>"101110100",
  19751=>"011101110",
  19752=>"100100101",
  19753=>"101000111",
  19754=>"111001100",
  19755=>"111010001",
  19756=>"100110100",
  19757=>"111110111",
  19758=>"000000001",
  19759=>"111111100",
  19760=>"111001100",
  19761=>"111101110",
  19762=>"101011010",
  19763=>"000101000",
  19764=>"100011101",
  19765=>"010111001",
  19766=>"000010000",
  19767=>"011001111",
  19768=>"110101011",
  19769=>"100000010",
  19770=>"000000011",
  19771=>"011110110",
  19772=>"111010010",
  19773=>"000010101",
  19774=>"000000101",
  19775=>"101011100",
  19776=>"010110110",
  19777=>"100010101",
  19778=>"011111111",
  19779=>"010001111",
  19780=>"101001011",
  19781=>"101010000",
  19782=>"110100111",
  19783=>"100011101",
  19784=>"000111101",
  19785=>"001101001",
  19786=>"000110100",
  19787=>"000111111",
  19788=>"101000101",
  19789=>"001010101",
  19790=>"100010000",
  19791=>"001010011",
  19792=>"011111110",
  19793=>"111100010",
  19794=>"011011001",
  19795=>"001101000",
  19796=>"000101111",
  19797=>"110000110",
  19798=>"110000010",
  19799=>"101110000",
  19800=>"110011110",
  19801=>"111001010",
  19802=>"010100101",
  19803=>"101101110",
  19804=>"111010011",
  19805=>"111000010",
  19806=>"110001000",
  19807=>"101001101",
  19808=>"000000100",
  19809=>"110001010",
  19810=>"000111101",
  19811=>"000011111",
  19812=>"100110001",
  19813=>"100000000",
  19814=>"110110111",
  19815=>"001111010",
  19816=>"010111111",
  19817=>"000000111",
  19818=>"010111010",
  19819=>"100010101",
  19820=>"011111110",
  19821=>"101001100",
  19822=>"111100110",
  19823=>"101101110",
  19824=>"001011000",
  19825=>"110001111",
  19826=>"000001001",
  19827=>"111101111",
  19828=>"101100100",
  19829=>"110011101",
  19830=>"001001010",
  19831=>"100010000",
  19832=>"101010010",
  19833=>"010100111",
  19834=>"111110101",
  19835=>"100010100",
  19836=>"101010000",
  19837=>"011101110",
  19838=>"001001011",
  19839=>"101100100",
  19840=>"100000000",
  19841=>"011111010",
  19842=>"100111111",
  19843=>"000001111",
  19844=>"010111000",
  19845=>"000001010",
  19846=>"111110011",
  19847=>"100011001",
  19848=>"000100111",
  19849=>"011110000",
  19850=>"101010010",
  19851=>"000101111",
  19852=>"010101111",
  19853=>"101100111",
  19854=>"010000100",
  19855=>"010001100",
  19856=>"010000100",
  19857=>"000110010",
  19858=>"011010111",
  19859=>"001101110",
  19860=>"011110000",
  19861=>"000111010",
  19862=>"100010011",
  19863=>"101000011",
  19864=>"011100000",
  19865=>"000011000",
  19866=>"101001111",
  19867=>"111000011",
  19868=>"001100111",
  19869=>"100110011",
  19870=>"000001110",
  19871=>"110010001",
  19872=>"000100101",
  19873=>"111000100",
  19874=>"111101110",
  19875=>"101001100",
  19876=>"011011001",
  19877=>"010100001",
  19878=>"010011000",
  19879=>"111000110",
  19880=>"010010101",
  19881=>"111010110",
  19882=>"000001000",
  19883=>"111111001",
  19884=>"010011111",
  19885=>"010111000",
  19886=>"100011001",
  19887=>"001011001",
  19888=>"011100011",
  19889=>"101111000",
  19890=>"100000000",
  19891=>"111010110",
  19892=>"011101100",
  19893=>"111010100",
  19894=>"110100011",
  19895=>"010111010",
  19896=>"111000101",
  19897=>"011011110",
  19898=>"111101110",
  19899=>"111011111",
  19900=>"001101110",
  19901=>"110010000",
  19902=>"101111110",
  19903=>"001111110",
  19904=>"001001111",
  19905=>"100111110",
  19906=>"011110111",
  19907=>"100110101",
  19908=>"100001011",
  19909=>"010011101",
  19910=>"110111111",
  19911=>"101011111",
  19912=>"011101100",
  19913=>"101000010",
  19914=>"011101111",
  19915=>"101101111",
  19916=>"011110110",
  19917=>"100101001",
  19918=>"111111101",
  19919=>"001000101",
  19920=>"111010001",
  19921=>"110101010",
  19922=>"111100001",
  19923=>"101101111",
  19924=>"110110111",
  19925=>"101111011",
  19926=>"000111111",
  19927=>"000000100",
  19928=>"001011101",
  19929=>"110000101",
  19930=>"011010010",
  19931=>"100001111",
  19932=>"101110001",
  19933=>"110000000",
  19934=>"011111110",
  19935=>"011100001",
  19936=>"100101101",
  19937=>"000000011",
  19938=>"111111110",
  19939=>"000111001",
  19940=>"101100011",
  19941=>"010000001",
  19942=>"110111011",
  19943=>"101100111",
  19944=>"100101100",
  19945=>"100100000",
  19946=>"110110100",
  19947=>"010110101",
  19948=>"101100111",
  19949=>"011010011",
  19950=>"001111100",
  19951=>"001011011",
  19952=>"100000011",
  19953=>"010101110",
  19954=>"000100010",
  19955=>"100001100",
  19956=>"101110011",
  19957=>"100010001",
  19958=>"001010000",
  19959=>"101000010",
  19960=>"101001001",
  19961=>"101111001",
  19962=>"110010011",
  19963=>"110100000",
  19964=>"010101011",
  19965=>"000001111",
  19966=>"110000011",
  19967=>"100001110",
  19968=>"101010110",
  19969=>"101100000",
  19970=>"111011000",
  19971=>"011000010",
  19972=>"000100001",
  19973=>"101111100",
  19974=>"100110111",
  19975=>"100001100",
  19976=>"011100100",
  19977=>"000010111",
  19978=>"101101110",
  19979=>"000110001",
  19980=>"010000110",
  19981=>"001000111",
  19982=>"110101000",
  19983=>"111101011",
  19984=>"000011110",
  19985=>"110101101",
  19986=>"001100000",
  19987=>"101110010",
  19988=>"111111101",
  19989=>"111010111",
  19990=>"011010001",
  19991=>"000100011",
  19992=>"011010010",
  19993=>"110011001",
  19994=>"100011101",
  19995=>"111101100",
  19996=>"000011001",
  19997=>"001000001",
  19998=>"110011101",
  19999=>"011010001",
  20000=>"010011111",
  20001=>"001101001",
  20002=>"111000110",
  20003=>"010000000",
  20004=>"101100100",
  20005=>"000000100",
  20006=>"001101101",
  20007=>"000101000",
  20008=>"010001100",
  20009=>"110001011",
  20010=>"100101110",
  20011=>"110101101",
  20012=>"100100010",
  20013=>"011001001",
  20014=>"100110100",
  20015=>"101100100",
  20016=>"110011110",
  20017=>"101001001",
  20018=>"000010101",
  20019=>"001111110",
  20020=>"110100100",
  20021=>"010000000",
  20022=>"100010000",
  20023=>"010100101",
  20024=>"111001110",
  20025=>"000001000",
  20026=>"100010001",
  20027=>"001101111",
  20028=>"000101000",
  20029=>"111011111",
  20030=>"110101001",
  20031=>"010000010",
  20032=>"011111010",
  20033=>"011101011",
  20034=>"001101000",
  20035=>"110000011",
  20036=>"011110001",
  20037=>"111111111",
  20038=>"100100010",
  20039=>"001011010",
  20040=>"101000100",
  20041=>"010011111",
  20042=>"010111000",
  20043=>"100011111",
  20044=>"001001110",
  20045=>"111101011",
  20046=>"101101011",
  20047=>"000000010",
  20048=>"111011011",
  20049=>"111000101",
  20050=>"101010011",
  20051=>"010111111",
  20052=>"001110011",
  20053=>"011110111",
  20054=>"101011100",
  20055=>"010110110",
  20056=>"010000101",
  20057=>"011111110",
  20058=>"001011111",
  20059=>"010110101",
  20060=>"100000011",
  20061=>"101000110",
  20062=>"000111001",
  20063=>"001110010",
  20064=>"011011000",
  20065=>"111000101",
  20066=>"100001000",
  20067=>"001001011",
  20068=>"001001011",
  20069=>"000010101",
  20070=>"001010001",
  20071=>"000101010",
  20072=>"101101011",
  20073=>"101100110",
  20074=>"100001000",
  20075=>"110010111",
  20076=>"110001000",
  20077=>"101001100",
  20078=>"110111110",
  20079=>"001001000",
  20080=>"011101011",
  20081=>"001010111",
  20082=>"110011001",
  20083=>"100011100",
  20084=>"110111001",
  20085=>"000111101",
  20086=>"001101000",
  20087=>"101010010",
  20088=>"110100110",
  20089=>"110100110",
  20090=>"111011011",
  20091=>"100110000",
  20092=>"010001011",
  20093=>"111111100",
  20094=>"010000000",
  20095=>"100001001",
  20096=>"110110110",
  20097=>"100001010",
  20098=>"000000000",
  20099=>"001101010",
  20100=>"101111100",
  20101=>"111110101",
  20102=>"101010000",
  20103=>"010000010",
  20104=>"110000000",
  20105=>"010001000",
  20106=>"001000111",
  20107=>"001010001",
  20108=>"100000111",
  20109=>"000100100",
  20110=>"110000010",
  20111=>"010000111",
  20112=>"001011010",
  20113=>"010010000",
  20114=>"100111100",
  20115=>"110101110",
  20116=>"100101001",
  20117=>"011100111",
  20118=>"100011110",
  20119=>"111001010",
  20120=>"111100100",
  20121=>"100100101",
  20122=>"111100001",
  20123=>"010000101",
  20124=>"111010100",
  20125=>"100111110",
  20126=>"111110001",
  20127=>"111001010",
  20128=>"101101011",
  20129=>"101001111",
  20130=>"010110111",
  20131=>"110101011",
  20132=>"000001000",
  20133=>"101001100",
  20134=>"011101000",
  20135=>"110100100",
  20136=>"000000011",
  20137=>"111111110",
  20138=>"100110111",
  20139=>"001000110",
  20140=>"001010010",
  20141=>"111101001",
  20142=>"101001110",
  20143=>"001011011",
  20144=>"011110111",
  20145=>"010101011",
  20146=>"100101111",
  20147=>"100110100",
  20148=>"111011110",
  20149=>"001011111",
  20150=>"111111110",
  20151=>"110001111",
  20152=>"100110010",
  20153=>"000110011",
  20154=>"100001010",
  20155=>"111001110",
  20156=>"000101011",
  20157=>"010011010",
  20158=>"001101011",
  20159=>"001100011",
  20160=>"100000101",
  20161=>"111111000",
  20162=>"001010001",
  20163=>"001101001",
  20164=>"010000101",
  20165=>"001010011",
  20166=>"000000101",
  20167=>"000011111",
  20168=>"001100110",
  20169=>"010100010",
  20170=>"001011011",
  20171=>"100000101",
  20172=>"000000011",
  20173=>"010101010",
  20174=>"001000011",
  20175=>"101010010",
  20176=>"001001000",
  20177=>"011000111",
  20178=>"010111101",
  20179=>"101101111",
  20180=>"111111111",
  20181=>"111011010",
  20182=>"010110010",
  20183=>"011000001",
  20184=>"010100000",
  20185=>"010011010",
  20186=>"110101101",
  20187=>"010011100",
  20188=>"101110111",
  20189=>"000111111",
  20190=>"000110111",
  20191=>"111110001",
  20192=>"011001000",
  20193=>"110000100",
  20194=>"111001001",
  20195=>"100110000",
  20196=>"100010001",
  20197=>"111111100",
  20198=>"101101011",
  20199=>"111101010",
  20200=>"000010111",
  20201=>"000100011",
  20202=>"110001000",
  20203=>"110110001",
  20204=>"011000010",
  20205=>"101011000",
  20206=>"001001010",
  20207=>"101110010",
  20208=>"110110100",
  20209=>"001100010",
  20210=>"000110100",
  20211=>"100010011",
  20212=>"100110101",
  20213=>"011100101",
  20214=>"100000000",
  20215=>"101110111",
  20216=>"000010000",
  20217=>"000011101",
  20218=>"010010000",
  20219=>"101001110",
  20220=>"111110001",
  20221=>"100000110",
  20222=>"001110011",
  20223=>"100111010",
  20224=>"011001111",
  20225=>"110001010",
  20226=>"010111101",
  20227=>"110101110",
  20228=>"001111001",
  20229=>"111010010",
  20230=>"011110001",
  20231=>"111100101",
  20232=>"011110010",
  20233=>"001111000",
  20234=>"100000011",
  20235=>"011100110",
  20236=>"111001010",
  20237=>"101111001",
  20238=>"001100110",
  20239=>"011010111",
  20240=>"100011101",
  20241=>"101101000",
  20242=>"111000000",
  20243=>"101010100",
  20244=>"110011000",
  20245=>"110110100",
  20246=>"111101111",
  20247=>"111001010",
  20248=>"101100101",
  20249=>"001010101",
  20250=>"010011011",
  20251=>"010111010",
  20252=>"101010011",
  20253=>"100001100",
  20254=>"100010111",
  20255=>"111101001",
  20256=>"111010001",
  20257=>"011101011",
  20258=>"111100010",
  20259=>"001101111",
  20260=>"011001111",
  20261=>"001000100",
  20262=>"000101100",
  20263=>"110000000",
  20264=>"001010111",
  20265=>"101010111",
  20266=>"010000010",
  20267=>"111111111",
  20268=>"010111111",
  20269=>"111110111",
  20270=>"001101100",
  20271=>"010111010",
  20272=>"101111011",
  20273=>"101001001",
  20274=>"010001000",
  20275=>"101001011",
  20276=>"110101111",
  20277=>"110110100",
  20278=>"100101111",
  20279=>"110001101",
  20280=>"001110110",
  20281=>"100011011",
  20282=>"110000001",
  20283=>"001010100",
  20284=>"001000001",
  20285=>"011110010",
  20286=>"001000011",
  20287=>"000000011",
  20288=>"101001000",
  20289=>"001111010",
  20290=>"011000000",
  20291=>"110100011",
  20292=>"100111000",
  20293=>"010100110",
  20294=>"111010010",
  20295=>"010000111",
  20296=>"010110000",
  20297=>"010000001",
  20298=>"111001110",
  20299=>"100110010",
  20300=>"011110101",
  20301=>"100100001",
  20302=>"101001111",
  20303=>"110000110",
  20304=>"110000100",
  20305=>"010101011",
  20306=>"000101001",
  20307=>"111000000",
  20308=>"011010110",
  20309=>"101000000",
  20310=>"111001001",
  20311=>"010100101",
  20312=>"100011100",
  20313=>"011100000",
  20314=>"011101001",
  20315=>"010011111",
  20316=>"111010110",
  20317=>"000001001",
  20318=>"111111110",
  20319=>"101000101",
  20320=>"000100111",
  20321=>"110010001",
  20322=>"110111100",
  20323=>"100100001",
  20324=>"111000001",
  20325=>"110000001",
  20326=>"111000110",
  20327=>"010000110",
  20328=>"110000110",
  20329=>"111101110",
  20330=>"111000101",
  20331=>"111111000",
  20332=>"100101100",
  20333=>"011011100",
  20334=>"011101100",
  20335=>"111101000",
  20336=>"100110010",
  20337=>"110001110",
  20338=>"111100011",
  20339=>"010100101",
  20340=>"011010010",
  20341=>"011011101",
  20342=>"011111100",
  20343=>"101100000",
  20344=>"100000111",
  20345=>"001010001",
  20346=>"110000100",
  20347=>"001001111",
  20348=>"100011100",
  20349=>"000100000",
  20350=>"101101110",
  20351=>"001000101",
  20352=>"101100000",
  20353=>"000101001",
  20354=>"011010010",
  20355=>"010001000",
  20356=>"001000101",
  20357=>"001111001",
  20358=>"111111000",
  20359=>"001101010",
  20360=>"000001110",
  20361=>"011001001",
  20362=>"001111010",
  20363=>"010000101",
  20364=>"110000101",
  20365=>"110001000",
  20366=>"001100111",
  20367=>"111111000",
  20368=>"011000010",
  20369=>"001100111",
  20370=>"001001011",
  20371=>"010000011",
  20372=>"111111111",
  20373=>"101111111",
  20374=>"000100110",
  20375=>"101010010",
  20376=>"011111100",
  20377=>"010000000",
  20378=>"010011111",
  20379=>"111110011",
  20380=>"001111110",
  20381=>"001001110",
  20382=>"001011110",
  20383=>"011011100",
  20384=>"001110011",
  20385=>"011101000",
  20386=>"101110100",
  20387=>"110111110",
  20388=>"100101011",
  20389=>"000101000",
  20390=>"010011111",
  20391=>"000101111",
  20392=>"010101101",
  20393=>"010011100",
  20394=>"010000100",
  20395=>"010011110",
  20396=>"100111101",
  20397=>"111001101",
  20398=>"000110110",
  20399=>"111100100",
  20400=>"100100000",
  20401=>"011000101",
  20402=>"111110101",
  20403=>"100000111",
  20404=>"001011111",
  20405=>"001101011",
  20406=>"100000000",
  20407=>"110001110",
  20408=>"110111111",
  20409=>"001010000",
  20410=>"001001000",
  20411=>"101011100",
  20412=>"010000010",
  20413=>"010111001",
  20414=>"111111101",
  20415=>"011001110",
  20416=>"000000010",
  20417=>"000101011",
  20418=>"101011000",
  20419=>"110010011",
  20420=>"000101101",
  20421=>"111100111",
  20422=>"111111001",
  20423=>"000011011",
  20424=>"010011100",
  20425=>"000010101",
  20426=>"110001101",
  20427=>"110110111",
  20428=>"010000000",
  20429=>"101010101",
  20430=>"010010100",
  20431=>"111101001",
  20432=>"001111100",
  20433=>"000010010",
  20434=>"000111000",
  20435=>"011101001",
  20436=>"011111011",
  20437=>"100110101",
  20438=>"110111100",
  20439=>"000010001",
  20440=>"011100101",
  20441=>"111000101",
  20442=>"100111100",
  20443=>"011110101",
  20444=>"111101100",
  20445=>"011001000",
  20446=>"101001000",
  20447=>"010010011",
  20448=>"001011110",
  20449=>"110010110",
  20450=>"100010011",
  20451=>"100101001",
  20452=>"011000111",
  20453=>"111111111",
  20454=>"000111011",
  20455=>"001010011",
  20456=>"000001011",
  20457=>"110011110",
  20458=>"001000011",
  20459=>"110101011",
  20460=>"010000110",
  20461=>"001101110",
  20462=>"100011110",
  20463=>"010001110",
  20464=>"010001100",
  20465=>"111001011",
  20466=>"001100111",
  20467=>"001101100",
  20468=>"000001010",
  20469=>"011101000",
  20470=>"111001001",
  20471=>"110100110",
  20472=>"011101010",
  20473=>"000011100",
  20474=>"100010000",
  20475=>"100010010",
  20476=>"100000011",
  20477=>"010000011",
  20478=>"000100000",
  20479=>"011101101",
  20480=>"011010001",
  20481=>"011110010",
  20482=>"010001100",
  20483=>"011000000",
  20484=>"100001001",
  20485=>"001111011",
  20486=>"110001110",
  20487=>"010010100",
  20488=>"101011000",
  20489=>"100000000",
  20490=>"000100101",
  20491=>"101010100",
  20492=>"101111000",
  20493=>"011101111",
  20494=>"100000000",
  20495=>"110100101",
  20496=>"100100010",
  20497=>"100101110",
  20498=>"001010010",
  20499=>"101011110",
  20500=>"100001010",
  20501=>"111011101",
  20502=>"111011111",
  20503=>"101111011",
  20504=>"100100100",
  20505=>"010111000",
  20506=>"010100000",
  20507=>"100101001",
  20508=>"011111111",
  20509=>"111001010",
  20510=>"101100110",
  20511=>"000001101",
  20512=>"100000010",
  20513=>"100010100",
  20514=>"100010011",
  20515=>"010100111",
  20516=>"111011001",
  20517=>"010010010",
  20518=>"100101010",
  20519=>"001001101",
  20520=>"101010010",
  20521=>"000000000",
  20522=>"001011110",
  20523=>"110001110",
  20524=>"000111111",
  20525=>"100100101",
  20526=>"101110101",
  20527=>"001110101",
  20528=>"101101100",
  20529=>"011101011",
  20530=>"101011100",
  20531=>"101110001",
  20532=>"011001111",
  20533=>"100001100",
  20534=>"100110110",
  20535=>"111011001",
  20536=>"101110100",
  20537=>"110000000",
  20538=>"000011101",
  20539=>"000011110",
  20540=>"100100000",
  20541=>"111011010",
  20542=>"011100000",
  20543=>"011000100",
  20544=>"101010001",
  20545=>"101111101",
  20546=>"100011000",
  20547=>"010011111",
  20548=>"011110111",
  20549=>"000001000",
  20550=>"001010100",
  20551=>"110001011",
  20552=>"010110001",
  20553=>"001000001",
  20554=>"101111101",
  20555=>"101000110",
  20556=>"000101110",
  20557=>"011011101",
  20558=>"111101110",
  20559=>"010010101",
  20560=>"100100001",
  20561=>"001001000",
  20562=>"111010000",
  20563=>"101010010",
  20564=>"101100010",
  20565=>"000011011",
  20566=>"001100011",
  20567=>"010101110",
  20568=>"101000111",
  20569=>"011000110",
  20570=>"000101110",
  20571=>"010010111",
  20572=>"000010110",
  20573=>"110011011",
  20574=>"001100110",
  20575=>"001010011",
  20576=>"001111110",
  20577=>"100001100",
  20578=>"101110011",
  20579=>"011001111",
  20580=>"110100011",
  20581=>"101110000",
  20582=>"001011111",
  20583=>"111001001",
  20584=>"000011010",
  20585=>"001100110",
  20586=>"001000001",
  20587=>"101111101",
  20588=>"100111000",
  20589=>"101100100",
  20590=>"000001111",
  20591=>"111110001",
  20592=>"000101100",
  20593=>"110001101",
  20594=>"001010101",
  20595=>"000010011",
  20596=>"111011111",
  20597=>"000000110",
  20598=>"111110010",
  20599=>"001101000",
  20600=>"101101010",
  20601=>"100101111",
  20602=>"000011001",
  20603=>"110010001",
  20604=>"000100101",
  20605=>"010111001",
  20606=>"001101000",
  20607=>"011000001",
  20608=>"111010110",
  20609=>"001100100",
  20610=>"101010111",
  20611=>"001101111",
  20612=>"001011010",
  20613=>"010111110",
  20614=>"010010010",
  20615=>"101000100",
  20616=>"001111101",
  20617=>"111100001",
  20618=>"001110101",
  20619=>"111000101",
  20620=>"001011101",
  20621=>"111100111",
  20622=>"110110010",
  20623=>"011001100",
  20624=>"101001001",
  20625=>"011110001",
  20626=>"001110010",
  20627=>"111100100",
  20628=>"001010110",
  20629=>"011011101",
  20630=>"000001000",
  20631=>"011100000",
  20632=>"001111110",
  20633=>"011110000",
  20634=>"011010011",
  20635=>"000001010",
  20636=>"000101001",
  20637=>"111100010",
  20638=>"111100111",
  20639=>"100011000",
  20640=>"111101100",
  20641=>"100000011",
  20642=>"010000110",
  20643=>"111010000",
  20644=>"111111110",
  20645=>"001101110",
  20646=>"011101110",
  20647=>"010100000",
  20648=>"000000010",
  20649=>"111000111",
  20650=>"010011100",
  20651=>"010010111",
  20652=>"101100101",
  20653=>"110101111",
  20654=>"110101011",
  20655=>"110011101",
  20656=>"111011100",
  20657=>"101001001",
  20658=>"000010111",
  20659=>"000001101",
  20660=>"100110101",
  20661=>"001011111",
  20662=>"000011010",
  20663=>"010101101",
  20664=>"001000111",
  20665=>"110111111",
  20666=>"111110111",
  20667=>"000010001",
  20668=>"001100010",
  20669=>"111111011",
  20670=>"100001100",
  20671=>"111110001",
  20672=>"100101010",
  20673=>"001011110",
  20674=>"001000011",
  20675=>"100011101",
  20676=>"011100101",
  20677=>"111011000",
  20678=>"010110110",
  20679=>"010000110",
  20680=>"110111011",
  20681=>"010000011",
  20682=>"101110100",
  20683=>"000000001",
  20684=>"111111110",
  20685=>"100111001",
  20686=>"101010010",
  20687=>"100111000",
  20688=>"000000010",
  20689=>"001111101",
  20690=>"110000010",
  20691=>"111011011",
  20692=>"001000100",
  20693=>"101000000",
  20694=>"111101100",
  20695=>"110101010",
  20696=>"010101011",
  20697=>"111000101",
  20698=>"110000100",
  20699=>"001010101",
  20700=>"010100110",
  20701=>"010010011",
  20702=>"010101110",
  20703=>"011010011",
  20704=>"011110010",
  20705=>"000011010",
  20706=>"001000100",
  20707=>"010001001",
  20708=>"101110100",
  20709=>"111011110",
  20710=>"111101111",
  20711=>"101110111",
  20712=>"111110111",
  20713=>"001111010",
  20714=>"110010010",
  20715=>"001001100",
  20716=>"011010100",
  20717=>"111000010",
  20718=>"000011011",
  20719=>"010111011",
  20720=>"110111111",
  20721=>"010001111",
  20722=>"001000010",
  20723=>"010010001",
  20724=>"101100101",
  20725=>"100011101",
  20726=>"111100001",
  20727=>"000101111",
  20728=>"010100100",
  20729=>"111011101",
  20730=>"100111010",
  20731=>"001001011",
  20732=>"111000111",
  20733=>"000011010",
  20734=>"011000010",
  20735=>"101101001",
  20736=>"100110110",
  20737=>"101011010",
  20738=>"000011011",
  20739=>"111100111",
  20740=>"010000000",
  20741=>"010110111",
  20742=>"000110101",
  20743=>"111110101",
  20744=>"010001011",
  20745=>"111011111",
  20746=>"110110000",
  20747=>"110110101",
  20748=>"100001101",
  20749=>"001100111",
  20750=>"100101111",
  20751=>"000001101",
  20752=>"100010101",
  20753=>"000011011",
  20754=>"001010000",
  20755=>"111101010",
  20756=>"011000001",
  20757=>"110100000",
  20758=>"001001001",
  20759=>"101010011",
  20760=>"001001111",
  20761=>"111110001",
  20762=>"101101010",
  20763=>"110000000",
  20764=>"000110100",
  20765=>"010111011",
  20766=>"110000110",
  20767=>"011010111",
  20768=>"010011000",
  20769=>"011110001",
  20770=>"010110100",
  20771=>"100101001",
  20772=>"011110001",
  20773=>"111001110",
  20774=>"111011000",
  20775=>"010010111",
  20776=>"110100111",
  20777=>"000101001",
  20778=>"111100000",
  20779=>"001010111",
  20780=>"100101111",
  20781=>"110010010",
  20782=>"100100110",
  20783=>"001001010",
  20784=>"000000011",
  20785=>"111011000",
  20786=>"001100000",
  20787=>"110011011",
  20788=>"001010111",
  20789=>"010100011",
  20790=>"001101101",
  20791=>"000011111",
  20792=>"111011101",
  20793=>"001101101",
  20794=>"011000011",
  20795=>"011111000",
  20796=>"010001110",
  20797=>"110111111",
  20798=>"111111111",
  20799=>"110110010",
  20800=>"100111010",
  20801=>"111110101",
  20802=>"101100111",
  20803=>"101010010",
  20804=>"100011100",
  20805=>"111110100",
  20806=>"110110001",
  20807=>"001111101",
  20808=>"001001001",
  20809=>"001001000",
  20810=>"110101011",
  20811=>"001011100",
  20812=>"000111101",
  20813=>"000101001",
  20814=>"111010011",
  20815=>"000011010",
  20816=>"100111101",
  20817=>"100000100",
  20818=>"111110100",
  20819=>"000100000",
  20820=>"100101010",
  20821=>"011011011",
  20822=>"001110101",
  20823=>"011000101",
  20824=>"100100110",
  20825=>"011000100",
  20826=>"011100101",
  20827=>"101101010",
  20828=>"111001010",
  20829=>"110110110",
  20830=>"010111101",
  20831=>"101101101",
  20832=>"001011111",
  20833=>"100111010",
  20834=>"001111110",
  20835=>"010001010",
  20836=>"000010010",
  20837=>"001101001",
  20838=>"010000000",
  20839=>"010100000",
  20840=>"010010000",
  20841=>"100100010",
  20842=>"010100111",
  20843=>"110001000",
  20844=>"001101100",
  20845=>"101001101",
  20846=>"010111110",
  20847=>"100011101",
  20848=>"110100101",
  20849=>"001100111",
  20850=>"111111010",
  20851=>"111100101",
  20852=>"110010110",
  20853=>"000001010",
  20854=>"100111011",
  20855=>"100001011",
  20856=>"011110110",
  20857=>"110010001",
  20858=>"100111011",
  20859=>"010001110",
  20860=>"100001000",
  20861=>"010011100",
  20862=>"110011110",
  20863=>"000101101",
  20864=>"101110001",
  20865=>"100011000",
  20866=>"011000010",
  20867=>"000110010",
  20868=>"010010001",
  20869=>"011111011",
  20870=>"101101001",
  20871=>"111100110",
  20872=>"011001010",
  20873=>"100011111",
  20874=>"110111100",
  20875=>"001001111",
  20876=>"010101111",
  20877=>"010010100",
  20878=>"100101000",
  20879=>"011100011",
  20880=>"111101010",
  20881=>"000010010",
  20882=>"001001000",
  20883=>"001001001",
  20884=>"111111111",
  20885=>"000111110",
  20886=>"110101110",
  20887=>"110001100",
  20888=>"111000101",
  20889=>"001011010",
  20890=>"001011001",
  20891=>"001011010",
  20892=>"010101000",
  20893=>"011000010",
  20894=>"101101110",
  20895=>"110101110",
  20896=>"001001011",
  20897=>"111101101",
  20898=>"011000110",
  20899=>"000001011",
  20900=>"110100000",
  20901=>"111100000",
  20902=>"101001111",
  20903=>"100010100",
  20904=>"111011101",
  20905=>"011101010",
  20906=>"110110010",
  20907=>"011001000",
  20908=>"000010100",
  20909=>"110101100",
  20910=>"000001011",
  20911=>"100100010",
  20912=>"111110011",
  20913=>"111011110",
  20914=>"011010111",
  20915=>"110000100",
  20916=>"000101000",
  20917=>"010001001",
  20918=>"000101110",
  20919=>"010110100",
  20920=>"111101111",
  20921=>"111000001",
  20922=>"010000111",
  20923=>"110001000",
  20924=>"101011001",
  20925=>"010000110",
  20926=>"100100111",
  20927=>"101101111",
  20928=>"000000010",
  20929=>"000100010",
  20930=>"010111100",
  20931=>"010000000",
  20932=>"011110110",
  20933=>"011110111",
  20934=>"000101101",
  20935=>"001011001",
  20936=>"000101010",
  20937=>"010000000",
  20938=>"111111010",
  20939=>"100011001",
  20940=>"111010011",
  20941=>"001111101",
  20942=>"101011000",
  20943=>"000010101",
  20944=>"001011011",
  20945=>"101100000",
  20946=>"010100000",
  20947=>"000011110",
  20948=>"111110000",
  20949=>"110110001",
  20950=>"100100011",
  20951=>"111000010",
  20952=>"100101100",
  20953=>"001011010",
  20954=>"101000111",
  20955=>"011000000",
  20956=>"000111011",
  20957=>"111101111",
  20958=>"100110111",
  20959=>"100010101",
  20960=>"000100011",
  20961=>"101010101",
  20962=>"110011000",
  20963=>"110111111",
  20964=>"011100111",
  20965=>"100110001",
  20966=>"111101010",
  20967=>"110011100",
  20968=>"011110101",
  20969=>"110101100",
  20970=>"001100110",
  20971=>"011010000",
  20972=>"101100110",
  20973=>"010110110",
  20974=>"000111011",
  20975=>"110100011",
  20976=>"000110001",
  20977=>"110111000",
  20978=>"001110111",
  20979=>"000110000",
  20980=>"010001111",
  20981=>"000111101",
  20982=>"000111010",
  20983=>"001010100",
  20984=>"111111101",
  20985=>"010111011",
  20986=>"110011000",
  20987=>"000110100",
  20988=>"100100000",
  20989=>"100000010",
  20990=>"110101000",
  20991=>"011001000",
  20992=>"100100011",
  20993=>"011010111",
  20994=>"111101110",
  20995=>"000111000",
  20996=>"000111010",
  20997=>"110011011",
  20998=>"111100011",
  20999=>"011100001",
  21000=>"001100110",
  21001=>"001111011",
  21002=>"101000011",
  21003=>"001000100",
  21004=>"010010010",
  21005=>"101011100",
  21006=>"001111000",
  21007=>"110110101",
  21008=>"001011001",
  21009=>"011000000",
  21010=>"000011011",
  21011=>"111010111",
  21012=>"100101100",
  21013=>"110111011",
  21014=>"110111001",
  21015=>"101111111",
  21016=>"101100101",
  21017=>"101000000",
  21018=>"010000110",
  21019=>"011010011",
  21020=>"011000000",
  21021=>"000000111",
  21022=>"101011111",
  21023=>"011000011",
  21024=>"011001100",
  21025=>"110010110",
  21026=>"111101010",
  21027=>"111111101",
  21028=>"100000011",
  21029=>"111101111",
  21030=>"001110010",
  21031=>"101101100",
  21032=>"111100111",
  21033=>"111111001",
  21034=>"011000000",
  21035=>"011010110",
  21036=>"000101111",
  21037=>"110011010",
  21038=>"000000000",
  21039=>"000111111",
  21040=>"001011011",
  21041=>"111001111",
  21042=>"000000111",
  21043=>"000110010",
  21044=>"100010100",
  21045=>"100000011",
  21046=>"100001101",
  21047=>"100000000",
  21048=>"011101111",
  21049=>"011100011",
  21050=>"001110010",
  21051=>"011100000",
  21052=>"001001100",
  21053=>"100001000",
  21054=>"001111000",
  21055=>"010110111",
  21056=>"011110101",
  21057=>"101101110",
  21058=>"111001110",
  21059=>"100000011",
  21060=>"111101000",
  21061=>"001100001",
  21062=>"100000000",
  21063=>"111001011",
  21064=>"100011101",
  21065=>"010011110",
  21066=>"011011000",
  21067=>"100100101",
  21068=>"110011000",
  21069=>"000101101",
  21070=>"100111111",
  21071=>"011101110",
  21072=>"101001110",
  21073=>"111101001",
  21074=>"000101000",
  21075=>"001111000",
  21076=>"110101000",
  21077=>"010111010",
  21078=>"000000010",
  21079=>"011110101",
  21080=>"000011100",
  21081=>"110110001",
  21082=>"000111001",
  21083=>"111101101",
  21084=>"010100110",
  21085=>"010001100",
  21086=>"111110000",
  21087=>"111100111",
  21088=>"011000011",
  21089=>"000101010",
  21090=>"010101110",
  21091=>"011111001",
  21092=>"011010000",
  21093=>"110001000",
  21094=>"010010011",
  21095=>"011001100",
  21096=>"111000011",
  21097=>"011101101",
  21098=>"110100100",
  21099=>"011000011",
  21100=>"100110001",
  21101=>"011111011",
  21102=>"001011000",
  21103=>"011001010",
  21104=>"101001110",
  21105=>"100111001",
  21106=>"001000011",
  21107=>"011001001",
  21108=>"101101010",
  21109=>"100000001",
  21110=>"110010110",
  21111=>"011000100",
  21112=>"111000110",
  21113=>"011000111",
  21114=>"111011100",
  21115=>"010010010",
  21116=>"000111110",
  21117=>"100011010",
  21118=>"110110100",
  21119=>"111000101",
  21120=>"010101100",
  21121=>"100101101",
  21122=>"110000110",
  21123=>"001010011",
  21124=>"011000100",
  21125=>"110011110",
  21126=>"100110010",
  21127=>"100111110",
  21128=>"100011101",
  21129=>"111101100",
  21130=>"110010000",
  21131=>"010010110",
  21132=>"101100100",
  21133=>"011110101",
  21134=>"110110101",
  21135=>"001010101",
  21136=>"101010110",
  21137=>"000001011",
  21138=>"000000001",
  21139=>"010111101",
  21140=>"000000100",
  21141=>"011110011",
  21142=>"011000100",
  21143=>"110011101",
  21144=>"010001010",
  21145=>"000110010",
  21146=>"100000101",
  21147=>"000000010",
  21148=>"000000101",
  21149=>"110100010",
  21150=>"010000111",
  21151=>"100100111",
  21152=>"111011010",
  21153=>"111001011",
  21154=>"100001111",
  21155=>"110110000",
  21156=>"011011010",
  21157=>"001000110",
  21158=>"100101011",
  21159=>"101101000",
  21160=>"010001011",
  21161=>"000000111",
  21162=>"110011010",
  21163=>"101100110",
  21164=>"001000110",
  21165=>"000100101",
  21166=>"010101000",
  21167=>"010100110",
  21168=>"000101011",
  21169=>"010001011",
  21170=>"101111010",
  21171=>"001110110",
  21172=>"110000000",
  21173=>"000010110",
  21174=>"111010110",
  21175=>"001001000",
  21176=>"010100000",
  21177=>"101010110",
  21178=>"010011001",
  21179=>"110000000",
  21180=>"100000100",
  21181=>"100101111",
  21182=>"000001110",
  21183=>"100001000",
  21184=>"100011001",
  21185=>"000001000",
  21186=>"111011010",
  21187=>"001001000",
  21188=>"111000100",
  21189=>"001001101",
  21190=>"110111000",
  21191=>"010010000",
  21192=>"100001000",
  21193=>"101000100",
  21194=>"111110000",
  21195=>"001101111",
  21196=>"110101011",
  21197=>"111000101",
  21198=>"010011110",
  21199=>"000001100",
  21200=>"110001100",
  21201=>"011000000",
  21202=>"001010000",
  21203=>"011100111",
  21204=>"101111111",
  21205=>"110110110",
  21206=>"100010100",
  21207=>"101000101",
  21208=>"111111101",
  21209=>"100100100",
  21210=>"110011111",
  21211=>"011000001",
  21212=>"011000010",
  21213=>"001001111",
  21214=>"000001111",
  21215=>"110001110",
  21216=>"001100101",
  21217=>"111100001",
  21218=>"000110011",
  21219=>"010001011",
  21220=>"110001000",
  21221=>"100001100",
  21222=>"010110000",
  21223=>"110101110",
  21224=>"100111000",
  21225=>"001101000",
  21226=>"001100111",
  21227=>"110010110",
  21228=>"010100101",
  21229=>"001110100",
  21230=>"000110001",
  21231=>"000100100",
  21232=>"100111010",
  21233=>"001101101",
  21234=>"101100111",
  21235=>"001101010",
  21236=>"011011110",
  21237=>"100001001",
  21238=>"000011110",
  21239=>"100000110",
  21240=>"100001111",
  21241=>"110000100",
  21242=>"101111000",
  21243=>"011010100",
  21244=>"011010001",
  21245=>"111100100",
  21246=>"100110010",
  21247=>"010001000",
  21248=>"101000011",
  21249=>"010101110",
  21250=>"000001011",
  21251=>"100111011",
  21252=>"100110101",
  21253=>"000101101",
  21254=>"111011100",
  21255=>"010110100",
  21256=>"100101111",
  21257=>"110001010",
  21258=>"001000100",
  21259=>"010010001",
  21260=>"000111100",
  21261=>"111011100",
  21262=>"000011111",
  21263=>"001110000",
  21264=>"000011101",
  21265=>"110000111",
  21266=>"101000001",
  21267=>"100110110",
  21268=>"110100111",
  21269=>"000101110",
  21270=>"110001100",
  21271=>"100001111",
  21272=>"011111011",
  21273=>"100100111",
  21274=>"101100100",
  21275=>"011001011",
  21276=>"110111001",
  21277=>"100110110",
  21278=>"111101111",
  21279=>"011110010",
  21280=>"100111101",
  21281=>"001111111",
  21282=>"001010110",
  21283=>"001011111",
  21284=>"110110010",
  21285=>"101110010",
  21286=>"101110100",
  21287=>"101110111",
  21288=>"000011110",
  21289=>"010011010",
  21290=>"001001111",
  21291=>"110100000",
  21292=>"111011011",
  21293=>"110001100",
  21294=>"000001011",
  21295=>"100001000",
  21296=>"001101001",
  21297=>"100011011",
  21298=>"001101011",
  21299=>"110011111",
  21300=>"110011000",
  21301=>"010110111",
  21302=>"001010010",
  21303=>"111101010",
  21304=>"111011010",
  21305=>"000010010",
  21306=>"100011010",
  21307=>"110100100",
  21308=>"010101110",
  21309=>"010000000",
  21310=>"011101000",
  21311=>"001111101",
  21312=>"001100001",
  21313=>"110111110",
  21314=>"011001110",
  21315=>"000010111",
  21316=>"111000110",
  21317=>"111011111",
  21318=>"001010111",
  21319=>"010011000",
  21320=>"110011110",
  21321=>"101111000",
  21322=>"011111000",
  21323=>"111011010",
  21324=>"110100110",
  21325=>"100101101",
  21326=>"000100001",
  21327=>"000100100",
  21328=>"100100010",
  21329=>"001111000",
  21330=>"011011110",
  21331=>"110111111",
  21332=>"011110010",
  21333=>"111000100",
  21334=>"111100100",
  21335=>"101000010",
  21336=>"111111011",
  21337=>"110100001",
  21338=>"111110100",
  21339=>"010001001",
  21340=>"011100001",
  21341=>"010000000",
  21342=>"010100100",
  21343=>"111110011",
  21344=>"011100011",
  21345=>"111101001",
  21346=>"100001011",
  21347=>"101011111",
  21348=>"100000001",
  21349=>"101100110",
  21350=>"110100000",
  21351=>"110110100",
  21352=>"001101110",
  21353=>"111010000",
  21354=>"111111100",
  21355=>"001000100",
  21356=>"110110011",
  21357=>"000011100",
  21358=>"001111000",
  21359=>"100010010",
  21360=>"100000100",
  21361=>"101010101",
  21362=>"101011110",
  21363=>"001001111",
  21364=>"010000100",
  21365=>"100101100",
  21366=>"101000110",
  21367=>"110000111",
  21368=>"011010100",
  21369=>"011001000",
  21370=>"111100111",
  21371=>"010010001",
  21372=>"011111001",
  21373=>"100110111",
  21374=>"010100001",
  21375=>"001111101",
  21376=>"001001001",
  21377=>"001001011",
  21378=>"100011110",
  21379=>"110000101",
  21380=>"110100000",
  21381=>"110000011",
  21382=>"110110101",
  21383=>"101001111",
  21384=>"101010100",
  21385=>"101101011",
  21386=>"010100111",
  21387=>"000101011",
  21388=>"101100000",
  21389=>"000110001",
  21390=>"000101011",
  21391=>"001111101",
  21392=>"111001000",
  21393=>"101011101",
  21394=>"011000101",
  21395=>"110011010",
  21396=>"000100011",
  21397=>"001010001",
  21398=>"011100101",
  21399=>"101111000",
  21400=>"001010111",
  21401=>"011111111",
  21402=>"000001110",
  21403=>"110101111",
  21404=>"111110111",
  21405=>"010101011",
  21406=>"101001001",
  21407=>"111011111",
  21408=>"000110101",
  21409=>"110011111",
  21410=>"010011001",
  21411=>"111001010",
  21412=>"010111000",
  21413=>"000000110",
  21414=>"101010110",
  21415=>"000001101",
  21416=>"001111000",
  21417=>"111010111",
  21418=>"011111100",
  21419=>"110000000",
  21420=>"100010001",
  21421=>"010000111",
  21422=>"110101100",
  21423=>"000000110",
  21424=>"000100010",
  21425=>"110101111",
  21426=>"010111100",
  21427=>"010010011",
  21428=>"111100011",
  21429=>"111100011",
  21430=>"011111100",
  21431=>"000111111",
  21432=>"111110000",
  21433=>"011010100",
  21434=>"101001000",
  21435=>"010111001",
  21436=>"110111111",
  21437=>"010000101",
  21438=>"111011010",
  21439=>"001100001",
  21440=>"101100111",
  21441=>"000001111",
  21442=>"100111110",
  21443=>"011110000",
  21444=>"101110111",
  21445=>"011001100",
  21446=>"000101110",
  21447=>"011000011",
  21448=>"101110011",
  21449=>"111010010",
  21450=>"010011000",
  21451=>"101000110",
  21452=>"011011011",
  21453=>"000001110",
  21454=>"000011100",
  21455=>"001001000",
  21456=>"100010111",
  21457=>"100011110",
  21458=>"010110101",
  21459=>"000100101",
  21460=>"010110111",
  21461=>"000011111",
  21462=>"010000110",
  21463=>"111101010",
  21464=>"101011101",
  21465=>"110000010",
  21466=>"100000010",
  21467=>"101010011",
  21468=>"101111000",
  21469=>"001100110",
  21470=>"110010101",
  21471=>"101101101",
  21472=>"101100011",
  21473=>"110100110",
  21474=>"000001111",
  21475=>"110100010",
  21476=>"100000101",
  21477=>"000011111",
  21478=>"000000010",
  21479=>"001110101",
  21480=>"000000110",
  21481=>"001110010",
  21482=>"101111111",
  21483=>"110001110",
  21484=>"001000101",
  21485=>"101110100",
  21486=>"101111101",
  21487=>"110110111",
  21488=>"110100101",
  21489=>"010010100",
  21490=>"000110111",
  21491=>"001000001",
  21492=>"110110011",
  21493=>"100110011",
  21494=>"010011001",
  21495=>"111111100",
  21496=>"100101111",
  21497=>"100100010",
  21498=>"100011100",
  21499=>"100111111",
  21500=>"101001110",
  21501=>"000010000",
  21502=>"100100000",
  21503=>"101010000",
  21504=>"000100001",
  21505=>"101101000",
  21506=>"101011010",
  21507=>"010000101",
  21508=>"101100111",
  21509=>"100011100",
  21510=>"001101101",
  21511=>"110011011",
  21512=>"001101000",
  21513=>"110001010",
  21514=>"100110111",
  21515=>"011101111",
  21516=>"000100010",
  21517=>"111010011",
  21518=>"101111111",
  21519=>"111110110",
  21520=>"101110101",
  21521=>"110101010",
  21522=>"010001011",
  21523=>"011001001",
  21524=>"001011111",
  21525=>"110000110",
  21526=>"000111100",
  21527=>"011011000",
  21528=>"111011111",
  21529=>"100001001",
  21530=>"011000100",
  21531=>"010101101",
  21532=>"100011101",
  21533=>"101001011",
  21534=>"010101011",
  21535=>"010111001",
  21536=>"001110011",
  21537=>"000001110",
  21538=>"010001100",
  21539=>"001001111",
  21540=>"010101110",
  21541=>"101111000",
  21542=>"100010101",
  21543=>"100001110",
  21544=>"011110010",
  21545=>"111100100",
  21546=>"000111111",
  21547=>"101011000",
  21548=>"111111101",
  21549=>"110010011",
  21550=>"011100110",
  21551=>"000010011",
  21552=>"101111110",
  21553=>"101000001",
  21554=>"110101111",
  21555=>"010001010",
  21556=>"100010010",
  21557=>"001001111",
  21558=>"111010111",
  21559=>"110000010",
  21560=>"011101111",
  21561=>"000011110",
  21562=>"100010011",
  21563=>"010101111",
  21564=>"000110001",
  21565=>"110011010",
  21566=>"011101101",
  21567=>"111000001",
  21568=>"101001100",
  21569=>"000111010",
  21570=>"111101011",
  21571=>"001010000",
  21572=>"010001001",
  21573=>"011100010",
  21574=>"100000011",
  21575=>"001100001",
  21576=>"001100000",
  21577=>"100111100",
  21578=>"111101110",
  21579=>"000101010",
  21580=>"000100000",
  21581=>"111011101",
  21582=>"111111001",
  21583=>"001110101",
  21584=>"010110011",
  21585=>"111010010",
  21586=>"000010101",
  21587=>"110110011",
  21588=>"011101110",
  21589=>"000100000",
  21590=>"000000100",
  21591=>"100110100",
  21592=>"110000101",
  21593=>"100110111",
  21594=>"101110000",
  21595=>"111011010",
  21596=>"100010001",
  21597=>"000100100",
  21598=>"111010001",
  21599=>"011001011",
  21600=>"100111000",
  21601=>"101001100",
  21602=>"110111110",
  21603=>"000010000",
  21604=>"010111111",
  21605=>"010111101",
  21606=>"110001001",
  21607=>"110100011",
  21608=>"100100101",
  21609=>"000011100",
  21610=>"110000010",
  21611=>"000000111",
  21612=>"011111111",
  21613=>"111110001",
  21614=>"111101111",
  21615=>"010010111",
  21616=>"111100100",
  21617=>"010100000",
  21618=>"110111111",
  21619=>"110001000",
  21620=>"111011000",
  21621=>"010111110",
  21622=>"101010101",
  21623=>"110011011",
  21624=>"000001101",
  21625=>"110110101",
  21626=>"100011000",
  21627=>"000000011",
  21628=>"000101000",
  21629=>"000001010",
  21630=>"000001110",
  21631=>"110111110",
  21632=>"010000111",
  21633=>"011101010",
  21634=>"011000100",
  21635=>"010010111",
  21636=>"101111100",
  21637=>"111111101",
  21638=>"111000000",
  21639=>"010111011",
  21640=>"000011000",
  21641=>"111011001",
  21642=>"011111011",
  21643=>"000110100",
  21644=>"001000101",
  21645=>"110001011",
  21646=>"100100100",
  21647=>"010000110",
  21648=>"011000000",
  21649=>"000100011",
  21650=>"101100111",
  21651=>"011100000",
  21652=>"001110100",
  21653=>"010110001",
  21654=>"101100010",
  21655=>"110101110",
  21656=>"111001010",
  21657=>"100011111",
  21658=>"110100000",
  21659=>"100100110",
  21660=>"110000010",
  21661=>"011001010",
  21662=>"111011000",
  21663=>"111111111",
  21664=>"101100111",
  21665=>"010000101",
  21666=>"010001110",
  21667=>"110110011",
  21668=>"111111010",
  21669=>"111101111",
  21670=>"001110001",
  21671=>"010001001",
  21672=>"101010000",
  21673=>"111100100",
  21674=>"000110000",
  21675=>"000100000",
  21676=>"101000111",
  21677=>"000100000",
  21678=>"111101101",
  21679=>"011110110",
  21680=>"111100110",
  21681=>"011111010",
  21682=>"111000001",
  21683=>"000000001",
  21684=>"100001111",
  21685=>"110001110",
  21686=>"110111000",
  21687=>"011111111",
  21688=>"111111010",
  21689=>"101101001",
  21690=>"110111000",
  21691=>"010000111",
  21692=>"110111111",
  21693=>"111010010",
  21694=>"011111100",
  21695=>"100111011",
  21696=>"011111011",
  21697=>"010000111",
  21698=>"111110000",
  21699=>"000110101",
  21700=>"000110100",
  21701=>"101111010",
  21702=>"111111010",
  21703=>"011110100",
  21704=>"000000010",
  21705=>"000110011",
  21706=>"111100110",
  21707=>"010011101",
  21708=>"110010000",
  21709=>"011001001",
  21710=>"000100110",
  21711=>"111010110",
  21712=>"001000010",
  21713=>"011101110",
  21714=>"001100110",
  21715=>"111011000",
  21716=>"010111110",
  21717=>"001011101",
  21718=>"110011011",
  21719=>"000011011",
  21720=>"100101101",
  21721=>"001101010",
  21722=>"101100111",
  21723=>"110000101",
  21724=>"011111110",
  21725=>"011010000",
  21726=>"000001100",
  21727=>"000101001",
  21728=>"000001011",
  21729=>"001011000",
  21730=>"111001000",
  21731=>"000100110",
  21732=>"111010001",
  21733=>"000000100",
  21734=>"010111000",
  21735=>"001000010",
  21736=>"011111110",
  21737=>"101010100",
  21738=>"111111011",
  21739=>"100000110",
  21740=>"001101000",
  21741=>"111100011",
  21742=>"000101010",
  21743=>"000010000",
  21744=>"001011111",
  21745=>"111010011",
  21746=>"111101011",
  21747=>"101001010",
  21748=>"111111110",
  21749=>"001011110",
  21750=>"110110011",
  21751=>"100001000",
  21752=>"010000010",
  21753=>"010010111",
  21754=>"110011111",
  21755=>"111001000",
  21756=>"101011000",
  21757=>"110010110",
  21758=>"111101000",
  21759=>"110001100",
  21760=>"011001010",
  21761=>"010001011",
  21762=>"010111100",
  21763=>"101100001",
  21764=>"000111110",
  21765=>"000000100",
  21766=>"010100000",
  21767=>"010011110",
  21768=>"000111100",
  21769=>"100101110",
  21770=>"000110010",
  21771=>"101001001",
  21772=>"101101111",
  21773=>"111111000",
  21774=>"011000001",
  21775=>"110100010",
  21776=>"110100011",
  21777=>"101110101",
  21778=>"101010111",
  21779=>"111010000",
  21780=>"000001100",
  21781=>"110011011",
  21782=>"110111010",
  21783=>"111000100",
  21784=>"110010101",
  21785=>"001000011",
  21786=>"100010001",
  21787=>"001101101",
  21788=>"001110110",
  21789=>"110110111",
  21790=>"101101011",
  21791=>"100000100",
  21792=>"101001010",
  21793=>"000100010",
  21794=>"011010111",
  21795=>"011001101",
  21796=>"010000000",
  21797=>"110100111",
  21798=>"001000010",
  21799=>"011001111",
  21800=>"101011111",
  21801=>"111110101",
  21802=>"110111100",
  21803=>"011101111",
  21804=>"010110011",
  21805=>"100111011",
  21806=>"010010111",
  21807=>"111010111",
  21808=>"110100110",
  21809=>"011100000",
  21810=>"111110110",
  21811=>"001001111",
  21812=>"100000100",
  21813=>"011011010",
  21814=>"011110000",
  21815=>"100000110",
  21816=>"100011100",
  21817=>"001101111",
  21818=>"000100101",
  21819=>"011010100",
  21820=>"111011111",
  21821=>"101010010",
  21822=>"010000010",
  21823=>"100000101",
  21824=>"001000101",
  21825=>"011001111",
  21826=>"111011011",
  21827=>"111111111",
  21828=>"110110000",
  21829=>"010110011",
  21830=>"101000000",
  21831=>"001000110",
  21832=>"001110101",
  21833=>"011100111",
  21834=>"000000100",
  21835=>"100101100",
  21836=>"100001011",
  21837=>"111011010",
  21838=>"010100001",
  21839=>"011001111",
  21840=>"111011110",
  21841=>"010101010",
  21842=>"101000111",
  21843=>"101100111",
  21844=>"000010000",
  21845=>"011010100",
  21846=>"000100011",
  21847=>"110010110",
  21848=>"101010010",
  21849=>"010101101",
  21850=>"110101000",
  21851=>"100100100",
  21852=>"100110000",
  21853=>"100001111",
  21854=>"010100000",
  21855=>"101101110",
  21856=>"101001100",
  21857=>"111001100",
  21858=>"101010110",
  21859=>"010010110",
  21860=>"111101110",
  21861=>"101001011",
  21862=>"000010101",
  21863=>"011110010",
  21864=>"010000100",
  21865=>"000011001",
  21866=>"111011011",
  21867=>"100101010",
  21868=>"011000001",
  21869=>"111101111",
  21870=>"010000000",
  21871=>"000110010",
  21872=>"110010010",
  21873=>"110011010",
  21874=>"000111010",
  21875=>"010100010",
  21876=>"011100010",
  21877=>"010001100",
  21878=>"111001010",
  21879=>"100111110",
  21880=>"111010000",
  21881=>"101010010",
  21882=>"000010110",
  21883=>"011110000",
  21884=>"001101110",
  21885=>"110010011",
  21886=>"110110000",
  21887=>"000111010",
  21888=>"000111010",
  21889=>"000011001",
  21890=>"101110011",
  21891=>"000000010",
  21892=>"100000111",
  21893=>"011100100",
  21894=>"111110110",
  21895=>"000001000",
  21896=>"100000010",
  21897=>"111100100",
  21898=>"010101011",
  21899=>"101000110",
  21900=>"001000101",
  21901=>"111001010",
  21902=>"111011011",
  21903=>"011010000",
  21904=>"101100000",
  21905=>"000110000",
  21906=>"101100010",
  21907=>"101001001",
  21908=>"101000011",
  21909=>"011010001",
  21910=>"110011011",
  21911=>"100110110",
  21912=>"100111000",
  21913=>"101101011",
  21914=>"110000000",
  21915=>"110000010",
  21916=>"100111111",
  21917=>"100011000",
  21918=>"111100010",
  21919=>"000000100",
  21920=>"001110011",
  21921=>"000111111",
  21922=>"110000010",
  21923=>"101111100",
  21924=>"100111010",
  21925=>"011111111",
  21926=>"110011100",
  21927=>"000101000",
  21928=>"000101110",
  21929=>"000101000",
  21930=>"101100000",
  21931=>"100010011",
  21932=>"001111010",
  21933=>"010000001",
  21934=>"000100010",
  21935=>"101010111",
  21936=>"110101010",
  21937=>"101110101",
  21938=>"011001101",
  21939=>"000110110",
  21940=>"101000011",
  21941=>"010011101",
  21942=>"101000111",
  21943=>"011010100",
  21944=>"100011010",
  21945=>"100000011",
  21946=>"000000000",
  21947=>"010000111",
  21948=>"011010000",
  21949=>"111011110",
  21950=>"011011000",
  21951=>"011011000",
  21952=>"111101000",
  21953=>"000101000",
  21954=>"001011111",
  21955=>"010101100",
  21956=>"100000011",
  21957=>"011000000",
  21958=>"100111111",
  21959=>"111100000",
  21960=>"110110111",
  21961=>"001011011",
  21962=>"010110100",
  21963=>"011111101",
  21964=>"011010000",
  21965=>"001101000",
  21966=>"000101101",
  21967=>"101000010",
  21968=>"010111010",
  21969=>"011001101",
  21970=>"110010110",
  21971=>"011001111",
  21972=>"100100010",
  21973=>"101111110",
  21974=>"111001110",
  21975=>"001000010",
  21976=>"111110010",
  21977=>"101001101",
  21978=>"100111101",
  21979=>"111011010",
  21980=>"001000001",
  21981=>"000110010",
  21982=>"010101011",
  21983=>"111101111",
  21984=>"000000000",
  21985=>"110111001",
  21986=>"011100001",
  21987=>"000000010",
  21988=>"010110101",
  21989=>"010011111",
  21990=>"000000000",
  21991=>"011000010",
  21992=>"100110100",
  21993=>"001000011",
  21994=>"100101011",
  21995=>"100110110",
  21996=>"110110001",
  21997=>"101001011",
  21998=>"000101001",
  21999=>"011001101",
  22000=>"011000110",
  22001=>"010000111",
  22002=>"000111110",
  22003=>"110011100",
  22004=>"001001011",
  22005=>"101010001",
  22006=>"111111101",
  22007=>"101101100",
  22008=>"010010100",
  22009=>"111101011",
  22010=>"000110111",
  22011=>"111001000",
  22012=>"001010011",
  22013=>"001001001",
  22014=>"000110110",
  22015=>"000111001",
  22016=>"000100000",
  22017=>"011001010",
  22018=>"010110010",
  22019=>"100001110",
  22020=>"101111011",
  22021=>"101010100",
  22022=>"111111101",
  22023=>"011010001",
  22024=>"001100110",
  22025=>"011101010",
  22026=>"011000010",
  22027=>"000001000",
  22028=>"100100011",
  22029=>"000011000",
  22030=>"111101010",
  22031=>"100011101",
  22032=>"111011000",
  22033=>"001011110",
  22034=>"111011101",
  22035=>"011001000",
  22036=>"100011101",
  22037=>"110111001",
  22038=>"111000011",
  22039=>"100111001",
  22040=>"101111101",
  22041=>"111101001",
  22042=>"101111111",
  22043=>"001111000",
  22044=>"101011001",
  22045=>"110111101",
  22046=>"000000111",
  22047=>"101000010",
  22048=>"110100001",
  22049=>"100111011",
  22050=>"111010000",
  22051=>"000001110",
  22052=>"100101111",
  22053=>"110100000",
  22054=>"100000011",
  22055=>"001001101",
  22056=>"110011100",
  22057=>"010001001",
  22058=>"100001110",
  22059=>"110000101",
  22060=>"111010011",
  22061=>"101100111",
  22062=>"001000111",
  22063=>"111100100",
  22064=>"010110111",
  22065=>"100101011",
  22066=>"111011110",
  22067=>"011000011",
  22068=>"111001100",
  22069=>"010101000",
  22070=>"001001101",
  22071=>"111100011",
  22072=>"001000000",
  22073=>"001001010",
  22074=>"011000001",
  22075=>"011111110",
  22076=>"100001000",
  22077=>"011001100",
  22078=>"100011011",
  22079=>"100111001",
  22080=>"100101101",
  22081=>"000000110",
  22082=>"111101101",
  22083=>"001111110",
  22084=>"010000011",
  22085=>"100111100",
  22086=>"000011100",
  22087=>"111100100",
  22088=>"001101101",
  22089=>"110001101",
  22090=>"001111001",
  22091=>"110111000",
  22092=>"101100001",
  22093=>"110001100",
  22094=>"011001100",
  22095=>"010101001",
  22096=>"100110100",
  22097=>"010001111",
  22098=>"110001010",
  22099=>"011001011",
  22100=>"001111100",
  22101=>"010011001",
  22102=>"001101010",
  22103=>"000011100",
  22104=>"000000100",
  22105=>"111101011",
  22106=>"001000110",
  22107=>"000000110",
  22108=>"011011111",
  22109=>"011001110",
  22110=>"000111001",
  22111=>"111111111",
  22112=>"011011101",
  22113=>"101010111",
  22114=>"011000100",
  22115=>"100111101",
  22116=>"010000010",
  22117=>"001101100",
  22118=>"011011111",
  22119=>"001010001",
  22120=>"101101111",
  22121=>"001001000",
  22122=>"001100111",
  22123=>"111111111",
  22124=>"110100101",
  22125=>"000100001",
  22126=>"101110111",
  22127=>"101101010",
  22128=>"100111100",
  22129=>"000010100",
  22130=>"010111101",
  22131=>"111110000",
  22132=>"100100000",
  22133=>"100000101",
  22134=>"010001000",
  22135=>"101100001",
  22136=>"000100010",
  22137=>"000001000",
  22138=>"010101110",
  22139=>"110001110",
  22140=>"000001011",
  22141=>"000101001",
  22142=>"111010001",
  22143=>"010101100",
  22144=>"011101110",
  22145=>"111110010",
  22146=>"000100011",
  22147=>"100101100",
  22148=>"101111010",
  22149=>"110000100",
  22150=>"010100001",
  22151=>"001001001",
  22152=>"110010011",
  22153=>"010111110",
  22154=>"010110101",
  22155=>"100110011",
  22156=>"001000011",
  22157=>"110110000",
  22158=>"100110010",
  22159=>"000010100",
  22160=>"001010110",
  22161=>"101010010",
  22162=>"111110000",
  22163=>"000100000",
  22164=>"010010011",
  22165=>"000111011",
  22166=>"001000100",
  22167=>"111001010",
  22168=>"000010000",
  22169=>"001001001",
  22170=>"011111010",
  22171=>"010011110",
  22172=>"000011010",
  22173=>"000100110",
  22174=>"000101010",
  22175=>"110111111",
  22176=>"111101111",
  22177=>"001010011",
  22178=>"110001100",
  22179=>"010100010",
  22180=>"110111010",
  22181=>"100011110",
  22182=>"101010111",
  22183=>"010001001",
  22184=>"011101111",
  22185=>"100011000",
  22186=>"001100001",
  22187=>"010011101",
  22188=>"100011111",
  22189=>"101100100",
  22190=>"011011010",
  22191=>"111110101",
  22192=>"101010111",
  22193=>"100001001",
  22194=>"001001110",
  22195=>"111111110",
  22196=>"011011010",
  22197=>"011010111",
  22198=>"011111010",
  22199=>"101001100",
  22200=>"110100101",
  22201=>"000100101",
  22202=>"011011010",
  22203=>"111101001",
  22204=>"001101000",
  22205=>"110110000",
  22206=>"100001100",
  22207=>"101001111",
  22208=>"100111101",
  22209=>"001001001",
  22210=>"001010110",
  22211=>"000000000",
  22212=>"010111001",
  22213=>"000111110",
  22214=>"001011101",
  22215=>"001010100",
  22216=>"100000100",
  22217=>"001100111",
  22218=>"010111000",
  22219=>"001101110",
  22220=>"001010011",
  22221=>"001001000",
  22222=>"111010100",
  22223=>"011000000",
  22224=>"101111011",
  22225=>"000001001",
  22226=>"001010000",
  22227=>"011000101",
  22228=>"000000011",
  22229=>"000100010",
  22230=>"111000001",
  22231=>"001110001",
  22232=>"100111111",
  22233=>"011010101",
  22234=>"101010010",
  22235=>"010111101",
  22236=>"000010100",
  22237=>"011110101",
  22238=>"001111010",
  22239=>"100111011",
  22240=>"101111001",
  22241=>"011010101",
  22242=>"111111000",
  22243=>"101110100",
  22244=>"011110000",
  22245=>"111101111",
  22246=>"001111110",
  22247=>"101110001",
  22248=>"100100000",
  22249=>"000010100",
  22250=>"011010111",
  22251=>"100001111",
  22252=>"001000010",
  22253=>"011101101",
  22254=>"100110000",
  22255=>"101101101",
  22256=>"011111001",
  22257=>"010010100",
  22258=>"011111001",
  22259=>"111100111",
  22260=>"110010111",
  22261=>"000000011",
  22262=>"100110110",
  22263=>"111111100",
  22264=>"111011101",
  22265=>"111101101",
  22266=>"101101110",
  22267=>"100000110",
  22268=>"011100101",
  22269=>"111010011",
  22270=>"101000000",
  22271=>"011010011",
  22272=>"010100001",
  22273=>"000001101",
  22274=>"101111101",
  22275=>"000010101",
  22276=>"101011111",
  22277=>"000100100",
  22278=>"001101010",
  22279=>"000110000",
  22280=>"000001001",
  22281=>"001100101",
  22282=>"000111100",
  22283=>"001101100",
  22284=>"001001010",
  22285=>"000111100",
  22286=>"000110101",
  22287=>"001000111",
  22288=>"110101010",
  22289=>"000101111",
  22290=>"011011100",
  22291=>"010111001",
  22292=>"101010110",
  22293=>"000111110",
  22294=>"111001010",
  22295=>"100100000",
  22296=>"000011011",
  22297=>"100000100",
  22298=>"000000101",
  22299=>"011100101",
  22300=>"001100000",
  22301=>"001110111",
  22302=>"010111110",
  22303=>"100110110",
  22304=>"101000011",
  22305=>"111110110",
  22306=>"001100001",
  22307=>"010110110",
  22308=>"100111000",
  22309=>"110011011",
  22310=>"111100111",
  22311=>"011001101",
  22312=>"111000011",
  22313=>"110100101",
  22314=>"111110000",
  22315=>"001110011",
  22316=>"001000110",
  22317=>"000000000",
  22318=>"001111010",
  22319=>"010001011",
  22320=>"000000100",
  22321=>"000111011",
  22322=>"010101110",
  22323=>"011000100",
  22324=>"001100111",
  22325=>"100100111",
  22326=>"111101111",
  22327=>"110001111",
  22328=>"111110101",
  22329=>"010100111",
  22330=>"001100100",
  22331=>"010001000",
  22332=>"101100101",
  22333=>"110101011",
  22334=>"101101010",
  22335=>"111001100",
  22336=>"110000110",
  22337=>"000010011",
  22338=>"010110001",
  22339=>"111010001",
  22340=>"111001011",
  22341=>"111010001",
  22342=>"111001001",
  22343=>"111111011",
  22344=>"010110001",
  22345=>"000011010",
  22346=>"011100100",
  22347=>"010011011",
  22348=>"101011110",
  22349=>"100000101",
  22350=>"110010010",
  22351=>"001011100",
  22352=>"001110000",
  22353=>"000010100",
  22354=>"010100000",
  22355=>"111111110",
  22356=>"110000010",
  22357=>"101101100",
  22358=>"000110011",
  22359=>"010000010",
  22360=>"100010011",
  22361=>"001001011",
  22362=>"101100011",
  22363=>"001001101",
  22364=>"010110010",
  22365=>"101000011",
  22366=>"110111010",
  22367=>"100000000",
  22368=>"101110100",
  22369=>"000111011",
  22370=>"100101010",
  22371=>"100100101",
  22372=>"001110110",
  22373=>"110011010",
  22374=>"101110111",
  22375=>"101110000",
  22376=>"100101101",
  22377=>"000100110",
  22378=>"110001010",
  22379=>"001001011",
  22380=>"101010100",
  22381=>"110011000",
  22382=>"001110011",
  22383=>"000111010",
  22384=>"111100010",
  22385=>"110110101",
  22386=>"010011101",
  22387=>"011000100",
  22388=>"000100000",
  22389=>"100000111",
  22390=>"100111000",
  22391=>"001111100",
  22392=>"111101010",
  22393=>"010000000",
  22394=>"000010101",
  22395=>"100101001",
  22396=>"000111110",
  22397=>"000010111",
  22398=>"111101111",
  22399=>"001110101",
  22400=>"111100101",
  22401=>"011010100",
  22402=>"001110111",
  22403=>"110001001",
  22404=>"010010001",
  22405=>"111110110",
  22406=>"100111100",
  22407=>"100111111",
  22408=>"101010010",
  22409=>"101011011",
  22410=>"101111000",
  22411=>"100101110",
  22412=>"001010001",
  22413=>"100001011",
  22414=>"001100010",
  22415=>"100010000",
  22416=>"000000110",
  22417=>"010110010",
  22418=>"010111110",
  22419=>"001000011",
  22420=>"000100100",
  22421=>"010101100",
  22422=>"000100100",
  22423=>"010100011",
  22424=>"011111100",
  22425=>"100011010",
  22426=>"101000100",
  22427=>"100011011",
  22428=>"011001111",
  22429=>"110111010",
  22430=>"111001010",
  22431=>"111010101",
  22432=>"000110011",
  22433=>"101110010",
  22434=>"100100100",
  22435=>"100011010",
  22436=>"001001111",
  22437=>"110010001",
  22438=>"100100101",
  22439=>"010100101",
  22440=>"100000101",
  22441=>"000110011",
  22442=>"011110011",
  22443=>"000010000",
  22444=>"111100100",
  22445=>"001010100",
  22446=>"101010010",
  22447=>"100000010",
  22448=>"011011110",
  22449=>"101000011",
  22450=>"011010010",
  22451=>"110001101",
  22452=>"010101010",
  22453=>"110001000",
  22454=>"110110010",
  22455=>"111000111",
  22456=>"111101011",
  22457=>"010011100",
  22458=>"010110000",
  22459=>"110101000",
  22460=>"011111100",
  22461=>"101010011",
  22462=>"101011100",
  22463=>"111100110",
  22464=>"010011111",
  22465=>"100110101",
  22466=>"100110110",
  22467=>"000100001",
  22468=>"001100011",
  22469=>"010000110",
  22470=>"111001010",
  22471=>"100001001",
  22472=>"011010000",
  22473=>"010110010",
  22474=>"100010111",
  22475=>"010010111",
  22476=>"100011101",
  22477=>"001101111",
  22478=>"001000110",
  22479=>"100100110",
  22480=>"110001100",
  22481=>"010001100",
  22482=>"111001001",
  22483=>"010000000",
  22484=>"101100001",
  22485=>"101111000",
  22486=>"000010010",
  22487=>"111100101",
  22488=>"000100100",
  22489=>"010010000",
  22490=>"001010110",
  22491=>"000011000",
  22492=>"010000100",
  22493=>"010001100",
  22494=>"000111100",
  22495=>"111100010",
  22496=>"111111111",
  22497=>"011000010",
  22498=>"011011101",
  22499=>"110011100",
  22500=>"111110001",
  22501=>"011110101",
  22502=>"000011111",
  22503=>"011001011",
  22504=>"011100000",
  22505=>"011101011",
  22506=>"110110100",
  22507=>"011111101",
  22508=>"010111010",
  22509=>"010100000",
  22510=>"010110011",
  22511=>"010101001",
  22512=>"010000001",
  22513=>"110111001",
  22514=>"001001001",
  22515=>"000100010",
  22516=>"000011010",
  22517=>"010101001",
  22518=>"010011110",
  22519=>"011101001",
  22520=>"110110011",
  22521=>"100110000",
  22522=>"111101101",
  22523=>"100110010",
  22524=>"001010000",
  22525=>"110100100",
  22526=>"010011101",
  22527=>"000010000",
  22528=>"110110001",
  22529=>"010111100",
  22530=>"001111001",
  22531=>"111101101",
  22532=>"101011001",
  22533=>"101000101",
  22534=>"100101101",
  22535=>"001100111",
  22536=>"000010110",
  22537=>"110101101",
  22538=>"011100101",
  22539=>"010100111",
  22540=>"111000111",
  22541=>"011011011",
  22542=>"011111111",
  22543=>"000001110",
  22544=>"000011011",
  22545=>"111110001",
  22546=>"101111010",
  22547=>"011010000",
  22548=>"011101010",
  22549=>"001001100",
  22550=>"000101010",
  22551=>"101100111",
  22552=>"101111000",
  22553=>"000101110",
  22554=>"001100110",
  22555=>"110000001",
  22556=>"011001011",
  22557=>"111000110",
  22558=>"010111000",
  22559=>"100101001",
  22560=>"011011011",
  22561=>"010011100",
  22562=>"111101111",
  22563=>"010001110",
  22564=>"111101111",
  22565=>"110001111",
  22566=>"000110010",
  22567=>"001111011",
  22568=>"000110100",
  22569=>"111010110",
  22570=>"111101111",
  22571=>"110010110",
  22572=>"100000100",
  22573=>"001011011",
  22574=>"010110000",
  22575=>"101010111",
  22576=>"010000010",
  22577=>"111101001",
  22578=>"001111000",
  22579=>"110000001",
  22580=>"000110000",
  22581=>"010111000",
  22582=>"110001111",
  22583=>"011100110",
  22584=>"101110001",
  22585=>"110100110",
  22586=>"010111100",
  22587=>"110100110",
  22588=>"010000101",
  22589=>"110010011",
  22590=>"000101101",
  22591=>"000111000",
  22592=>"100001111",
  22593=>"001000000",
  22594=>"001111111",
  22595=>"100110100",
  22596=>"101100101",
  22597=>"100010100",
  22598=>"100001011",
  22599=>"011110111",
  22600=>"100001011",
  22601=>"100011011",
  22602=>"100000000",
  22603=>"000010101",
  22604=>"000100100",
  22605=>"011100011",
  22606=>"111001111",
  22607=>"010101001",
  22608=>"110100101",
  22609=>"110010001",
  22610=>"011111101",
  22611=>"011001110",
  22612=>"101000100",
  22613=>"001110110",
  22614=>"101110000",
  22615=>"000001011",
  22616=>"010010001",
  22617=>"011101001",
  22618=>"000100011",
  22619=>"101100110",
  22620=>"111100011",
  22621=>"110101100",
  22622=>"000000111",
  22623=>"101101001",
  22624=>"001101011",
  22625=>"010110100",
  22626=>"010000100",
  22627=>"000001001",
  22628=>"111100100",
  22629=>"000000000",
  22630=>"101110011",
  22631=>"100110001",
  22632=>"001101111",
  22633=>"000111110",
  22634=>"111110111",
  22635=>"100000111",
  22636=>"010010101",
  22637=>"011101110",
  22638=>"001011011",
  22639=>"110001101",
  22640=>"111101010",
  22641=>"001001011",
  22642=>"110110000",
  22643=>"010110111",
  22644=>"000001110",
  22645=>"101011110",
  22646=>"100010100",
  22647=>"010100101",
  22648=>"110101110",
  22649=>"001001100",
  22650=>"010110100",
  22651=>"001111011",
  22652=>"110010000",
  22653=>"101110000",
  22654=>"000000000",
  22655=>"001000000",
  22656=>"111100001",
  22657=>"110100001",
  22658=>"100111100",
  22659=>"000111110",
  22660=>"100111110",
  22661=>"010001101",
  22662=>"010011111",
  22663=>"001111000",
  22664=>"101001001",
  22665=>"111011110",
  22666=>"100010111",
  22667=>"110010010",
  22668=>"011011000",
  22669=>"100011001",
  22670=>"110011010",
  22671=>"110101101",
  22672=>"000100110",
  22673=>"100011111",
  22674=>"000111011",
  22675=>"000001010",
  22676=>"011001010",
  22677=>"000001110",
  22678=>"100000101",
  22679=>"101100101",
  22680=>"101101011",
  22681=>"101010000",
  22682=>"011001001",
  22683=>"110101101",
  22684=>"000001101",
  22685=>"101100000",
  22686=>"000100001",
  22687=>"001010110",
  22688=>"001000010",
  22689=>"101000100",
  22690=>"001111011",
  22691=>"010101000",
  22692=>"111011110",
  22693=>"010010000",
  22694=>"001101011",
  22695=>"000001100",
  22696=>"100101010",
  22697=>"010001011",
  22698=>"001100100",
  22699=>"101001011",
  22700=>"101001011",
  22701=>"001101001",
  22702=>"101111111",
  22703=>"101001000",
  22704=>"110010101",
  22705=>"001111001",
  22706=>"001010000",
  22707=>"010001101",
  22708=>"010111111",
  22709=>"101000010",
  22710=>"011110100",
  22711=>"000000010",
  22712=>"101011000",
  22713=>"011111001",
  22714=>"010000100",
  22715=>"110101111",
  22716=>"111111110",
  22717=>"111011101",
  22718=>"111011001",
  22719=>"101110111",
  22720=>"100010100",
  22721=>"010100101",
  22722=>"010011100",
  22723=>"111100011",
  22724=>"000010111",
  22725=>"011000001",
  22726=>"001001010",
  22727=>"001011000",
  22728=>"100100000",
  22729=>"010000000",
  22730=>"111000111",
  22731=>"111111010",
  22732=>"001011011",
  22733=>"000000000",
  22734=>"001110110",
  22735=>"110100011",
  22736=>"101110110",
  22737=>"101011111",
  22738=>"000110101",
  22739=>"110111100",
  22740=>"100000101",
  22741=>"110101010",
  22742=>"000000111",
  22743=>"000000010",
  22744=>"110000110",
  22745=>"011001101",
  22746=>"111100100",
  22747=>"011000110",
  22748=>"100000100",
  22749=>"111111101",
  22750=>"110101110",
  22751=>"111111101",
  22752=>"010001011",
  22753=>"110101111",
  22754=>"001000011",
  22755=>"110110001",
  22756=>"001000010",
  22757=>"110101011",
  22758=>"010000010",
  22759=>"100010110",
  22760=>"100111111",
  22761=>"110011110",
  22762=>"101010111",
  22763=>"100001000",
  22764=>"101011010",
  22765=>"000000011",
  22766=>"000100001",
  22767=>"000110101",
  22768=>"011111110",
  22769=>"101101110",
  22770=>"100101101",
  22771=>"111100000",
  22772=>"010110011",
  22773=>"010010101",
  22774=>"110110010",
  22775=>"100110101",
  22776=>"000000101",
  22777=>"010010001",
  22778=>"011101001",
  22779=>"011011000",
  22780=>"101100101",
  22781=>"000011001",
  22782=>"001011001",
  22783=>"000001111",
  22784=>"100111100",
  22785=>"000011001",
  22786=>"011010110",
  22787=>"011100011",
  22788=>"110001010",
  22789=>"001110010",
  22790=>"011000001",
  22791=>"001001011",
  22792=>"110011000",
  22793=>"000011010",
  22794=>"101100101",
  22795=>"101111011",
  22796=>"010101110",
  22797=>"100000111",
  22798=>"001101001",
  22799=>"000011001",
  22800=>"101010000",
  22801=>"110011001",
  22802=>"100001010",
  22803=>"110111111",
  22804=>"000110110",
  22805=>"011001010",
  22806=>"111100000",
  22807=>"110110001",
  22808=>"101111100",
  22809=>"000100101",
  22810=>"101011010",
  22811=>"101010011",
  22812=>"011110101",
  22813=>"110011001",
  22814=>"111001011",
  22815=>"000010100",
  22816=>"011100100",
  22817=>"000101011",
  22818=>"100000101",
  22819=>"001001000",
  22820=>"110101101",
  22821=>"010110001",
  22822=>"110011010",
  22823=>"111001110",
  22824=>"010101000",
  22825=>"101010100",
  22826=>"111110111",
  22827=>"000010111",
  22828=>"101010101",
  22829=>"100011000",
  22830=>"011110000",
  22831=>"000110110",
  22832=>"101100001",
  22833=>"111100111",
  22834=>"010100101",
  22835=>"000111011",
  22836=>"010000000",
  22837=>"001011000",
  22838=>"100110000",
  22839=>"001000000",
  22840=>"000111010",
  22841=>"000101110",
  22842=>"000000010",
  22843=>"111100101",
  22844=>"111010000",
  22845=>"001100010",
  22846=>"001001110",
  22847=>"000001101",
  22848=>"000010000",
  22849=>"000100110",
  22850=>"110110011",
  22851=>"110101100",
  22852=>"111011111",
  22853=>"000101100",
  22854=>"001010111",
  22855=>"001111001",
  22856=>"010111111",
  22857=>"001110010",
  22858=>"111111101",
  22859=>"001110110",
  22860=>"100110100",
  22861=>"100111010",
  22862=>"101010001",
  22863=>"111000011",
  22864=>"101111101",
  22865=>"110101110",
  22866=>"101000100",
  22867=>"100000000",
  22868=>"011111110",
  22869=>"000111111",
  22870=>"111010000",
  22871=>"101011100",
  22872=>"011101110",
  22873=>"100000011",
  22874=>"000001100",
  22875=>"111100111",
  22876=>"010101100",
  22877=>"101110111",
  22878=>"010000100",
  22879=>"000111000",
  22880=>"100110100",
  22881=>"010000010",
  22882=>"000000000",
  22883=>"000110010",
  22884=>"111111101",
  22885=>"100011100",
  22886=>"000000110",
  22887=>"011000011",
  22888=>"111101111",
  22889=>"001110111",
  22890=>"110110101",
  22891=>"111100001",
  22892=>"000111100",
  22893=>"101001000",
  22894=>"101010000",
  22895=>"011011000",
  22896=>"111110100",
  22897=>"011100000",
  22898=>"101010110",
  22899=>"101100010",
  22900=>"110101000",
  22901=>"011101111",
  22902=>"010011110",
  22903=>"111000011",
  22904=>"001111101",
  22905=>"111111001",
  22906=>"111111011",
  22907=>"000000011",
  22908=>"111101001",
  22909=>"011010101",
  22910=>"001110001",
  22911=>"101000011",
  22912=>"000101000",
  22913=>"100100100",
  22914=>"100001111",
  22915=>"011101110",
  22916=>"101111010",
  22917=>"100111001",
  22918=>"110010010",
  22919=>"111000101",
  22920=>"000000000",
  22921=>"111100110",
  22922=>"011010011",
  22923=>"001010110",
  22924=>"000001100",
  22925=>"011011101",
  22926=>"001100000",
  22927=>"111110001",
  22928=>"001001101",
  22929=>"001001100",
  22930=>"010000100",
  22931=>"010111101",
  22932=>"010100100",
  22933=>"001000110",
  22934=>"000000100",
  22935=>"000010010",
  22936=>"001101000",
  22937=>"010101011",
  22938=>"000111011",
  22939=>"110001110",
  22940=>"100100000",
  22941=>"011100001",
  22942=>"001101001",
  22943=>"001111110",
  22944=>"110001100",
  22945=>"000011101",
  22946=>"100111000",
  22947=>"001011100",
  22948=>"000100101",
  22949=>"100110101",
  22950=>"000100000",
  22951=>"000010111",
  22952=>"001000011",
  22953=>"101000110",
  22954=>"001001000",
  22955=>"010110111",
  22956=>"110111011",
  22957=>"001110101",
  22958=>"111001010",
  22959=>"101000010",
  22960=>"001010000",
  22961=>"000010100",
  22962=>"011001001",
  22963=>"111100111",
  22964=>"011101101",
  22965=>"101000011",
  22966=>"010011010",
  22967=>"001011000",
  22968=>"010110001",
  22969=>"101011100",
  22970=>"000110110",
  22971=>"101101111",
  22972=>"001001010",
  22973=>"100011010",
  22974=>"100010100",
  22975=>"000111001",
  22976=>"100011100",
  22977=>"111110110",
  22978=>"000111110",
  22979=>"011101111",
  22980=>"000011010",
  22981=>"010011111",
  22982=>"110011011",
  22983=>"100111101",
  22984=>"000110100",
  22985=>"111010000",
  22986=>"001110010",
  22987=>"110101011",
  22988=>"011001000",
  22989=>"010010010",
  22990=>"011011101",
  22991=>"000001110",
  22992=>"010001110",
  22993=>"100010101",
  22994=>"010001001",
  22995=>"000010101",
  22996=>"010111011",
  22997=>"010000000",
  22998=>"011110101",
  22999=>"011100000",
  23000=>"001010010",
  23001=>"010101101",
  23002=>"111110001",
  23003=>"100111010",
  23004=>"011101111",
  23005=>"001010101",
  23006=>"000100010",
  23007=>"001000011",
  23008=>"101000010",
  23009=>"011001010",
  23010=>"101100110",
  23011=>"110100001",
  23012=>"101101011",
  23013=>"000011010",
  23014=>"000110111",
  23015=>"001010111",
  23016=>"010010000",
  23017=>"001101111",
  23018=>"110101000",
  23019=>"001011111",
  23020=>"101111100",
  23021=>"011000100",
  23022=>"011000111",
  23023=>"011111000",
  23024=>"000010011",
  23025=>"100011000",
  23026=>"111110010",
  23027=>"101001010",
  23028=>"100011000",
  23029=>"011111101",
  23030=>"100001100",
  23031=>"111001011",
  23032=>"000110101",
  23033=>"010110010",
  23034=>"111000101",
  23035=>"110101010",
  23036=>"001011011",
  23037=>"100001100",
  23038=>"001010010",
  23039=>"010111001",
  23040=>"000010000",
  23041=>"011001101",
  23042=>"000000101",
  23043=>"010100000",
  23044=>"110010101",
  23045=>"000100010",
  23046=>"001011001",
  23047=>"010101101",
  23048=>"010000000",
  23049=>"000000111",
  23050=>"110101111",
  23051=>"110101110",
  23052=>"110000010",
  23053=>"011101011",
  23054=>"111110101",
  23055=>"110111110",
  23056=>"011010100",
  23057=>"111000111",
  23058=>"010111100",
  23059=>"010101111",
  23060=>"101010101",
  23061=>"001001001",
  23062=>"101011000",
  23063=>"010111101",
  23064=>"011101111",
  23065=>"110011010",
  23066=>"000000100",
  23067=>"010010100",
  23068=>"101111010",
  23069=>"100100001",
  23070=>"111100101",
  23071=>"111001110",
  23072=>"111100100",
  23073=>"000110101",
  23074=>"010111011",
  23075=>"111001011",
  23076=>"010010111",
  23077=>"110010111",
  23078=>"111110001",
  23079=>"100100110",
  23080=>"001100011",
  23081=>"000000010",
  23082=>"100011111",
  23083=>"001001001",
  23084=>"110000100",
  23085=>"000110000",
  23086=>"111110001",
  23087=>"100111001",
  23088=>"100001010",
  23089=>"111010110",
  23090=>"000011000",
  23091=>"010000001",
  23092=>"011100001",
  23093=>"101111011",
  23094=>"100101101",
  23095=>"011110001",
  23096=>"101111011",
  23097=>"010100001",
  23098=>"101000001",
  23099=>"011100111",
  23100=>"101011110",
  23101=>"110000011",
  23102=>"010101100",
  23103=>"101110001",
  23104=>"001000011",
  23105=>"100101101",
  23106=>"110110110",
  23107=>"010001100",
  23108=>"010110111",
  23109=>"001101001",
  23110=>"010110100",
  23111=>"100010011",
  23112=>"110001101",
  23113=>"111001011",
  23114=>"011011110",
  23115=>"101111110",
  23116=>"111110111",
  23117=>"000100110",
  23118=>"010100010",
  23119=>"011011100",
  23120=>"010100100",
  23121=>"011000111",
  23122=>"101100100",
  23123=>"000100110",
  23124=>"110000010",
  23125=>"000110110",
  23126=>"000011000",
  23127=>"001111111",
  23128=>"111001001",
  23129=>"010010110",
  23130=>"101111101",
  23131=>"101110111",
  23132=>"011001000",
  23133=>"100011100",
  23134=>"000100010",
  23135=>"100000000",
  23136=>"110011010",
  23137=>"111001010",
  23138=>"100001000",
  23139=>"000100001",
  23140=>"111010010",
  23141=>"000001101",
  23142=>"010100111",
  23143=>"010111111",
  23144=>"110011000",
  23145=>"001100100",
  23146=>"010000011",
  23147=>"000100010",
  23148=>"001101000",
  23149=>"110000110",
  23150=>"100011100",
  23151=>"011100010",
  23152=>"110000001",
  23153=>"010111110",
  23154=>"110100110",
  23155=>"111111011",
  23156=>"100010111",
  23157=>"011010110",
  23158=>"101101001",
  23159=>"001110001",
  23160=>"110011101",
  23161=>"010111101",
  23162=>"100000100",
  23163=>"101110000",
  23164=>"111010101",
  23165=>"110100110",
  23166=>"001100011",
  23167=>"010010100",
  23168=>"010010000",
  23169=>"110001111",
  23170=>"111111011",
  23171=>"111101100",
  23172=>"010100101",
  23173=>"100000000",
  23174=>"001111101",
  23175=>"000101010",
  23176=>"111000110",
  23177=>"101101000",
  23178=>"010000111",
  23179=>"001110001",
  23180=>"011101001",
  23181=>"110000000",
  23182=>"110100010",
  23183=>"010101000",
  23184=>"111101001",
  23185=>"000101111",
  23186=>"011001011",
  23187=>"100101100",
  23188=>"010000000",
  23189=>"011000100",
  23190=>"001101001",
  23191=>"110010011",
  23192=>"001101001",
  23193=>"111010110",
  23194=>"111110110",
  23195=>"110000010",
  23196=>"101110100",
  23197=>"011110101",
  23198=>"011001011",
  23199=>"101001110",
  23200=>"110110000",
  23201=>"101100011",
  23202=>"101011110",
  23203=>"001001100",
  23204=>"111101011",
  23205=>"111001101",
  23206=>"101101110",
  23207=>"110100011",
  23208=>"101110011",
  23209=>"011111000",
  23210=>"001000101",
  23211=>"101001100",
  23212=>"001000001",
  23213=>"000000011",
  23214=>"011011111",
  23215=>"011111010",
  23216=>"101000111",
  23217=>"010000101",
  23218=>"111000100",
  23219=>"110101110",
  23220=>"100011111",
  23221=>"111101101",
  23222=>"100111101",
  23223=>"100101100",
  23224=>"100010001",
  23225=>"000010001",
  23226=>"111011111",
  23227=>"000010001",
  23228=>"110110111",
  23229=>"011101000",
  23230=>"010110101",
  23231=>"010001001",
  23232=>"000000011",
  23233=>"110110110",
  23234=>"100101100",
  23235=>"100011011",
  23236=>"011000101",
  23237=>"111001110",
  23238=>"011100011",
  23239=>"011100001",
  23240=>"101100001",
  23241=>"110101000",
  23242=>"010011000",
  23243=>"010001101",
  23244=>"000011111",
  23245=>"100011001",
  23246=>"101101000",
  23247=>"010010010",
  23248=>"010010010",
  23249=>"110011110",
  23250=>"000100110",
  23251=>"011010011",
  23252=>"111110011",
  23253=>"010001110",
  23254=>"110011101",
  23255=>"001101010",
  23256=>"000001010",
  23257=>"111001011",
  23258=>"001110100",
  23259=>"000110010",
  23260=>"010111110",
  23261=>"001100000",
  23262=>"111000010",
  23263=>"001111101",
  23264=>"110101100",
  23265=>"110000001",
  23266=>"110100100",
  23267=>"010100011",
  23268=>"101111001",
  23269=>"100110000",
  23270=>"100100000",
  23271=>"001111101",
  23272=>"001011111",
  23273=>"100010101",
  23274=>"011010011",
  23275=>"000011101",
  23276=>"111101110",
  23277=>"101110111",
  23278=>"000011111",
  23279=>"101100011",
  23280=>"101100010",
  23281=>"001110001",
  23282=>"001100010",
  23283=>"100110001",
  23284=>"111010110",
  23285=>"001001111",
  23286=>"110111100",
  23287=>"001000101",
  23288=>"001001101",
  23289=>"010000001",
  23290=>"110000100",
  23291=>"000001111",
  23292=>"110000110",
  23293=>"011010011",
  23294=>"010100001",
  23295=>"000010010",
  23296=>"000110011",
  23297=>"111101000",
  23298=>"100110011",
  23299=>"011000000",
  23300=>"101101110",
  23301=>"110111010",
  23302=>"110110000",
  23303=>"000011010",
  23304=>"111000001",
  23305=>"001111101",
  23306=>"101010101",
  23307=>"111100111",
  23308=>"111011101",
  23309=>"011110100",
  23310=>"110101100",
  23311=>"001101000",
  23312=>"001111110",
  23313=>"110000101",
  23314=>"111010001",
  23315=>"111010111",
  23316=>"001100000",
  23317=>"111001000",
  23318=>"111100100",
  23319=>"001010100",
  23320=>"110010101",
  23321=>"000010011",
  23322=>"001111110",
  23323=>"101101000",
  23324=>"100001010",
  23325=>"100011100",
  23326=>"110010100",
  23327=>"010010111",
  23328=>"011101111",
  23329=>"011101100",
  23330=>"011101110",
  23331=>"000011011",
  23332=>"110001001",
  23333=>"011101010",
  23334=>"011100111",
  23335=>"111001101",
  23336=>"001101011",
  23337=>"101100000",
  23338=>"100111000",
  23339=>"110011100",
  23340=>"110001010",
  23341=>"000100101",
  23342=>"011000010",
  23343=>"110000011",
  23344=>"111100110",
  23345=>"011011000",
  23346=>"111100010",
  23347=>"100110010",
  23348=>"111110100",
  23349=>"001011110",
  23350=>"001100011",
  23351=>"010001001",
  23352=>"101101101",
  23353=>"001001000",
  23354=>"001001110",
  23355=>"010010111",
  23356=>"101101110",
  23357=>"010101011",
  23358=>"111100010",
  23359=>"000001100",
  23360=>"111101010",
  23361=>"101010111",
  23362=>"100111001",
  23363=>"101111111",
  23364=>"111101011",
  23365=>"111011000",
  23366=>"101101100",
  23367=>"101011001",
  23368=>"101000000",
  23369=>"011010100",
  23370=>"000100100",
  23371=>"111110000",
  23372=>"101110010",
  23373=>"010100011",
  23374=>"001100011",
  23375=>"000111000",
  23376=>"110110011",
  23377=>"100101001",
  23378=>"111101110",
  23379=>"000010000",
  23380=>"111001000",
  23381=>"101100110",
  23382=>"100001111",
  23383=>"010001101",
  23384=>"100001101",
  23385=>"010001101",
  23386=>"000100101",
  23387=>"101000101",
  23388=>"101101010",
  23389=>"100111000",
  23390=>"101011011",
  23391=>"110000101",
  23392=>"100101011",
  23393=>"011000111",
  23394=>"111101101",
  23395=>"000110010",
  23396=>"010100001",
  23397=>"100011001",
  23398=>"100100101",
  23399=>"000000110",
  23400=>"101011101",
  23401=>"110100111",
  23402=>"111011100",
  23403=>"100001111",
  23404=>"101010001",
  23405=>"011100011",
  23406=>"011100001",
  23407=>"100010001",
  23408=>"110011100",
  23409=>"000101101",
  23410=>"000110100",
  23411=>"100101100",
  23412=>"110110011",
  23413=>"001010100",
  23414=>"100001010",
  23415=>"111110111",
  23416=>"100011000",
  23417=>"000001101",
  23418=>"101000111",
  23419=>"110111111",
  23420=>"011101001",
  23421=>"101100100",
  23422=>"010110010",
  23423=>"001001111",
  23424=>"110100111",
  23425=>"111110010",
  23426=>"111100100",
  23427=>"001111110",
  23428=>"001100010",
  23429=>"101100111",
  23430=>"001011001",
  23431=>"001001101",
  23432=>"011000000",
  23433=>"110011100",
  23434=>"111110001",
  23435=>"011001011",
  23436=>"001010100",
  23437=>"111111011",
  23438=>"100000000",
  23439=>"111011001",
  23440=>"111001110",
  23441=>"111111010",
  23442=>"111010000",
  23443=>"100110010",
  23444=>"111101100",
  23445=>"111101101",
  23446=>"101111011",
  23447=>"000010110",
  23448=>"111101100",
  23449=>"111111001",
  23450=>"100010110",
  23451=>"011100000",
  23452=>"001010101",
  23453=>"000101010",
  23454=>"010010001",
  23455=>"101110111",
  23456=>"100000101",
  23457=>"101110011",
  23458=>"000111110",
  23459=>"101100011",
  23460=>"111100101",
  23461=>"101111100",
  23462=>"101100110",
  23463=>"101011001",
  23464=>"010110001",
  23465=>"001010000",
  23466=>"111110111",
  23467=>"001001000",
  23468=>"111000011",
  23469=>"000010011",
  23470=>"001011000",
  23471=>"000110010",
  23472=>"100001010",
  23473=>"010101100",
  23474=>"010111001",
  23475=>"111001100",
  23476=>"101001100",
  23477=>"000100001",
  23478=>"001101001",
  23479=>"011010001",
  23480=>"110000101",
  23481=>"000010001",
  23482=>"111101000",
  23483=>"110110110",
  23484=>"100011000",
  23485=>"011101001",
  23486=>"111100111",
  23487=>"101001001",
  23488=>"011010011",
  23489=>"101100010",
  23490=>"000111011",
  23491=>"000100010",
  23492=>"111111010",
  23493=>"111111011",
  23494=>"100101110",
  23495=>"011011101",
  23496=>"100110010",
  23497=>"011101000",
  23498=>"011001100",
  23499=>"100011110",
  23500=>"110001110",
  23501=>"100100000",
  23502=>"001001101",
  23503=>"010110110",
  23504=>"111010101",
  23505=>"110000000",
  23506=>"101011001",
  23507=>"001101100",
  23508=>"110010100",
  23509=>"001100101",
  23510=>"110000010",
  23511=>"000100001",
  23512=>"100100000",
  23513=>"111011100",
  23514=>"111100100",
  23515=>"110110100",
  23516=>"111111111",
  23517=>"110111111",
  23518=>"000000000",
  23519=>"111010101",
  23520=>"010010001",
  23521=>"101101011",
  23522=>"011011101",
  23523=>"010101000",
  23524=>"101001110",
  23525=>"110101100",
  23526=>"100000101",
  23527=>"100110001",
  23528=>"011110101",
  23529=>"110101011",
  23530=>"101010110",
  23531=>"000100011",
  23532=>"110010011",
  23533=>"101101111",
  23534=>"000000010",
  23535=>"100111111",
  23536=>"100001111",
  23537=>"101011011",
  23538=>"011011000",
  23539=>"000001111",
  23540=>"110101000",
  23541=>"111111011",
  23542=>"111001001",
  23543=>"100011100",
  23544=>"111100001",
  23545=>"000001001",
  23546=>"110010100",
  23547=>"101110000",
  23548=>"011000000",
  23549=>"011001010",
  23550=>"100101010",
  23551=>"101111101",
  23552=>"110111110",
  23553=>"000101100",
  23554=>"100110110",
  23555=>"000111000",
  23556=>"101011101",
  23557=>"001000001",
  23558=>"101101001",
  23559=>"000101100",
  23560=>"110100110",
  23561=>"101111111",
  23562=>"001101110",
  23563=>"010100011",
  23564=>"100100000",
  23565=>"110010001",
  23566=>"000011110",
  23567=>"010101010",
  23568=>"100011011",
  23569=>"100000110",
  23570=>"111111111",
  23571=>"011001100",
  23572=>"010010100",
  23573=>"111110100",
  23574=>"011101111",
  23575=>"100000100",
  23576=>"011011110",
  23577=>"000000101",
  23578=>"000011110",
  23579=>"000100001",
  23580=>"101101100",
  23581=>"000110111",
  23582=>"010110111",
  23583=>"001100010",
  23584=>"011011100",
  23585=>"010001101",
  23586=>"001100110",
  23587=>"100011111",
  23588=>"101011010",
  23589=>"000010110",
  23590=>"010011010",
  23591=>"000111110",
  23592=>"101000101",
  23593=>"010011001",
  23594=>"110011011",
  23595=>"101111100",
  23596=>"111011110",
  23597=>"001001101",
  23598=>"011101100",
  23599=>"010110101",
  23600=>"011011010",
  23601=>"000110010",
  23602=>"100010010",
  23603=>"001000110",
  23604=>"000101000",
  23605=>"010101001",
  23606=>"110100001",
  23607=>"010010011",
  23608=>"010101100",
  23609=>"000110010",
  23610=>"001011100",
  23611=>"101110101",
  23612=>"011000001",
  23613=>"001101011",
  23614=>"101100011",
  23615=>"000101010",
  23616=>"110111010",
  23617=>"001100010",
  23618=>"101111001",
  23619=>"000110001",
  23620=>"111010010",
  23621=>"000111001",
  23622=>"100110001",
  23623=>"011010101",
  23624=>"100111010",
  23625=>"101000011",
  23626=>"101000100",
  23627=>"000101010",
  23628=>"110000011",
  23629=>"101001101",
  23630=>"111111011",
  23631=>"101000011",
  23632=>"010000110",
  23633=>"000010100",
  23634=>"010010110",
  23635=>"111001101",
  23636=>"001010100",
  23637=>"111111100",
  23638=>"001011000",
  23639=>"000010111",
  23640=>"100110110",
  23641=>"101111101",
  23642=>"001011010",
  23643=>"001100001",
  23644=>"010001000",
  23645=>"001011011",
  23646=>"001101000",
  23647=>"000000111",
  23648=>"110010001",
  23649=>"011011111",
  23650=>"100110100",
  23651=>"000111001",
  23652=>"000100000",
  23653=>"001000011",
  23654=>"110100000",
  23655=>"000000000",
  23656=>"111110101",
  23657=>"101110011",
  23658=>"000000001",
  23659=>"011011001",
  23660=>"101011010",
  23661=>"100000001",
  23662=>"010111100",
  23663=>"001111001",
  23664=>"001100000",
  23665=>"010110110",
  23666=>"100001111",
  23667=>"000010111",
  23668=>"011000010",
  23669=>"011010110",
  23670=>"010000101",
  23671=>"101111111",
  23672=>"001011100",
  23673=>"010101000",
  23674=>"000001100",
  23675=>"101000110",
  23676=>"000000110",
  23677=>"101101101",
  23678=>"010010000",
  23679=>"111000110",
  23680=>"000000000",
  23681=>"000110010",
  23682=>"000010000",
  23683=>"000010100",
  23684=>"000101000",
  23685=>"000000110",
  23686=>"111111000",
  23687=>"100101110",
  23688=>"101010010",
  23689=>"100011100",
  23690=>"011001111",
  23691=>"011110110",
  23692=>"110111010",
  23693=>"011111001",
  23694=>"001011110",
  23695=>"101001110",
  23696=>"001000000",
  23697=>"111100000",
  23698=>"001000011",
  23699=>"011100011",
  23700=>"101101011",
  23701=>"001110100",
  23702=>"000111100",
  23703=>"000000011",
  23704=>"000010001",
  23705=>"101001110",
  23706=>"010101100",
  23707=>"000111101",
  23708=>"000010111",
  23709=>"100001110",
  23710=>"111011011",
  23711=>"110101100",
  23712=>"011110111",
  23713=>"100111011",
  23714=>"001010010",
  23715=>"111110001",
  23716=>"101011000",
  23717=>"110010010",
  23718=>"011100011",
  23719=>"110100001",
  23720=>"110000101",
  23721=>"001011110",
  23722=>"000111110",
  23723=>"111110100",
  23724=>"001000111",
  23725=>"100011101",
  23726=>"000010110",
  23727=>"111011111",
  23728=>"000001010",
  23729=>"100001000",
  23730=>"000111011",
  23731=>"100100011",
  23732=>"110100100",
  23733=>"111011101",
  23734=>"000101000",
  23735=>"011111100",
  23736=>"001111110",
  23737=>"010111010",
  23738=>"100001101",
  23739=>"111101100",
  23740=>"010110100",
  23741=>"000000101",
  23742=>"100000011",
  23743=>"001001111",
  23744=>"111110010",
  23745=>"001100110",
  23746=>"000010000",
  23747=>"111000000",
  23748=>"101000100",
  23749=>"001101100",
  23750=>"001001010",
  23751=>"110010110",
  23752=>"111011001",
  23753=>"101000010",
  23754=>"101011111",
  23755=>"111110010",
  23756=>"111111010",
  23757=>"100100001",
  23758=>"000000000",
  23759=>"111011100",
  23760=>"001100100",
  23761=>"100111000",
  23762=>"011011110",
  23763=>"100101110",
  23764=>"111110111",
  23765=>"001100101",
  23766=>"000011110",
  23767=>"100101101",
  23768=>"010010011",
  23769=>"110011100",
  23770=>"100110111",
  23771=>"100001111",
  23772=>"001111100",
  23773=>"010100100",
  23774=>"000011001",
  23775=>"011111010",
  23776=>"101010111",
  23777=>"011001011",
  23778=>"100100101",
  23779=>"000000110",
  23780=>"011101001",
  23781=>"000001000",
  23782=>"000010101",
  23783=>"010111010",
  23784=>"100101000",
  23785=>"011011011",
  23786=>"100111000",
  23787=>"100000111",
  23788=>"001001111",
  23789=>"100100111",
  23790=>"111010010",
  23791=>"000100000",
  23792=>"001101000",
  23793=>"001010000",
  23794=>"000110110",
  23795=>"011000011",
  23796=>"000000000",
  23797=>"110000010",
  23798=>"001111101",
  23799=>"000011000",
  23800=>"001010011",
  23801=>"100101100",
  23802=>"001010110",
  23803=>"000010011",
  23804=>"101011011",
  23805=>"100111000",
  23806=>"111110100",
  23807=>"111100100",
  23808=>"111000010",
  23809=>"100110011",
  23810=>"001000110",
  23811=>"000110101",
  23812=>"100010101",
  23813=>"101100111",
  23814=>"100011110",
  23815=>"110011100",
  23816=>"100110000",
  23817=>"100000001",
  23818=>"110111010",
  23819=>"100000000",
  23820=>"001101100",
  23821=>"000000101",
  23822=>"100011100",
  23823=>"100110110",
  23824=>"011010110",
  23825=>"101001101",
  23826=>"111010100",
  23827=>"111110001",
  23828=>"010111111",
  23829=>"011101100",
  23830=>"011000100",
  23831=>"010111011",
  23832=>"011010011",
  23833=>"111011000",
  23834=>"110101101",
  23835=>"111100001",
  23836=>"001100000",
  23837=>"010000100",
  23838=>"100110110",
  23839=>"110111011",
  23840=>"110110011",
  23841=>"011101111",
  23842=>"000001011",
  23843=>"001001001",
  23844=>"000101000",
  23845=>"000001101",
  23846=>"111010110",
  23847=>"100001101",
  23848=>"110100000",
  23849=>"100011111",
  23850=>"110110011",
  23851=>"011100100",
  23852=>"111111010",
  23853=>"010100101",
  23854=>"101000011",
  23855=>"100001100",
  23856=>"100011000",
  23857=>"111111100",
  23858=>"011000010",
  23859=>"100011010",
  23860=>"001011110",
  23861=>"100100011",
  23862=>"100001100",
  23863=>"101100110",
  23864=>"000000000",
  23865=>"101100101",
  23866=>"100110101",
  23867=>"100110111",
  23868=>"010010111",
  23869=>"011101100",
  23870=>"101111110",
  23871=>"101111111",
  23872=>"010111001",
  23873=>"000000000",
  23874=>"101100011",
  23875=>"111000010",
  23876=>"000111001",
  23877=>"100001111",
  23878=>"011000000",
  23879=>"100100001",
  23880=>"001001101",
  23881=>"000100000",
  23882=>"100100010",
  23883=>"001000000",
  23884=>"001001100",
  23885=>"111010000",
  23886=>"001100101",
  23887=>"011111010",
  23888=>"000011011",
  23889=>"001101010",
  23890=>"110011000",
  23891=>"001000010",
  23892=>"000100000",
  23893=>"010000000",
  23894=>"010010001",
  23895=>"110111000",
  23896=>"000111100",
  23897=>"101101111",
  23898=>"000111010",
  23899=>"110101111",
  23900=>"110010111",
  23901=>"100111111",
  23902=>"011010101",
  23903=>"000011111",
  23904=>"010101000",
  23905=>"111010000",
  23906=>"010101010",
  23907=>"000111000",
  23908=>"100001111",
  23909=>"010000101",
  23910=>"101100001",
  23911=>"101100000",
  23912=>"000011110",
  23913=>"100110111",
  23914=>"011110010",
  23915=>"000111111",
  23916=>"111110001",
  23917=>"100000010",
  23918=>"010000010",
  23919=>"011001000",
  23920=>"000011001",
  23921=>"000000011",
  23922=>"101110111",
  23923=>"111001101",
  23924=>"011010001",
  23925=>"110101000",
  23926=>"010000001",
  23927=>"110101101",
  23928=>"110011101",
  23929=>"001111000",
  23930=>"000001011",
  23931=>"001111000",
  23932=>"010101101",
  23933=>"101111010",
  23934=>"110011010",
  23935=>"110010111",
  23936=>"011101110",
  23937=>"010101101",
  23938=>"000100000",
  23939=>"110010010",
  23940=>"010100110",
  23941=>"111101101",
  23942=>"000101111",
  23943=>"011001111",
  23944=>"111000001",
  23945=>"001000000",
  23946=>"001100000",
  23947=>"000010111",
  23948=>"011101110",
  23949=>"010100010",
  23950=>"101111000",
  23951=>"001010111",
  23952=>"100010110",
  23953=>"100000001",
  23954=>"100011110",
  23955=>"111000100",
  23956=>"111010010",
  23957=>"100111011",
  23958=>"100111100",
  23959=>"111010111",
  23960=>"101100011",
  23961=>"000101101",
  23962=>"110010111",
  23963=>"100111111",
  23964=>"101100011",
  23965=>"011010010",
  23966=>"011001001",
  23967=>"011111101",
  23968=>"111101100",
  23969=>"000111010",
  23970=>"000000001",
  23971=>"000010000",
  23972=>"110100100",
  23973=>"011011000",
  23974=>"110100000",
  23975=>"011011101",
  23976=>"010001111",
  23977=>"001001111",
  23978=>"010111000",
  23979=>"110110100",
  23980=>"111100100",
  23981=>"000011001",
  23982=>"100000000",
  23983=>"100110110",
  23984=>"001010110",
  23985=>"000111100",
  23986=>"010000010",
  23987=>"010111100",
  23988=>"011001111",
  23989=>"010110010",
  23990=>"001011010",
  23991=>"000110011",
  23992=>"111100010",
  23993=>"000010010",
  23994=>"000000010",
  23995=>"000001111",
  23996=>"011011000",
  23997=>"101100110",
  23998=>"100011101",
  23999=>"000100110",
  24000=>"010011000",
  24001=>"000111001",
  24002=>"100000100",
  24003=>"111011101",
  24004=>"010101001",
  24005=>"000010010",
  24006=>"000000010",
  24007=>"001100101",
  24008=>"001010011",
  24009=>"110010101",
  24010=>"010010000",
  24011=>"100111100",
  24012=>"111011111",
  24013=>"111010000",
  24014=>"000101111",
  24015=>"111101110",
  24016=>"110001010",
  24017=>"001100000",
  24018=>"001100010",
  24019=>"011110111",
  24020=>"110011110",
  24021=>"001100100",
  24022=>"110000010",
  24023=>"110000111",
  24024=>"000110111",
  24025=>"101011011",
  24026=>"111101001",
  24027=>"000101010",
  24028=>"111111010",
  24029=>"001010111",
  24030=>"010110111",
  24031=>"101000111",
  24032=>"110111000",
  24033=>"110110101",
  24034=>"001100000",
  24035=>"101001111",
  24036=>"011001100",
  24037=>"111110000",
  24038=>"110001001",
  24039=>"010000010",
  24040=>"110111100",
  24041=>"101100100",
  24042=>"000100001",
  24043=>"101101110",
  24044=>"011101011",
  24045=>"000111001",
  24046=>"110110100",
  24047=>"001110001",
  24048=>"100100110",
  24049=>"111111011",
  24050=>"100010101",
  24051=>"101001100",
  24052=>"001011110",
  24053=>"000001111",
  24054=>"101000110",
  24055=>"101101111",
  24056=>"001110001",
  24057=>"110001001",
  24058=>"000111010",
  24059=>"001101001",
  24060=>"000110000",
  24061=>"101101110",
  24062=>"101101010",
  24063=>"100110010",
  24064=>"110100010",
  24065=>"111001110",
  24066=>"110110001",
  24067=>"011000100",
  24068=>"100101010",
  24069=>"101111110",
  24070=>"011101111",
  24071=>"011110001",
  24072=>"001000001",
  24073=>"101101011",
  24074=>"001000101",
  24075=>"001100100",
  24076=>"110110111",
  24077=>"000001100",
  24078=>"111011000",
  24079=>"011100000",
  24080=>"100101100",
  24081=>"101010010",
  24082=>"101100101",
  24083=>"100010001",
  24084=>"000100100",
  24085=>"010010001",
  24086=>"111011111",
  24087=>"101010010",
  24088=>"001000011",
  24089=>"010110011",
  24090=>"000101101",
  24091=>"111010011",
  24092=>"111000011",
  24093=>"100001111",
  24094=>"000100000",
  24095=>"111001010",
  24096=>"101011101",
  24097=>"111010101",
  24098=>"000011011",
  24099=>"010000110",
  24100=>"110100011",
  24101=>"111010011",
  24102=>"001101000",
  24103=>"111101010",
  24104=>"000011111",
  24105=>"111101000",
  24106=>"101101101",
  24107=>"101111011",
  24108=>"110010011",
  24109=>"111001100",
  24110=>"000111000",
  24111=>"000100011",
  24112=>"101000101",
  24113=>"111100111",
  24114=>"110111110",
  24115=>"100110010",
  24116=>"000011000",
  24117=>"001100010",
  24118=>"110110011",
  24119=>"011000100",
  24120=>"101101000",
  24121=>"101001000",
  24122=>"101001011",
  24123=>"101110000",
  24124=>"011011110",
  24125=>"100010100",
  24126=>"111000011",
  24127=>"100101100",
  24128=>"101110001",
  24129=>"110011111",
  24130=>"000101001",
  24131=>"010100110",
  24132=>"000010011",
  24133=>"011111010",
  24134=>"110110010",
  24135=>"010110001",
  24136=>"001001100",
  24137=>"100100000",
  24138=>"001110100",
  24139=>"100111100",
  24140=>"011110011",
  24141=>"011100011",
  24142=>"010111101",
  24143=>"111001100",
  24144=>"011100110",
  24145=>"110111000",
  24146=>"101010001",
  24147=>"100100111",
  24148=>"011000100",
  24149=>"000111000",
  24150=>"000000000",
  24151=>"010100111",
  24152=>"100000110",
  24153=>"010111111",
  24154=>"000100000",
  24155=>"000001011",
  24156=>"011111100",
  24157=>"000011111",
  24158=>"101001010",
  24159=>"000101110",
  24160=>"011111100",
  24161=>"001110110",
  24162=>"001100100",
  24163=>"010100111",
  24164=>"011011010",
  24165=>"110100111",
  24166=>"110001110",
  24167=>"010011001",
  24168=>"000100001",
  24169=>"110010110",
  24170=>"001111101",
  24171=>"011100001",
  24172=>"101011100",
  24173=>"110101110",
  24174=>"101011001",
  24175=>"101101001",
  24176=>"000010100",
  24177=>"001100100",
  24178=>"111101010",
  24179=>"111111100",
  24180=>"100001001",
  24181=>"010111000",
  24182=>"000001110",
  24183=>"010000111",
  24184=>"111011000",
  24185=>"010111111",
  24186=>"001000101",
  24187=>"011100100",
  24188=>"001000111",
  24189=>"111011110",
  24190=>"010010100",
  24191=>"001111100",
  24192=>"110101010",
  24193=>"010111111",
  24194=>"110001100",
  24195=>"000100101",
  24196=>"000111001",
  24197=>"010111010",
  24198=>"111100101",
  24199=>"010101001",
  24200=>"011111000",
  24201=>"110000011",
  24202=>"010011010",
  24203=>"011100010",
  24204=>"011000100",
  24205=>"011011010",
  24206=>"110010000",
  24207=>"110001110",
  24208=>"110001100",
  24209=>"111101010",
  24210=>"000000000",
  24211=>"000111100",
  24212=>"010000001",
  24213=>"010111101",
  24214=>"100010000",
  24215=>"000010111",
  24216=>"111000110",
  24217=>"111001001",
  24218=>"000001111",
  24219=>"100110110",
  24220=>"111001101",
  24221=>"111110011",
  24222=>"010111010",
  24223=>"001101011",
  24224=>"111001010",
  24225=>"111011010",
  24226=>"101100111",
  24227=>"011100111",
  24228=>"111101111",
  24229=>"100110101",
  24230=>"100111010",
  24231=>"001000001",
  24232=>"010001000",
  24233=>"101000100",
  24234=>"110111011",
  24235=>"101010101",
  24236=>"000100110",
  24237=>"101100010",
  24238=>"110110100",
  24239=>"011110100",
  24240=>"000001011",
  24241=>"111011000",
  24242=>"100100001",
  24243=>"100101011",
  24244=>"101111110",
  24245=>"010110011",
  24246=>"101111110",
  24247=>"111011110",
  24248=>"000110011",
  24249=>"000011100",
  24250=>"101101110",
  24251=>"111001111",
  24252=>"101111010",
  24253=>"111010101",
  24254=>"100000111",
  24255=>"010011110",
  24256=>"111011011",
  24257=>"011101011",
  24258=>"100010111",
  24259=>"011001000",
  24260=>"000110001",
  24261=>"110100111",
  24262=>"011000101",
  24263=>"000101111",
  24264=>"111111000",
  24265=>"111110000",
  24266=>"101111001",
  24267=>"100000000",
  24268=>"100111110",
  24269=>"001100010",
  24270=>"111111001",
  24271=>"000010010",
  24272=>"000001011",
  24273=>"001101010",
  24274=>"001001111",
  24275=>"000101111",
  24276=>"011011111",
  24277=>"000111011",
  24278=>"100101000",
  24279=>"010001000",
  24280=>"100100000",
  24281=>"101100011",
  24282=>"001011101",
  24283=>"110100011",
  24284=>"111110111",
  24285=>"110001000",
  24286=>"000111010",
  24287=>"010001001",
  24288=>"010000010",
  24289=>"000000100",
  24290=>"111010001",
  24291=>"001110011",
  24292=>"001000110",
  24293=>"011010010",
  24294=>"100000110",
  24295=>"000100111",
  24296=>"001001111",
  24297=>"111101011",
  24298=>"111111110",
  24299=>"001000001",
  24300=>"000100101",
  24301=>"001010110",
  24302=>"111110110",
  24303=>"101000110",
  24304=>"100101010",
  24305=>"110101101",
  24306=>"100000011",
  24307=>"111101100",
  24308=>"000101110",
  24309=>"101001101",
  24310=>"110101010",
  24311=>"110001110",
  24312=>"011101000",
  24313=>"010110011",
  24314=>"010001111",
  24315=>"101100101",
  24316=>"100110000",
  24317=>"011010011",
  24318=>"010001100",
  24319=>"010101101",
  24320=>"000111010",
  24321=>"100110000",
  24322=>"000110000",
  24323=>"001001101",
  24324=>"111111011",
  24325=>"000101001",
  24326=>"001100111",
  24327=>"110110011",
  24328=>"110100011",
  24329=>"101010100",
  24330=>"110101101",
  24331=>"110010001",
  24332=>"000001101",
  24333=>"110000000",
  24334=>"011110001",
  24335=>"110101001",
  24336=>"100001100",
  24337=>"110010001",
  24338=>"111011001",
  24339=>"111111111",
  24340=>"100001111",
  24341=>"110100000",
  24342=>"011110001",
  24343=>"111000101",
  24344=>"001010111",
  24345=>"100010101",
  24346=>"000110100",
  24347=>"010010100",
  24348=>"001000000",
  24349=>"101001100",
  24350=>"101000000",
  24351=>"110101100",
  24352=>"100101000",
  24353=>"011001010",
  24354=>"010100101",
  24355=>"001001111",
  24356=>"101001010",
  24357=>"111001010",
  24358=>"100111111",
  24359=>"010111101",
  24360=>"101101101",
  24361=>"111011000",
  24362=>"100101011",
  24363=>"111100110",
  24364=>"011100100",
  24365=>"010101101",
  24366=>"100110010",
  24367=>"100101000",
  24368=>"000000110",
  24369=>"110010100",
  24370=>"010100001",
  24371=>"000011000",
  24372=>"110111101",
  24373=>"010000001",
  24374=>"000000110",
  24375=>"011000101",
  24376=>"011001000",
  24377=>"111001011",
  24378=>"101000111",
  24379=>"101111111",
  24380=>"000001110",
  24381=>"001001100",
  24382=>"000000111",
  24383=>"101111100",
  24384=>"000001011",
  24385=>"111010010",
  24386=>"110111000",
  24387=>"100011000",
  24388=>"110111111",
  24389=>"111011000",
  24390=>"100001001",
  24391=>"100011000",
  24392=>"011111010",
  24393=>"110011010",
  24394=>"111110101",
  24395=>"001111010",
  24396=>"111011011",
  24397=>"111011011",
  24398=>"111000010",
  24399=>"000000000",
  24400=>"011001011",
  24401=>"010100011",
  24402=>"111101111",
  24403=>"101110100",
  24404=>"110011000",
  24405=>"011001101",
  24406=>"000000110",
  24407=>"011111010",
  24408=>"001110101",
  24409=>"010100100",
  24410=>"001101011",
  24411=>"101000010",
  24412=>"100001110",
  24413=>"110100111",
  24414=>"101101000",
  24415=>"110100000",
  24416=>"101100001",
  24417=>"100111001",
  24418=>"000100111",
  24419=>"010111000",
  24420=>"110000101",
  24421=>"001111011",
  24422=>"110110011",
  24423=>"111011101",
  24424=>"111000011",
  24425=>"101111110",
  24426=>"010111101",
  24427=>"011011001",
  24428=>"111101101",
  24429=>"100011000",
  24430=>"010001011",
  24431=>"111110011",
  24432=>"001101010",
  24433=>"000100111",
  24434=>"100000100",
  24435=>"111111110",
  24436=>"011011000",
  24437=>"011110011",
  24438=>"011110001",
  24439=>"010001000",
  24440=>"011111000",
  24441=>"100111000",
  24442=>"111110001",
  24443=>"000110001",
  24444=>"000000000",
  24445=>"011010011",
  24446=>"010111000",
  24447=>"010110101",
  24448=>"011101010",
  24449=>"111101101",
  24450=>"000001000",
  24451=>"011000001",
  24452=>"100000010",
  24453=>"110110101",
  24454=>"011001001",
  24455=>"101010110",
  24456=>"101011111",
  24457=>"100000010",
  24458=>"110111100",
  24459=>"010110110",
  24460=>"101011101",
  24461=>"011011000",
  24462=>"100000111",
  24463=>"011101010",
  24464=>"011110001",
  24465=>"010000011",
  24466=>"100000000",
  24467=>"110000011",
  24468=>"101000000",
  24469=>"001110011",
  24470=>"010110100",
  24471=>"000010111",
  24472=>"010111101",
  24473=>"110010001",
  24474=>"100110101",
  24475=>"001010100",
  24476=>"110111111",
  24477=>"001110111",
  24478=>"010001110",
  24479=>"000000100",
  24480=>"100001111",
  24481=>"010111110",
  24482=>"010101110",
  24483=>"000100100",
  24484=>"000000110",
  24485=>"101111101",
  24486=>"100101001",
  24487=>"011101100",
  24488=>"011110010",
  24489=>"000111000",
  24490=>"000110101",
  24491=>"111100100",
  24492=>"110110010",
  24493=>"101001000",
  24494=>"000000110",
  24495=>"001101111",
  24496=>"001000100",
  24497=>"111010110",
  24498=>"000101011",
  24499=>"001100110",
  24500=>"111000101",
  24501=>"010000111",
  24502=>"001001000",
  24503=>"110101001",
  24504=>"100000010",
  24505=>"111011001",
  24506=>"110001010",
  24507=>"010101010",
  24508=>"011010000",
  24509=>"101101111",
  24510=>"100000000",
  24511=>"101101110",
  24512=>"110111100",
  24513=>"001101010",
  24514=>"010111110",
  24515=>"101011111",
  24516=>"100111001",
  24517=>"110100111",
  24518=>"001010000",
  24519=>"110011010",
  24520=>"101011111",
  24521=>"100001000",
  24522=>"000000001",
  24523=>"011101011",
  24524=>"110110011",
  24525=>"000000110",
  24526=>"101000010",
  24527=>"111011110",
  24528=>"000010011",
  24529=>"010100011",
  24530=>"110010101",
  24531=>"100101100",
  24532=>"000111010",
  24533=>"100100111",
  24534=>"000000111",
  24535=>"010100010",
  24536=>"001110100",
  24537=>"101110110",
  24538=>"010010000",
  24539=>"000110001",
  24540=>"110111100",
  24541=>"100101100",
  24542=>"110010001",
  24543=>"010001010",
  24544=>"001000100",
  24545=>"001111100",
  24546=>"000101101",
  24547=>"111001011",
  24548=>"001110100",
  24549=>"001100000",
  24550=>"000011000",
  24551=>"011000010",
  24552=>"110101100",
  24553=>"100011011",
  24554=>"011000011",
  24555=>"000100110",
  24556=>"100101000",
  24557=>"101001011",
  24558=>"011000111",
  24559=>"011101001",
  24560=>"100010101",
  24561=>"000010110",
  24562=>"001100011",
  24563=>"001010010",
  24564=>"110001000",
  24565=>"000111101",
  24566=>"011101001",
  24567=>"111101001",
  24568=>"110010001",
  24569=>"110100010",
  24570=>"010101000",
  24571=>"011100100",
  24572=>"010100000",
  24573=>"000010011",
  24574=>"001000011",
  24575=>"010011010",
  24576=>"100000111",
  24577=>"110001001",
  24578=>"010010001",
  24579=>"111111000",
  24580=>"011011001",
  24581=>"100011101",
  24582=>"111101000",
  24583=>"100100100",
  24584=>"110001100",
  24585=>"110111000",
  24586=>"010111101",
  24587=>"010001001",
  24588=>"111011100",
  24589=>"101110000",
  24590=>"001110111",
  24591=>"101001010",
  24592=>"111001101",
  24593=>"000101001",
  24594=>"101101110",
  24595=>"011000100",
  24596=>"111000110",
  24597=>"101001111",
  24598=>"100100101",
  24599=>"110000011",
  24600=>"000101110",
  24601=>"001000110",
  24602=>"101000000",
  24603=>"010101111",
  24604=>"000011001",
  24605=>"111010110",
  24606=>"101111101",
  24607=>"011010101",
  24608=>"111011000",
  24609=>"011100100",
  24610=>"011000110",
  24611=>"110101011",
  24612=>"111100111",
  24613=>"101011101",
  24614=>"010010100",
  24615=>"100001011",
  24616=>"001000000",
  24617=>"100101010",
  24618=>"001101101",
  24619=>"001010100",
  24620=>"000001000",
  24621=>"001100000",
  24622=>"011001101",
  24623=>"001000101",
  24624=>"011010011",
  24625=>"101111011",
  24626=>"011110100",
  24627=>"100110000",
  24628=>"100010111",
  24629=>"011101111",
  24630=>"101001100",
  24631=>"000101101",
  24632=>"000001001",
  24633=>"101000101",
  24634=>"101000000",
  24635=>"011101100",
  24636=>"101101001",
  24637=>"100110011",
  24638=>"100000100",
  24639=>"101010110",
  24640=>"100100110",
  24641=>"110111111",
  24642=>"000100110",
  24643=>"011100000",
  24644=>"101111000",
  24645=>"111010011",
  24646=>"110111100",
  24647=>"010000100",
  24648=>"101010111",
  24649=>"111110110",
  24650=>"111110101",
  24651=>"001010111",
  24652=>"011111011",
  24653=>"111000111",
  24654=>"110110101",
  24655=>"111111010",
  24656=>"010011111",
  24657=>"001011010",
  24658=>"010010100",
  24659=>"110001000",
  24660=>"111100100",
  24661=>"001111110",
  24662=>"011000100",
  24663=>"000101001",
  24664=>"001000011",
  24665=>"110101010",
  24666=>"100111000",
  24667=>"000000011",
  24668=>"011101000",
  24669=>"001000110",
  24670=>"100110001",
  24671=>"100000001",
  24672=>"011111000",
  24673=>"110100100",
  24674=>"000011100",
  24675=>"111000010",
  24676=>"000111011",
  24677=>"101011011",
  24678=>"001001100",
  24679=>"000101101",
  24680=>"000001000",
  24681=>"000111110",
  24682=>"110101011",
  24683=>"111010000",
  24684=>"100000101",
  24685=>"000011010",
  24686=>"001110110",
  24687=>"010111000",
  24688=>"011101001",
  24689=>"011111010",
  24690=>"010011101",
  24691=>"000100101",
  24692=>"111111011",
  24693=>"010100111",
  24694=>"100011110",
  24695=>"001100110",
  24696=>"011100010",
  24697=>"000010000",
  24698=>"010011011",
  24699=>"100100100",
  24700=>"110100100",
  24701=>"111000110",
  24702=>"010001100",
  24703=>"111010000",
  24704=>"101001111",
  24705=>"110100101",
  24706=>"011110000",
  24707=>"010111111",
  24708=>"000000100",
  24709=>"110100100",
  24710=>"001000100",
  24711=>"111000100",
  24712=>"110100001",
  24713=>"011110000",
  24714=>"100110100",
  24715=>"111010101",
  24716=>"101110100",
  24717=>"100000110",
  24718=>"100011111",
  24719=>"101000001",
  24720=>"110110010",
  24721=>"110100000",
  24722=>"001111000",
  24723=>"010001011",
  24724=>"100010010",
  24725=>"010010100",
  24726=>"111110000",
  24727=>"000110000",
  24728=>"010111011",
  24729=>"100101101",
  24730=>"101100001",
  24731=>"100011010",
  24732=>"010011001",
  24733=>"011011011",
  24734=>"000001010",
  24735=>"100000011",
  24736=>"100000000",
  24737=>"001010011",
  24738=>"110011100",
  24739=>"101001100",
  24740=>"111010001",
  24741=>"101100010",
  24742=>"110010100",
  24743=>"111010110",
  24744=>"001011100",
  24745=>"011111110",
  24746=>"000100101",
  24747=>"101100101",
  24748=>"110100011",
  24749=>"000111110",
  24750=>"011001000",
  24751=>"010000011",
  24752=>"010000010",
  24753=>"011010110",
  24754=>"110100000",
  24755=>"101010011",
  24756=>"001000010",
  24757=>"111101001",
  24758=>"011100000",
  24759=>"100010001",
  24760=>"011000001",
  24761=>"101110011",
  24762=>"111110110",
  24763=>"001100110",
  24764=>"111111001",
  24765=>"010111100",
  24766=>"000111011",
  24767=>"000100000",
  24768=>"011110011",
  24769=>"010111001",
  24770=>"101111001",
  24771=>"100101101",
  24772=>"000010101",
  24773=>"111000011",
  24774=>"111101110",
  24775=>"011110011",
  24776=>"000110110",
  24777=>"111111001",
  24778=>"111010101",
  24779=>"100111011",
  24780=>"000001110",
  24781=>"010011111",
  24782=>"101100001",
  24783=>"100010000",
  24784=>"111010010",
  24785=>"001100110",
  24786=>"110011010",
  24787=>"111000010",
  24788=>"110101001",
  24789=>"011111100",
  24790=>"101011100",
  24791=>"001001110",
  24792=>"000010001",
  24793=>"100111100",
  24794=>"101101011",
  24795=>"101111010",
  24796=>"011000100",
  24797=>"000010100",
  24798=>"100100001",
  24799=>"100010101",
  24800=>"010010000",
  24801=>"001100000",
  24802=>"011100111",
  24803=>"000001001",
  24804=>"010000100",
  24805=>"001110001",
  24806=>"110101101",
  24807=>"000010010",
  24808=>"110010101",
  24809=>"010101110",
  24810=>"100011110",
  24811=>"110001011",
  24812=>"110101100",
  24813=>"101111001",
  24814=>"100010001",
  24815=>"000101010",
  24816=>"110111110",
  24817=>"001111001",
  24818=>"111010110",
  24819=>"000000101",
  24820=>"011101111",
  24821=>"111000000",
  24822=>"111100011",
  24823=>"000011010",
  24824=>"101110100",
  24825=>"101110110",
  24826=>"111000011",
  24827=>"001101011",
  24828=>"101001111",
  24829=>"100010000",
  24830=>"001111100",
  24831=>"001000100",
  24832=>"110010100",
  24833=>"100001100",
  24834=>"110101100",
  24835=>"101001010",
  24836=>"101001110",
  24837=>"101110011",
  24838=>"000010000",
  24839=>"101100000",
  24840=>"001011101",
  24841=>"010001000",
  24842=>"001100110",
  24843=>"001001100",
  24844=>"101010110",
  24845=>"000011111",
  24846=>"100011111",
  24847=>"000001101",
  24848=>"001111110",
  24849=>"011000001",
  24850=>"001000110",
  24851=>"111001011",
  24852=>"110100101",
  24853=>"000001110",
  24854=>"001001111",
  24855=>"100000101",
  24856=>"110000101",
  24857=>"000001011",
  24858=>"000000001",
  24859=>"111011001",
  24860=>"110001000",
  24861=>"001101110",
  24862=>"000000100",
  24863=>"000001101",
  24864=>"010001110",
  24865=>"110101001",
  24866=>"101111111",
  24867=>"101011001",
  24868=>"001011011",
  24869=>"100010010",
  24870=>"111000000",
  24871=>"100100100",
  24872=>"010000010",
  24873=>"001001101",
  24874=>"011010000",
  24875=>"111100101",
  24876=>"001111011",
  24877=>"100010000",
  24878=>"111011101",
  24879=>"101110001",
  24880=>"000100100",
  24881=>"110101011",
  24882=>"001100110",
  24883=>"101101000",
  24884=>"000000101",
  24885=>"110001011",
  24886=>"011111101",
  24887=>"101110001",
  24888=>"000001111",
  24889=>"101101010",
  24890=>"010001001",
  24891=>"101111110",
  24892=>"100110100",
  24893=>"010001011",
  24894=>"001110111",
  24895=>"001011001",
  24896=>"100101001",
  24897=>"111111101",
  24898=>"110101011",
  24899=>"010101101",
  24900=>"000000011",
  24901=>"000110000",
  24902=>"001100001",
  24903=>"101010100",
  24904=>"100101100",
  24905=>"110001010",
  24906=>"101010011",
  24907=>"010100100",
  24908=>"101101001",
  24909=>"000100000",
  24910=>"010001010",
  24911=>"011001101",
  24912=>"000101101",
  24913=>"110101011",
  24914=>"101000101",
  24915=>"111101111",
  24916=>"101000011",
  24917=>"010010100",
  24918=>"010110000",
  24919=>"101010110",
  24920=>"000100100",
  24921=>"000000101",
  24922=>"100000101",
  24923=>"001101010",
  24924=>"011111101",
  24925=>"010010010",
  24926=>"011011011",
  24927=>"011000010",
  24928=>"010101100",
  24929=>"101010100",
  24930=>"000110110",
  24931=>"010011001",
  24932=>"000101001",
  24933=>"101010001",
  24934=>"010100101",
  24935=>"100110110",
  24936=>"001111011",
  24937=>"001111010",
  24938=>"000101011",
  24939=>"111111000",
  24940=>"010001000",
  24941=>"001000000",
  24942=>"000111000",
  24943=>"011101101",
  24944=>"010110110",
  24945=>"100101100",
  24946=>"011110101",
  24947=>"011000011",
  24948=>"000010111",
  24949=>"000110010",
  24950=>"100010100",
  24951=>"010101000",
  24952=>"110101010",
  24953=>"000011100",
  24954=>"101000000",
  24955=>"101000111",
  24956=>"010100110",
  24957=>"000110001",
  24958=>"011111001",
  24959=>"111111111",
  24960=>"000010010",
  24961=>"111000111",
  24962=>"101111111",
  24963=>"101000101",
  24964=>"011100000",
  24965=>"100010000",
  24966=>"101001111",
  24967=>"110101000",
  24968=>"101001010",
  24969=>"101100101",
  24970=>"001001011",
  24971=>"001010100",
  24972=>"100000000",
  24973=>"011001101",
  24974=>"000000100",
  24975=>"000101110",
  24976=>"110100000",
  24977=>"000100011",
  24978=>"100011101",
  24979=>"111111011",
  24980=>"100100111",
  24981=>"010111010",
  24982=>"001001000",
  24983=>"110100100",
  24984=>"000101001",
  24985=>"100111010",
  24986=>"111110000",
  24987=>"001101000",
  24988=>"100010100",
  24989=>"111111011",
  24990=>"000111011",
  24991=>"011101111",
  24992=>"010011010",
  24993=>"010100000",
  24994=>"110010011",
  24995=>"100000101",
  24996=>"111111110",
  24997=>"000101111",
  24998=>"010111110",
  24999=>"111110011",
  25000=>"101101101",
  25001=>"101001100",
  25002=>"011111101",
  25003=>"100110100",
  25004=>"111001111",
  25005=>"001110100",
  25006=>"011111111",
  25007=>"000011110",
  25008=>"011110110",
  25009=>"100100010",
  25010=>"000001011",
  25011=>"101100100",
  25012=>"001001100",
  25013=>"101110111",
  25014=>"011110010",
  25015=>"000110000",
  25016=>"111110010",
  25017=>"010100111",
  25018=>"100100001",
  25019=>"011000111",
  25020=>"010001010",
  25021=>"111011000",
  25022=>"001010001",
  25023=>"010110000",
  25024=>"000000101",
  25025=>"101000101",
  25026=>"000100000",
  25027=>"000111010",
  25028=>"010101100",
  25029=>"001101001",
  25030=>"000111010",
  25031=>"001011001",
  25032=>"010110011",
  25033=>"110111111",
  25034=>"110101100",
  25035=>"010000110",
  25036=>"111100000",
  25037=>"101011011",
  25038=>"110100000",
  25039=>"101111010",
  25040=>"011001011",
  25041=>"001011011",
  25042=>"100110100",
  25043=>"110111101",
  25044=>"110010010",
  25045=>"101101011",
  25046=>"111100000",
  25047=>"111100110",
  25048=>"010111011",
  25049=>"111000001",
  25050=>"001101111",
  25051=>"000010110",
  25052=>"011111001",
  25053=>"001111111",
  25054=>"010111110",
  25055=>"111001000",
  25056=>"100011100",
  25057=>"100001100",
  25058=>"011111110",
  25059=>"111101010",
  25060=>"110010101",
  25061=>"110000100",
  25062=>"011101001",
  25063=>"110000011",
  25064=>"101101000",
  25065=>"110000101",
  25066=>"000100000",
  25067=>"110001101",
  25068=>"101001111",
  25069=>"111110100",
  25070=>"011100100",
  25071=>"000011000",
  25072=>"101110101",
  25073=>"100100000",
  25074=>"010101000",
  25075=>"001101111",
  25076=>"110101001",
  25077=>"111111111",
  25078=>"010101001",
  25079=>"010011001",
  25080=>"110111101",
  25081=>"011001011",
  25082=>"101001000",
  25083=>"111100100",
  25084=>"000110111",
  25085=>"001001010",
  25086=>"111010011",
  25087=>"101100000",
  25088=>"110001101",
  25089=>"100100111",
  25090=>"010101100",
  25091=>"001001111",
  25092=>"010101101",
  25093=>"010011011",
  25094=>"010001010",
  25095=>"011111101",
  25096=>"010111011",
  25097=>"101100111",
  25098=>"000010011",
  25099=>"100111110",
  25100=>"001001100",
  25101=>"000101010",
  25102=>"001011000",
  25103=>"000101010",
  25104=>"000110011",
  25105=>"101011101",
  25106=>"111011000",
  25107=>"100101001",
  25108=>"101101100",
  25109=>"000110100",
  25110=>"111101110",
  25111=>"100110011",
  25112=>"101001101",
  25113=>"110110100",
  25114=>"000000101",
  25115=>"001101110",
  25116=>"100000101",
  25117=>"110001000",
  25118=>"000011010",
  25119=>"101110010",
  25120=>"111001101",
  25121=>"111101010",
  25122=>"111000100",
  25123=>"111100010",
  25124=>"101111011",
  25125=>"110010010",
  25126=>"001000110",
  25127=>"100010000",
  25128=>"111110000",
  25129=>"001000001",
  25130=>"111101001",
  25131=>"110100110",
  25132=>"110010101",
  25133=>"000111100",
  25134=>"011000101",
  25135=>"010000010",
  25136=>"001010011",
  25137=>"001010101",
  25138=>"011100101",
  25139=>"000111010",
  25140=>"000010100",
  25141=>"000100110",
  25142=>"111101111",
  25143=>"111000001",
  25144=>"100010101",
  25145=>"011110011",
  25146=>"010111110",
  25147=>"100110111",
  25148=>"100001100",
  25149=>"000000100",
  25150=>"010111101",
  25151=>"011010101",
  25152=>"111111000",
  25153=>"001111100",
  25154=>"110101010",
  25155=>"011101111",
  25156=>"001101011",
  25157=>"101000111",
  25158=>"011000100",
  25159=>"010110111",
  25160=>"110011101",
  25161=>"101011011",
  25162=>"001110110",
  25163=>"000101111",
  25164=>"110000111",
  25165=>"010011101",
  25166=>"000101111",
  25167=>"110000000",
  25168=>"101111110",
  25169=>"100111111",
  25170=>"000001110",
  25171=>"000101111",
  25172=>"000001000",
  25173=>"110000100",
  25174=>"100111111",
  25175=>"100000110",
  25176=>"101011000",
  25177=>"010001010",
  25178=>"011101110",
  25179=>"001001001",
  25180=>"010001110",
  25181=>"011001111",
  25182=>"101000110",
  25183=>"101100101",
  25184=>"110110110",
  25185=>"111010110",
  25186=>"100000110",
  25187=>"010000101",
  25188=>"111111110",
  25189=>"110010001",
  25190=>"101100001",
  25191=>"011001001",
  25192=>"010000000",
  25193=>"110100000",
  25194=>"111101101",
  25195=>"111001100",
  25196=>"100100110",
  25197=>"001100110",
  25198=>"011000001",
  25199=>"111010011",
  25200=>"000101001",
  25201=>"011100100",
  25202=>"001101111",
  25203=>"010110010",
  25204=>"011000100",
  25205=>"010100011",
  25206=>"110111111",
  25207=>"010000101",
  25208=>"111001111",
  25209=>"001010011",
  25210=>"011000101",
  25211=>"101000011",
  25212=>"000111110",
  25213=>"101110000",
  25214=>"010110100",
  25215=>"000110101",
  25216=>"011011001",
  25217=>"111011010",
  25218=>"100111100",
  25219=>"011101000",
  25220=>"111100010",
  25221=>"110101000",
  25222=>"010010010",
  25223=>"101000101",
  25224=>"011001100",
  25225=>"011010101",
  25226=>"100011101",
  25227=>"110111101",
  25228=>"010111011",
  25229=>"001100000",
  25230=>"110010001",
  25231=>"010011110",
  25232=>"011010111",
  25233=>"011011101",
  25234=>"110111111",
  25235=>"000011011",
  25236=>"110110001",
  25237=>"000011011",
  25238=>"101110101",
  25239=>"111100110",
  25240=>"001011000",
  25241=>"001100111",
  25242=>"101000011",
  25243=>"011110010",
  25244=>"100011001",
  25245=>"011010101",
  25246=>"000110111",
  25247=>"001101100",
  25248=>"011001100",
  25249=>"011101001",
  25250=>"110001110",
  25251=>"111000110",
  25252=>"000010011",
  25253=>"001110011",
  25254=>"100100101",
  25255=>"100001111",
  25256=>"011101010",
  25257=>"101010111",
  25258=>"100100110",
  25259=>"100100000",
  25260=>"010000000",
  25261=>"100001011",
  25262=>"111001100",
  25263=>"000100000",
  25264=>"111111001",
  25265=>"111000000",
  25266=>"000011101",
  25267=>"101001000",
  25268=>"100110010",
  25269=>"111110001",
  25270=>"000100111",
  25271=>"001100000",
  25272=>"011101100",
  25273=>"111100100",
  25274=>"011100101",
  25275=>"010010001",
  25276=>"100010000",
  25277=>"000100001",
  25278=>"111001110",
  25279=>"110100110",
  25280=>"011011101",
  25281=>"110101110",
  25282=>"011110100",
  25283=>"001001011",
  25284=>"101100110",
  25285=>"101101111",
  25286=>"000101111",
  25287=>"011000001",
  25288=>"001001000",
  25289=>"111100101",
  25290=>"110111010",
  25291=>"001000010",
  25292=>"011111111",
  25293=>"101010101",
  25294=>"000000000",
  25295=>"010111010",
  25296=>"101010001",
  25297=>"000000010",
  25298=>"111000011",
  25299=>"011110010",
  25300=>"110111110",
  25301=>"001101101",
  25302=>"001011101",
  25303=>"001000110",
  25304=>"010011101",
  25305=>"111010011",
  25306=>"011000001",
  25307=>"011010101",
  25308=>"010100100",
  25309=>"100010000",
  25310=>"101010100",
  25311=>"000011000",
  25312=>"110101001",
  25313=>"000101010",
  25314=>"101010111",
  25315=>"011011101",
  25316=>"110010000",
  25317=>"110011011",
  25318=>"010010001",
  25319=>"000011111",
  25320=>"000100101",
  25321=>"001001111",
  25322=>"101111001",
  25323=>"011111011",
  25324=>"000100001",
  25325=>"101001011",
  25326=>"001101011",
  25327=>"100011001",
  25328=>"101000011",
  25329=>"011101111",
  25330=>"001110011",
  25331=>"101111011",
  25332=>"110010010",
  25333=>"100111010",
  25334=>"110111000",
  25335=>"000000111",
  25336=>"111011010",
  25337=>"111001010",
  25338=>"010101000",
  25339=>"011011111",
  25340=>"110110110",
  25341=>"000011100",
  25342=>"011101010",
  25343=>"001101101",
  25344=>"111011000",
  25345=>"010101010",
  25346=>"011011001",
  25347=>"011101101",
  25348=>"011101110",
  25349=>"101101111",
  25350=>"111010010",
  25351=>"001100101",
  25352=>"000111010",
  25353=>"101011001",
  25354=>"111111100",
  25355=>"110001110",
  25356=>"101100100",
  25357=>"110000101",
  25358=>"011111001",
  25359=>"101011110",
  25360=>"000110101",
  25361=>"010000001",
  25362=>"100110111",
  25363=>"010001110",
  25364=>"000010010",
  25365=>"011011010",
  25366=>"000000110",
  25367=>"010001000",
  25368=>"110100000",
  25369=>"101011100",
  25370=>"101001111",
  25371=>"000101101",
  25372=>"110101010",
  25373=>"111100111",
  25374=>"011011100",
  25375=>"101110101",
  25376=>"100001100",
  25377=>"110101111",
  25378=>"100100001",
  25379=>"000111000",
  25380=>"010011100",
  25381=>"011000001",
  25382=>"010011110",
  25383=>"000100111",
  25384=>"001111000",
  25385=>"001010000",
  25386=>"111010000",
  25387=>"001010100",
  25388=>"000000100",
  25389=>"100101101",
  25390=>"110000000",
  25391=>"010000101",
  25392=>"000010011",
  25393=>"110001010",
  25394=>"111000110",
  25395=>"001001000",
  25396=>"010101100",
  25397=>"110011000",
  25398=>"110001010",
  25399=>"000000001",
  25400=>"000100001",
  25401=>"011111010",
  25402=>"010011110",
  25403=>"000001101",
  25404=>"111000001",
  25405=>"011011110",
  25406=>"010100010",
  25407=>"100010001",
  25408=>"011000010",
  25409=>"110001110",
  25410=>"101000010",
  25411=>"111001011",
  25412=>"100100110",
  25413=>"100000100",
  25414=>"011001111",
  25415=>"010010110",
  25416=>"111011010",
  25417=>"110011010",
  25418=>"111011000",
  25419=>"110101100",
  25420=>"110101110",
  25421=>"100101101",
  25422=>"000100100",
  25423=>"111000001",
  25424=>"100001001",
  25425=>"010001100",
  25426=>"000110011",
  25427=>"100000100",
  25428=>"110110110",
  25429=>"000010110",
  25430=>"000110000",
  25431=>"001110101",
  25432=>"011011101",
  25433=>"110110010",
  25434=>"001101000",
  25435=>"000001101",
  25436=>"010111011",
  25437=>"111101111",
  25438=>"110000111",
  25439=>"000010011",
  25440=>"011000010",
  25441=>"100010110",
  25442=>"001010011",
  25443=>"011110100",
  25444=>"100010000",
  25445=>"000100101",
  25446=>"101100000",
  25447=>"010110100",
  25448=>"110101010",
  25449=>"000000001",
  25450=>"000111101",
  25451=>"000010110",
  25452=>"100101000",
  25453=>"000100100",
  25454=>"111001011",
  25455=>"001111110",
  25456=>"010010111",
  25457=>"011001011",
  25458=>"110101011",
  25459=>"100110000",
  25460=>"111000001",
  25461=>"111101010",
  25462=>"111111101",
  25463=>"101101001",
  25464=>"010011110",
  25465=>"110111100",
  25466=>"010111110",
  25467=>"000010111",
  25468=>"110000001",
  25469=>"110000111",
  25470=>"001110101",
  25471=>"010100011",
  25472=>"110110110",
  25473=>"101110011",
  25474=>"000111111",
  25475=>"010101000",
  25476=>"010100100",
  25477=>"100111110",
  25478=>"101011000",
  25479=>"100010000",
  25480=>"100011011",
  25481=>"110000001",
  25482=>"011000110",
  25483=>"100011101",
  25484=>"101010100",
  25485=>"101000011",
  25486=>"101001101",
  25487=>"101110000",
  25488=>"010111101",
  25489=>"111111010",
  25490=>"010010000",
  25491=>"001010000",
  25492=>"001000110",
  25493=>"100111001",
  25494=>"100011111",
  25495=>"010010100",
  25496=>"000010010",
  25497=>"000110101",
  25498=>"111001011",
  25499=>"111111101",
  25500=>"111011000",
  25501=>"111101101",
  25502=>"011100111",
  25503=>"011100001",
  25504=>"100011111",
  25505=>"001010100",
  25506=>"110010010",
  25507=>"001110001",
  25508=>"101011000",
  25509=>"110000011",
  25510=>"011101101",
  25511=>"100110011",
  25512=>"110001000",
  25513=>"010100010",
  25514=>"000101111",
  25515=>"011101111",
  25516=>"000010000",
  25517=>"011110010",
  25518=>"110011000",
  25519=>"110100010",
  25520=>"010000000",
  25521=>"001100010",
  25522=>"101011010",
  25523=>"001101110",
  25524=>"010011101",
  25525=>"001101111",
  25526=>"110000111",
  25527=>"110110011",
  25528=>"110100101",
  25529=>"000110010",
  25530=>"010000011",
  25531=>"111011001",
  25532=>"110101110",
  25533=>"100000101",
  25534=>"111000000",
  25535=>"111111011",
  25536=>"110000010",
  25537=>"100110000",
  25538=>"111100001",
  25539=>"100001100",
  25540=>"101010111",
  25541=>"100011110",
  25542=>"010111000",
  25543=>"001011101",
  25544=>"110100010",
  25545=>"100110000",
  25546=>"010010000",
  25547=>"110110010",
  25548=>"011110000",
  25549=>"000101011",
  25550=>"010110000",
  25551=>"110001110",
  25552=>"011001001",
  25553=>"001011110",
  25554=>"000101101",
  25555=>"100000011",
  25556=>"100100110",
  25557=>"010101101",
  25558=>"110110001",
  25559=>"101110001",
  25560=>"111110110",
  25561=>"110100110",
  25562=>"010010111",
  25563=>"001000100",
  25564=>"101010000",
  25565=>"110100001",
  25566=>"101000011",
  25567=>"111111110",
  25568=>"000100000",
  25569=>"110000101",
  25570=>"100010011",
  25571=>"101000110",
  25572=>"101010000",
  25573=>"011100011",
  25574=>"010011110",
  25575=>"111000000",
  25576=>"010110011",
  25577=>"111010111",
  25578=>"111110001",
  25579=>"001101101",
  25580=>"100010101",
  25581=>"111101000",
  25582=>"000010001",
  25583=>"100101000",
  25584=>"000010001",
  25585=>"111100000",
  25586=>"011011101",
  25587=>"100000100",
  25588=>"110100100",
  25589=>"001011110",
  25590=>"100101101",
  25591=>"000001110",
  25592=>"010110011",
  25593=>"101100010",
  25594=>"010110000",
  25595=>"000101110",
  25596=>"100100010",
  25597=>"000101001",
  25598=>"000101111",
  25599=>"101010100",
  25600=>"110010010",
  25601=>"001001010",
  25602=>"111111100",
  25603=>"111100010",
  25604=>"010100000",
  25605=>"000000101",
  25606=>"111011110",
  25607=>"111001011",
  25608=>"001100011",
  25609=>"011000000",
  25610=>"111010100",
  25611=>"100110111",
  25612=>"010111011",
  25613=>"110110010",
  25614=>"110110000",
  25615=>"111001000",
  25616=>"010011001",
  25617=>"110100100",
  25618=>"000010010",
  25619=>"101011011",
  25620=>"001100010",
  25621=>"110111010",
  25622=>"000111101",
  25623=>"111011011",
  25624=>"111110001",
  25625=>"111001101",
  25626=>"110010110",
  25627=>"111101000",
  25628=>"001110101",
  25629=>"001000001",
  25630=>"100010100",
  25631=>"000000000",
  25632=>"101010000",
  25633=>"000001110",
  25634=>"101110111",
  25635=>"001110001",
  25636=>"000111110",
  25637=>"110010111",
  25638=>"101001010",
  25639=>"010000011",
  25640=>"011100101",
  25641=>"000101001",
  25642=>"011101011",
  25643=>"011010010",
  25644=>"000000100",
  25645=>"001111111",
  25646=>"000010100",
  25647=>"111101010",
  25648=>"010001011",
  25649=>"100100100",
  25650=>"001000101",
  25651=>"000111101",
  25652=>"101011010",
  25653=>"111010010",
  25654=>"111000011",
  25655=>"101001001",
  25656=>"101000011",
  25657=>"010000110",
  25658=>"100101011",
  25659=>"011100010",
  25660=>"101000100",
  25661=>"011100100",
  25662=>"001010011",
  25663=>"101000010",
  25664=>"111010001",
  25665=>"101000101",
  25666=>"011011000",
  25667=>"100101111",
  25668=>"110111010",
  25669=>"111100100",
  25670=>"011010111",
  25671=>"000001110",
  25672=>"000001111",
  25673=>"000101010",
  25674=>"101010000",
  25675=>"011010110",
  25676=>"110110111",
  25677=>"101010001",
  25678=>"011011000",
  25679=>"001111110",
  25680=>"001001101",
  25681=>"111101111",
  25682=>"011011001",
  25683=>"111010110",
  25684=>"100101101",
  25685=>"010011001",
  25686=>"101001000",
  25687=>"111111011",
  25688=>"101111010",
  25689=>"010111101",
  25690=>"001011011",
  25691=>"010101100",
  25692=>"010111111",
  25693=>"101110001",
  25694=>"011111010",
  25695=>"111001011",
  25696=>"010100010",
  25697=>"010000011",
  25698=>"100000000",
  25699=>"101001111",
  25700=>"100110000",
  25701=>"100000000",
  25702=>"111101110",
  25703=>"001000101",
  25704=>"010001111",
  25705=>"000101000",
  25706=>"011001010",
  25707=>"011010011",
  25708=>"111110010",
  25709=>"100100111",
  25710=>"111100001",
  25711=>"111110010",
  25712=>"111011000",
  25713=>"001111001",
  25714=>"110110001",
  25715=>"110100011",
  25716=>"000001000",
  25717=>"111101111",
  25718=>"111100011",
  25719=>"001001110",
  25720=>"010011000",
  25721=>"001101101",
  25722=>"011111111",
  25723=>"000010100",
  25724=>"100111101",
  25725=>"111010111",
  25726=>"111010001",
  25727=>"101101001",
  25728=>"111101110",
  25729=>"000001111",
  25730=>"110100000",
  25731=>"100000010",
  25732=>"000010111",
  25733=>"010000001",
  25734=>"110111011",
  25735=>"001001011",
  25736=>"101101010",
  25737=>"000001010",
  25738=>"100100001",
  25739=>"111001101",
  25740=>"000000111",
  25741=>"100000010",
  25742=>"110101100",
  25743=>"001011101",
  25744=>"010110000",
  25745=>"000001110",
  25746=>"110101000",
  25747=>"101000000",
  25748=>"100101111",
  25749=>"101110011",
  25750=>"110110111",
  25751=>"000001111",
  25752=>"111111011",
  25753=>"011011001",
  25754=>"101100111",
  25755=>"111010110",
  25756=>"010001000",
  25757=>"101001000",
  25758=>"010000000",
  25759=>"000000011",
  25760=>"110010000",
  25761=>"111111010",
  25762=>"001111010",
  25763=>"011111010",
  25764=>"101011100",
  25765=>"110111010",
  25766=>"011011001",
  25767=>"100000001",
  25768=>"101000000",
  25769=>"011000011",
  25770=>"111110110",
  25771=>"111011000",
  25772=>"111110001",
  25773=>"101110001",
  25774=>"101010111",
  25775=>"011101100",
  25776=>"110001010",
  25777=>"000010010",
  25778=>"101010001",
  25779=>"000011111",
  25780=>"010000110",
  25781=>"010001010",
  25782=>"010001010",
  25783=>"001001001",
  25784=>"110110001",
  25785=>"111110110",
  25786=>"011010000",
  25787=>"110111011",
  25788=>"010011101",
  25789=>"001111110",
  25790=>"111111100",
  25791=>"101111111",
  25792=>"110010010",
  25793=>"000110111",
  25794=>"000110110",
  25795=>"010001011",
  25796=>"000111111",
  25797=>"110111100",
  25798=>"010001000",
  25799=>"101000101",
  25800=>"010111100",
  25801=>"010110100",
  25802=>"111111101",
  25803=>"111001010",
  25804=>"011101001",
  25805=>"101010100",
  25806=>"110000100",
  25807=>"110000111",
  25808=>"101001100",
  25809=>"011000110",
  25810=>"010110010",
  25811=>"000100101",
  25812=>"111000100",
  25813=>"010001100",
  25814=>"101110010",
  25815=>"111000111",
  25816=>"111010101",
  25817=>"010000000",
  25818=>"001100001",
  25819=>"101100010",
  25820=>"101110101",
  25821=>"010001101",
  25822=>"010110001",
  25823=>"100111000",
  25824=>"111010010",
  25825=>"111101101",
  25826=>"101001101",
  25827=>"011011110",
  25828=>"100110100",
  25829=>"110001010",
  25830=>"111111000",
  25831=>"010110100",
  25832=>"011001100",
  25833=>"110111000",
  25834=>"001101010",
  25835=>"000010101",
  25836=>"010100000",
  25837=>"111111001",
  25838=>"000010000",
  25839=>"110110001",
  25840=>"000000011",
  25841=>"110011101",
  25842=>"001011100",
  25843=>"101010100",
  25844=>"100101010",
  25845=>"000110110",
  25846=>"000101000",
  25847=>"001100100",
  25848=>"111110001",
  25849=>"010101001",
  25850=>"101011000",
  25851=>"000111100",
  25852=>"111001000",
  25853=>"010101010",
  25854=>"010101100",
  25855=>"111011000",
  25856=>"101000101",
  25857=>"111001110",
  25858=>"010000011",
  25859=>"010010011",
  25860=>"001100101",
  25861=>"010011100",
  25862=>"111100110",
  25863=>"010100010",
  25864=>"100010100",
  25865=>"101100010",
  25866=>"010010011",
  25867=>"100101010",
  25868=>"100100001",
  25869=>"111010010",
  25870=>"101000000",
  25871=>"111000100",
  25872=>"011000101",
  25873=>"010000000",
  25874=>"110100110",
  25875=>"000110010",
  25876=>"011011101",
  25877=>"011000101",
  25878=>"111111100",
  25879=>"111000101",
  25880=>"111011001",
  25881=>"100101111",
  25882=>"010010011",
  25883=>"111011101",
  25884=>"001001110",
  25885=>"010101100",
  25886=>"100110111",
  25887=>"011100111",
  25888=>"111001000",
  25889=>"000011001",
  25890=>"010010010",
  25891=>"111111010",
  25892=>"000000000",
  25893=>"010100000",
  25894=>"011101100",
  25895=>"111100000",
  25896=>"011001111",
  25897=>"000011110",
  25898=>"101101011",
  25899=>"111101111",
  25900=>"011010011",
  25901=>"110101001",
  25902=>"101110011",
  25903=>"011001000",
  25904=>"010100100",
  25905=>"011100010",
  25906=>"100001111",
  25907=>"010110000",
  25908=>"001110111",
  25909=>"000111101",
  25910=>"100110100",
  25911=>"110110111",
  25912=>"100000000",
  25913=>"001110101",
  25914=>"000000110",
  25915=>"001000001",
  25916=>"100000010",
  25917=>"011011111",
  25918=>"111101111",
  25919=>"010110100",
  25920=>"010001010",
  25921=>"110101111",
  25922=>"111001001",
  25923=>"001101100",
  25924=>"001101101",
  25925=>"011010111",
  25926=>"001100001",
  25927=>"011000110",
  25928=>"100110110",
  25929=>"111010011",
  25930=>"000000010",
  25931=>"011100011",
  25932=>"001010011",
  25933=>"111101110",
  25934=>"111111110",
  25935=>"111000011",
  25936=>"001111110",
  25937=>"000111111",
  25938=>"000010000",
  25939=>"110101111",
  25940=>"001000001",
  25941=>"011101011",
  25942=>"100001111",
  25943=>"110011110",
  25944=>"011011011",
  25945=>"100011001",
  25946=>"001010110",
  25947=>"011001010",
  25948=>"101111001",
  25949=>"011111111",
  25950=>"100000111",
  25951=>"001101010",
  25952=>"111010011",
  25953=>"111110111",
  25954=>"100010010",
  25955=>"001011000",
  25956=>"111000011",
  25957=>"010111100",
  25958=>"000000000",
  25959=>"111010100",
  25960=>"100001100",
  25961=>"001111110",
  25962=>"100111001",
  25963=>"001100111",
  25964=>"101010000",
  25965=>"010100001",
  25966=>"011111111",
  25967=>"110111010",
  25968=>"010100100",
  25969=>"100111010",
  25970=>"101111100",
  25971=>"010011110",
  25972=>"101001110",
  25973=>"101111101",
  25974=>"011100100",
  25975=>"100000111",
  25976=>"110010110",
  25977=>"100101011",
  25978=>"110001000",
  25979=>"011000100",
  25980=>"001001110",
  25981=>"111011111",
  25982=>"100100101",
  25983=>"010001011",
  25984=>"101110100",
  25985=>"000010010",
  25986=>"111111101",
  25987=>"100100000",
  25988=>"100010000",
  25989=>"110011001",
  25990=>"101101010",
  25991=>"000110111",
  25992=>"001011000",
  25993=>"101111011",
  25994=>"011101111",
  25995=>"001001010",
  25996=>"111111001",
  25997=>"010011011",
  25998=>"101111000",
  25999=>"000111111",
  26000=>"100011111",
  26001=>"011011001",
  26002=>"011111100",
  26003=>"110000110",
  26004=>"100001000",
  26005=>"001110101",
  26006=>"100010000",
  26007=>"000100111",
  26008=>"110110011",
  26009=>"000011001",
  26010=>"000111001",
  26011=>"100011001",
  26012=>"110111011",
  26013=>"101111110",
  26014=>"011101000",
  26015=>"001100000",
  26016=>"000110101",
  26017=>"100000100",
  26018=>"101100001",
  26019=>"111110110",
  26020=>"000000001",
  26021=>"000110011",
  26022=>"111101000",
  26023=>"111100000",
  26024=>"101100101",
  26025=>"011110101",
  26026=>"010100100",
  26027=>"111010001",
  26028=>"001100101",
  26029=>"010000101",
  26030=>"010101110",
  26031=>"011100000",
  26032=>"010010001",
  26033=>"101001100",
  26034=>"000101100",
  26035=>"100011000",
  26036=>"111111100",
  26037=>"011000001",
  26038=>"001011011",
  26039=>"010111101",
  26040=>"111001111",
  26041=>"110000111",
  26042=>"001001001",
  26043=>"010110110",
  26044=>"001001000",
  26045=>"001010101",
  26046=>"111011010",
  26047=>"111110010",
  26048=>"101100110",
  26049=>"101010001",
  26050=>"101000110",
  26051=>"000000010",
  26052=>"111000111",
  26053=>"111110101",
  26054=>"100100100",
  26055=>"100000000",
  26056=>"010011111",
  26057=>"001110010",
  26058=>"000000110",
  26059=>"001011100",
  26060=>"010010110",
  26061=>"111000011",
  26062=>"110011101",
  26063=>"010101001",
  26064=>"001100011",
  26065=>"110001101",
  26066=>"000000011",
  26067=>"011101001",
  26068=>"100010010",
  26069=>"011101000",
  26070=>"101100111",
  26071=>"010010111",
  26072=>"110111101",
  26073=>"110111111",
  26074=>"001100001",
  26075=>"010001101",
  26076=>"100110100",
  26077=>"101000111",
  26078=>"001111100",
  26079=>"111110101",
  26080=>"100010110",
  26081=>"010110110",
  26082=>"110100101",
  26083=>"101000101",
  26084=>"101010000",
  26085=>"111000000",
  26086=>"000011100",
  26087=>"011010000",
  26088=>"110001100",
  26089=>"111101000",
  26090=>"101001110",
  26091=>"010001001",
  26092=>"001011001",
  26093=>"110000100",
  26094=>"001111010",
  26095=>"010010000",
  26096=>"000100000",
  26097=>"000111000",
  26098=>"011011100",
  26099=>"011011111",
  26100=>"011100111",
  26101=>"100000101",
  26102=>"001001110",
  26103=>"000001010",
  26104=>"001000111",
  26105=>"100100110",
  26106=>"011001101",
  26107=>"111110101",
  26108=>"000011000",
  26109=>"000100000",
  26110=>"001010100",
  26111=>"011111111",
  26112=>"110110110",
  26113=>"001100101",
  26114=>"010111000",
  26115=>"111000000",
  26116=>"100100101",
  26117=>"100111111",
  26118=>"111111100",
  26119=>"010000001",
  26120=>"000100001",
  26121=>"011101000",
  26122=>"010000111",
  26123=>"000000001",
  26124=>"000001011",
  26125=>"111110000",
  26126=>"010000000",
  26127=>"111100010",
  26128=>"100001000",
  26129=>"000010010",
  26130=>"111000001",
  26131=>"010011110",
  26132=>"000110010",
  26133=>"101111000",
  26134=>"100000110",
  26135=>"100110111",
  26136=>"101001111",
  26137=>"101011101",
  26138=>"100000000",
  26139=>"111111011",
  26140=>"011111111",
  26141=>"000110100",
  26142=>"000100011",
  26143=>"010000101",
  26144=>"111100111",
  26145=>"100000010",
  26146=>"000010110",
  26147=>"110000000",
  26148=>"001001001",
  26149=>"100011111",
  26150=>"101011100",
  26151=>"000010011",
  26152=>"101000101",
  26153=>"001000100",
  26154=>"100011010",
  26155=>"110100010",
  26156=>"110100000",
  26157=>"101111111",
  26158=>"010100001",
  26159=>"111000010",
  26160=>"111110001",
  26161=>"000110111",
  26162=>"001000111",
  26163=>"011100110",
  26164=>"101101010",
  26165=>"010011101",
  26166=>"010001011",
  26167=>"001101110",
  26168=>"111001001",
  26169=>"101111001",
  26170=>"000111101",
  26171=>"101111100",
  26172=>"110011001",
  26173=>"101000110",
  26174=>"000000001",
  26175=>"010010001",
  26176=>"001010001",
  26177=>"010000101",
  26178=>"011111111",
  26179=>"101101001",
  26180=>"001111001",
  26181=>"100101101",
  26182=>"111010100",
  26183=>"100011011",
  26184=>"010010011",
  26185=>"001010110",
  26186=>"110011101",
  26187=>"101011011",
  26188=>"000111010",
  26189=>"110001011",
  26190=>"001111000",
  26191=>"000011010",
  26192=>"000101000",
  26193=>"101010000",
  26194=>"010101111",
  26195=>"100001001",
  26196=>"001110100",
  26197=>"000010101",
  26198=>"000111101",
  26199=>"111001001",
  26200=>"110111000",
  26201=>"000101001",
  26202=>"101111111",
  26203=>"001001101",
  26204=>"011100100",
  26205=>"000000010",
  26206=>"101110100",
  26207=>"110000000",
  26208=>"110100001",
  26209=>"001101011",
  26210=>"100010001",
  26211=>"001010011",
  26212=>"111000010",
  26213=>"001110000",
  26214=>"110010100",
  26215=>"010111101",
  26216=>"101000100",
  26217=>"000001001",
  26218=>"100011001",
  26219=>"111110010",
  26220=>"111110100",
  26221=>"101001100",
  26222=>"110011010",
  26223=>"000111001",
  26224=>"011110001",
  26225=>"000010000",
  26226=>"001001001",
  26227=>"001111101",
  26228=>"001001010",
  26229=>"101011010",
  26230=>"000111010",
  26231=>"000101010",
  26232=>"000001000",
  26233=>"100011101",
  26234=>"010011100",
  26235=>"011111001",
  26236=>"110011010",
  26237=>"000001001",
  26238=>"111100101",
  26239=>"101001100",
  26240=>"001111111",
  26241=>"110111110",
  26242=>"000010000",
  26243=>"010111011",
  26244=>"011101100",
  26245=>"101110111",
  26246=>"011101011",
  26247=>"001001000",
  26248=>"100011100",
  26249=>"100010010",
  26250=>"100011001",
  26251=>"001001101",
  26252=>"100001111",
  26253=>"100010001",
  26254=>"001110110",
  26255=>"011011011",
  26256=>"010111010",
  26257=>"001000000",
  26258=>"100110111",
  26259=>"001110001",
  26260=>"111001100",
  26261=>"110010101",
  26262=>"111100001",
  26263=>"100101001",
  26264=>"010110110",
  26265=>"111111101",
  26266=>"111101101",
  26267=>"101001110",
  26268=>"000111101",
  26269=>"000001011",
  26270=>"010101101",
  26271=>"001011110",
  26272=>"001001001",
  26273=>"000110010",
  26274=>"100011101",
  26275=>"000000100",
  26276=>"011010100",
  26277=>"001101100",
  26278=>"100011011",
  26279=>"000111111",
  26280=>"110010000",
  26281=>"101110100",
  26282=>"001010110",
  26283=>"001001100",
  26284=>"111001110",
  26285=>"101010000",
  26286=>"011010011",
  26287=>"010111011",
  26288=>"100001111",
  26289=>"111100111",
  26290=>"101001010",
  26291=>"110111110",
  26292=>"111100001",
  26293=>"110110011",
  26294=>"100100011",
  26295=>"100110110",
  26296=>"001111100",
  26297=>"011100010",
  26298=>"101010110",
  26299=>"101000010",
  26300=>"111101111",
  26301=>"101101001",
  26302=>"101101100",
  26303=>"110101010",
  26304=>"111100011",
  26305=>"010010111",
  26306=>"000001101",
  26307=>"111100110",
  26308=>"110001000",
  26309=>"000100110",
  26310=>"001001001",
  26311=>"010000010",
  26312=>"011010001",
  26313=>"001111010",
  26314=>"110001111",
  26315=>"101000011",
  26316=>"000000010",
  26317=>"101111011",
  26318=>"000001010",
  26319=>"010000001",
  26320=>"111111100",
  26321=>"000101100",
  26322=>"001100001",
  26323=>"110000011",
  26324=>"110011110",
  26325=>"100111001",
  26326=>"010101101",
  26327=>"101110111",
  26328=>"010110101",
  26329=>"011110011",
  26330=>"011011101",
  26331=>"010100001",
  26332=>"100100000",
  26333=>"000100001",
  26334=>"001101001",
  26335=>"010010000",
  26336=>"011111010",
  26337=>"101100101",
  26338=>"001111110",
  26339=>"001011101",
  26340=>"100001111",
  26341=>"101000001",
  26342=>"011001100",
  26343=>"110101101",
  26344=>"001011100",
  26345=>"010110000",
  26346=>"011110000",
  26347=>"100101011",
  26348=>"000101000",
  26349=>"010010111",
  26350=>"110000100",
  26351=>"000101111",
  26352=>"110001101",
  26353=>"000011010",
  26354=>"010111111",
  26355=>"011011111",
  26356=>"011011101",
  26357=>"111011111",
  26358=>"010100111",
  26359=>"001110100",
  26360=>"101110001",
  26361=>"111011111",
  26362=>"000101101",
  26363=>"011001101",
  26364=>"111100010",
  26365=>"000110011",
  26366=>"100000001",
  26367=>"000001000",
  26368=>"110001011",
  26369=>"100110011",
  26370=>"010001010",
  26371=>"011111111",
  26372=>"000011010",
  26373=>"010001000",
  26374=>"011110001",
  26375=>"100101000",
  26376=>"100011000",
  26377=>"000010001",
  26378=>"111000110",
  26379=>"010111110",
  26380=>"101100011",
  26381=>"010101110",
  26382=>"100010101",
  26383=>"011111001",
  26384=>"110010111",
  26385=>"100001010",
  26386=>"101010000",
  26387=>"011100001",
  26388=>"010011010",
  26389=>"000111000",
  26390=>"001011110",
  26391=>"000110011",
  26392=>"000011100",
  26393=>"100000110",
  26394=>"011000000",
  26395=>"001000110",
  26396=>"100100101",
  26397=>"000101011",
  26398=>"110110101",
  26399=>"000111111",
  26400=>"110110111",
  26401=>"110011111",
  26402=>"100111101",
  26403=>"101111111",
  26404=>"110000111",
  26405=>"100001011",
  26406=>"100100010",
  26407=>"001100000",
  26408=>"001110000",
  26409=>"001100110",
  26410=>"000000101",
  26411=>"001001001",
  26412=>"011101011",
  26413=>"111001000",
  26414=>"110001010",
  26415=>"010100110",
  26416=>"011000011",
  26417=>"001000111",
  26418=>"000010101",
  26419=>"011100010",
  26420=>"000101101",
  26421=>"010111110",
  26422=>"111011000",
  26423=>"000111111",
  26424=>"011111011",
  26425=>"001100110",
  26426=>"000111001",
  26427=>"010000001",
  26428=>"100100000",
  26429=>"001001000",
  26430=>"100010110",
  26431=>"100100111",
  26432=>"011001010",
  26433=>"110011001",
  26434=>"000010000",
  26435=>"110010000",
  26436=>"000000010",
  26437=>"110000000",
  26438=>"111011110",
  26439=>"000101000",
  26440=>"011101001",
  26441=>"110110111",
  26442=>"000011000",
  26443=>"011110000",
  26444=>"010000011",
  26445=>"011010111",
  26446=>"000100001",
  26447=>"010011000",
  26448=>"111101010",
  26449=>"000000000",
  26450=>"100110001",
  26451=>"000010011",
  26452=>"111100101",
  26453=>"011110010",
  26454=>"110011110",
  26455=>"101001000",
  26456=>"000101100",
  26457=>"010001111",
  26458=>"100101110",
  26459=>"101100001",
  26460=>"001100111",
  26461=>"111001101",
  26462=>"001111011",
  26463=>"000000101",
  26464=>"010011111",
  26465=>"001100010",
  26466=>"011100000",
  26467=>"000011110",
  26468=>"101001000",
  26469=>"010010111",
  26470=>"101010111",
  26471=>"001010001",
  26472=>"100111101",
  26473=>"111101111",
  26474=>"001110000",
  26475=>"100000100",
  26476=>"110000101",
  26477=>"111000011",
  26478=>"100101011",
  26479=>"101011110",
  26480=>"110110001",
  26481=>"101011100",
  26482=>"011101101",
  26483=>"010010010",
  26484=>"010011010",
  26485=>"000001100",
  26486=>"110110001",
  26487=>"100100101",
  26488=>"011010111",
  26489=>"111101000",
  26490=>"001100000",
  26491=>"111000111",
  26492=>"000100010",
  26493=>"000101100",
  26494=>"000000011",
  26495=>"110111001",
  26496=>"011111110",
  26497=>"100011001",
  26498=>"010101111",
  26499=>"111010001",
  26500=>"001011111",
  26501=>"010001110",
  26502=>"001100010",
  26503=>"011011101",
  26504=>"110000010",
  26505=>"010111100",
  26506=>"000010100",
  26507=>"111010111",
  26508=>"011000101",
  26509=>"010001101",
  26510=>"100100111",
  26511=>"101001011",
  26512=>"001001011",
  26513=>"011100001",
  26514=>"011010111",
  26515=>"100011100",
  26516=>"100111001",
  26517=>"010111100",
  26518=>"000011110",
  26519=>"111110101",
  26520=>"100100110",
  26521=>"111101111",
  26522=>"001111110",
  26523=>"110000011",
  26524=>"111010010",
  26525=>"101110110",
  26526=>"001011101",
  26527=>"001000010",
  26528=>"010110011",
  26529=>"100000011",
  26530=>"110111000",
  26531=>"001000111",
  26532=>"100101101",
  26533=>"111010010",
  26534=>"100100100",
  26535=>"101100110",
  26536=>"010000000",
  26537=>"000100000",
  26538=>"001000010",
  26539=>"110100010",
  26540=>"001110000",
  26541=>"110111101",
  26542=>"100000110",
  26543=>"101010110",
  26544=>"101111110",
  26545=>"100101011",
  26546=>"001101110",
  26547=>"001101110",
  26548=>"001100010",
  26549=>"101110011",
  26550=>"110011111",
  26551=>"101011001",
  26552=>"011111101",
  26553=>"100101100",
  26554=>"110001110",
  26555=>"110111100",
  26556=>"000011000",
  26557=>"001110001",
  26558=>"110001011",
  26559=>"000000000",
  26560=>"011010010",
  26561=>"000001000",
  26562=>"011111010",
  26563=>"101100110",
  26564=>"101100000",
  26565=>"010011110",
  26566=>"010110001",
  26567=>"001011010",
  26568=>"111110001",
  26569=>"100000101",
  26570=>"100110001",
  26571=>"110100000",
  26572=>"100000111",
  26573=>"101110101",
  26574=>"110101000",
  26575=>"110000111",
  26576=>"100100110",
  26577=>"100110000",
  26578=>"010000000",
  26579=>"111110111",
  26580=>"001000101",
  26581=>"100001110",
  26582=>"011110100",
  26583=>"101000010",
  26584=>"111011011",
  26585=>"010010110",
  26586=>"010011001",
  26587=>"001111110",
  26588=>"100000101",
  26589=>"010010001",
  26590=>"100110001",
  26591=>"001111101",
  26592=>"111111101",
  26593=>"011010000",
  26594=>"101001000",
  26595=>"010100100",
  26596=>"101001001",
  26597=>"111101000",
  26598=>"100001101",
  26599=>"010100011",
  26600=>"011011111",
  26601=>"010010111",
  26602=>"011110001",
  26603=>"101010011",
  26604=>"100001111",
  26605=>"000011011",
  26606=>"010011110",
  26607=>"000010001",
  26608=>"000101110",
  26609=>"111001100",
  26610=>"011110111",
  26611=>"100110001",
  26612=>"100011101",
  26613=>"000111100",
  26614=>"110111110",
  26615=>"111101101",
  26616=>"101110010",
  26617=>"000010000",
  26618=>"001010001",
  26619=>"000111101",
  26620=>"101010110",
  26621=>"101011100",
  26622=>"001000001",
  26623=>"111010000",
  26624=>"000001100",
  26625=>"100011011",
  26626=>"100011000",
  26627=>"101010100",
  26628=>"010011110",
  26629=>"010010010",
  26630=>"000110000",
  26631=>"010101100",
  26632=>"000110101",
  26633=>"111110101",
  26634=>"010001010",
  26635=>"001011101",
  26636=>"101111110",
  26637=>"101110100",
  26638=>"111100000",
  26639=>"010000000",
  26640=>"101010110",
  26641=>"111001110",
  26642=>"000001111",
  26643=>"010000000",
  26644=>"111110010",
  26645=>"110100000",
  26646=>"001100111",
  26647=>"000011101",
  26648=>"011111101",
  26649=>"000110000",
  26650=>"100001101",
  26651=>"000011100",
  26652=>"101001000",
  26653=>"101100010",
  26654=>"101010111",
  26655=>"010100010",
  26656=>"000001010",
  26657=>"011111010",
  26658=>"110000011",
  26659=>"010111000",
  26660=>"101100011",
  26661=>"111000011",
  26662=>"000110111",
  26663=>"001001110",
  26664=>"011011010",
  26665=>"111001110",
  26666=>"110110110",
  26667=>"110110101",
  26668=>"000001101",
  26669=>"101000001",
  26670=>"111100110",
  26671=>"000001111",
  26672=>"110101111",
  26673=>"111101011",
  26674=>"011010110",
  26675=>"101110011",
  26676=>"101111101",
  26677=>"011001011",
  26678=>"110101000",
  26679=>"100100010",
  26680=>"011100101",
  26681=>"110001100",
  26682=>"000100000",
  26683=>"011100000",
  26684=>"100111100",
  26685=>"101000001",
  26686=>"111010101",
  26687=>"011011101",
  26688=>"101000100",
  26689=>"011100000",
  26690=>"101100010",
  26691=>"110111110",
  26692=>"110010111",
  26693=>"001001010",
  26694=>"100101011",
  26695=>"000010010",
  26696=>"111100000",
  26697=>"000110111",
  26698=>"110011111",
  26699=>"001000010",
  26700=>"001100100",
  26701=>"010100011",
  26702=>"101000110",
  26703=>"011101000",
  26704=>"101100001",
  26705=>"100111010",
  26706=>"011111000",
  26707=>"011100011",
  26708=>"111001111",
  26709=>"011001110",
  26710=>"111101010",
  26711=>"101101001",
  26712=>"101011111",
  26713=>"011000001",
  26714=>"001001010",
  26715=>"100111110",
  26716=>"001101111",
  26717=>"100111000",
  26718=>"000100011",
  26719=>"001100101",
  26720=>"010000100",
  26721=>"000110111",
  26722=>"100101101",
  26723=>"101010101",
  26724=>"010011000",
  26725=>"111011110",
  26726=>"010001111",
  26727=>"101010010",
  26728=>"101001110",
  26729=>"100011110",
  26730=>"110000000",
  26731=>"110111011",
  26732=>"110011100",
  26733=>"010101110",
  26734=>"101111110",
  26735=>"100100111",
  26736=>"101001001",
  26737=>"011101011",
  26738=>"111000100",
  26739=>"100110100",
  26740=>"000010000",
  26741=>"000100100",
  26742=>"111010100",
  26743=>"110101000",
  26744=>"110111011",
  26745=>"001001010",
  26746=>"010010010",
  26747=>"110000011",
  26748=>"000101101",
  26749=>"010010101",
  26750=>"000000001",
  26751=>"010000001",
  26752=>"100001100",
  26753=>"111101010",
  26754=>"001101011",
  26755=>"000111010",
  26756=>"100101101",
  26757=>"111011101",
  26758=>"110010110",
  26759=>"001011110",
  26760=>"010000101",
  26761=>"100000010",
  26762=>"000000010",
  26763=>"011011111",
  26764=>"110100010",
  26765=>"000110101",
  26766=>"000001111",
  26767=>"110100101",
  26768=>"101111101",
  26769=>"001000101",
  26770=>"000011000",
  26771=>"110010001",
  26772=>"010110010",
  26773=>"100011010",
  26774=>"000001000",
  26775=>"111110100",
  26776=>"010011110",
  26777=>"010101001",
  26778=>"110001010",
  26779=>"111111000",
  26780=>"011000001",
  26781=>"111101111",
  26782=>"010010100",
  26783=>"100101000",
  26784=>"111110011",
  26785=>"100010111",
  26786=>"010000001",
  26787=>"011101010",
  26788=>"000010000",
  26789=>"010001100",
  26790=>"000001111",
  26791=>"011001001",
  26792=>"111001011",
  26793=>"011010110",
  26794=>"110111000",
  26795=>"000100100",
  26796=>"110110110",
  26797=>"101111000",
  26798=>"110011011",
  26799=>"110101110",
  26800=>"011101001",
  26801=>"101001100",
  26802=>"011101101",
  26803=>"001100110",
  26804=>"000001011",
  26805=>"101101101",
  26806=>"001011100",
  26807=>"100010111",
  26808=>"010110000",
  26809=>"001001100",
  26810=>"111001000",
  26811=>"101111100",
  26812=>"101010111",
  26813=>"110111100",
  26814=>"001000010",
  26815=>"101000101",
  26816=>"001111011",
  26817=>"011000000",
  26818=>"001100000",
  26819=>"001001001",
  26820=>"000100010",
  26821=>"110000001",
  26822=>"000000111",
  26823=>"101000010",
  26824=>"000000100",
  26825=>"000011010",
  26826=>"111001010",
  26827=>"011100111",
  26828=>"111000010",
  26829=>"000011000",
  26830=>"001001010",
  26831=>"011001100",
  26832=>"011011111",
  26833=>"001101110",
  26834=>"001010010",
  26835=>"111000111",
  26836=>"101011100",
  26837=>"110111111",
  26838=>"001101001",
  26839=>"101110101",
  26840=>"001001000",
  26841=>"000100110",
  26842=>"101001011",
  26843=>"111000011",
  26844=>"110000000",
  26845=>"110001011",
  26846=>"111001101",
  26847=>"101101101",
  26848=>"111000111",
  26849=>"010010001",
  26850=>"111000110",
  26851=>"001100001",
  26852=>"101001110",
  26853=>"111000001",
  26854=>"101000110",
  26855=>"001111110",
  26856=>"011101011",
  26857=>"100100000",
  26858=>"000100001",
  26859=>"111101110",
  26860=>"001000000",
  26861=>"010110111",
  26862=>"111001011",
  26863=>"011010001",
  26864=>"001000111",
  26865=>"000100110",
  26866=>"011000000",
  26867=>"100010101",
  26868=>"110111010",
  26869=>"001111001",
  26870=>"000011000",
  26871=>"110000100",
  26872=>"100111110",
  26873=>"010001111",
  26874=>"001010001",
  26875=>"010100100",
  26876=>"111101011",
  26877=>"100101011",
  26878=>"101000100",
  26879=>"000010000",
  26880=>"110110001",
  26881=>"001111000",
  26882=>"001001010",
  26883=>"001110110",
  26884=>"010010100",
  26885=>"110111000",
  26886=>"010110010",
  26887=>"111110011",
  26888=>"010101001",
  26889=>"001000101",
  26890=>"010001100",
  26891=>"100110100",
  26892=>"110000011",
  26893=>"111000101",
  26894=>"001001001",
  26895=>"011111001",
  26896=>"001011001",
  26897=>"010100001",
  26898=>"001101100",
  26899=>"111101001",
  26900=>"001101100",
  26901=>"101011011",
  26902=>"101000110",
  26903=>"101101000",
  26904=>"001111110",
  26905=>"111010110",
  26906=>"010110111",
  26907=>"001111100",
  26908=>"101011010",
  26909=>"010110101",
  26910=>"101001100",
  26911=>"111001010",
  26912=>"110000111",
  26913=>"011101001",
  26914=>"011111010",
  26915=>"011110010",
  26916=>"010011101",
  26917=>"010010001",
  26918=>"110100111",
  26919=>"111010010",
  26920=>"010010011",
  26921=>"010000000",
  26922=>"100110000",
  26923=>"110100000",
  26924=>"010000101",
  26925=>"110011000",
  26926=>"101000000",
  26927=>"001111111",
  26928=>"101100010",
  26929=>"000111001",
  26930=>"111110101",
  26931=>"011110011",
  26932=>"111111010",
  26933=>"110101100",
  26934=>"111101010",
  26935=>"100001001",
  26936=>"100000010",
  26937=>"011101001",
  26938=>"001000110",
  26939=>"011101000",
  26940=>"011101110",
  26941=>"000000101",
  26942=>"010010110",
  26943=>"110101100",
  26944=>"111100101",
  26945=>"001101010",
  26946=>"110010011",
  26947=>"001010011",
  26948=>"101100101",
  26949=>"011100011",
  26950=>"010101011",
  26951=>"101111011",
  26952=>"110111010",
  26953=>"011001111",
  26954=>"100001011",
  26955=>"000011101",
  26956=>"101110101",
  26957=>"001011110",
  26958=>"111001111",
  26959=>"101110010",
  26960=>"110110110",
  26961=>"111100100",
  26962=>"001110101",
  26963=>"001010101",
  26964=>"101111110",
  26965=>"101111110",
  26966=>"111110010",
  26967=>"100110110",
  26968=>"001001101",
  26969=>"100001110",
  26970=>"000010000",
  26971=>"100011111",
  26972=>"111001111",
  26973=>"111110110",
  26974=>"011011010",
  26975=>"100100100",
  26976=>"000011110",
  26977=>"010011010",
  26978=>"101000110",
  26979=>"101000000",
  26980=>"111010011",
  26981=>"011011001",
  26982=>"111010011",
  26983=>"000001001",
  26984=>"110100000",
  26985=>"111100001",
  26986=>"010001111",
  26987=>"111000100",
  26988=>"001101010",
  26989=>"101111110",
  26990=>"100110001",
  26991=>"010100011",
  26992=>"111000100",
  26993=>"000111011",
  26994=>"101011001",
  26995=>"110110011",
  26996=>"101011011",
  26997=>"000111110",
  26998=>"100001110",
  26999=>"001100110",
  27000=>"000100001",
  27001=>"110101101",
  27002=>"110010110",
  27003=>"001111100",
  27004=>"010100000",
  27005=>"110011111",
  27006=>"010001111",
  27007=>"111110011",
  27008=>"010000100",
  27009=>"111011101",
  27010=>"111000000",
  27011=>"111011110",
  27012=>"100110100",
  27013=>"000101100",
  27014=>"101110110",
  27015=>"010101110",
  27016=>"001010010",
  27017=>"001000001",
  27018=>"011011111",
  27019=>"111010010",
  27020=>"000101111",
  27021=>"111101001",
  27022=>"101010101",
  27023=>"001011001",
  27024=>"111011011",
  27025=>"001110100",
  27026=>"000001110",
  27027=>"100110001",
  27028=>"100011100",
  27029=>"000100001",
  27030=>"101111000",
  27031=>"111001100",
  27032=>"001101100",
  27033=>"001000000",
  27034=>"100001100",
  27035=>"110100011",
  27036=>"010010101",
  27037=>"000001111",
  27038=>"110111000",
  27039=>"101110110",
  27040=>"100111111",
  27041=>"110100101",
  27042=>"111110111",
  27043=>"100001111",
  27044=>"010100011",
  27045=>"010000100",
  27046=>"111111100",
  27047=>"111000101",
  27048=>"101010011",
  27049=>"010110000",
  27050=>"010000101",
  27051=>"000101000",
  27052=>"100100011",
  27053=>"001100000",
  27054=>"101010011",
  27055=>"000101101",
  27056=>"100110001",
  27057=>"111100101",
  27058=>"000110100",
  27059=>"101001011",
  27060=>"110011011",
  27061=>"010011011",
  27062=>"110100100",
  27063=>"000100111",
  27064=>"111000100",
  27065=>"001000001",
  27066=>"001110111",
  27067=>"111101000",
  27068=>"000000010",
  27069=>"100111000",
  27070=>"111111100",
  27071=>"111111000",
  27072=>"010110101",
  27073=>"010100011",
  27074=>"011001101",
  27075=>"111101010",
  27076=>"000000000",
  27077=>"110001000",
  27078=>"011101101",
  27079=>"001000001",
  27080=>"001101101",
  27081=>"110010000",
  27082=>"010000111",
  27083=>"010101000",
  27084=>"101110011",
  27085=>"100010110",
  27086=>"011001111",
  27087=>"001101101",
  27088=>"001001000",
  27089=>"100010010",
  27090=>"100000010",
  27091=>"111101001",
  27092=>"100110111",
  27093=>"000011100",
  27094=>"100011101",
  27095=>"110100010",
  27096=>"110010100",
  27097=>"000101101",
  27098=>"001010011",
  27099=>"111100000",
  27100=>"001110100",
  27101=>"010100010",
  27102=>"110111000",
  27103=>"011110101",
  27104=>"100101011",
  27105=>"100100111",
  27106=>"111110010",
  27107=>"101011111",
  27108=>"010101011",
  27109=>"011000100",
  27110=>"111001111",
  27111=>"000000000",
  27112=>"110110101",
  27113=>"010011110",
  27114=>"110101100",
  27115=>"011011101",
  27116=>"101101111",
  27117=>"000101110",
  27118=>"101100010",
  27119=>"001001010",
  27120=>"100011000",
  27121=>"011100000",
  27122=>"110111100",
  27123=>"101100001",
  27124=>"000010100",
  27125=>"000000101",
  27126=>"010011001",
  27127=>"001000110",
  27128=>"110011100",
  27129=>"111000001",
  27130=>"010111100",
  27131=>"001010100",
  27132=>"100110000",
  27133=>"111110110",
  27134=>"000110000",
  27135=>"010001100",
  27136=>"011110001",
  27137=>"100111000",
  27138=>"010110101",
  27139=>"100000001",
  27140=>"001000011",
  27141=>"010001101",
  27142=>"000110001",
  27143=>"001110110",
  27144=>"100110111",
  27145=>"001001011",
  27146=>"111100111",
  27147=>"110001011",
  27148=>"111000101",
  27149=>"110011001",
  27150=>"011000010",
  27151=>"001010110",
  27152=>"101001100",
  27153=>"110101110",
  27154=>"001101110",
  27155=>"100001111",
  27156=>"100111000",
  27157=>"011101001",
  27158=>"010101110",
  27159=>"011100001",
  27160=>"000010110",
  27161=>"010001111",
  27162=>"100110011",
  27163=>"011000000",
  27164=>"101100011",
  27165=>"011100001",
  27166=>"100001111",
  27167=>"000010110",
  27168=>"101001100",
  27169=>"100111000",
  27170=>"101100110",
  27171=>"001000000",
  27172=>"111011001",
  27173=>"010000010",
  27174=>"011011001",
  27175=>"100101000",
  27176=>"110011000",
  27177=>"100111101",
  27178=>"101010110",
  27179=>"101110000",
  27180=>"010101100",
  27181=>"100111101",
  27182=>"111111001",
  27183=>"111100111",
  27184=>"010100101",
  27185=>"111001110",
  27186=>"011000111",
  27187=>"110001010",
  27188=>"011000011",
  27189=>"100111010",
  27190=>"110001000",
  27191=>"011111010",
  27192=>"001110111",
  27193=>"101100000",
  27194=>"011000000",
  27195=>"100110000",
  27196=>"111100000",
  27197=>"001101010",
  27198=>"110001000",
  27199=>"110111101",
  27200=>"101010101",
  27201=>"010001100",
  27202=>"010000111",
  27203=>"101101100",
  27204=>"101110001",
  27205=>"000001110",
  27206=>"001100000",
  27207=>"000101000",
  27208=>"000101110",
  27209=>"111110100",
  27210=>"001110000",
  27211=>"101010100",
  27212=>"000000000",
  27213=>"101101110",
  27214=>"111011011",
  27215=>"010101111",
  27216=>"000010110",
  27217=>"111011101",
  27218=>"100000010",
  27219=>"111111111",
  27220=>"100100101",
  27221=>"101011111",
  27222=>"001011000",
  27223=>"001110010",
  27224=>"111011010",
  27225=>"010111000",
  27226=>"000000000",
  27227=>"110101010",
  27228=>"100000100",
  27229=>"000101000",
  27230=>"000010101",
  27231=>"011111000",
  27232=>"110101111",
  27233=>"101101011",
  27234=>"000010111",
  27235=>"101100001",
  27236=>"011111000",
  27237=>"010101001",
  27238=>"000010010",
  27239=>"100100001",
  27240=>"000001000",
  27241=>"000111001",
  27242=>"100001011",
  27243=>"001100011",
  27244=>"001000100",
  27245=>"011111011",
  27246=>"010001001",
  27247=>"000100101",
  27248=>"000011100",
  27249=>"010010110",
  27250=>"010000001",
  27251=>"110111100",
  27252=>"101111111",
  27253=>"110101001",
  27254=>"111111111",
  27255=>"111100001",
  27256=>"001110010",
  27257=>"111110100",
  27258=>"011100110",
  27259=>"101100011",
  27260=>"101100010",
  27261=>"100110110",
  27262=>"110011001",
  27263=>"001011111",
  27264=>"001010011",
  27265=>"010111110",
  27266=>"101011111",
  27267=>"111111101",
  27268=>"011010000",
  27269=>"010100000",
  27270=>"001011100",
  27271=>"000010111",
  27272=>"001110010",
  27273=>"100101010",
  27274=>"011010110",
  27275=>"101110000",
  27276=>"101010100",
  27277=>"010100000",
  27278=>"110110101",
  27279=>"011010000",
  27280=>"001011011",
  27281=>"001011100",
  27282=>"111010000",
  27283=>"011010011",
  27284=>"101001000",
  27285=>"111011111",
  27286=>"101100000",
  27287=>"110100010",
  27288=>"111011110",
  27289=>"000100101",
  27290=>"100001000",
  27291=>"010001011",
  27292=>"100111101",
  27293=>"011110110",
  27294=>"100001010",
  27295=>"001110101",
  27296=>"100000011",
  27297=>"001000001",
  27298=>"100011000",
  27299=>"001111001",
  27300=>"010001001",
  27301=>"000101000",
  27302=>"100101000",
  27303=>"101000110",
  27304=>"010110101",
  27305=>"101101110",
  27306=>"001011010",
  27307=>"001001110",
  27308=>"100011100",
  27309=>"100010001",
  27310=>"001110101",
  27311=>"011110111",
  27312=>"110010010",
  27313=>"000011011",
  27314=>"111000011",
  27315=>"001001011",
  27316=>"110101011",
  27317=>"011101000",
  27318=>"100000000",
  27319=>"011111001",
  27320=>"010010101",
  27321=>"010101110",
  27322=>"111111111",
  27323=>"011011111",
  27324=>"111001011",
  27325=>"010010100",
  27326=>"100001001",
  27327=>"111011101",
  27328=>"011111010",
  27329=>"111011010",
  27330=>"011011000",
  27331=>"110010011",
  27332=>"101000100",
  27333=>"010010101",
  27334=>"100110001",
  27335=>"011001100",
  27336=>"100110101",
  27337=>"100110000",
  27338=>"010110100",
  27339=>"000110000",
  27340=>"000000011",
  27341=>"010101101",
  27342=>"010100101",
  27343=>"001000010",
  27344=>"000000100",
  27345=>"100001010",
  27346=>"000001010",
  27347=>"011000011",
  27348=>"001000000",
  27349=>"111100111",
  27350=>"010111000",
  27351=>"111000000",
  27352=>"001111111",
  27353=>"110011011",
  27354=>"001011001",
  27355=>"110001010",
  27356=>"001100100",
  27357=>"111011001",
  27358=>"100001100",
  27359=>"001000011",
  27360=>"010100011",
  27361=>"000110110",
  27362=>"111111100",
  27363=>"110001110",
  27364=>"000000000",
  27365=>"011110011",
  27366=>"000001110",
  27367=>"111111010",
  27368=>"000000101",
  27369=>"110111001",
  27370=>"011000010",
  27371=>"010000011",
  27372=>"111001001",
  27373=>"000011110",
  27374=>"011101000",
  27375=>"111000101",
  27376=>"010001011",
  27377=>"000110110",
  27378=>"011010100",
  27379=>"011000011",
  27380=>"001110110",
  27381=>"000100000",
  27382=>"000100011",
  27383=>"101000000",
  27384=>"101101010",
  27385=>"010001100",
  27386=>"001001110",
  27387=>"100011011",
  27388=>"011001111",
  27389=>"001010011",
  27390=>"110001110",
  27391=>"000010110",
  27392=>"010110111",
  27393=>"001001110",
  27394=>"000111110",
  27395=>"110011011",
  27396=>"100100001",
  27397=>"010101111",
  27398=>"000001010",
  27399=>"101110101",
  27400=>"101100010",
  27401=>"000111110",
  27402=>"110110100",
  27403=>"110001101",
  27404=>"011110001",
  27405=>"000010110",
  27406=>"100100001",
  27407=>"010111010",
  27408=>"011110000",
  27409=>"111110010",
  27410=>"000111100",
  27411=>"001100100",
  27412=>"100111111",
  27413=>"110011111",
  27414=>"001010010",
  27415=>"100011111",
  27416=>"100100100",
  27417=>"111100011",
  27418=>"011101001",
  27419=>"111111101",
  27420=>"100010100",
  27421=>"101110111",
  27422=>"011011110",
  27423=>"011111110",
  27424=>"100001101",
  27425=>"000010011",
  27426=>"011110011",
  27427=>"100001101",
  27428=>"111010110",
  27429=>"000101110",
  27430=>"111110111",
  27431=>"000010001",
  27432=>"111101011",
  27433=>"110000011",
  27434=>"011101011",
  27435=>"111011011",
  27436=>"011000000",
  27437=>"100011111",
  27438=>"110100110",
  27439=>"010000001",
  27440=>"111100110",
  27441=>"011111001",
  27442=>"111101001",
  27443=>"111010110",
  27444=>"010111000",
  27445=>"110111000",
  27446=>"111010110",
  27447=>"111001010",
  27448=>"001011110",
  27449=>"100111001",
  27450=>"111011001",
  27451=>"110010000",
  27452=>"110000110",
  27453=>"100001100",
  27454=>"001000000",
  27455=>"110001010",
  27456=>"100110110",
  27457=>"110001001",
  27458=>"110111001",
  27459=>"010101100",
  27460=>"011001001",
  27461=>"100101101",
  27462=>"101101010",
  27463=>"110111010",
  27464=>"011010001",
  27465=>"001000001",
  27466=>"111100111",
  27467=>"100100110",
  27468=>"011101000",
  27469=>"101000110",
  27470=>"100100011",
  27471=>"011110001",
  27472=>"110101101",
  27473=>"110011000",
  27474=>"100010000",
  27475=>"000000010",
  27476=>"000100101",
  27477=>"100111100",
  27478=>"001000110",
  27479=>"010010011",
  27480=>"001100110",
  27481=>"111110000",
  27482=>"101100001",
  27483=>"000001011",
  27484=>"011100110",
  27485=>"111000110",
  27486=>"111000011",
  27487=>"111100101",
  27488=>"110001111",
  27489=>"101011110",
  27490=>"001101001",
  27491=>"110001010",
  27492=>"111011010",
  27493=>"110010111",
  27494=>"001011100",
  27495=>"001100101",
  27496=>"011000000",
  27497=>"100110100",
  27498=>"000001001",
  27499=>"000001000",
  27500=>"110111001",
  27501=>"001001110",
  27502=>"010001001",
  27503=>"100100000",
  27504=>"101001010",
  27505=>"100010111",
  27506=>"111010110",
  27507=>"000000100",
  27508=>"100000000",
  27509=>"001111111",
  27510=>"100100100",
  27511=>"011101011",
  27512=>"100101101",
  27513=>"010100001",
  27514=>"010101111",
  27515=>"011010100",
  27516=>"001110000",
  27517=>"100010011",
  27518=>"100110011",
  27519=>"000110011",
  27520=>"011100001",
  27521=>"110011101",
  27522=>"101110001",
  27523=>"110001010",
  27524=>"011100011",
  27525=>"000101100",
  27526=>"101001001",
  27527=>"010010111",
  27528=>"011001000",
  27529=>"010000000",
  27530=>"110001101",
  27531=>"010110100",
  27532=>"110111010",
  27533=>"101100100",
  27534=>"001100101",
  27535=>"111001111",
  27536=>"111110100",
  27537=>"011001011",
  27538=>"011111111",
  27539=>"001011001",
  27540=>"011101011",
  27541=>"100100101",
  27542=>"000111000",
  27543=>"000110100",
  27544=>"001000011",
  27545=>"100011101",
  27546=>"001110011",
  27547=>"001110011",
  27548=>"100110100",
  27549=>"110001000",
  27550=>"001110101",
  27551=>"011001011",
  27552=>"011001100",
  27553=>"110110111",
  27554=>"111110001",
  27555=>"011000000",
  27556=>"110111010",
  27557=>"000011101",
  27558=>"101010000",
  27559=>"001000000",
  27560=>"000100010",
  27561=>"000101111",
  27562=>"010100110",
  27563=>"010000101",
  27564=>"100111010",
  27565=>"011001000",
  27566=>"011001101",
  27567=>"011110011",
  27568=>"011001100",
  27569=>"100100010",
  27570=>"110110010",
  27571=>"111111001",
  27572=>"011000000",
  27573=>"011110000",
  27574=>"011011001",
  27575=>"111111110",
  27576=>"101000111",
  27577=>"011001010",
  27578=>"110111000",
  27579=>"000111000",
  27580=>"000100110",
  27581=>"000001111",
  27582=>"100110000",
  27583=>"101111111",
  27584=>"111001010",
  27585=>"110111100",
  27586=>"011100111",
  27587=>"111010000",
  27588=>"010101000",
  27589=>"111111001",
  27590=>"001011100",
  27591=>"000110100",
  27592=>"111100100",
  27593=>"001011001",
  27594=>"101110001",
  27595=>"111100000",
  27596=>"011101001",
  27597=>"111000101",
  27598=>"011101110",
  27599=>"010000011",
  27600=>"100111111",
  27601=>"110111011",
  27602=>"110111000",
  27603=>"011000000",
  27604=>"111111100",
  27605=>"000001000",
  27606=>"010101000",
  27607=>"011111110",
  27608=>"100010011",
  27609=>"101100111",
  27610=>"011011110",
  27611=>"100100000",
  27612=>"111101100",
  27613=>"011111100",
  27614=>"011010110",
  27615=>"000001010",
  27616=>"100100100",
  27617=>"010010001",
  27618=>"111111100",
  27619=>"001100010",
  27620=>"011011001",
  27621=>"111111000",
  27622=>"101111001",
  27623=>"111011011",
  27624=>"101011101",
  27625=>"110001111",
  27626=>"111100111",
  27627=>"011101011",
  27628=>"010001001",
  27629=>"101000010",
  27630=>"111101011",
  27631=>"011110010",
  27632=>"101010100",
  27633=>"100001111",
  27634=>"001000100",
  27635=>"001011001",
  27636=>"010111111",
  27637=>"000011001",
  27638=>"100100110",
  27639=>"100000111",
  27640=>"000111000",
  27641=>"111111110",
  27642=>"000110101",
  27643=>"000101101",
  27644=>"110101101",
  27645=>"000100100",
  27646=>"111010111",
  27647=>"001110111",
  27648=>"000010000",
  27649=>"101000000",
  27650=>"010101111",
  27651=>"000101111",
  27652=>"010110001",
  27653=>"000110000",
  27654=>"101000000",
  27655=>"101111100",
  27656=>"000111011",
  27657=>"010000111",
  27658=>"111011111",
  27659=>"100010011",
  27660=>"110101110",
  27661=>"011101011",
  27662=>"110111010",
  27663=>"000010000",
  27664=>"001000001",
  27665=>"010100100",
  27666=>"000010011",
  27667=>"010000001",
  27668=>"001001101",
  27669=>"001100011",
  27670=>"111101111",
  27671=>"010100110",
  27672=>"000101010",
  27673=>"101000000",
  27674=>"110110010",
  27675=>"010001111",
  27676=>"000011000",
  27677=>"110111100",
  27678=>"010010100",
  27679=>"110000100",
  27680=>"011100001",
  27681=>"000101111",
  27682=>"001011001",
  27683=>"010101000",
  27684=>"011011001",
  27685=>"000100010",
  27686=>"110101110",
  27687=>"100011110",
  27688=>"000000110",
  27689=>"101100111",
  27690=>"100111010",
  27691=>"110100000",
  27692=>"010010110",
  27693=>"010100110",
  27694=>"101001011",
  27695=>"010110100",
  27696=>"110111111",
  27697=>"110110101",
  27698=>"110100101",
  27699=>"000001001",
  27700=>"010110100",
  27701=>"100111001",
  27702=>"011000000",
  27703=>"011011110",
  27704=>"001010111",
  27705=>"000110100",
  27706=>"110000101",
  27707=>"000100111",
  27708=>"011000000",
  27709=>"111110010",
  27710=>"001111000",
  27711=>"000010100",
  27712=>"000110000",
  27713=>"101000001",
  27714=>"000001100",
  27715=>"100111111",
  27716=>"111110001",
  27717=>"100100111",
  27718=>"010111010",
  27719=>"000101001",
  27720=>"011010000",
  27721=>"110111101",
  27722=>"000001000",
  27723=>"010110011",
  27724=>"001011000",
  27725=>"101111010",
  27726=>"011010100",
  27727=>"101011011",
  27728=>"101010001",
  27729=>"111011100",
  27730=>"010010100",
  27731=>"111011111",
  27732=>"101100100",
  27733=>"011101111",
  27734=>"111100101",
  27735=>"001001001",
  27736=>"000110000",
  27737=>"110010111",
  27738=>"011100010",
  27739=>"010001010",
  27740=>"101011000",
  27741=>"110011111",
  27742=>"101001010",
  27743=>"000110101",
  27744=>"010100000",
  27745=>"101100101",
  27746=>"111101111",
  27747=>"011001111",
  27748=>"100011011",
  27749=>"000111000",
  27750=>"010111101",
  27751=>"011111101",
  27752=>"000100100",
  27753=>"101111010",
  27754=>"101111011",
  27755=>"100010111",
  27756=>"111010111",
  27757=>"010100011",
  27758=>"111000010",
  27759=>"001101110",
  27760=>"101100010",
  27761=>"110110011",
  27762=>"000100011",
  27763=>"110000111",
  27764=>"000100011",
  27765=>"010100111",
  27766=>"001000011",
  27767=>"000001000",
  27768=>"101001010",
  27769=>"110101001",
  27770=>"000010100",
  27771=>"100000111",
  27772=>"100000000",
  27773=>"101111100",
  27774=>"000010010",
  27775=>"010111011",
  27776=>"000000010",
  27777=>"110000010",
  27778=>"100001111",
  27779=>"001110100",
  27780=>"000100100",
  27781=>"011001100",
  27782=>"110000011",
  27783=>"010100111",
  27784=>"011000111",
  27785=>"100010010",
  27786=>"000000011",
  27787=>"111010100",
  27788=>"001111010",
  27789=>"110000101",
  27790=>"101011111",
  27791=>"011111111",
  27792=>"010111111",
  27793=>"110111110",
  27794=>"000101011",
  27795=>"100110001",
  27796=>"101001001",
  27797=>"110011001",
  27798=>"001101010",
  27799=>"010000010",
  27800=>"101101000",
  27801=>"101000100",
  27802=>"000001000",
  27803=>"110100101",
  27804=>"101111111",
  27805=>"000111101",
  27806=>"010011000",
  27807=>"010100000",
  27808=>"000011101",
  27809=>"001001100",
  27810=>"101111011",
  27811=>"110011001",
  27812=>"010000001",
  27813=>"101110010",
  27814=>"111011011",
  27815=>"100101111",
  27816=>"000101100",
  27817=>"011011001",
  27818=>"000011000",
  27819=>"101101001",
  27820=>"110011000",
  27821=>"000111011",
  27822=>"010010111",
  27823=>"111110110",
  27824=>"100000101",
  27825=>"100000000",
  27826=>"010100010",
  27827=>"110000111",
  27828=>"011010101",
  27829=>"000001110",
  27830=>"000100111",
  27831=>"011001110",
  27832=>"011111000",
  27833=>"110101111",
  27834=>"111100001",
  27835=>"111100001",
  27836=>"110101110",
  27837=>"010101001",
  27838=>"100010111",
  27839=>"000011010",
  27840=>"011000011",
  27841=>"101111001",
  27842=>"001111001",
  27843=>"011110000",
  27844=>"100100000",
  27845=>"101111100",
  27846=>"101111001",
  27847=>"010111100",
  27848=>"010101101",
  27849=>"001011001",
  27850=>"110000110",
  27851=>"110101100",
  27852=>"101001011",
  27853=>"011101101",
  27854=>"001001000",
  27855=>"000010011",
  27856=>"010001011",
  27857=>"100000011",
  27858=>"000010000",
  27859=>"101011011",
  27860=>"111111111",
  27861=>"011111101",
  27862=>"000000000",
  27863=>"110100101",
  27864=>"010111011",
  27865=>"001100010",
  27866=>"010111110",
  27867=>"010100000",
  27868=>"011110111",
  27869=>"111001110",
  27870=>"111110111",
  27871=>"010011111",
  27872=>"110000000",
  27873=>"000110000",
  27874=>"101101111",
  27875=>"000110011",
  27876=>"111110001",
  27877=>"111111100",
  27878=>"100111000",
  27879=>"010100111",
  27880=>"100111000",
  27881=>"100100011",
  27882=>"010011010",
  27883=>"001000011",
  27884=>"111110010",
  27885=>"101010100",
  27886=>"001000011",
  27887=>"010010110",
  27888=>"010000001",
  27889=>"011101110",
  27890=>"001111001",
  27891=>"100101110",
  27892=>"000111111",
  27893=>"001110000",
  27894=>"110100001",
  27895=>"100000010",
  27896=>"001010001",
  27897=>"010011010",
  27898=>"111011010",
  27899=>"101100001",
  27900=>"110011000",
  27901=>"001000000",
  27902=>"011000001",
  27903=>"100010011",
  27904=>"100001011",
  27905=>"100011010",
  27906=>"010001111",
  27907=>"111101101",
  27908=>"001000101",
  27909=>"001111111",
  27910=>"111101011",
  27911=>"110101100",
  27912=>"110001011",
  27913=>"001010000",
  27914=>"100101011",
  27915=>"100100000",
  27916=>"000111001",
  27917=>"001111111",
  27918=>"110110011",
  27919=>"011100001",
  27920=>"010100010",
  27921=>"010110011",
  27922=>"011001101",
  27923=>"001000000",
  27924=>"010010101",
  27925=>"010001101",
  27926=>"001100101",
  27927=>"010011101",
  27928=>"100011011",
  27929=>"010010010",
  27930=>"110011001",
  27931=>"101010001",
  27932=>"101100110",
  27933=>"100101010",
  27934=>"001111111",
  27935=>"011011100",
  27936=>"010110101",
  27937=>"010111011",
  27938=>"101011010",
  27939=>"010110101",
  27940=>"110101011",
  27941=>"011110100",
  27942=>"001000110",
  27943=>"000000100",
  27944=>"110010001",
  27945=>"001010010",
  27946=>"101110101",
  27947=>"010100110",
  27948=>"011100110",
  27949=>"000010001",
  27950=>"001100101",
  27951=>"110000101",
  27952=>"111001100",
  27953=>"100010011",
  27954=>"101011011",
  27955=>"001001111",
  27956=>"000001101",
  27957=>"000000000",
  27958=>"111110111",
  27959=>"110101011",
  27960=>"100011101",
  27961=>"000011111",
  27962=>"001100001",
  27963=>"100110101",
  27964=>"111111101",
  27965=>"101001111",
  27966=>"011111001",
  27967=>"001110100",
  27968=>"110110110",
  27969=>"000001011",
  27970=>"010010111",
  27971=>"110010101",
  27972=>"110001011",
  27973=>"101101111",
  27974=>"101110000",
  27975=>"010010011",
  27976=>"111111101",
  27977=>"111010010",
  27978=>"011100000",
  27979=>"001000100",
  27980=>"100110110",
  27981=>"001011101",
  27982=>"000000000",
  27983=>"101111010",
  27984=>"111111111",
  27985=>"110101001",
  27986=>"001011000",
  27987=>"100011011",
  27988=>"111010101",
  27989=>"101000000",
  27990=>"001000100",
  27991=>"101011101",
  27992=>"101000111",
  27993=>"000010000",
  27994=>"010001010",
  27995=>"110001010",
  27996=>"110111100",
  27997=>"111111111",
  27998=>"011110011",
  27999=>"100010000",
  28000=>"110111110",
  28001=>"110110001",
  28002=>"000110011",
  28003=>"011111000",
  28004=>"011100111",
  28005=>"100100101",
  28006=>"100011110",
  28007=>"110101111",
  28008=>"000000110",
  28009=>"011010000",
  28010=>"011011001",
  28011=>"010100100",
  28012=>"010110011",
  28013=>"011001100",
  28014=>"000011101",
  28015=>"100100011",
  28016=>"001000001",
  28017=>"101001011",
  28018=>"100100001",
  28019=>"111011000",
  28020=>"000001100",
  28021=>"101000001",
  28022=>"100111101",
  28023=>"101100010",
  28024=>"000001101",
  28025=>"010111110",
  28026=>"011001010",
  28027=>"001010010",
  28028=>"011010100",
  28029=>"000111011",
  28030=>"101101110",
  28031=>"100111001",
  28032=>"110000010",
  28033=>"010110111",
  28034=>"000011001",
  28035=>"011001010",
  28036=>"101001101",
  28037=>"010110111",
  28038=>"010101101",
  28039=>"000000011",
  28040=>"000001001",
  28041=>"110111101",
  28042=>"111000000",
  28043=>"110011000",
  28044=>"111111101",
  28045=>"100000000",
  28046=>"101010000",
  28047=>"110001110",
  28048=>"101010100",
  28049=>"010111000",
  28050=>"001001101",
  28051=>"001111111",
  28052=>"100110001",
  28053=>"110000011",
  28054=>"101110111",
  28055=>"001111111",
  28056=>"110110100",
  28057=>"000101111",
  28058=>"100110011",
  28059=>"000000001",
  28060=>"011100000",
  28061=>"110010101",
  28062=>"111101001",
  28063=>"010010001",
  28064=>"101100110",
  28065=>"011100001",
  28066=>"001010100",
  28067=>"111011101",
  28068=>"001100001",
  28069=>"111111111",
  28070=>"001110010",
  28071=>"101111100",
  28072=>"011100100",
  28073=>"111001111",
  28074=>"001010110",
  28075=>"111001101",
  28076=>"010111010",
  28077=>"111010011",
  28078=>"011011110",
  28079=>"111110101",
  28080=>"001100011",
  28081=>"101111100",
  28082=>"100011101",
  28083=>"101010000",
  28084=>"000010001",
  28085=>"100010010",
  28086=>"111000111",
  28087=>"011001100",
  28088=>"011001011",
  28089=>"100111010",
  28090=>"101101001",
  28091=>"000001111",
  28092=>"101011110",
  28093=>"100101110",
  28094=>"101101110",
  28095=>"011010111",
  28096=>"101000010",
  28097=>"010000000",
  28098=>"111001100",
  28099=>"011100110",
  28100=>"100001100",
  28101=>"011000011",
  28102=>"010000001",
  28103=>"001000000",
  28104=>"001000111",
  28105=>"100101100",
  28106=>"000000100",
  28107=>"111001000",
  28108=>"111010110",
  28109=>"000101000",
  28110=>"000100010",
  28111=>"101011011",
  28112=>"001010000",
  28113=>"011100011",
  28114=>"010110110",
  28115=>"010111011",
  28116=>"000111100",
  28117=>"011110010",
  28118=>"110111111",
  28119=>"001010010",
  28120=>"001000010",
  28121=>"101011001",
  28122=>"010100111",
  28123=>"111100000",
  28124=>"101001001",
  28125=>"110011011",
  28126=>"000111110",
  28127=>"111100101",
  28128=>"001010000",
  28129=>"001101100",
  28130=>"100110110",
  28131=>"111001001",
  28132=>"100010111",
  28133=>"100000000",
  28134=>"010111001",
  28135=>"011000011",
  28136=>"111001000",
  28137=>"111111100",
  28138=>"000010000",
  28139=>"001111011",
  28140=>"000111011",
  28141=>"111100000",
  28142=>"110110100",
  28143=>"111100100",
  28144=>"110001111",
  28145=>"000001000",
  28146=>"100110101",
  28147=>"000000000",
  28148=>"001100010",
  28149=>"101000101",
  28150=>"010101111",
  28151=>"100001001",
  28152=>"001111111",
  28153=>"010010010",
  28154=>"111000100",
  28155=>"010011101",
  28156=>"101110100",
  28157=>"111100111",
  28158=>"101000101",
  28159=>"001111000",
  28160=>"000110010",
  28161=>"011101010",
  28162=>"101101101",
  28163=>"100010101",
  28164=>"101010111",
  28165=>"100101110",
  28166=>"111001011",
  28167=>"001000000",
  28168=>"011000010",
  28169=>"000011101",
  28170=>"111101010",
  28171=>"010000001",
  28172=>"010101000",
  28173=>"111100110",
  28174=>"111000011",
  28175=>"101111011",
  28176=>"000111101",
  28177=>"000110100",
  28178=>"101011000",
  28179=>"111011011",
  28180=>"101001111",
  28181=>"111001001",
  28182=>"111010101",
  28183=>"100100010",
  28184=>"101100001",
  28185=>"011111111",
  28186=>"011110101",
  28187=>"010010100",
  28188=>"011010111",
  28189=>"110010000",
  28190=>"111000001",
  28191=>"100001110",
  28192=>"100011100",
  28193=>"011000100",
  28194=>"111100100",
  28195=>"100010000",
  28196=>"001100111",
  28197=>"011101100",
  28198=>"100011001",
  28199=>"000010010",
  28200=>"011111101",
  28201=>"010001110",
  28202=>"101010010",
  28203=>"101110101",
  28204=>"011001000",
  28205=>"101010001",
  28206=>"011001100",
  28207=>"011101101",
  28208=>"011011101",
  28209=>"001101111",
  28210=>"010110010",
  28211=>"101000101",
  28212=>"001001000",
  28213=>"001000000",
  28214=>"101110000",
  28215=>"011000110",
  28216=>"111001111",
  28217=>"001111111",
  28218=>"101011010",
  28219=>"011100011",
  28220=>"010101111",
  28221=>"000000011",
  28222=>"011001010",
  28223=>"100100000",
  28224=>"100011010",
  28225=>"100101010",
  28226=>"101101110",
  28227=>"111011010",
  28228=>"010001000",
  28229=>"010010000",
  28230=>"101000000",
  28231=>"111111100",
  28232=>"001000110",
  28233=>"111011001",
  28234=>"100101111",
  28235=>"111101011",
  28236=>"010100000",
  28237=>"111101100",
  28238=>"000011110",
  28239=>"101010101",
  28240=>"111110010",
  28241=>"001000101",
  28242=>"101101111",
  28243=>"110111101",
  28244=>"000010000",
  28245=>"010000110",
  28246=>"100001101",
  28247=>"010101111",
  28248=>"111111001",
  28249=>"101000010",
  28250=>"101101101",
  28251=>"001000000",
  28252=>"111001101",
  28253=>"000000010",
  28254=>"101101010",
  28255=>"000011110",
  28256=>"011110100",
  28257=>"100101011",
  28258=>"111001000",
  28259=>"000000100",
  28260=>"000001110",
  28261=>"001001111",
  28262=>"000100001",
  28263=>"111001111",
  28264=>"110000111",
  28265=>"001011000",
  28266=>"110011000",
  28267=>"010010110",
  28268=>"111100001",
  28269=>"011001111",
  28270=>"111101001",
  28271=>"010001000",
  28272=>"000000101",
  28273=>"100010110",
  28274=>"011110001",
  28275=>"011000101",
  28276=>"100111100",
  28277=>"001111111",
  28278=>"011011111",
  28279=>"010100010",
  28280=>"111101101",
  28281=>"110000001",
  28282=>"101000101",
  28283=>"001011000",
  28284=>"100110110",
  28285=>"110110101",
  28286=>"111111101",
  28287=>"000000110",
  28288=>"110010111",
  28289=>"000111110",
  28290=>"000111000",
  28291=>"110111110",
  28292=>"001101001",
  28293=>"100010010",
  28294=>"101110101",
  28295=>"100100101",
  28296=>"101000010",
  28297=>"001100111",
  28298=>"011001110",
  28299=>"010101110",
  28300=>"001100000",
  28301=>"010001101",
  28302=>"111111111",
  28303=>"101010111",
  28304=>"011101011",
  28305=>"111000011",
  28306=>"011010011",
  28307=>"011000110",
  28308=>"111010000",
  28309=>"100100010",
  28310=>"011010110",
  28311=>"010100000",
  28312=>"001101111",
  28313=>"001010101",
  28314=>"001100000",
  28315=>"101111101",
  28316=>"001101001",
  28317=>"001110100",
  28318=>"011000101",
  28319=>"001111000",
  28320=>"011111111",
  28321=>"100111000",
  28322=>"010101111",
  28323=>"101100000",
  28324=>"000000111",
  28325=>"110101100",
  28326=>"111010111",
  28327=>"101001110",
  28328=>"101110100",
  28329=>"000000000",
  28330=>"001101100",
  28331=>"011000010",
  28332=>"111000000",
  28333=>"001010000",
  28334=>"010010000",
  28335=>"000111111",
  28336=>"111101110",
  28337=>"110100111",
  28338=>"101000111",
  28339=>"101100001",
  28340=>"110000010",
  28341=>"111111101",
  28342=>"111110110",
  28343=>"000011111",
  28344=>"101000011",
  28345=>"001101000",
  28346=>"111111100",
  28347=>"011000010",
  28348=>"011000101",
  28349=>"111101100",
  28350=>"101010001",
  28351=>"011111011",
  28352=>"111001000",
  28353=>"110000111",
  28354=>"111010000",
  28355=>"110100110",
  28356=>"000001100",
  28357=>"010001001",
  28358=>"100001011",
  28359=>"101111011",
  28360=>"010111100",
  28361=>"111010100",
  28362=>"010000101",
  28363=>"000010001",
  28364=>"100000110",
  28365=>"010110100",
  28366=>"010111101",
  28367=>"110111110",
  28368=>"010111001",
  28369=>"001001000",
  28370=>"010100011",
  28371=>"111100110",
  28372=>"111000011",
  28373=>"110001110",
  28374=>"110110000",
  28375=>"000111101",
  28376=>"100000100",
  28377=>"011001000",
  28378=>"111011111",
  28379=>"101001111",
  28380=>"000111110",
  28381=>"000001101",
  28382=>"110111011",
  28383=>"000101011",
  28384=>"111110110",
  28385=>"100100011",
  28386=>"111101101",
  28387=>"111001011",
  28388=>"010111011",
  28389=>"000000111",
  28390=>"110101110",
  28391=>"111001111",
  28392=>"000011101",
  28393=>"101010110",
  28394=>"010000010",
  28395=>"101010110",
  28396=>"000011101",
  28397=>"010101100",
  28398=>"011011111",
  28399=>"001110011",
  28400=>"111001111",
  28401=>"111011110",
  28402=>"111000101",
  28403=>"001100111",
  28404=>"111010010",
  28405=>"110100111",
  28406=>"001000100",
  28407=>"100111011",
  28408=>"110011001",
  28409=>"110010111",
  28410=>"101000011",
  28411=>"010010011",
  28412=>"100011100",
  28413=>"000011101",
  28414=>"111000000",
  28415=>"000000000",
  28416=>"110010010",
  28417=>"011110000",
  28418=>"110011001",
  28419=>"110001101",
  28420=>"001001000",
  28421=>"010011111",
  28422=>"011100100",
  28423=>"101101010",
  28424=>"100111101",
  28425=>"110101010",
  28426=>"110001110",
  28427=>"101100011",
  28428=>"011001001",
  28429=>"101100001",
  28430=>"001011010",
  28431=>"011111100",
  28432=>"110111011",
  28433=>"000000100",
  28434=>"111111110",
  28435=>"000110100",
  28436=>"000011100",
  28437=>"011110001",
  28438=>"110101011",
  28439=>"000001111",
  28440=>"001001100",
  28441=>"000100001",
  28442=>"000000101",
  28443=>"000100011",
  28444=>"011010110",
  28445=>"000111001",
  28446=>"110010011",
  28447=>"101100110",
  28448=>"010110110",
  28449=>"100101000",
  28450=>"110001100",
  28451=>"000001111",
  28452=>"111001011",
  28453=>"010101010",
  28454=>"111001010",
  28455=>"001100000",
  28456=>"010110000",
  28457=>"111010010",
  28458=>"001000001",
  28459=>"111111000",
  28460=>"101001010",
  28461=>"111101101",
  28462=>"100001000",
  28463=>"100011101",
  28464=>"101001111",
  28465=>"000101001",
  28466=>"101100010",
  28467=>"000001001",
  28468=>"010011011",
  28469=>"010011100",
  28470=>"000010001",
  28471=>"001111010",
  28472=>"010100101",
  28473=>"100001001",
  28474=>"011110011",
  28475=>"110010010",
  28476=>"111001101",
  28477=>"010111111",
  28478=>"110010111",
  28479=>"100000101",
  28480=>"001001101",
  28481=>"010100000",
  28482=>"000011111",
  28483=>"111001101",
  28484=>"010110011",
  28485=>"110100101",
  28486=>"001111111",
  28487=>"111101111",
  28488=>"100000010",
  28489=>"010001010",
  28490=>"100010010",
  28491=>"100000000",
  28492=>"010001101",
  28493=>"111010010",
  28494=>"001110100",
  28495=>"001010010",
  28496=>"010111000",
  28497=>"000001111",
  28498=>"000001010",
  28499=>"100110101",
  28500=>"101000000",
  28501=>"000111010",
  28502=>"010111011",
  28503=>"000100110",
  28504=>"000100101",
  28505=>"100010100",
  28506=>"010011110",
  28507=>"000010101",
  28508=>"110001100",
  28509=>"100011110",
  28510=>"111111110",
  28511=>"001000010",
  28512=>"011001111",
  28513=>"000001010",
  28514=>"110011100",
  28515=>"111011001",
  28516=>"010111001",
  28517=>"001000100",
  28518=>"000101000",
  28519=>"111100110",
  28520=>"100101011",
  28521=>"100110100",
  28522=>"011110011",
  28523=>"101101111",
  28524=>"100101110",
  28525=>"001011011",
  28526=>"100100011",
  28527=>"011101010",
  28528=>"000011101",
  28529=>"000001110",
  28530=>"001100100",
  28531=>"110111100",
  28532=>"101010110",
  28533=>"000000011",
  28534=>"101110001",
  28535=>"100011000",
  28536=>"110000011",
  28537=>"110111000",
  28538=>"111101100",
  28539=>"011100000",
  28540=>"111111101",
  28541=>"101000100",
  28542=>"100000101",
  28543=>"110111111",
  28544=>"010100010",
  28545=>"111100101",
  28546=>"110110101",
  28547=>"011100011",
  28548=>"100010010",
  28549=>"001001010",
  28550=>"001111011",
  28551=>"101010100",
  28552=>"111010110",
  28553=>"011100111",
  28554=>"111101000",
  28555=>"000000000",
  28556=>"011001101",
  28557=>"110101001",
  28558=>"110010101",
  28559=>"101111000",
  28560=>"100001110",
  28561=>"011111010",
  28562=>"100101100",
  28563=>"011011110",
  28564=>"001100001",
  28565=>"110111001",
  28566=>"010001010",
  28567=>"000001100",
  28568=>"011100001",
  28569=>"110011101",
  28570=>"101100001",
  28571=>"100111010",
  28572=>"111010111",
  28573=>"001010111",
  28574=>"000001100",
  28575=>"101111000",
  28576=>"010101110",
  28577=>"001110010",
  28578=>"101111101",
  28579=>"010001011",
  28580=>"100111110",
  28581=>"110111000",
  28582=>"011111001",
  28583=>"110100000",
  28584=>"000000000",
  28585=>"000001111",
  28586=>"111010101",
  28587=>"011100111",
  28588=>"001000100",
  28589=>"001011000",
  28590=>"111001010",
  28591=>"100010000",
  28592=>"010000010",
  28593=>"010100110",
  28594=>"011010110",
  28595=>"001100101",
  28596=>"001010101",
  28597=>"101101110",
  28598=>"000010101",
  28599=>"111010110",
  28600=>"011001100",
  28601=>"010100111",
  28602=>"000111000",
  28603=>"110100001",
  28604=>"001011101",
  28605=>"000001000",
  28606=>"011001011",
  28607=>"101001000",
  28608=>"100110001",
  28609=>"111110011",
  28610=>"101011001",
  28611=>"110110000",
  28612=>"110110100",
  28613=>"001100011",
  28614=>"100100001",
  28615=>"100000111",
  28616=>"001010000",
  28617=>"010010101",
  28618=>"111101001",
  28619=>"001010110",
  28620=>"010001000",
  28621=>"000010010",
  28622=>"011001100",
  28623=>"001001110",
  28624=>"101111011",
  28625=>"000000111",
  28626=>"010110101",
  28627=>"110100000",
  28628=>"010011000",
  28629=>"111111101",
  28630=>"111101100",
  28631=>"011001001",
  28632=>"111111100",
  28633=>"001100001",
  28634=>"000110000",
  28635=>"001101111",
  28636=>"110000110",
  28637=>"001011111",
  28638=>"100001101",
  28639=>"101000100",
  28640=>"110011110",
  28641=>"000010011",
  28642=>"111010000",
  28643=>"001100101",
  28644=>"101111001",
  28645=>"111111100",
  28646=>"001001011",
  28647=>"110100000",
  28648=>"101011100",
  28649=>"100100101",
  28650=>"011010001",
  28651=>"101010111",
  28652=>"010000001",
  28653=>"111010101",
  28654=>"000101100",
  28655=>"110110100",
  28656=>"000101101",
  28657=>"101100100",
  28658=>"000100010",
  28659=>"010111101",
  28660=>"111010011",
  28661=>"001010110",
  28662=>"010111000",
  28663=>"101000000",
  28664=>"101010111",
  28665=>"000000110",
  28666=>"111101111",
  28667=>"001111110",
  28668=>"111110000",
  28669=>"000000000",
  28670=>"110001010",
  28671=>"010000011",
  28672=>"110100011",
  28673=>"000100010",
  28674=>"110011101",
  28675=>"101111011",
  28676=>"011001011",
  28677=>"110010001",
  28678=>"001000110",
  28679=>"100110100",
  28680=>"110101111",
  28681=>"110101101",
  28682=>"001001111",
  28683=>"111000001",
  28684=>"010010111",
  28685=>"001101111",
  28686=>"100001100",
  28687=>"000100010",
  28688=>"010011110",
  28689=>"101010010",
  28690=>"010110111",
  28691=>"010010110",
  28692=>"001100011",
  28693=>"001100000",
  28694=>"111101001",
  28695=>"000011100",
  28696=>"011100100",
  28697=>"100000011",
  28698=>"010010101",
  28699=>"000100001",
  28700=>"110100000",
  28701=>"110111101",
  28702=>"111100011",
  28703=>"111011010",
  28704=>"110101110",
  28705=>"000010011",
  28706=>"011100000",
  28707=>"100011001",
  28708=>"000010010",
  28709=>"100001001",
  28710=>"000010000",
  28711=>"110001111",
  28712=>"110000111",
  28713=>"111011001",
  28714=>"110100000",
  28715=>"111101111",
  28716=>"010000100",
  28717=>"110001101",
  28718=>"100101001",
  28719=>"100100000",
  28720=>"001001010",
  28721=>"011110010",
  28722=>"001100011",
  28723=>"011100111",
  28724=>"010101011",
  28725=>"000000010",
  28726=>"000101000",
  28727=>"100000000",
  28728=>"000100111",
  28729=>"100010001",
  28730=>"000011010",
  28731=>"100000010",
  28732=>"111110000",
  28733=>"101111101",
  28734=>"011000000",
  28735=>"000001100",
  28736=>"000100111",
  28737=>"110001001",
  28738=>"100110111",
  28739=>"111000100",
  28740=>"100110000",
  28741=>"111101101",
  28742=>"111011111",
  28743=>"010000100",
  28744=>"101000101",
  28745=>"000001110",
  28746=>"010011100",
  28747=>"010000011",
  28748=>"101001100",
  28749=>"001110110",
  28750=>"000101100",
  28751=>"110101101",
  28752=>"001010000",
  28753=>"000000011",
  28754=>"111010011",
  28755=>"101000111",
  28756=>"111000011",
  28757=>"001010010",
  28758=>"111010000",
  28759=>"111000101",
  28760=>"111000011",
  28761=>"101101111",
  28762=>"111001000",
  28763=>"101100110",
  28764=>"111100100",
  28765=>"000000011",
  28766=>"110100010",
  28767=>"111100101",
  28768=>"100010111",
  28769=>"010111111",
  28770=>"010000001",
  28771=>"100100100",
  28772=>"011111100",
  28773=>"101101110",
  28774=>"101111111",
  28775=>"001001001",
  28776=>"110110101",
  28777=>"111111001",
  28778=>"010100101",
  28779=>"000001000",
  28780=>"001001001",
  28781=>"000111001",
  28782=>"100011111",
  28783=>"000100000",
  28784=>"101110110",
  28785=>"001000100",
  28786=>"001111001",
  28787=>"110011111",
  28788=>"110010000",
  28789=>"100111100",
  28790=>"011100010",
  28791=>"010101110",
  28792=>"100001010",
  28793=>"100000100",
  28794=>"110111100",
  28795=>"000101011",
  28796=>"101111000",
  28797=>"010111000",
  28798=>"010000110",
  28799=>"100010111",
  28800=>"101010100",
  28801=>"111010101",
  28802=>"111000100",
  28803=>"010110010",
  28804=>"010100001",
  28805=>"110001110",
  28806=>"110101100",
  28807=>"000010111",
  28808=>"110101110",
  28809=>"100000000",
  28810=>"100001001",
  28811=>"110010101",
  28812=>"001111001",
  28813=>"000101101",
  28814=>"100010101",
  28815=>"000011011",
  28816=>"011001110",
  28817=>"011001100",
  28818=>"101101001",
  28819=>"111010001",
  28820=>"010001101",
  28821=>"010110000",
  28822=>"010100110",
  28823=>"010001000",
  28824=>"111100111",
  28825=>"110111011",
  28826=>"001011011",
  28827=>"101011111",
  28828=>"000110010",
  28829=>"100100000",
  28830=>"110000010",
  28831=>"111110011",
  28832=>"011111100",
  28833=>"001000111",
  28834=>"110111001",
  28835=>"110000010",
  28836=>"001010101",
  28837=>"010100000",
  28838=>"011100010",
  28839=>"011100111",
  28840=>"101000001",
  28841=>"111110010",
  28842=>"001011110",
  28843=>"000111100",
  28844=>"010100001",
  28845=>"101101110",
  28846=>"101110110",
  28847=>"100000100",
  28848=>"110101001",
  28849=>"010001000",
  28850=>"101100101",
  28851=>"111001111",
  28852=>"000000001",
  28853=>"011110000",
  28854=>"111111100",
  28855=>"001010010",
  28856=>"001100011",
  28857=>"111101011",
  28858=>"000001001",
  28859=>"010000100",
  28860=>"010011001",
  28861=>"011001010",
  28862=>"111101111",
  28863=>"001111000",
  28864=>"001111011",
  28865=>"000011101",
  28866=>"100001101",
  28867=>"001100100",
  28868=>"011101101",
  28869=>"101011111",
  28870=>"110001111",
  28871=>"110110110",
  28872=>"110011101",
  28873=>"101110000",
  28874=>"011011000",
  28875=>"000011110",
  28876=>"111101011",
  28877=>"000001000",
  28878=>"011011001",
  28879=>"010111010",
  28880=>"001110111",
  28881=>"111101111",
  28882=>"011111010",
  28883=>"010010111",
  28884=>"111000011",
  28885=>"000110000",
  28886=>"101011111",
  28887=>"111011010",
  28888=>"001101010",
  28889=>"001000000",
  28890=>"011100011",
  28891=>"111100111",
  28892=>"010101101",
  28893=>"011001001",
  28894=>"111001011",
  28895=>"000110001",
  28896=>"101000011",
  28897=>"100011011",
  28898=>"111001101",
  28899=>"110101010",
  28900=>"000010001",
  28901=>"110000100",
  28902=>"001010100",
  28903=>"000010101",
  28904=>"100000010",
  28905=>"100010001",
  28906=>"000100110",
  28907=>"101111000",
  28908=>"111010000",
  28909=>"001101100",
  28910=>"001100000",
  28911=>"100101000",
  28912=>"000101010",
  28913=>"010101110",
  28914=>"001100100",
  28915=>"110010100",
  28916=>"000110010",
  28917=>"010010000",
  28918=>"110110110",
  28919=>"100000000",
  28920=>"100011111",
  28921=>"010101010",
  28922=>"010010101",
  28923=>"010000111",
  28924=>"101000000",
  28925=>"110100110",
  28926=>"000001001",
  28927=>"010010001",
  28928=>"010100110",
  28929=>"111110111",
  28930=>"011001100",
  28931=>"000110110",
  28932=>"001001011",
  28933=>"110000111",
  28934=>"000101001",
  28935=>"011000000",
  28936=>"110001010",
  28937=>"101001110",
  28938=>"010000100",
  28939=>"111110101",
  28940=>"101000110",
  28941=>"101101000",
  28942=>"101110011",
  28943=>"110010110",
  28944=>"101011110",
  28945=>"111111001",
  28946=>"010010000",
  28947=>"100010110",
  28948=>"110100101",
  28949=>"011011001",
  28950=>"001011001",
  28951=>"110010111",
  28952=>"000111111",
  28953=>"110011111",
  28954=>"111010110",
  28955=>"001011000",
  28956=>"111001000",
  28957=>"101010011",
  28958=>"111111101",
  28959=>"010111000",
  28960=>"001110001",
  28961=>"111101001",
  28962=>"001010110",
  28963=>"000101011",
  28964=>"101010001",
  28965=>"101001011",
  28966=>"000100011",
  28967=>"101111101",
  28968=>"100001010",
  28969=>"111010100",
  28970=>"110001010",
  28971=>"100001100",
  28972=>"100100011",
  28973=>"111101011",
  28974=>"100000010",
  28975=>"111100001",
  28976=>"111000100",
  28977=>"101001000",
  28978=>"111011101",
  28979=>"000011000",
  28980=>"001110110",
  28981=>"000010011",
  28982=>"010000100",
  28983=>"000100000",
  28984=>"110110100",
  28985=>"000011000",
  28986=>"010101001",
  28987=>"111101000",
  28988=>"011111101",
  28989=>"001110101",
  28990=>"101000010",
  28991=>"010101011",
  28992=>"011100011",
  28993=>"110111101",
  28994=>"011010001",
  28995=>"011011011",
  28996=>"001110101",
  28997=>"100001100",
  28998=>"011010100",
  28999=>"000000011",
  29000=>"111111101",
  29001=>"010001001",
  29002=>"001011100",
  29003=>"110111111",
  29004=>"111101101",
  29005=>"011000011",
  29006=>"000001011",
  29007=>"000111001",
  29008=>"111101001",
  29009=>"000101101",
  29010=>"010010000",
  29011=>"010111111",
  29012=>"100010111",
  29013=>"110011101",
  29014=>"000001101",
  29015=>"000010001",
  29016=>"001010100",
  29017=>"000000000",
  29018=>"010101000",
  29019=>"111101011",
  29020=>"100110110",
  29021=>"001001100",
  29022=>"000001010",
  29023=>"001010011",
  29024=>"101010110",
  29025=>"111110000",
  29026=>"111111011",
  29027=>"000011110",
  29028=>"110111110",
  29029=>"101000011",
  29030=>"001010101",
  29031=>"010000000",
  29032=>"101000100",
  29033=>"111101111",
  29034=>"000000010",
  29035=>"000100100",
  29036=>"011010011",
  29037=>"101111100",
  29038=>"000010010",
  29039=>"010110100",
  29040=>"101100011",
  29041=>"011011001",
  29042=>"000110001",
  29043=>"101100110",
  29044=>"100001011",
  29045=>"011100000",
  29046=>"000111110",
  29047=>"110000010",
  29048=>"010100101",
  29049=>"101111011",
  29050=>"000001000",
  29051=>"110110001",
  29052=>"011110011",
  29053=>"000100001",
  29054=>"001010111",
  29055=>"010101111",
  29056=>"101111101",
  29057=>"011111001",
  29058=>"110101111",
  29059=>"101000010",
  29060=>"111011000",
  29061=>"011111101",
  29062=>"100101110",
  29063=>"110011000",
  29064=>"100000101",
  29065=>"010010001",
  29066=>"001011100",
  29067=>"000011011",
  29068=>"011001000",
  29069=>"011111001",
  29070=>"001000111",
  29071=>"101001011",
  29072=>"010111111",
  29073=>"100000011",
  29074=>"111101010",
  29075=>"001001101",
  29076=>"000011100",
  29077=>"010101000",
  29078=>"010010001",
  29079=>"111000011",
  29080=>"000001000",
  29081=>"010101111",
  29082=>"111001011",
  29083=>"010000001",
  29084=>"010001000",
  29085=>"001101111",
  29086=>"011100100",
  29087=>"001111011",
  29088=>"000011001",
  29089=>"100100001",
  29090=>"100001100",
  29091=>"100001111",
  29092=>"010010101",
  29093=>"110000011",
  29094=>"000101000",
  29095=>"101111110",
  29096=>"001000111",
  29097=>"100101100",
  29098=>"000011010",
  29099=>"101110101",
  29100=>"100111110",
  29101=>"101101111",
  29102=>"010011010",
  29103=>"111010100",
  29104=>"101101100",
  29105=>"011001000",
  29106=>"111000010",
  29107=>"011010010",
  29108=>"101100000",
  29109=>"011011100",
  29110=>"000110011",
  29111=>"110010111",
  29112=>"000100110",
  29113=>"100111010",
  29114=>"101111101",
  29115=>"000110011",
  29116=>"010001010",
  29117=>"001001001",
  29118=>"100000000",
  29119=>"101010111",
  29120=>"100000111",
  29121=>"111111100",
  29122=>"010000011",
  29123=>"011111110",
  29124=>"011001110",
  29125=>"111100001",
  29126=>"000010101",
  29127=>"101110111",
  29128=>"010100101",
  29129=>"001011010",
  29130=>"001000001",
  29131=>"111001100",
  29132=>"000101111",
  29133=>"010001011",
  29134=>"011001010",
  29135=>"110110010",
  29136=>"001001010",
  29137=>"101101001",
  29138=>"100101011",
  29139=>"000101000",
  29140=>"010000010",
  29141=>"001110011",
  29142=>"110010101",
  29143=>"110001111",
  29144=>"111001001",
  29145=>"000000010",
  29146=>"000100000",
  29147=>"011111011",
  29148=>"111001100",
  29149=>"111110011",
  29150=>"110111100",
  29151=>"011100110",
  29152=>"100100101",
  29153=>"000100101",
  29154=>"110111010",
  29155=>"110111000",
  29156=>"110001111",
  29157=>"110101001",
  29158=>"011111111",
  29159=>"000010100",
  29160=>"110111110",
  29161=>"111010101",
  29162=>"000010000",
  29163=>"110001011",
  29164=>"100001101",
  29165=>"101100000",
  29166=>"110110000",
  29167=>"011110010",
  29168=>"001101001",
  29169=>"010011110",
  29170=>"110011011",
  29171=>"010011010",
  29172=>"111100111",
  29173=>"100000000",
  29174=>"001101010",
  29175=>"100011100",
  29176=>"101100110",
  29177=>"001001101",
  29178=>"000010010",
  29179=>"101000010",
  29180=>"010110010",
  29181=>"010001100",
  29182=>"000001100",
  29183=>"001011111",
  29184=>"000100011",
  29185=>"101010111",
  29186=>"010010000",
  29187=>"111001100",
  29188=>"001100111",
  29189=>"101000010",
  29190=>"110110101",
  29191=>"011011001",
  29192=>"111001110",
  29193=>"000010011",
  29194=>"001100110",
  29195=>"011011110",
  29196=>"001110001",
  29197=>"001111111",
  29198=>"000110011",
  29199=>"011000100",
  29200=>"100101010",
  29201=>"101111000",
  29202=>"010010111",
  29203=>"011010110",
  29204=>"010111101",
  29205=>"000111111",
  29206=>"011011010",
  29207=>"011011010",
  29208=>"000111111",
  29209=>"110001000",
  29210=>"111111011",
  29211=>"100100100",
  29212=>"011101001",
  29213=>"101000011",
  29214=>"000110110",
  29215=>"000000001",
  29216=>"111010011",
  29217=>"001101111",
  29218=>"110000110",
  29219=>"011110111",
  29220=>"011101110",
  29221=>"001101001",
  29222=>"100100111",
  29223=>"000010011",
  29224=>"110111110",
  29225=>"101111101",
  29226=>"111101011",
  29227=>"110011111",
  29228=>"011101110",
  29229=>"110010001",
  29230=>"110000010",
  29231=>"010111010",
  29232=>"101111000",
  29233=>"111010001",
  29234=>"001110010",
  29235=>"101001001",
  29236=>"100111111",
  29237=>"101110010",
  29238=>"010110010",
  29239=>"110001101",
  29240=>"001110111",
  29241=>"010101010",
  29242=>"010110101",
  29243=>"111000000",
  29244=>"101001001",
  29245=>"001111100",
  29246=>"101101111",
  29247=>"010000000",
  29248=>"111011001",
  29249=>"100100111",
  29250=>"010001010",
  29251=>"011001101",
  29252=>"111001100",
  29253=>"110000001",
  29254=>"100100010",
  29255=>"000101111",
  29256=>"011111011",
  29257=>"101011100",
  29258=>"111010000",
  29259=>"010000011",
  29260=>"011000001",
  29261=>"100011110",
  29262=>"101111100",
  29263=>"100110111",
  29264=>"110110011",
  29265=>"111001001",
  29266=>"010010000",
  29267=>"001001001",
  29268=>"000000010",
  29269=>"000000000",
  29270=>"111100111",
  29271=>"011100000",
  29272=>"111111111",
  29273=>"100100100",
  29274=>"110001101",
  29275=>"000010110",
  29276=>"000000001",
  29277=>"011000111",
  29278=>"000011101",
  29279=>"100111111",
  29280=>"001100011",
  29281=>"011100110",
  29282=>"100011010",
  29283=>"100010101",
  29284=>"011100101",
  29285=>"101100010",
  29286=>"101010101",
  29287=>"100001101",
  29288=>"110110111",
  29289=>"110010110",
  29290=>"010100110",
  29291=>"111110111",
  29292=>"100000101",
  29293=>"101100001",
  29294=>"010110011",
  29295=>"111010100",
  29296=>"111101110",
  29297=>"010100001",
  29298=>"001010100",
  29299=>"110011011",
  29300=>"100100000",
  29301=>"000101110",
  29302=>"101101010",
  29303=>"110111111",
  29304=>"010010111",
  29305=>"000001100",
  29306=>"100001010",
  29307=>"110111001",
  29308=>"010001101",
  29309=>"100110111",
  29310=>"100000001",
  29311=>"000011110",
  29312=>"011000001",
  29313=>"001010000",
  29314=>"000001000",
  29315=>"001110100",
  29316=>"010000100",
  29317=>"010001111",
  29318=>"100010111",
  29319=>"110011110",
  29320=>"010010001",
  29321=>"000010000",
  29322=>"111010110",
  29323=>"001001100",
  29324=>"000101100",
  29325=>"111011000",
  29326=>"010100111",
  29327=>"000000001",
  29328=>"100110011",
  29329=>"100011001",
  29330=>"010001110",
  29331=>"110010100",
  29332=>"000001001",
  29333=>"000111010",
  29334=>"001001101",
  29335=>"011001110",
  29336=>"000000001",
  29337=>"111100111",
  29338=>"011111010",
  29339=>"011001111",
  29340=>"101110001",
  29341=>"111111100",
  29342=>"011011001",
  29343=>"100101111",
  29344=>"000011110",
  29345=>"010010000",
  29346=>"100101100",
  29347=>"100001111",
  29348=>"100011111",
  29349=>"101010011",
  29350=>"001010101",
  29351=>"011010111",
  29352=>"100001000",
  29353=>"010101101",
  29354=>"110011001",
  29355=>"000000101",
  29356=>"111011111",
  29357=>"100000000",
  29358=>"101110011",
  29359=>"101101010",
  29360=>"111111111",
  29361=>"101111100",
  29362=>"110011111",
  29363=>"010110111",
  29364=>"010100010",
  29365=>"000010101",
  29366=>"001001100",
  29367=>"010101101",
  29368=>"011010101",
  29369=>"000110111",
  29370=>"101011001",
  29371=>"100111011",
  29372=>"010010010",
  29373=>"001100000",
  29374=>"111101110",
  29375=>"110000100",
  29376=>"011101000",
  29377=>"110000011",
  29378=>"010010001",
  29379=>"000011000",
  29380=>"000110110",
  29381=>"000111111",
  29382=>"101100111",
  29383=>"101010111",
  29384=>"100110100",
  29385=>"110011011",
  29386=>"001000000",
  29387=>"111001000",
  29388=>"100010001",
  29389=>"101111100",
  29390=>"011110101",
  29391=>"110100000",
  29392=>"011011010",
  29393=>"001010110",
  29394=>"110111100",
  29395=>"000110010",
  29396=>"001000001",
  29397=>"111111100",
  29398=>"101011101",
  29399=>"000010100",
  29400=>"000000000",
  29401=>"001011110",
  29402=>"110011000",
  29403=>"010111010",
  29404=>"110001000",
  29405=>"000001101",
  29406=>"000001010",
  29407=>"000001111",
  29408=>"010110000",
  29409=>"101110110",
  29410=>"100100010",
  29411=>"001000100",
  29412=>"000000010",
  29413=>"011101010",
  29414=>"101001110",
  29415=>"000000110",
  29416=>"001100010",
  29417=>"001000001",
  29418=>"000001001",
  29419=>"111001011",
  29420=>"001001101",
  29421=>"010110111",
  29422=>"100000111",
  29423=>"111011111",
  29424=>"111111110",
  29425=>"100000100",
  29426=>"000010011",
  29427=>"011001001",
  29428=>"110111101",
  29429=>"000100010",
  29430=>"010110100",
  29431=>"101001000",
  29432=>"001100001",
  29433=>"101101000",
  29434=>"010101111",
  29435=>"000100000",
  29436=>"101011010",
  29437=>"010000100",
  29438=>"110110111",
  29439=>"011110011",
  29440=>"010000001",
  29441=>"101010110",
  29442=>"100101000",
  29443=>"110110001",
  29444=>"011001101",
  29445=>"000110011",
  29446=>"011100111",
  29447=>"010001101",
  29448=>"101110111",
  29449=>"101000011",
  29450=>"010011010",
  29451=>"010111100",
  29452=>"011011111",
  29453=>"000111111",
  29454=>"101100100",
  29455=>"111101100",
  29456=>"010011111",
  29457=>"000010101",
  29458=>"100110000",
  29459=>"100110010",
  29460=>"001001010",
  29461=>"111001111",
  29462=>"000111011",
  29463=>"011001000",
  29464=>"111010001",
  29465=>"011100111",
  29466=>"010010101",
  29467=>"010110011",
  29468=>"111111101",
  29469=>"100110010",
  29470=>"100010000",
  29471=>"110001001",
  29472=>"110111000",
  29473=>"001100111",
  29474=>"011100111",
  29475=>"110111110",
  29476=>"011001001",
  29477=>"000000110",
  29478=>"000000010",
  29479=>"011111011",
  29480=>"010111011",
  29481=>"111101001",
  29482=>"101011011",
  29483=>"111110011",
  29484=>"110110010",
  29485=>"101000000",
  29486=>"000100001",
  29487=>"111000000",
  29488=>"110010101",
  29489=>"011000110",
  29490=>"010000110",
  29491=>"111000001",
  29492=>"101111011",
  29493=>"010110011",
  29494=>"011101001",
  29495=>"011100110",
  29496=>"110000111",
  29497=>"001110000",
  29498=>"001011011",
  29499=>"011101011",
  29500=>"011111110",
  29501=>"101010010",
  29502=>"111100011",
  29503=>"010110111",
  29504=>"001001111",
  29505=>"011100101",
  29506=>"100111101",
  29507=>"111100101",
  29508=>"000011100",
  29509=>"010011100",
  29510=>"101001010",
  29511=>"000001000",
  29512=>"011110001",
  29513=>"110000010",
  29514=>"110101001",
  29515=>"011011010",
  29516=>"011011000",
  29517=>"001111110",
  29518=>"110100110",
  29519=>"001010000",
  29520=>"110010000",
  29521=>"111101011",
  29522=>"100101011",
  29523=>"101101011",
  29524=>"100100100",
  29525=>"110101010",
  29526=>"101000000",
  29527=>"001110000",
  29528=>"101010111",
  29529=>"000000111",
  29530=>"001101000",
  29531=>"011111000",
  29532=>"100111010",
  29533=>"101010100",
  29534=>"100111001",
  29535=>"000000000",
  29536=>"001011000",
  29537=>"010000000",
  29538=>"010111010",
  29539=>"000100110",
  29540=>"000000010",
  29541=>"101100000",
  29542=>"001010010",
  29543=>"001110001",
  29544=>"010110011",
  29545=>"001000000",
  29546=>"110101001",
  29547=>"110001011",
  29548=>"100001011",
  29549=>"110101110",
  29550=>"101011011",
  29551=>"001110001",
  29552=>"100011111",
  29553=>"101011011",
  29554=>"001101011",
  29555=>"101011110",
  29556=>"010010110",
  29557=>"110110001",
  29558=>"011101011",
  29559=>"011111000",
  29560=>"000001011",
  29561=>"010101010",
  29562=>"101100010",
  29563=>"101010110",
  29564=>"000011010",
  29565=>"011001011",
  29566=>"101000100",
  29567=>"101011011",
  29568=>"000001010",
  29569=>"110111010",
  29570=>"110010110",
  29571=>"100000111",
  29572=>"010110101",
  29573=>"000101100",
  29574=>"000010000",
  29575=>"101000100",
  29576=>"111000110",
  29577=>"111001000",
  29578=>"010000011",
  29579=>"001101001",
  29580=>"111011111",
  29581=>"100011000",
  29582=>"001010110",
  29583=>"101001100",
  29584=>"001010101",
  29585=>"101101001",
  29586=>"111010110",
  29587=>"111000001",
  29588=>"100011101",
  29589=>"111000000",
  29590=>"000010011",
  29591=>"010000011",
  29592=>"001011101",
  29593=>"100101011",
  29594=>"000010000",
  29595=>"001011110",
  29596=>"011011110",
  29597=>"011000110",
  29598=>"010100100",
  29599=>"010100001",
  29600=>"010010010",
  29601=>"111111111",
  29602=>"111101111",
  29603=>"110010101",
  29604=>"100011100",
  29605=>"000010100",
  29606=>"010100110",
  29607=>"010111011",
  29608=>"111001100",
  29609=>"000101110",
  29610=>"000011001",
  29611=>"001101111",
  29612=>"100111101",
  29613=>"100001000",
  29614=>"011010101",
  29615=>"010001001",
  29616=>"001100000",
  29617=>"111000010",
  29618=>"001100011",
  29619=>"111000010",
  29620=>"000000001",
  29621=>"000110010",
  29622=>"000110100",
  29623=>"101100010",
  29624=>"101010010",
  29625=>"111010001",
  29626=>"101111110",
  29627=>"110100011",
  29628=>"010001010",
  29629=>"010111000",
  29630=>"011101111",
  29631=>"000000011",
  29632=>"000110101",
  29633=>"001011111",
  29634=>"000111000",
  29635=>"111010000",
  29636=>"000000011",
  29637=>"111010111",
  29638=>"010000000",
  29639=>"111111110",
  29640=>"000001110",
  29641=>"100111100",
  29642=>"001111000",
  29643=>"000100110",
  29644=>"010111100",
  29645=>"101011001",
  29646=>"111000111",
  29647=>"110001000",
  29648=>"111011011",
  29649=>"000111100",
  29650=>"110111110",
  29651=>"011010010",
  29652=>"010100110",
  29653=>"110111001",
  29654=>"110000111",
  29655=>"000001000",
  29656=>"110111110",
  29657=>"010010001",
  29658=>"110111000",
  29659=>"011011001",
  29660=>"101011110",
  29661=>"100000110",
  29662=>"000111011",
  29663=>"100010101",
  29664=>"011111010",
  29665=>"011100010",
  29666=>"000010000",
  29667=>"010001110",
  29668=>"010000010",
  29669=>"110110111",
  29670=>"010001000",
  29671=>"011011101",
  29672=>"111010011",
  29673=>"110010000",
  29674=>"010010010",
  29675=>"011010011",
  29676=>"010001010",
  29677=>"111101110",
  29678=>"100101010",
  29679=>"011001100",
  29680=>"001111100",
  29681=>"111000000",
  29682=>"100001111",
  29683=>"101110110",
  29684=>"110101110",
  29685=>"111010010",
  29686=>"011110110",
  29687=>"110010111",
  29688=>"001111001",
  29689=>"000100100",
  29690=>"101011011",
  29691=>"101111101",
  29692=>"001110101",
  29693=>"010011110",
  29694=>"100100001",
  29695=>"011000110",
  29696=>"001010000",
  29697=>"100001000",
  29698=>"111110010",
  29699=>"010001001",
  29700=>"100000100",
  29701=>"110011101",
  29702=>"011100001",
  29703=>"101000111",
  29704=>"110001100",
  29705=>"111000010",
  29706=>"011010100",
  29707=>"101010000",
  29708=>"011000011",
  29709=>"011101101",
  29710=>"101111101",
  29711=>"101001000",
  29712=>"100011010",
  29713=>"101011000",
  29714=>"000111100",
  29715=>"100011001",
  29716=>"100001111",
  29717=>"000110010",
  29718=>"011101001",
  29719=>"001100000",
  29720=>"001100001",
  29721=>"010011100",
  29722=>"111000000",
  29723=>"001111010",
  29724=>"111000110",
  29725=>"111001101",
  29726=>"101000110",
  29727=>"101011000",
  29728=>"001010010",
  29729=>"011000111",
  29730=>"000001010",
  29731=>"011001101",
  29732=>"011011011",
  29733=>"110001010",
  29734=>"110011000",
  29735=>"110111101",
  29736=>"011101011",
  29737=>"010110000",
  29738=>"000100100",
  29739=>"110110011",
  29740=>"100000111",
  29741=>"100110111",
  29742=>"101000010",
  29743=>"111011010",
  29744=>"001000010",
  29745=>"111110010",
  29746=>"100110001",
  29747=>"011010000",
  29748=>"110101110",
  29749=>"100011011",
  29750=>"001100000",
  29751=>"010101100",
  29752=>"110010000",
  29753=>"001110010",
  29754=>"000111010",
  29755=>"110011011",
  29756=>"101100111",
  29757=>"110001000",
  29758=>"000011111",
  29759=>"010001101",
  29760=>"010110011",
  29761=>"111000001",
  29762=>"100110010",
  29763=>"010000011",
  29764=>"110010010",
  29765=>"101000011",
  29766=>"011101011",
  29767=>"101110000",
  29768=>"100011101",
  29769=>"010100101",
  29770=>"010001110",
  29771=>"001111011",
  29772=>"111010001",
  29773=>"101010111",
  29774=>"011101111",
  29775=>"000011010",
  29776=>"111101100",
  29777=>"000100100",
  29778=>"110000110",
  29779=>"111110100",
  29780=>"111011010",
  29781=>"011100110",
  29782=>"011011010",
  29783=>"101010010",
  29784=>"100011110",
  29785=>"110111101",
  29786=>"001000100",
  29787=>"000000110",
  29788=>"001110010",
  29789=>"000111010",
  29790=>"110111000",
  29791=>"100110110",
  29792=>"011010111",
  29793=>"101100000",
  29794=>"001011110",
  29795=>"111110110",
  29796=>"110111000",
  29797=>"110111101",
  29798=>"010111000",
  29799=>"100000011",
  29800=>"001011010",
  29801=>"011101011",
  29802=>"000011101",
  29803=>"111010000",
  29804=>"111001011",
  29805=>"000100010",
  29806=>"101101100",
  29807=>"010011001",
  29808=>"111100110",
  29809=>"000101001",
  29810=>"010111111",
  29811=>"101111101",
  29812=>"111011101",
  29813=>"010101111",
  29814=>"111101011",
  29815=>"111101011",
  29816=>"011001011",
  29817=>"110101010",
  29818=>"001100110",
  29819=>"011001001",
  29820=>"101000111",
  29821=>"101111100",
  29822=>"111111001",
  29823=>"010000110",
  29824=>"010100001",
  29825=>"100101011",
  29826=>"011011011",
  29827=>"011111110",
  29828=>"001011001",
  29829=>"010100101",
  29830=>"001011010",
  29831=>"010111010",
  29832=>"110100110",
  29833=>"111100101",
  29834=>"010011100",
  29835=>"100111000",
  29836=>"101011111",
  29837=>"100100010",
  29838=>"110000000",
  29839=>"011011011",
  29840=>"100110000",
  29841=>"000000001",
  29842=>"110001110",
  29843=>"010110100",
  29844=>"101110110",
  29845=>"001110111",
  29846=>"100011010",
  29847=>"000100011",
  29848=>"111111111",
  29849=>"101100100",
  29850=>"111100011",
  29851=>"111101001",
  29852=>"000101111",
  29853=>"110100111",
  29854=>"010100101",
  29855=>"010110010",
  29856=>"101111010",
  29857=>"011010011",
  29858=>"100011010",
  29859=>"011110101",
  29860=>"011111011",
  29861=>"101110100",
  29862=>"011101110",
  29863=>"010011001",
  29864=>"011001111",
  29865=>"100011110",
  29866=>"110101010",
  29867=>"001100001",
  29868=>"001000101",
  29869=>"100110111",
  29870=>"000101000",
  29871=>"101100000",
  29872=>"001011111",
  29873=>"011101010",
  29874=>"100001011",
  29875=>"000001111",
  29876=>"110110000",
  29877=>"001000010",
  29878=>"010010011",
  29879=>"011100000",
  29880=>"000001011",
  29881=>"001101000",
  29882=>"010001011",
  29883=>"110101010",
  29884=>"001010110",
  29885=>"011001111",
  29886=>"010111001",
  29887=>"010011000",
  29888=>"111001101",
  29889=>"110000101",
  29890=>"000111010",
  29891=>"001111011",
  29892=>"010110010",
  29893=>"111011100",
  29894=>"010110100",
  29895=>"110110110",
  29896=>"000010101",
  29897=>"010010011",
  29898=>"100000111",
  29899=>"011111100",
  29900=>"010010000",
  29901=>"011000100",
  29902=>"010001001",
  29903=>"101000110",
  29904=>"110101000",
  29905=>"101011000",
  29906=>"000111110",
  29907=>"100100011",
  29908=>"000000001",
  29909=>"110110010",
  29910=>"110111011",
  29911=>"111010100",
  29912=>"101101100",
  29913=>"000100111",
  29914=>"000000111",
  29915=>"000001111",
  29916=>"011110000",
  29917=>"010010011",
  29918=>"001001101",
  29919=>"010011001",
  29920=>"000100010",
  29921=>"001000111",
  29922=>"111110010",
  29923=>"010010001",
  29924=>"001110100",
  29925=>"011101100",
  29926=>"100111011",
  29927=>"100100100",
  29928=>"100100100",
  29929=>"011010011",
  29930=>"001011010",
  29931=>"100111010",
  29932=>"110110001",
  29933=>"010000100",
  29934=>"011111011",
  29935=>"100001111",
  29936=>"001001011",
  29937=>"100010101",
  29938=>"110001111",
  29939=>"011001000",
  29940=>"010001100",
  29941=>"100011000",
  29942=>"011001110",
  29943=>"011010010",
  29944=>"100111100",
  29945=>"111000101",
  29946=>"000110110",
  29947=>"010001011",
  29948=>"011011111",
  29949=>"001100001",
  29950=>"110110010",
  29951=>"000001111",
  29952=>"110010011",
  29953=>"000110011",
  29954=>"011101100",
  29955=>"011010010",
  29956=>"101001100",
  29957=>"101110000",
  29958=>"000010010",
  29959=>"111101010",
  29960=>"010111101",
  29961=>"111001101",
  29962=>"110100001",
  29963=>"000000101",
  29964=>"000000010",
  29965=>"001101110",
  29966=>"010100000",
  29967=>"100011000",
  29968=>"001110000",
  29969=>"100001001",
  29970=>"110110110",
  29971=>"101101011",
  29972=>"101000000",
  29973=>"001000011",
  29974=>"111001010",
  29975=>"000110100",
  29976=>"111011111",
  29977=>"101110110",
  29978=>"100110110",
  29979=>"100000101",
  29980=>"011011111",
  29981=>"001010010",
  29982=>"111100010",
  29983=>"000110110",
  29984=>"110111000",
  29985=>"110100111",
  29986=>"010001101",
  29987=>"010100110",
  29988=>"000100100",
  29989=>"010000110",
  29990=>"010111010",
  29991=>"010111101",
  29992=>"101001101",
  29993=>"110011011",
  29994=>"000111000",
  29995=>"101011000",
  29996=>"110110111",
  29997=>"010001011",
  29998=>"011111011",
  29999=>"001001110",
  30000=>"101100001",
  30001=>"110010001",
  30002=>"000011101",
  30003=>"011010000",
  30004=>"100001110",
  30005=>"100001111",
  30006=>"101011100",
  30007=>"100111000",
  30008=>"111001101",
  30009=>"101001011",
  30010=>"101000101",
  30011=>"110111110",
  30012=>"011000111",
  30013=>"110011010",
  30014=>"001010001",
  30015=>"011011001",
  30016=>"001111000",
  30017=>"100010100",
  30018=>"000010110",
  30019=>"010000000",
  30020=>"100000001",
  30021=>"111000101",
  30022=>"101100010",
  30023=>"011111111",
  30024=>"100100100",
  30025=>"010110001",
  30026=>"101011100",
  30027=>"010010011",
  30028=>"001001000",
  30029=>"110001100",
  30030=>"010000000",
  30031=>"101000011",
  30032=>"001011111",
  30033=>"010110110",
  30034=>"010011001",
  30035=>"011111110",
  30036=>"000011101",
  30037=>"100001001",
  30038=>"111110110",
  30039=>"001110100",
  30040=>"111110111",
  30041=>"100111110",
  30042=>"001010000",
  30043=>"101111010",
  30044=>"000000000",
  30045=>"011010001",
  30046=>"101101111",
  30047=>"010011010",
  30048=>"000001011",
  30049=>"001011011",
  30050=>"101100100",
  30051=>"111001110",
  30052=>"011101111",
  30053=>"111111100",
  30054=>"001011111",
  30055=>"001111001",
  30056=>"001010001",
  30057=>"010110110",
  30058=>"100111001",
  30059=>"110111010",
  30060=>"110000000",
  30061=>"111101011",
  30062=>"110111101",
  30063=>"011000000",
  30064=>"011110011",
  30065=>"000100001",
  30066=>"100001011",
  30067=>"100010101",
  30068=>"110110010",
  30069=>"010011100",
  30070=>"001010001",
  30071=>"010011000",
  30072=>"101011000",
  30073=>"010001001",
  30074=>"011101100",
  30075=>"101111100",
  30076=>"111110000",
  30077=>"101110111",
  30078=>"010101010",
  30079=>"101001010",
  30080=>"011110110",
  30081=>"101011101",
  30082=>"101000110",
  30083=>"010100100",
  30084=>"111010110",
  30085=>"010111110",
  30086=>"111101100",
  30087=>"010011110",
  30088=>"010001000",
  30089=>"000000000",
  30090=>"000000000",
  30091=>"010101101",
  30092=>"100010000",
  30093=>"000111001",
  30094=>"001111111",
  30095=>"000110110",
  30096=>"000111011",
  30097=>"000100110",
  30098=>"111101111",
  30099=>"000001110",
  30100=>"101001101",
  30101=>"000000111",
  30102=>"010111001",
  30103=>"111001001",
  30104=>"101101100",
  30105=>"010100000",
  30106=>"100000111",
  30107=>"011011001",
  30108=>"110111101",
  30109=>"001100000",
  30110=>"001101110",
  30111=>"000001011",
  30112=>"000011010",
  30113=>"001110100",
  30114=>"001100011",
  30115=>"000000111",
  30116=>"110100001",
  30117=>"010101001",
  30118=>"001011101",
  30119=>"110000110",
  30120=>"101110000",
  30121=>"001010111",
  30122=>"101011000",
  30123=>"100110111",
  30124=>"111000100",
  30125=>"111100110",
  30126=>"101111111",
  30127=>"100111010",
  30128=>"110110001",
  30129=>"100110000",
  30130=>"011111101",
  30131=>"011100000",
  30132=>"111101000",
  30133=>"010110001",
  30134=>"000110111",
  30135=>"010000110",
  30136=>"010110111",
  30137=>"111001000",
  30138=>"000010111",
  30139=>"101110111",
  30140=>"111001111",
  30141=>"111011010",
  30142=>"000001101",
  30143=>"111101100",
  30144=>"110010010",
  30145=>"000111111",
  30146=>"111000000",
  30147=>"010000011",
  30148=>"011000110",
  30149=>"010111010",
  30150=>"000100011",
  30151=>"000011010",
  30152=>"110111100",
  30153=>"100111010",
  30154=>"010111010",
  30155=>"110101100",
  30156=>"100001101",
  30157=>"000110100",
  30158=>"001111010",
  30159=>"111110010",
  30160=>"110000011",
  30161=>"000110110",
  30162=>"111101100",
  30163=>"100101011",
  30164=>"111110111",
  30165=>"001110101",
  30166=>"101011111",
  30167=>"011010000",
  30168=>"001100011",
  30169=>"010110011",
  30170=>"100110001",
  30171=>"100000000",
  30172=>"011011110",
  30173=>"010011100",
  30174=>"110111101",
  30175=>"110011000",
  30176=>"111000000",
  30177=>"011001111",
  30178=>"001000010",
  30179=>"110010100",
  30180=>"110111000",
  30181=>"010101000",
  30182=>"101100000",
  30183=>"000111011",
  30184=>"001001111",
  30185=>"011000110",
  30186=>"001011101",
  30187=>"000000110",
  30188=>"000111011",
  30189=>"111101000",
  30190=>"001011010",
  30191=>"001100011",
  30192=>"101111011",
  30193=>"000111011",
  30194=>"000000011",
  30195=>"011010000",
  30196=>"100110111",
  30197=>"011010000",
  30198=>"010000101",
  30199=>"010001110",
  30200=>"010101101",
  30201=>"010011111",
  30202=>"110110101",
  30203=>"101101101",
  30204=>"111111100",
  30205=>"001110110",
  30206=>"111010011",
  30207=>"111111101",
  30208=>"111010111",
  30209=>"001010101",
  30210=>"001000101",
  30211=>"001010011",
  30212=>"000001111",
  30213=>"111100100",
  30214=>"000101110",
  30215=>"111110011",
  30216=>"000100010",
  30217=>"110111111",
  30218=>"000100110",
  30219=>"000101010",
  30220=>"101110011",
  30221=>"100111000",
  30222=>"000100100",
  30223=>"110110111",
  30224=>"011001110",
  30225=>"111000101",
  30226=>"100010010",
  30227=>"000001110",
  30228=>"100000011",
  30229=>"101101101",
  30230=>"000101110",
  30231=>"110010011",
  30232=>"000001111",
  30233=>"100100011",
  30234=>"011010011",
  30235=>"101010100",
  30236=>"100101110",
  30237=>"011101101",
  30238=>"110000011",
  30239=>"000001101",
  30240=>"000100000",
  30241=>"001110000",
  30242=>"000011010",
  30243=>"011100001",
  30244=>"100011010",
  30245=>"110011001",
  30246=>"011010001",
  30247=>"010010111",
  30248=>"010000000",
  30249=>"100110010",
  30250=>"100000000",
  30251=>"101100000",
  30252=>"010001000",
  30253=>"100110001",
  30254=>"000100010",
  30255=>"111000101",
  30256=>"001100111",
  30257=>"110001101",
  30258=>"111001110",
  30259=>"100001001",
  30260=>"010110101",
  30261=>"111111010",
  30262=>"010000111",
  30263=>"111011111",
  30264=>"001101111",
  30265=>"000111110",
  30266=>"011100101",
  30267=>"000101111",
  30268=>"000101000",
  30269=>"110011101",
  30270=>"100100011",
  30271=>"010101010",
  30272=>"000000100",
  30273=>"011010111",
  30274=>"110000100",
  30275=>"010010101",
  30276=>"111011000",
  30277=>"110110010",
  30278=>"010111001",
  30279=>"001110100",
  30280=>"000111100",
  30281=>"010001101",
  30282=>"100010000",
  30283=>"000010111",
  30284=>"000000011",
  30285=>"101000011",
  30286=>"110101010",
  30287=>"001000111",
  30288=>"110010010",
  30289=>"000000100",
  30290=>"100011010",
  30291=>"001101001",
  30292=>"010100001",
  30293=>"001100001",
  30294=>"100110000",
  30295=>"011101101",
  30296=>"000111111",
  30297=>"110111011",
  30298=>"000010011",
  30299=>"111110011",
  30300=>"011001111",
  30301=>"010001010",
  30302=>"111110011",
  30303=>"000001111",
  30304=>"011100110",
  30305=>"001111100",
  30306=>"011111101",
  30307=>"000100010",
  30308=>"010100110",
  30309=>"111010000",
  30310=>"101111101",
  30311=>"011100100",
  30312=>"000011001",
  30313=>"000101011",
  30314=>"100111101",
  30315=>"010000100",
  30316=>"110011011",
  30317=>"000100110",
  30318=>"110010100",
  30319=>"111100010",
  30320=>"111000010",
  30321=>"110101010",
  30322=>"000100000",
  30323=>"001001001",
  30324=>"011010001",
  30325=>"010011101",
  30326=>"111110100",
  30327=>"011010111",
  30328=>"000100010",
  30329=>"100111111",
  30330=>"101111010",
  30331=>"111111010",
  30332=>"011010100",
  30333=>"101000101",
  30334=>"111000101",
  30335=>"100110011",
  30336=>"011000000",
  30337=>"101100010",
  30338=>"111001000",
  30339=>"000101010",
  30340=>"100011100",
  30341=>"111000110",
  30342=>"110100000",
  30343=>"010010110",
  30344=>"000010011",
  30345=>"110100110",
  30346=>"101000101",
  30347=>"010000110",
  30348=>"100111111",
  30349=>"001111011",
  30350=>"000100111",
  30351=>"010011010",
  30352=>"010111000",
  30353=>"001010000",
  30354=>"101010111",
  30355=>"101111110",
  30356=>"110111100",
  30357=>"001000001",
  30358=>"001010011",
  30359=>"100100010",
  30360=>"010111101",
  30361=>"000010011",
  30362=>"011001001",
  30363=>"111100110",
  30364=>"010110001",
  30365=>"000000010",
  30366=>"001010100",
  30367=>"010011111",
  30368=>"111001100",
  30369=>"110010101",
  30370=>"111000010",
  30371=>"000010000",
  30372=>"011010110",
  30373=>"100000010",
  30374=>"011101101",
  30375=>"110011100",
  30376=>"110001111",
  30377=>"110100010",
  30378=>"011111010",
  30379=>"010110111",
  30380=>"000100000",
  30381=>"010110111",
  30382=>"011110001",
  30383=>"011101000",
  30384=>"000011101",
  30385=>"000101100",
  30386=>"101101000",
  30387=>"010100110",
  30388=>"111011010",
  30389=>"000001000",
  30390=>"111000000",
  30391=>"100000101",
  30392=>"111000111",
  30393=>"001101001",
  30394=>"110011111",
  30395=>"100100100",
  30396=>"111000011",
  30397=>"010001010",
  30398=>"101000110",
  30399=>"100110100",
  30400=>"000111110",
  30401=>"100011111",
  30402=>"011001101",
  30403=>"001100111",
  30404=>"111011111",
  30405=>"000110000",
  30406=>"010100110",
  30407=>"100100001",
  30408=>"011010010",
  30409=>"001101111",
  30410=>"011101100",
  30411=>"010010110",
  30412=>"001011011",
  30413=>"111010000",
  30414=>"101100001",
  30415=>"011101010",
  30416=>"010000100",
  30417=>"001001101",
  30418=>"100010000",
  30419=>"110001000",
  30420=>"001001011",
  30421=>"101100110",
  30422=>"101010101",
  30423=>"001101010",
  30424=>"001011100",
  30425=>"001001111",
  30426=>"001110011",
  30427=>"001111011",
  30428=>"000111101",
  30429=>"011100100",
  30430=>"010011001",
  30431=>"010101010",
  30432=>"100100110",
  30433=>"101010001",
  30434=>"100011010",
  30435=>"010111100",
  30436=>"001100000",
  30437=>"100101100",
  30438=>"110010001",
  30439=>"100100000",
  30440=>"111101001",
  30441=>"000101000",
  30442=>"101010110",
  30443=>"001100000",
  30444=>"100101111",
  30445=>"100000010",
  30446=>"000100101",
  30447=>"001000111",
  30448=>"110000110",
  30449=>"011100111",
  30450=>"000111011",
  30451=>"110001110",
  30452=>"101011111",
  30453=>"011110011",
  30454=>"111111011",
  30455=>"010000011",
  30456=>"101111001",
  30457=>"100000000",
  30458=>"100001010",
  30459=>"101000011",
  30460=>"100011000",
  30461=>"010001101",
  30462=>"000111100",
  30463=>"110001111",
  30464=>"001000100",
  30465=>"001011110",
  30466=>"101100011",
  30467=>"101100111",
  30468=>"000100011",
  30469=>"101011011",
  30470=>"010100001",
  30471=>"111001111",
  30472=>"110111011",
  30473=>"010100011",
  30474=>"101011001",
  30475=>"110111110",
  30476=>"111011111",
  30477=>"111111111",
  30478=>"110010000",
  30479=>"101110100",
  30480=>"010001110",
  30481=>"110110101",
  30482=>"000000100",
  30483=>"010000100",
  30484=>"000100011",
  30485=>"010011100",
  30486=>"010111000",
  30487=>"001001000",
  30488=>"001001011",
  30489=>"101111001",
  30490=>"100000001",
  30491=>"011101110",
  30492=>"010101100",
  30493=>"001100101",
  30494=>"011000110",
  30495=>"101000001",
  30496=>"101001100",
  30497=>"100000011",
  30498=>"000100000",
  30499=>"101001100",
  30500=>"101000110",
  30501=>"000001101",
  30502=>"010100111",
  30503=>"000100011",
  30504=>"100100000",
  30505=>"001010001",
  30506=>"110110101",
  30507=>"011001000",
  30508=>"111111010",
  30509=>"010000111",
  30510=>"001111010",
  30511=>"010110011",
  30512=>"010010100",
  30513=>"101100101",
  30514=>"111111110",
  30515=>"111111000",
  30516=>"010010001",
  30517=>"001010000",
  30518=>"000010110",
  30519=>"000101011",
  30520=>"110111000",
  30521=>"010110000",
  30522=>"111000111",
  30523=>"101011001",
  30524=>"010001011",
  30525=>"100111110",
  30526=>"101010100",
  30527=>"110110101",
  30528=>"100100111",
  30529=>"101101111",
  30530=>"100100010",
  30531=>"110011111",
  30532=>"001000110",
  30533=>"101100000",
  30534=>"000010100",
  30535=>"001001110",
  30536=>"110011100",
  30537=>"001111111",
  30538=>"100110110",
  30539=>"110111110",
  30540=>"000001000",
  30541=>"011010010",
  30542=>"001011000",
  30543=>"011100111",
  30544=>"001110100",
  30545=>"001000001",
  30546=>"100110000",
  30547=>"000110110",
  30548=>"110111101",
  30549=>"001100100",
  30550=>"011010011",
  30551=>"111100001",
  30552=>"111110110",
  30553=>"011111000",
  30554=>"000001101",
  30555=>"110101101",
  30556=>"011011110",
  30557=>"010111100",
  30558=>"010011010",
  30559=>"000011010",
  30560=>"011100110",
  30561=>"010110000",
  30562=>"011110001",
  30563=>"101011111",
  30564=>"101110000",
  30565=>"111110111",
  30566=>"111010011",
  30567=>"111101000",
  30568=>"101000010",
  30569=>"101010000",
  30570=>"001000010",
  30571=>"010011011",
  30572=>"001110101",
  30573=>"101011011",
  30574=>"100000111",
  30575=>"011001000",
  30576=>"011001001",
  30577=>"001101001",
  30578=>"011101010",
  30579=>"110011110",
  30580=>"100111101",
  30581=>"100111000",
  30582=>"111111000",
  30583=>"010111101",
  30584=>"001100111",
  30585=>"110011001",
  30586=>"111001000",
  30587=>"011101000",
  30588=>"100000001",
  30589=>"000111010",
  30590=>"000110001",
  30591=>"111001000",
  30592=>"010111011",
  30593=>"101001111",
  30594=>"101010001",
  30595=>"000011111",
  30596=>"010010111",
  30597=>"100000110",
  30598=>"010101001",
  30599=>"100110111",
  30600=>"000111111",
  30601=>"100111111",
  30602=>"101111101",
  30603=>"101000001",
  30604=>"111010001",
  30605=>"100010001",
  30606=>"001001010",
  30607=>"010011101",
  30608=>"001001101",
  30609=>"100111011",
  30610=>"001111110",
  30611=>"111101010",
  30612=>"000001011",
  30613=>"000011100",
  30614=>"001100011",
  30615=>"000011110",
  30616=>"000101110",
  30617=>"000011011",
  30618=>"010001000",
  30619=>"001011100",
  30620=>"001001111",
  30621=>"010000101",
  30622=>"110110001",
  30623=>"011011001",
  30624=>"110001110",
  30625=>"111000110",
  30626=>"000000111",
  30627=>"000101101",
  30628=>"000100010",
  30629=>"101101101",
  30630=>"001001010",
  30631=>"110101000",
  30632=>"000110001",
  30633=>"100101101",
  30634=>"100100100",
  30635=>"101011000",
  30636=>"111000100",
  30637=>"001000100",
  30638=>"101011101",
  30639=>"110101110",
  30640=>"111001000",
  30641=>"010110100",
  30642=>"010001000",
  30643=>"011010100",
  30644=>"000000100",
  30645=>"010000101",
  30646=>"111110100",
  30647=>"110000011",
  30648=>"100000010",
  30649=>"111000100",
  30650=>"010010101",
  30651=>"100110011",
  30652=>"011001000",
  30653=>"000100000",
  30654=>"010010010",
  30655=>"010011001",
  30656=>"000010011",
  30657=>"011101101",
  30658=>"100111011",
  30659=>"000110010",
  30660=>"011101111",
  30661=>"011010111",
  30662=>"101000010",
  30663=>"001000110",
  30664=>"101100010",
  30665=>"100110010",
  30666=>"000000111",
  30667=>"001101010",
  30668=>"101010101",
  30669=>"110001111",
  30670=>"010110101",
  30671=>"010011001",
  30672=>"010111000",
  30673=>"001100000",
  30674=>"011001110",
  30675=>"011000010",
  30676=>"000010011",
  30677=>"001101111",
  30678=>"000000000",
  30679=>"010011111",
  30680=>"110000000",
  30681=>"111101010",
  30682=>"111110100",
  30683=>"110011101",
  30684=>"001101111",
  30685=>"100110101",
  30686=>"100110111",
  30687=>"101110100",
  30688=>"010001000",
  30689=>"000001101",
  30690=>"110000001",
  30691=>"111101001",
  30692=>"001111000",
  30693=>"110011100",
  30694=>"000011010",
  30695=>"100010000",
  30696=>"110010011",
  30697=>"011010110",
  30698=>"101001000",
  30699=>"011111111",
  30700=>"001000110",
  30701=>"010000011",
  30702=>"111110101",
  30703=>"101111110",
  30704=>"110010010",
  30705=>"110011001",
  30706=>"010111011",
  30707=>"110010101",
  30708=>"111000010",
  30709=>"010000111",
  30710=>"100110010",
  30711=>"010011110",
  30712=>"101111011",
  30713=>"000011010",
  30714=>"000011010",
  30715=>"010000010",
  30716=>"011100001",
  30717=>"101111100",
  30718=>"110010110",
  30719=>"011011011",
  30720=>"010011000",
  30721=>"100001001",
  30722=>"010001001",
  30723=>"001011000",
  30724=>"101010001",
  30725=>"110011001",
  30726=>"010011101",
  30727=>"011100110",
  30728=>"100001000",
  30729=>"001010110",
  30730=>"110111010",
  30731=>"011001011",
  30732=>"100111000",
  30733=>"100011111",
  30734=>"111111000",
  30735=>"100101000",
  30736=>"011111110",
  30737=>"110001111",
  30738=>"111010010",
  30739=>"100101111",
  30740=>"000101001",
  30741=>"000000000",
  30742=>"010110110",
  30743=>"001100000",
  30744=>"111101100",
  30745=>"000011011",
  30746=>"110111010",
  30747=>"110111001",
  30748=>"000011110",
  30749=>"001000010",
  30750=>"100010001",
  30751=>"110100111",
  30752=>"001010010",
  30753=>"100100100",
  30754=>"001100011",
  30755=>"111100110",
  30756=>"001001011",
  30757=>"011010110",
  30758=>"110000000",
  30759=>"110111111",
  30760=>"001000001",
  30761=>"010110100",
  30762=>"101000110",
  30763=>"001100000",
  30764=>"011000010",
  30765=>"000101111",
  30766=>"001111010",
  30767=>"001010011",
  30768=>"000110011",
  30769=>"011010100",
  30770=>"101111101",
  30771=>"000110110",
  30772=>"110001000",
  30773=>"000001010",
  30774=>"010110100",
  30775=>"100111011",
  30776=>"100110000",
  30777=>"101100101",
  30778=>"000011110",
  30779=>"011010100",
  30780=>"010101000",
  30781=>"011011111",
  30782=>"010100001",
  30783=>"101100111",
  30784=>"101001100",
  30785=>"101010110",
  30786=>"011101000",
  30787=>"100010101",
  30788=>"000110110",
  30789=>"011011011",
  30790=>"010001000",
  30791=>"101100111",
  30792=>"011110001",
  30793=>"111111010",
  30794=>"101001011",
  30795=>"011001011",
  30796=>"111110001",
  30797=>"101110001",
  30798=>"111110000",
  30799=>"001110101",
  30800=>"100110100",
  30801=>"000000001",
  30802=>"011111011",
  30803=>"101101101",
  30804=>"001000101",
  30805=>"101100010",
  30806=>"010000101",
  30807=>"011010001",
  30808=>"011011010",
  30809=>"101000010",
  30810=>"100110001",
  30811=>"101001011",
  30812=>"010000111",
  30813=>"000011000",
  30814=>"111111010",
  30815=>"001101000",
  30816=>"000010110",
  30817=>"011100000",
  30818=>"010000000",
  30819=>"001111000",
  30820=>"110101011",
  30821=>"000000010",
  30822=>"001100010",
  30823=>"000101011",
  30824=>"011010111",
  30825=>"101111110",
  30826=>"110100100",
  30827=>"101110011",
  30828=>"101001010",
  30829=>"101011001",
  30830=>"100010101",
  30831=>"100100010",
  30832=>"010111111",
  30833=>"000000010",
  30834=>"001101001",
  30835=>"111111100",
  30836=>"010100100",
  30837=>"111100001",
  30838=>"101010011",
  30839=>"101101101",
  30840=>"000010001",
  30841=>"001100110",
  30842=>"110110111",
  30843=>"001000010",
  30844=>"111000101",
  30845=>"010000010",
  30846=>"101001100",
  30847=>"111001001",
  30848=>"101001100",
  30849=>"011110010",
  30850=>"111110101",
  30851=>"000000000",
  30852=>"111110111",
  30853=>"110010101",
  30854=>"001110010",
  30855=>"011110110",
  30856=>"100111000",
  30857=>"011011110",
  30858=>"010100100",
  30859=>"101101001",
  30860=>"001111111",
  30861=>"100101010",
  30862=>"000100010",
  30863=>"001011000",
  30864=>"001010010",
  30865=>"001010000",
  30866=>"010101101",
  30867=>"101110110",
  30868=>"100000000",
  30869=>"011100100",
  30870=>"001101100",
  30871=>"010110111",
  30872=>"010000101",
  30873=>"001111001",
  30874=>"101001011",
  30875=>"111111111",
  30876=>"011011100",
  30877=>"001001000",
  30878=>"111110001",
  30879=>"001000010",
  30880=>"100010100",
  30881=>"100000110",
  30882=>"101011110",
  30883=>"011011101",
  30884=>"101000100",
  30885=>"111100111",
  30886=>"001011111",
  30887=>"111010000",
  30888=>"100110101",
  30889=>"110111000",
  30890=>"100011001",
  30891=>"010101001",
  30892=>"011110000",
  30893=>"100101011",
  30894=>"000111000",
  30895=>"000100000",
  30896=>"110101000",
  30897=>"000111010",
  30898=>"010010000",
  30899=>"100101011",
  30900=>"100011110",
  30901=>"011011010",
  30902=>"000001011",
  30903=>"111110101",
  30904=>"110110111",
  30905=>"001010110",
  30906=>"110111111",
  30907=>"101110010",
  30908=>"000011000",
  30909=>"101111110",
  30910=>"111010111",
  30911=>"011100010",
  30912=>"110100101",
  30913=>"010100000",
  30914=>"001010001",
  30915=>"111110111",
  30916=>"101110001",
  30917=>"110100100",
  30918=>"010001101",
  30919=>"000101011",
  30920=>"101011011",
  30921=>"110101000",
  30922=>"000101010",
  30923=>"011101011",
  30924=>"111110010",
  30925=>"111111111",
  30926=>"001100011",
  30927=>"100110111",
  30928=>"010010111",
  30929=>"101001010",
  30930=>"011010000",
  30931=>"010110000",
  30932=>"001010111",
  30933=>"000110000",
  30934=>"100110011",
  30935=>"010010010",
  30936=>"011000010",
  30937=>"000010110",
  30938=>"100000011",
  30939=>"101111110",
  30940=>"000001010",
  30941=>"100110001",
  30942=>"111001000",
  30943=>"011010011",
  30944=>"101001100",
  30945=>"011100010",
  30946=>"001010001",
  30947=>"110011101",
  30948=>"110011111",
  30949=>"001000001",
  30950=>"001101010",
  30951=>"111101111",
  30952=>"000001010",
  30953=>"011101100",
  30954=>"111101000",
  30955=>"001000111",
  30956=>"110000010",
  30957=>"101100100",
  30958=>"111111100",
  30959=>"100000100",
  30960=>"010111001",
  30961=>"001110110",
  30962=>"010011001",
  30963=>"110001010",
  30964=>"100101000",
  30965=>"010111100",
  30966=>"110111110",
  30967=>"101101010",
  30968=>"111100011",
  30969=>"110101111",
  30970=>"100111001",
  30971=>"010101000",
  30972=>"001010000",
  30973=>"000101111",
  30974=>"000011111",
  30975=>"010000010",
  30976=>"011100000",
  30977=>"010100100",
  30978=>"111001010",
  30979=>"111001001",
  30980=>"101111001",
  30981=>"100001100",
  30982=>"111111011",
  30983=>"001110111",
  30984=>"000010010",
  30985=>"011110001",
  30986=>"111110110",
  30987=>"110000100",
  30988=>"000111001",
  30989=>"100000011",
  30990=>"001100111",
  30991=>"110010001",
  30992=>"011000110",
  30993=>"110100111",
  30994=>"000101101",
  30995=>"100101101",
  30996=>"011110100",
  30997=>"001100111",
  30998=>"001001000",
  30999=>"010100011",
  31000=>"111010001",
  31001=>"000111000",
  31002=>"000101101",
  31003=>"011100001",
  31004=>"010000011",
  31005=>"101110001",
  31006=>"001111100",
  31007=>"100011101",
  31008=>"100101110",
  31009=>"101001000",
  31010=>"010101101",
  31011=>"111010110",
  31012=>"100000010",
  31013=>"100010110",
  31014=>"111101000",
  31015=>"100101100",
  31016=>"000001111",
  31017=>"100111011",
  31018=>"110010100",
  31019=>"100000011",
  31020=>"000111001",
  31021=>"000110001",
  31022=>"100011011",
  31023=>"100111000",
  31024=>"010011111",
  31025=>"001111011",
  31026=>"100010111",
  31027=>"000100010",
  31028=>"101101100",
  31029=>"000000010",
  31030=>"100110001",
  31031=>"011111100",
  31032=>"011100000",
  31033=>"110010000",
  31034=>"110000110",
  31035=>"100000100",
  31036=>"111100111",
  31037=>"000111101",
  31038=>"000011111",
  31039=>"000000011",
  31040=>"010010100",
  31041=>"000110010",
  31042=>"111111101",
  31043=>"101001111",
  31044=>"101010001",
  31045=>"101110100",
  31046=>"010110101",
  31047=>"010110110",
  31048=>"100111000",
  31049=>"100100100",
  31050=>"010000110",
  31051=>"111001100",
  31052=>"110100010",
  31053=>"110011110",
  31054=>"011001010",
  31055=>"000110110",
  31056=>"100111001",
  31057=>"011010001",
  31058=>"100001110",
  31059=>"100100000",
  31060=>"100110010",
  31061=>"110010111",
  31062=>"100001000",
  31063=>"000101011",
  31064=>"000010000",
  31065=>"101000100",
  31066=>"110111111",
  31067=>"110011100",
  31068=>"111011110",
  31069=>"011111100",
  31070=>"111001110",
  31071=>"011110101",
  31072=>"011101111",
  31073=>"010100101",
  31074=>"000100001",
  31075=>"001011010",
  31076=>"111001101",
  31077=>"100000010",
  31078=>"000010111",
  31079=>"111100111",
  31080=>"101101100",
  31081=>"111110001",
  31082=>"000010001",
  31083=>"111111101",
  31084=>"110110101",
  31085=>"101000100",
  31086=>"011011110",
  31087=>"011111000",
  31088=>"000011101",
  31089=>"100100111",
  31090=>"000000001",
  31091=>"110110001",
  31092=>"110000011",
  31093=>"100001111",
  31094=>"011101101",
  31095=>"001111100",
  31096=>"000101101",
  31097=>"000000000",
  31098=>"111111111",
  31099=>"010011101",
  31100=>"100000100",
  31101=>"110000110",
  31102=>"100101100",
  31103=>"111011000",
  31104=>"000100001",
  31105=>"101101000",
  31106=>"111000110",
  31107=>"110101001",
  31108=>"110110001",
  31109=>"001001000",
  31110=>"001101010",
  31111=>"110110101",
  31112=>"011110100",
  31113=>"011100110",
  31114=>"000100011",
  31115=>"101111100",
  31116=>"100011011",
  31117=>"001001011",
  31118=>"101001011",
  31119=>"111000111",
  31120=>"010010001",
  31121=>"001111100",
  31122=>"000101100",
  31123=>"111000110",
  31124=>"011111111",
  31125=>"001100000",
  31126=>"101010101",
  31127=>"000100101",
  31128=>"111001100",
  31129=>"100000100",
  31130=>"000110000",
  31131=>"000010100",
  31132=>"111110101",
  31133=>"000101100",
  31134=>"001000011",
  31135=>"011110101",
  31136=>"101001110",
  31137=>"000111110",
  31138=>"110000001",
  31139=>"011000010",
  31140=>"010001011",
  31141=>"010000100",
  31142=>"011001101",
  31143=>"000111010",
  31144=>"000101010",
  31145=>"111001000",
  31146=>"000001000",
  31147=>"100101101",
  31148=>"111111011",
  31149=>"000110011",
  31150=>"000000111",
  31151=>"000011011",
  31152=>"000000010",
  31153=>"000000001",
  31154=>"100111100",
  31155=>"000010010",
  31156=>"101001001",
  31157=>"110011101",
  31158=>"001110110",
  31159=>"000100001",
  31160=>"101011100",
  31161=>"011101001",
  31162=>"101001001",
  31163=>"110010000",
  31164=>"111000011",
  31165=>"011101111",
  31166=>"011001000",
  31167=>"100001111",
  31168=>"111010011",
  31169=>"110111010",
  31170=>"100001001",
  31171=>"010010000",
  31172=>"101110110",
  31173=>"101110000",
  31174=>"111100111",
  31175=>"111101011",
  31176=>"011011000",
  31177=>"000110000",
  31178=>"010110011",
  31179=>"001100001",
  31180=>"001110011",
  31181=>"010100011",
  31182=>"100000100",
  31183=>"001110100",
  31184=>"111101010",
  31185=>"011100001",
  31186=>"011101111",
  31187=>"110011010",
  31188=>"111111111",
  31189=>"011101001",
  31190=>"111011000",
  31191=>"101101110",
  31192=>"010100110",
  31193=>"000010011",
  31194=>"101111011",
  31195=>"011111111",
  31196=>"100010011",
  31197=>"011101001",
  31198=>"001110000",
  31199=>"101001000",
  31200=>"010000101",
  31201=>"101100101",
  31202=>"010001111",
  31203=>"110011011",
  31204=>"111110001",
  31205=>"000000100",
  31206=>"000010010",
  31207=>"000111101",
  31208=>"110100010",
  31209=>"101001001",
  31210=>"110111111",
  31211=>"100001110",
  31212=>"100111011",
  31213=>"001111000",
  31214=>"100111101",
  31215=>"011010001",
  31216=>"011011001",
  31217=>"110110110",
  31218=>"110010010",
  31219=>"010001100",
  31220=>"101100101",
  31221=>"001010010",
  31222=>"110101001",
  31223=>"101100000",
  31224=>"100111110",
  31225=>"001001010",
  31226=>"010111101",
  31227=>"010111010",
  31228=>"001000000",
  31229=>"010010011",
  31230=>"110010110",
  31231=>"001000000",
  31232=>"010110111",
  31233=>"011011011",
  31234=>"110010111",
  31235=>"101000100",
  31236=>"100101000",
  31237=>"010011010",
  31238=>"010100111",
  31239=>"010001100",
  31240=>"011011100",
  31241=>"010111110",
  31242=>"001100011",
  31243=>"001011100",
  31244=>"111101010",
  31245=>"010010010",
  31246=>"101000001",
  31247=>"101011110",
  31248=>"011111100",
  31249=>"000110010",
  31250=>"110000000",
  31251=>"101101001",
  31252=>"000001000",
  31253=>"111111110",
  31254=>"011110000",
  31255=>"010110001",
  31256=>"011100101",
  31257=>"011100010",
  31258=>"101001001",
  31259=>"101111010",
  31260=>"101111001",
  31261=>"111011001",
  31262=>"101001011",
  31263=>"010010000",
  31264=>"101100001",
  31265=>"000111000",
  31266=>"111111101",
  31267=>"100110100",
  31268=>"100101101",
  31269=>"001101100",
  31270=>"100000000",
  31271=>"110110000",
  31272=>"100100111",
  31273=>"011000111",
  31274=>"111000000",
  31275=>"001101010",
  31276=>"110011000",
  31277=>"111001110",
  31278=>"100100001",
  31279=>"000010101",
  31280=>"001010000",
  31281=>"101101100",
  31282=>"010000100",
  31283=>"111101111",
  31284=>"111001100",
  31285=>"101011011",
  31286=>"001001110",
  31287=>"101111101",
  31288=>"000100111",
  31289=>"001100100",
  31290=>"100111000",
  31291=>"110101100",
  31292=>"011011111",
  31293=>"100010000",
  31294=>"011000010",
  31295=>"011010110",
  31296=>"001000010",
  31297=>"111100101",
  31298=>"011110011",
  31299=>"111000011",
  31300=>"010100010",
  31301=>"101001110",
  31302=>"100111010",
  31303=>"010000111",
  31304=>"000000001",
  31305=>"100001001",
  31306=>"000100010",
  31307=>"000001011",
  31308=>"110111110",
  31309=>"000101011",
  31310=>"010001100",
  31311=>"011010000",
  31312=>"010000000",
  31313=>"011000011",
  31314=>"101101110",
  31315=>"011101101",
  31316=>"110010110",
  31317=>"001100010",
  31318=>"010110000",
  31319=>"100111000",
  31320=>"010111101",
  31321=>"101011000",
  31322=>"011010001",
  31323=>"111101011",
  31324=>"101101000",
  31325=>"111010000",
  31326=>"011100100",
  31327=>"110011101",
  31328=>"100011101",
  31329=>"100100000",
  31330=>"101000011",
  31331=>"111110010",
  31332=>"010100011",
  31333=>"010110010",
  31334=>"111010010",
  31335=>"011010101",
  31336=>"011010100",
  31337=>"000100100",
  31338=>"001010000",
  31339=>"100101000",
  31340=>"111000110",
  31341=>"001010101",
  31342=>"110100100",
  31343=>"111010110",
  31344=>"000011111",
  31345=>"011000001",
  31346=>"101011110",
  31347=>"110111011",
  31348=>"111100000",
  31349=>"000100000",
  31350=>"011001000",
  31351=>"100100000",
  31352=>"000011101",
  31353=>"011111001",
  31354=>"100000111",
  31355=>"101100110",
  31356=>"010000110",
  31357=>"100000111",
  31358=>"111001110",
  31359=>"010000100",
  31360=>"100111100",
  31361=>"111000101",
  31362=>"001101111",
  31363=>"000000001",
  31364=>"101010010",
  31365=>"111001110",
  31366=>"101100100",
  31367=>"110011010",
  31368=>"111111101",
  31369=>"000111000",
  31370=>"101000111",
  31371=>"010000000",
  31372=>"110001010",
  31373=>"001110110",
  31374=>"001110101",
  31375=>"001010100",
  31376=>"111110111",
  31377=>"001001100",
  31378=>"000001111",
  31379=>"101011010",
  31380=>"010011000",
  31381=>"100010111",
  31382=>"101001001",
  31383=>"110010000",
  31384=>"110101110",
  31385=>"001111000",
  31386=>"111110011",
  31387=>"000111111",
  31388=>"000011000",
  31389=>"101100101",
  31390=>"100111100",
  31391=>"000010101",
  31392=>"000100001",
  31393=>"111000111",
  31394=>"110010100",
  31395=>"101111000",
  31396=>"111100101",
  31397=>"000101011",
  31398=>"100010101",
  31399=>"111000000",
  31400=>"101000100",
  31401=>"111001011",
  31402=>"000000001",
  31403=>"110101111",
  31404=>"100100011",
  31405=>"110100010",
  31406=>"011000100",
  31407=>"010010101",
  31408=>"010011010",
  31409=>"110000111",
  31410=>"101001000",
  31411=>"001101011",
  31412=>"110010110",
  31413=>"001101101",
  31414=>"110110011",
  31415=>"010010101",
  31416=>"011000010",
  31417=>"111001100",
  31418=>"110110001",
  31419=>"111001001",
  31420=>"011100111",
  31421=>"000001011",
  31422=>"100011000",
  31423=>"000110100",
  31424=>"001000010",
  31425=>"100010000",
  31426=>"010011000",
  31427=>"110011001",
  31428=>"011100101",
  31429=>"010000111",
  31430=>"101010000",
  31431=>"000010100",
  31432=>"110100000",
  31433=>"000010100",
  31434=>"010111110",
  31435=>"000001100",
  31436=>"001100101",
  31437=>"100001110",
  31438=>"011010001",
  31439=>"011001110",
  31440=>"111111110",
  31441=>"100100100",
  31442=>"110100010",
  31443=>"011011000",
  31444=>"101010111",
  31445=>"101101111",
  31446=>"111000011",
  31447=>"101101101",
  31448=>"010101111",
  31449=>"010110110",
  31450=>"111100101",
  31451=>"011011001",
  31452=>"111011000",
  31453=>"110101000",
  31454=>"100010010",
  31455=>"111100101",
  31456=>"011101100",
  31457=>"101011101",
  31458=>"000010110",
  31459=>"101011010",
  31460=>"100011111",
  31461=>"001001111",
  31462=>"100001101",
  31463=>"110110110",
  31464=>"000100001",
  31465=>"111110010",
  31466=>"011100001",
  31467=>"110111101",
  31468=>"010010001",
  31469=>"000100101",
  31470=>"010110010",
  31471=>"001111000",
  31472=>"010101010",
  31473=>"010111011",
  31474=>"010100000",
  31475=>"100101000",
  31476=>"011001110",
  31477=>"101111101",
  31478=>"111111110",
  31479=>"011010000",
  31480=>"110011100",
  31481=>"011010111",
  31482=>"100110001",
  31483=>"100000111",
  31484=>"101011111",
  31485=>"000011010",
  31486=>"100111100",
  31487=>"101001010",
  31488=>"111010101",
  31489=>"101001011",
  31490=>"011101010",
  31491=>"111011110",
  31492=>"100101000",
  31493=>"011000010",
  31494=>"111110111",
  31495=>"011011100",
  31496=>"110101100",
  31497=>"111101101",
  31498=>"010110001",
  31499=>"001011111",
  31500=>"110111101",
  31501=>"000101001",
  31502=>"111001001",
  31503=>"100110101",
  31504=>"010100010",
  31505=>"000111110",
  31506=>"110010100",
  31507=>"100110000",
  31508=>"110010010",
  31509=>"000000101",
  31510=>"000001110",
  31511=>"010000010",
  31512=>"001110110",
  31513=>"101111001",
  31514=>"111101100",
  31515=>"111100111",
  31516=>"110100100",
  31517=>"001011111",
  31518=>"111101111",
  31519=>"100011010",
  31520=>"101011111",
  31521=>"111000100",
  31522=>"100000110",
  31523=>"011110011",
  31524=>"001100101",
  31525=>"100010010",
  31526=>"000100101",
  31527=>"001100001",
  31528=>"111110111",
  31529=>"011001001",
  31530=>"011010011",
  31531=>"101100110",
  31532=>"011001101",
  31533=>"000011101",
  31534=>"101011111",
  31535=>"011010011",
  31536=>"110101101",
  31537=>"100000000",
  31538=>"001011110",
  31539=>"100011101",
  31540=>"000011001",
  31541=>"101100101",
  31542=>"000110000",
  31543=>"010101001",
  31544=>"111000001",
  31545=>"011100000",
  31546=>"000110010",
  31547=>"011100011",
  31548=>"010010100",
  31549=>"100111011",
  31550=>"000100000",
  31551=>"110011111",
  31552=>"011110000",
  31553=>"010100111",
  31554=>"100100110",
  31555=>"011111110",
  31556=>"011010000",
  31557=>"110110101",
  31558=>"000011110",
  31559=>"011010000",
  31560=>"011111100",
  31561=>"000101101",
  31562=>"100101010",
  31563=>"111000001",
  31564=>"101101100",
  31565=>"000010011",
  31566=>"010110010",
  31567=>"111101100",
  31568=>"011100101",
  31569=>"011011110",
  31570=>"001111100",
  31571=>"100110100",
  31572=>"101110010",
  31573=>"101111111",
  31574=>"101011010",
  31575=>"110100011",
  31576=>"101110010",
  31577=>"111010011",
  31578=>"101110110",
  31579=>"000110000",
  31580=>"000110001",
  31581=>"000011010",
  31582=>"001001001",
  31583=>"110000011",
  31584=>"001101011",
  31585=>"010100011",
  31586=>"001101001",
  31587=>"000100101",
  31588=>"111011001",
  31589=>"110001011",
  31590=>"110001000",
  31591=>"111000110",
  31592=>"011011010",
  31593=>"101100111",
  31594=>"011000001",
  31595=>"111010011",
  31596=>"000101011",
  31597=>"101000100",
  31598=>"111010100",
  31599=>"101110010",
  31600=>"001110000",
  31601=>"111111011",
  31602=>"111100111",
  31603=>"101001001",
  31604=>"001110101",
  31605=>"011011101",
  31606=>"111111010",
  31607=>"100011000",
  31608=>"100010111",
  31609=>"001000101",
  31610=>"101000111",
  31611=>"001111110",
  31612=>"100011110",
  31613=>"010011111",
  31614=>"101101001",
  31615=>"110111111",
  31616=>"011100000",
  31617=>"100111111",
  31618=>"011000110",
  31619=>"001001001",
  31620=>"101101101",
  31621=>"111011110",
  31622=>"000100010",
  31623=>"110001010",
  31624=>"010100001",
  31625=>"110111000",
  31626=>"111111111",
  31627=>"100100111",
  31628=>"001100000",
  31629=>"101110110",
  31630=>"111100110",
  31631=>"011111100",
  31632=>"111001101",
  31633=>"000001011",
  31634=>"011011001",
  31635=>"000111000",
  31636=>"011101111",
  31637=>"110101111",
  31638=>"001101001",
  31639=>"111101010",
  31640=>"001010010",
  31641=>"000100101",
  31642=>"100100100",
  31643=>"111111000",
  31644=>"110010111",
  31645=>"011000110",
  31646=>"100111101",
  31647=>"000101100",
  31648=>"000111010",
  31649=>"000001100",
  31650=>"111110100",
  31651=>"011101011",
  31652=>"000101111",
  31653=>"011001100",
  31654=>"110000100",
  31655=>"101011000",
  31656=>"100100111",
  31657=>"001101110",
  31658=>"100011001",
  31659=>"000000110",
  31660=>"101010001",
  31661=>"110110010",
  31662=>"111111101",
  31663=>"111010101",
  31664=>"011101100",
  31665=>"001001111",
  31666=>"010000000",
  31667=>"001101100",
  31668=>"010111100",
  31669=>"010101010",
  31670=>"111010111",
  31671=>"111110000",
  31672=>"000100100",
  31673=>"111010100",
  31674=>"011010111",
  31675=>"001111110",
  31676=>"110000101",
  31677=>"001001000",
  31678=>"100110101",
  31679=>"010000100",
  31680=>"100100001",
  31681=>"001111100",
  31682=>"011110001",
  31683=>"100000001",
  31684=>"110100000",
  31685=>"111001111",
  31686=>"100011101",
  31687=>"100101110",
  31688=>"010110010",
  31689=>"010110010",
  31690=>"100001001",
  31691=>"001010000",
  31692=>"001111111",
  31693=>"111101011",
  31694=>"100100011",
  31695=>"100111101",
  31696=>"010011010",
  31697=>"001010001",
  31698=>"000000100",
  31699=>"100011111",
  31700=>"010101110",
  31701=>"111000001",
  31702=>"110111000",
  31703=>"011101110",
  31704=>"000100011",
  31705=>"101111110",
  31706=>"000111110",
  31707=>"011100101",
  31708=>"111101011",
  31709=>"111011000",
  31710=>"110001001",
  31711=>"110010011",
  31712=>"110111101",
  31713=>"111101011",
  31714=>"110100010",
  31715=>"111110100",
  31716=>"010011011",
  31717=>"010110101",
  31718=>"110110000",
  31719=>"101010110",
  31720=>"001010000",
  31721=>"000010110",
  31722=>"101011101",
  31723=>"011011011",
  31724=>"110100110",
  31725=>"001111001",
  31726=>"111001110",
  31727=>"110001000",
  31728=>"101111101",
  31729=>"101101101",
  31730=>"000010100",
  31731=>"110101011",
  31732=>"111000100",
  31733=>"010011001",
  31734=>"001110101",
  31735=>"101010001",
  31736=>"110011101",
  31737=>"100000010",
  31738=>"110011011",
  31739=>"001111110",
  31740=>"010001110",
  31741=>"000111101",
  31742=>"101011100",
  31743=>"110100010",
  31744=>"110000000",
  31745=>"011101101",
  31746=>"001111011",
  31747=>"111110110",
  31748=>"001001111",
  31749=>"100000000",
  31750=>"100111011",
  31751=>"001001111",
  31752=>"000100010",
  31753=>"110000010",
  31754=>"011101111",
  31755=>"000000100",
  31756=>"101000000",
  31757=>"111110110",
  31758=>"011100001",
  31759=>"100101100",
  31760=>"001110100",
  31761=>"100010010",
  31762=>"011000000",
  31763=>"010000110",
  31764=>"111010110",
  31765=>"011101100",
  31766=>"110110000",
  31767=>"010011000",
  31768=>"011111001",
  31769=>"100010111",
  31770=>"000101011",
  31771=>"111001010",
  31772=>"111111101",
  31773=>"010001011",
  31774=>"001111111",
  31775=>"101111111",
  31776=>"101011111",
  31777=>"011011101",
  31778=>"000011100",
  31779=>"101010100",
  31780=>"001110000",
  31781=>"010101010",
  31782=>"010101011",
  31783=>"001100110",
  31784=>"000000101",
  31785=>"011111001",
  31786=>"010111011",
  31787=>"111111001",
  31788=>"110011110",
  31789=>"011110100",
  31790=>"111110010",
  31791=>"101100101",
  31792=>"010100111",
  31793=>"110100011",
  31794=>"100011011",
  31795=>"010000100",
  31796=>"111001101",
  31797=>"011111011",
  31798=>"000101001",
  31799=>"000011000",
  31800=>"000101100",
  31801=>"101101101",
  31802=>"000110100",
  31803=>"100000001",
  31804=>"001100001",
  31805=>"000010110",
  31806=>"000011100",
  31807=>"011000010",
  31808=>"011010001",
  31809=>"001110001",
  31810=>"110000000",
  31811=>"001101100",
  31812=>"110100011",
  31813=>"111111101",
  31814=>"100000111",
  31815=>"010101000",
  31816=>"110111001",
  31817=>"001010010",
  31818=>"010011010",
  31819=>"000110111",
  31820=>"101001100",
  31821=>"010011001",
  31822=>"011001010",
  31823=>"100000100",
  31824=>"101001011",
  31825=>"001000101",
  31826=>"111111111",
  31827=>"110000111",
  31828=>"100111111",
  31829=>"010100010",
  31830=>"010011000",
  31831=>"001010101",
  31832=>"101111111",
  31833=>"111011100",
  31834=>"100110101",
  31835=>"000110100",
  31836=>"101000110",
  31837=>"000101001",
  31838=>"111010010",
  31839=>"010011111",
  31840=>"010100010",
  31841=>"101101111",
  31842=>"010001101",
  31843=>"101001001",
  31844=>"101111100",
  31845=>"000110100",
  31846=>"101111110",
  31847=>"000010110",
  31848=>"111111101",
  31849=>"100100010",
  31850=>"001000100",
  31851=>"000101000",
  31852=>"010100000",
  31853=>"110111101",
  31854=>"110010111",
  31855=>"011010011",
  31856=>"101110111",
  31857=>"101100100",
  31858=>"011101100",
  31859=>"000010111",
  31860=>"000111101",
  31861=>"000100000",
  31862=>"001011001",
  31863=>"100100010",
  31864=>"111111010",
  31865=>"001100000",
  31866=>"010110101",
  31867=>"100101111",
  31868=>"000100001",
  31869=>"000110100",
  31870=>"010111111",
  31871=>"101001000",
  31872=>"111100011",
  31873=>"011111010",
  31874=>"100100101",
  31875=>"101000010",
  31876=>"000101011",
  31877=>"000010011",
  31878=>"110000010",
  31879=>"110100011",
  31880=>"101111101",
  31881=>"011101010",
  31882=>"000110010",
  31883=>"010101110",
  31884=>"010011011",
  31885=>"111101101",
  31886=>"111011011",
  31887=>"101100000",
  31888=>"000101010",
  31889=>"010010011",
  31890=>"101110110",
  31891=>"010101100",
  31892=>"111110010",
  31893=>"000000110",
  31894=>"110101010",
  31895=>"011000001",
  31896=>"100110101",
  31897=>"011010000",
  31898=>"010101001",
  31899=>"001100001",
  31900=>"101101010",
  31901=>"101011001",
  31902=>"110111011",
  31903=>"011010100",
  31904=>"111100101",
  31905=>"011010011",
  31906=>"100100101",
  31907=>"101010000",
  31908=>"001100001",
  31909=>"111011010",
  31910=>"000101110",
  31911=>"110010110",
  31912=>"111101101",
  31913=>"010001000",
  31914=>"011100110",
  31915=>"011001011",
  31916=>"010001111",
  31917=>"001111110",
  31918=>"100011110",
  31919=>"011001111",
  31920=>"000001010",
  31921=>"011110111",
  31922=>"111100010",
  31923=>"100010001",
  31924=>"110010100",
  31925=>"100111000",
  31926=>"011110100",
  31927=>"001100000",
  31928=>"011111101",
  31929=>"101000000",
  31930=>"101101011",
  31931=>"011111111",
  31932=>"110011010",
  31933=>"010101000",
  31934=>"000111111",
  31935=>"100001001",
  31936=>"010000001",
  31937=>"101000011",
  31938=>"001100010",
  31939=>"000011110",
  31940=>"100001100",
  31941=>"101000000",
  31942=>"011100101",
  31943=>"000100101",
  31944=>"111001010",
  31945=>"011011011",
  31946=>"101010001",
  31947=>"101000100",
  31948=>"101001111",
  31949=>"000111010",
  31950=>"100001001",
  31951=>"000101101",
  31952=>"111010111",
  31953=>"100101011",
  31954=>"110100010",
  31955=>"111111111",
  31956=>"101111110",
  31957=>"101000111",
  31958=>"001100100",
  31959=>"010101001",
  31960=>"000001111",
  31961=>"010010011",
  31962=>"101000101",
  31963=>"001010000",
  31964=>"010101111",
  31965=>"010011110",
  31966=>"010101101",
  31967=>"000111000",
  31968=>"011101101",
  31969=>"000110010",
  31970=>"000111101",
  31971=>"001101001",
  31972=>"010100100",
  31973=>"000110000",
  31974=>"110001100",
  31975=>"010000011",
  31976=>"111100010",
  31977=>"010010111",
  31978=>"010001101",
  31979=>"111010010",
  31980=>"100100011",
  31981=>"001011001",
  31982=>"010101101",
  31983=>"000010001",
  31984=>"111001000",
  31985=>"010010010",
  31986=>"110011101",
  31987=>"000011101",
  31988=>"000100000",
  31989=>"101111001",
  31990=>"011001001",
  31991=>"011100000",
  31992=>"011011000",
  31993=>"111100100",
  31994=>"111011011",
  31995=>"010111100",
  31996=>"001101011",
  31997=>"110011101",
  31998=>"000101101",
  31999=>"110011011",
  32000=>"111110110",
  32001=>"100001100",
  32002=>"010010011",
  32003=>"100110010",
  32004=>"001000010",
  32005=>"100110000",
  32006=>"110000101",
  32007=>"110101110",
  32008=>"100111111",
  32009=>"111011001",
  32010=>"010000001",
  32011=>"001001000",
  32012=>"010100011",
  32013=>"011011100",
  32014=>"010011101",
  32015=>"010000011",
  32016=>"100100010",
  32017=>"010111111",
  32018=>"111101001",
  32019=>"111001010",
  32020=>"101101010",
  32021=>"110001000",
  32022=>"001110010",
  32023=>"010100011",
  32024=>"001010100",
  32025=>"111111110",
  32026=>"000101111",
  32027=>"000101001",
  32028=>"111000011",
  32029=>"000000101",
  32030=>"001100111",
  32031=>"001110001",
  32032=>"000000011",
  32033=>"111110001",
  32034=>"010111101",
  32035=>"001101000",
  32036=>"100011100",
  32037=>"100000101",
  32038=>"101010100",
  32039=>"001110101",
  32040=>"110111000",
  32041=>"101010011",
  32042=>"111101111",
  32043=>"111101001",
  32044=>"100010010",
  32045=>"010000100",
  32046=>"100000000",
  32047=>"000001111",
  32048=>"100110101",
  32049=>"110011111",
  32050=>"100010111",
  32051=>"101110010",
  32052=>"110000101",
  32053=>"000001000",
  32054=>"111001000",
  32055=>"000010000",
  32056=>"111100110",
  32057=>"110110010",
  32058=>"111101011",
  32059=>"001111111",
  32060=>"110100001",
  32061=>"010100000",
  32062=>"100001001",
  32063=>"110111110",
  32064=>"011101011",
  32065=>"011001000",
  32066=>"101111000",
  32067=>"101111111",
  32068=>"100110001",
  32069=>"100101110",
  32070=>"000011011",
  32071=>"101000111",
  32072=>"101111110",
  32073=>"110110110",
  32074=>"111011001",
  32075=>"011011001",
  32076=>"100011000",
  32077=>"001011000",
  32078=>"011100010",
  32079=>"011111010",
  32080=>"111001010",
  32081=>"111001010",
  32082=>"100110000",
  32083=>"010100000",
  32084=>"000100100",
  32085=>"010010110",
  32086=>"000100100",
  32087=>"000010000",
  32088=>"111101110",
  32089=>"010010101",
  32090=>"101010110",
  32091=>"010100001",
  32092=>"110100011",
  32093=>"000001100",
  32094=>"001001111",
  32095=>"001111011",
  32096=>"010001001",
  32097=>"001001100",
  32098=>"001101010",
  32099=>"011101011",
  32100=>"111011111",
  32101=>"110101101",
  32102=>"110110001",
  32103=>"110001101",
  32104=>"001111111",
  32105=>"101111000",
  32106=>"101010011",
  32107=>"011001110",
  32108=>"011001001",
  32109=>"000000000",
  32110=>"100000110",
  32111=>"000111100",
  32112=>"010011001",
  32113=>"100010101",
  32114=>"110001000",
  32115=>"011010000",
  32116=>"100100110",
  32117=>"011101001",
  32118=>"100000011",
  32119=>"111010001",
  32120=>"101010111",
  32121=>"011010011",
  32122=>"101110101",
  32123=>"010011000",
  32124=>"111000101",
  32125=>"001111001",
  32126=>"000000110",
  32127=>"000000110",
  32128=>"111011011",
  32129=>"111101010",
  32130=>"110010001",
  32131=>"101110010",
  32132=>"011110101",
  32133=>"111110110",
  32134=>"101111010",
  32135=>"100101001",
  32136=>"100001000",
  32137=>"100110000",
  32138=>"111001010",
  32139=>"000011000",
  32140=>"000100101",
  32141=>"101101001",
  32142=>"011100001",
  32143=>"111110101",
  32144=>"010101100",
  32145=>"001011001",
  32146=>"000100110",
  32147=>"100010111",
  32148=>"100110011",
  32149=>"000111101",
  32150=>"000110100",
  32151=>"111000001",
  32152=>"101100001",
  32153=>"001100001",
  32154=>"101111111",
  32155=>"000000000",
  32156=>"010110111",
  32157=>"100110100",
  32158=>"101001000",
  32159=>"110101110",
  32160=>"010000001",
  32161=>"000000111",
  32162=>"100011101",
  32163=>"011000000",
  32164=>"010011001",
  32165=>"100010101",
  32166=>"110101000",
  32167=>"000001011",
  32168=>"001001011",
  32169=>"101100100",
  32170=>"101111000",
  32171=>"111101000",
  32172=>"001000000",
  32173=>"101010110",
  32174=>"101000101",
  32175=>"111110101",
  32176=>"101011111",
  32177=>"010000000",
  32178=>"000001101",
  32179=>"011111110",
  32180=>"110011010",
  32181=>"100101110",
  32182=>"110011010",
  32183=>"101011000",
  32184=>"000001010",
  32185=>"011010111",
  32186=>"101011101",
  32187=>"001110100",
  32188=>"101110000",
  32189=>"110000111",
  32190=>"100011100",
  32191=>"100111111",
  32192=>"001001111",
  32193=>"101011100",
  32194=>"110010011",
  32195=>"100110001",
  32196=>"100101011",
  32197=>"101001000",
  32198=>"001000111",
  32199=>"011011111",
  32200=>"011101110",
  32201=>"110011000",
  32202=>"001011111",
  32203=>"010011010",
  32204=>"001000100",
  32205=>"111111010",
  32206=>"110000100",
  32207=>"100110010",
  32208=>"111100110",
  32209=>"101101101",
  32210=>"011100101",
  32211=>"101000001",
  32212=>"000000001",
  32213=>"110100000",
  32214=>"000001011",
  32215=>"111000001",
  32216=>"010110100",
  32217=>"000001110",
  32218=>"011110100",
  32219=>"011011111",
  32220=>"101101101",
  32221=>"010110010",
  32222=>"010100000",
  32223=>"011100100",
  32224=>"011100010",
  32225=>"110100010",
  32226=>"000001000",
  32227=>"010111111",
  32228=>"101101100",
  32229=>"101110010",
  32230=>"000000010",
  32231=>"100000001",
  32232=>"101101101",
  32233=>"100000101",
  32234=>"000001011",
  32235=>"110001101",
  32236=>"101001110",
  32237=>"001001100",
  32238=>"111001110",
  32239=>"010101111",
  32240=>"110111101",
  32241=>"111110111",
  32242=>"111110111",
  32243=>"010001100",
  32244=>"111001110",
  32245=>"111000110",
  32246=>"100010110",
  32247=>"001010000",
  32248=>"100101111",
  32249=>"011101011",
  32250=>"100111000",
  32251=>"101110011",
  32252=>"110111010",
  32253=>"001000000",
  32254=>"010111000",
  32255=>"001000100",
  32256=>"011111000",
  32257=>"111111110",
  32258=>"011010001",
  32259=>"100101101",
  32260=>"010101011",
  32261=>"100111101",
  32262=>"000100011",
  32263=>"111111101",
  32264=>"001000100",
  32265=>"100101101",
  32266=>"001000010",
  32267=>"110100010",
  32268=>"000100101",
  32269=>"111101111",
  32270=>"000111001",
  32271=>"001110000",
  32272=>"000010100",
  32273=>"011000011",
  32274=>"101100101",
  32275=>"111011101",
  32276=>"110001111",
  32277=>"011011110",
  32278=>"010111011",
  32279=>"001111100",
  32280=>"011001000",
  32281=>"001001101",
  32282=>"001010010",
  32283=>"100110111",
  32284=>"111111101",
  32285=>"010101110",
  32286=>"101101011",
  32287=>"010101001",
  32288=>"011001001",
  32289=>"111011111",
  32290=>"111000111",
  32291=>"101001000",
  32292=>"110111110",
  32293=>"001110101",
  32294=>"011111110",
  32295=>"000010100",
  32296=>"010110110",
  32297=>"001101100",
  32298=>"000010111",
  32299=>"110000101",
  32300=>"011111010",
  32301=>"001111111",
  32302=>"001111100",
  32303=>"010011110",
  32304=>"100001100",
  32305=>"110010000",
  32306=>"101100100",
  32307=>"101010011",
  32308=>"111001111",
  32309=>"111110100",
  32310=>"001111111",
  32311=>"110011000",
  32312=>"001110101",
  32313=>"101001001",
  32314=>"110100010",
  32315=>"111011111",
  32316=>"111000011",
  32317=>"010010001",
  32318=>"100001001",
  32319=>"010010101",
  32320=>"111101001",
  32321=>"011100101",
  32322=>"011001011",
  32323=>"001101011",
  32324=>"001100101",
  32325=>"111011010",
  32326=>"101000001",
  32327=>"001101100",
  32328=>"010101111",
  32329=>"010111100",
  32330=>"000001100",
  32331=>"100100001",
  32332=>"111100010",
  32333=>"000000001",
  32334=>"000000011",
  32335=>"101011100",
  32336=>"011111110",
  32337=>"111111000",
  32338=>"100010000",
  32339=>"100010100",
  32340=>"111111000",
  32341=>"001011011",
  32342=>"111011110",
  32343=>"010001000",
  32344=>"110111010",
  32345=>"001001011",
  32346=>"111010110",
  32347=>"111101000",
  32348=>"000010011",
  32349=>"001110000",
  32350=>"010101000",
  32351=>"110011101",
  32352=>"100100000",
  32353=>"011110101",
  32354=>"110111101",
  32355=>"011110001",
  32356=>"101100010",
  32357=>"011001000",
  32358=>"110101000",
  32359=>"000110001",
  32360=>"111000101",
  32361=>"011011110",
  32362=>"100100000",
  32363=>"111010111",
  32364=>"011110111",
  32365=>"110101001",
  32366=>"000110110",
  32367=>"101000001",
  32368=>"001111111",
  32369=>"101100101",
  32370=>"011010001",
  32371=>"100000010",
  32372=>"111100010",
  32373=>"001010011",
  32374=>"011000011",
  32375=>"111110011",
  32376=>"000111101",
  32377=>"100011010",
  32378=>"011101010",
  32379=>"100010100",
  32380=>"011100101",
  32381=>"100110111",
  32382=>"100110011",
  32383=>"100101101",
  32384=>"101001101",
  32385=>"111000111",
  32386=>"110000101",
  32387=>"000000100",
  32388=>"111111001",
  32389=>"001111010",
  32390=>"110101100",
  32391=>"110101001",
  32392=>"101111100",
  32393=>"000101111",
  32394=>"101110010",
  32395=>"011110111",
  32396=>"000010000",
  32397=>"001000100",
  32398=>"001101101",
  32399=>"111110101",
  32400=>"100101001",
  32401=>"101110000",
  32402=>"000010011",
  32403=>"010000001",
  32404=>"110101110",
  32405=>"001111001",
  32406=>"000000001",
  32407=>"111010100",
  32408=>"011000001",
  32409=>"111110010",
  32410=>"001101000",
  32411=>"101111100",
  32412=>"110111100",
  32413=>"111001100",
  32414=>"010100100",
  32415=>"000001010",
  32416=>"010000101",
  32417=>"000101100",
  32418=>"100011011",
  32419=>"000001010",
  32420=>"101111110",
  32421=>"100001000",
  32422=>"110111001",
  32423=>"101001110",
  32424=>"100101000",
  32425=>"001111111",
  32426=>"000010111",
  32427=>"110110100",
  32428=>"111111000",
  32429=>"100011111",
  32430=>"111101010",
  32431=>"011001111",
  32432=>"111000000",
  32433=>"100101011",
  32434=>"111100010",
  32435=>"100011000",
  32436=>"111110110",
  32437=>"100100011",
  32438=>"111111111",
  32439=>"001110111",
  32440=>"111001101",
  32441=>"101100101",
  32442=>"110010100",
  32443=>"001100011",
  32444=>"001100010",
  32445=>"011100001",
  32446=>"001101000",
  32447=>"111101100",
  32448=>"101110011",
  32449=>"111100110",
  32450=>"100101110",
  32451=>"101111011",
  32452=>"010101101",
  32453=>"000101001",
  32454=>"111001101",
  32455=>"011010010",
  32456=>"001010110",
  32457=>"111111010",
  32458=>"010000000",
  32459=>"111100101",
  32460=>"101100000",
  32461=>"101000011",
  32462=>"111101101",
  32463=>"000001011",
  32464=>"011110111",
  32465=>"000101110",
  32466=>"001011101",
  32467=>"000010010",
  32468=>"100000011",
  32469=>"000111010",
  32470=>"100010100",
  32471=>"101111110",
  32472=>"001000101",
  32473=>"011000110",
  32474=>"100100110",
  32475=>"010000010",
  32476=>"011000101",
  32477=>"110110011",
  32478=>"110110100",
  32479=>"101000101",
  32480=>"001101000",
  32481=>"101111001",
  32482=>"011000110",
  32483=>"011010010",
  32484=>"110000100",
  32485=>"000100101",
  32486=>"101010000",
  32487=>"001011100",
  32488=>"000010111",
  32489=>"100101011",
  32490=>"111101011",
  32491=>"111011110",
  32492=>"101100101",
  32493=>"000010101",
  32494=>"000001111",
  32495=>"101110101",
  32496=>"010111011",
  32497=>"000010011",
  32498=>"011100101",
  32499=>"111001110",
  32500=>"101011111",
  32501=>"000110110",
  32502=>"101101011",
  32503=>"101101101",
  32504=>"101101101",
  32505=>"111011100",
  32506=>"101111011",
  32507=>"010100011",
  32508=>"011101010",
  32509=>"010011111",
  32510=>"101000100",
  32511=>"000111100",
  32512=>"011110000",
  32513=>"111001110",
  32514=>"100001010",
  32515=>"011010110",
  32516=>"011000101",
  32517=>"100111001",
  32518=>"101110110",
  32519=>"101010111",
  32520=>"010100000",
  32521=>"110101100",
  32522=>"011000101",
  32523=>"000101100",
  32524=>"001001000",
  32525=>"110101001",
  32526=>"100001101",
  32527=>"111011111",
  32528=>"010000100",
  32529=>"010001110",
  32530=>"010011010",
  32531=>"001010100",
  32532=>"100000011",
  32533=>"001010111",
  32534=>"101010101",
  32535=>"111111110",
  32536=>"011110100",
  32537=>"110010011",
  32538=>"011001110",
  32539=>"000010111",
  32540=>"010010001",
  32541=>"110011000",
  32542=>"011111000",
  32543=>"001000011",
  32544=>"000011011",
  32545=>"001000010",
  32546=>"001001010",
  32547=>"000000101",
  32548=>"011101111",
  32549=>"010011000",
  32550=>"001011000",
  32551=>"101100100",
  32552=>"010010100",
  32553=>"111110100",
  32554=>"100101101",
  32555=>"110111101",
  32556=>"011111010",
  32557=>"100111010",
  32558=>"100101110",
  32559=>"100000010",
  32560=>"000110111",
  32561=>"001100111",
  32562=>"011100001",
  32563=>"000011001",
  32564=>"010001111",
  32565=>"011010010",
  32566=>"001101001",
  32567=>"011011010",
  32568=>"110101001",
  32569=>"101101100",
  32570=>"011101110",
  32571=>"011110100",
  32572=>"111010111",
  32573=>"000100100",
  32574=>"000011001",
  32575=>"100110111",
  32576=>"100011100",
  32577=>"010111101",
  32578=>"100000011",
  32579=>"100001110",
  32580=>"000010000",
  32581=>"100001010",
  32582=>"100011101",
  32583=>"010000111",
  32584=>"111010100",
  32585=>"010110000",
  32586=>"110000001",
  32587=>"110010011",
  32588=>"001101110",
  32589=>"010010111",
  32590=>"001111101",
  32591=>"001000000",
  32592=>"010010001",
  32593=>"101001000",
  32594=>"011000101",
  32595=>"011111101",
  32596=>"111001010",
  32597=>"010101111",
  32598=>"100101001",
  32599=>"010111001",
  32600=>"011010101",
  32601=>"101100011",
  32602=>"010110101",
  32603=>"010011010",
  32604=>"111010000",
  32605=>"100100100",
  32606=>"111101100",
  32607=>"000001010",
  32608=>"001010011",
  32609=>"010110001",
  32610=>"101111111",
  32611=>"110010100",
  32612=>"111001110",
  32613=>"110000011",
  32614=>"111000010",
  32615=>"101100110",
  32616=>"001010000",
  32617=>"111110111",
  32618=>"100110010",
  32619=>"101100111",
  32620=>"001101000",
  32621=>"001000001",
  32622=>"111101000",
  32623=>"000000011",
  32624=>"111100011",
  32625=>"111000111",
  32626=>"011001001",
  32627=>"000000111",
  32628=>"101011110",
  32629=>"111101011",
  32630=>"011101111",
  32631=>"100100110",
  32632=>"100001100",
  32633=>"110110110",
  32634=>"101100010",
  32635=>"111110110",
  32636=>"111001110",
  32637=>"010100010",
  32638=>"110000000",
  32639=>"101111111",
  32640=>"100011001",
  32641=>"001011100",
  32642=>"000100000",
  32643=>"011110001",
  32644=>"100110101",
  32645=>"010001001",
  32646=>"011011011",
  32647=>"000101101",
  32648=>"111100011",
  32649=>"101001000",
  32650=>"000001000",
  32651=>"101001011",
  32652=>"110101111",
  32653=>"000101110",
  32654=>"111010000",
  32655=>"110110011",
  32656=>"101101011",
  32657=>"111101111",
  32658=>"010110011",
  32659=>"000101011",
  32660=>"111111100",
  32661=>"011001111",
  32662=>"010000110",
  32663=>"110010011",
  32664=>"111111100",
  32665=>"000001000",
  32666=>"001111101",
  32667=>"010000000",
  32668=>"100111111",
  32669=>"111001101",
  32670=>"100001110",
  32671=>"101001000",
  32672=>"001001101",
  32673=>"101101011",
  32674=>"000001000",
  32675=>"111001110",
  32676=>"000010000",
  32677=>"011111000",
  32678=>"000100110",
  32679=>"011011001",
  32680=>"111000110",
  32681=>"100111001",
  32682=>"011111000",
  32683=>"011111011",
  32684=>"111111000",
  32685=>"011111100",
  32686=>"110110111",
  32687=>"000010111",
  32688=>"101000101",
  32689=>"010110010",
  32690=>"100000100",
  32691=>"100010001",
  32692=>"000000100",
  32693=>"111001000",
  32694=>"111100110",
  32695=>"010110101",
  32696=>"111000110",
  32697=>"100011011",
  32698=>"011010000",
  32699=>"110011001",
  32700=>"010110110",
  32701=>"001011110",
  32702=>"111101111",
  32703=>"111001011",
  32704=>"110000101",
  32705=>"010010001",
  32706=>"010101000",
  32707=>"111101001",
  32708=>"000110010",
  32709=>"000110100",
  32710=>"111101100",
  32711=>"100000101",
  32712=>"101101000",
  32713=>"010110101",
  32714=>"001000000",
  32715=>"001100111",
  32716=>"000000000",
  32717=>"000000010",
  32718=>"001100100",
  32719=>"110000111",
  32720=>"000111100",
  32721=>"000100101",
  32722=>"101101000",
  32723=>"100000100",
  32724=>"010000011",
  32725=>"101010010",
  32726=>"101111110",
  32727=>"010000110",
  32728=>"001101111",
  32729=>"101001100",
  32730=>"101100110",
  32731=>"111110100",
  32732=>"011001010",
  32733=>"011101111",
  32734=>"111010011",
  32735=>"000100101",
  32736=>"111110001",
  32737=>"010010110",
  32738=>"011000010",
  32739=>"001110010",
  32740=>"000110001",
  32741=>"111111111",
  32742=>"100000000",
  32743=>"110100001",
  32744=>"001000001",
  32745=>"101011101",
  32746=>"101011010",
  32747=>"111100000",
  32748=>"000000100",
  32749=>"110011110",
  32750=>"101011110",
  32751=>"000001011",
  32752=>"110111110",
  32753=>"000010010",
  32754=>"011110001",
  32755=>"110101110",
  32756=>"111101110",
  32757=>"000111101",
  32758=>"111000000",
  32759=>"011001011",
  32760=>"110101111",
  32761=>"101011110",
  32762=>"100101111",
  32763=>"001110010",
  32764=>"000000001",
  32765=>"001100101",
  32766=>"110101000",
  32767=>"101010010",
  32768=>"001010010",
  32769=>"110000111",
  32770=>"001011000",
  32771=>"100011001",
  32772=>"000011110",
  32773=>"110011000",
  32774=>"100011010",
  32775=>"010001101",
  32776=>"101100111",
  32777=>"011101011",
  32778=>"001101111",
  32779=>"111010100",
  32780=>"101110001",
  32781=>"111111000",
  32782=>"111001010",
  32783=>"010000001",
  32784=>"000001000",
  32785=>"100010011",
  32786=>"111001111",
  32787=>"110111100",
  32788=>"010110010",
  32789=>"011101001",
  32790=>"110000000",
  32791=>"011001101",
  32792=>"100101100",
  32793=>"001000001",
  32794=>"100001010",
  32795=>"100010101",
  32796=>"100010111",
  32797=>"011011000",
  32798=>"011101011",
  32799=>"111000011",
  32800=>"100010001",
  32801=>"011000110",
  32802=>"111100111",
  32803=>"100110110",
  32804=>"101100001",
  32805=>"101111011",
  32806=>"011101101",
  32807=>"111111101",
  32808=>"111100011",
  32809=>"000001000",
  32810=>"000110001",
  32811=>"110011000",
  32812=>"000010001",
  32813=>"010010111",
  32814=>"110011101",
  32815=>"111101101",
  32816=>"110110101",
  32817=>"010100011",
  32818=>"011101011",
  32819=>"001110100",
  32820=>"100100001",
  32821=>"000100110",
  32822=>"000101111",
  32823=>"011011110",
  32824=>"000111111",
  32825=>"111011001",
  32826=>"001100100",
  32827=>"110110011",
  32828=>"101101100",
  32829=>"111001000",
  32830=>"001011011",
  32831=>"000001001",
  32832=>"110010001",
  32833=>"101010111",
  32834=>"101011101",
  32835=>"111001100",
  32836=>"111101101",
  32837=>"100111000",
  32838=>"111101100",
  32839=>"110111000",
  32840=>"001111101",
  32841=>"001100001",
  32842=>"000011111",
  32843=>"100100010",
  32844=>"000100101",
  32845=>"010100110",
  32846=>"100110111",
  32847=>"000101100",
  32848=>"011010010",
  32849=>"111010100",
  32850=>"101011011",
  32851=>"111111101",
  32852=>"110010011",
  32853=>"001010111",
  32854=>"101110110",
  32855=>"000010101",
  32856=>"001000101",
  32857=>"111000001",
  32858=>"111101001",
  32859=>"011000000",
  32860=>"100100011",
  32861=>"100111000",
  32862=>"111100111",
  32863=>"001100100",
  32864=>"011100110",
  32865=>"001110001",
  32866=>"110010001",
  32867=>"000011001",
  32868=>"011000101",
  32869=>"010111000",
  32870=>"001010101",
  32871=>"000011011",
  32872=>"110001000",
  32873=>"101111111",
  32874=>"111111111",
  32875=>"001001001",
  32876=>"000010111",
  32877=>"000010111",
  32878=>"001010000",
  32879=>"100110000",
  32880=>"110101001",
  32881=>"010001110",
  32882=>"010111111",
  32883=>"011101101",
  32884=>"110111110",
  32885=>"111111011",
  32886=>"100101111",
  32887=>"011100100",
  32888=>"111101101",
  32889=>"000110011",
  32890=>"100010000",
  32891=>"101100101",
  32892=>"011101000",
  32893=>"000110001",
  32894=>"100010000",
  32895=>"110010110",
  32896=>"010001000",
  32897=>"110101100",
  32898=>"010000111",
  32899=>"111001001",
  32900=>"111011101",
  32901=>"010110100",
  32902=>"110111101",
  32903=>"110011010",
  32904=>"110101111",
  32905=>"100001001",
  32906=>"001100111",
  32907=>"110110000",
  32908=>"101000011",
  32909=>"101000001",
  32910=>"000110011",
  32911=>"001000000",
  32912=>"011101110",
  32913=>"110010111",
  32914=>"110000001",
  32915=>"001100100",
  32916=>"110111111",
  32917=>"011101011",
  32918=>"001010010",
  32919=>"010110101",
  32920=>"111111001",
  32921=>"111001111",
  32922=>"111100011",
  32923=>"110111111",
  32924=>"110110001",
  32925=>"000100010",
  32926=>"010100011",
  32927=>"000000111",
  32928=>"101000000",
  32929=>"100110011",
  32930=>"011001111",
  32931=>"101110101",
  32932=>"111000101",
  32933=>"100110110",
  32934=>"101101011",
  32935=>"101011111",
  32936=>"101100110",
  32937=>"110000100",
  32938=>"110101101",
  32939=>"001000110",
  32940=>"110001010",
  32941=>"110001000",
  32942=>"110101001",
  32943=>"000110101",
  32944=>"010011110",
  32945=>"011111110",
  32946=>"101001111",
  32947=>"101001100",
  32948=>"110101010",
  32949=>"111001110",
  32950=>"110000010",
  32951=>"110000001",
  32952=>"111011010",
  32953=>"011111111",
  32954=>"111110010",
  32955=>"101110101",
  32956=>"101101101",
  32957=>"110010001",
  32958=>"001011111",
  32959=>"111111111",
  32960=>"100010011",
  32961=>"110111000",
  32962=>"101101010",
  32963=>"011000111",
  32964=>"010000011",
  32965=>"000010010",
  32966=>"110010001",
  32967=>"000100100",
  32968=>"110110100",
  32969=>"100001101",
  32970=>"100010110",
  32971=>"011111001",
  32972=>"111010001",
  32973=>"011010011",
  32974=>"100000000",
  32975=>"001001000",
  32976=>"011111100",
  32977=>"011001110",
  32978=>"001001000",
  32979=>"111010110",
  32980=>"010111110",
  32981=>"001110010",
  32982=>"111010110",
  32983=>"110111000",
  32984=>"011010101",
  32985=>"001001000",
  32986=>"110010001",
  32987=>"101011110",
  32988=>"011010100",
  32989=>"101011000",
  32990=>"111110111",
  32991=>"101111011",
  32992=>"001100101",
  32993=>"000100100",
  32994=>"110110001",
  32995=>"100011011",
  32996=>"000011011",
  32997=>"100101000",
  32998=>"101110011",
  32999=>"101111111",
  33000=>"100011011",
  33001=>"000111111",
  33002=>"110100000",
  33003=>"001000001",
  33004=>"110110110",
  33005=>"101110011",
  33006=>"110100001",
  33007=>"010010000",
  33008=>"011000100",
  33009=>"101110111",
  33010=>"000110101",
  33011=>"011010000",
  33012=>"010111011",
  33013=>"101011001",
  33014=>"101001101",
  33015=>"100011101",
  33016=>"110001100",
  33017=>"110010111",
  33018=>"011000000",
  33019=>"000110110",
  33020=>"110001000",
  33021=>"110001000",
  33022=>"100011100",
  33023=>"100111011",
  33024=>"100001010",
  33025=>"001010111",
  33026=>"001100110",
  33027=>"110100111",
  33028=>"100101111",
  33029=>"110001111",
  33030=>"111101100",
  33031=>"111000101",
  33032=>"010110001",
  33033=>"010010101",
  33034=>"001111100",
  33035=>"110100000",
  33036=>"001001110",
  33037=>"011100110",
  33038=>"100100010",
  33039=>"111101000",
  33040=>"111010110",
  33041=>"010101111",
  33042=>"011000101",
  33043=>"100100100",
  33044=>"101001011",
  33045=>"111111100",
  33046=>"100010000",
  33047=>"101101100",
  33048=>"000001000",
  33049=>"100010000",
  33050=>"111011010",
  33051=>"011110000",
  33052=>"001001100",
  33053=>"010000011",
  33054=>"001000111",
  33055=>"101100000",
  33056=>"101001110",
  33057=>"110110001",
  33058=>"010000000",
  33059=>"011110110",
  33060=>"001011010",
  33061=>"110010011",
  33062=>"111101101",
  33063=>"110000000",
  33064=>"111001100",
  33065=>"111101101",
  33066=>"011111110",
  33067=>"100001000",
  33068=>"101000111",
  33069=>"011000100",
  33070=>"000100110",
  33071=>"111111111",
  33072=>"111101101",
  33073=>"001000000",
  33074=>"001100101",
  33075=>"010010100",
  33076=>"011001010",
  33077=>"110011011",
  33078=>"101111000",
  33079=>"010111000",
  33080=>"010010110",
  33081=>"001001001",
  33082=>"001111111",
  33083=>"110100101",
  33084=>"101001110",
  33085=>"110001010",
  33086=>"110101100",
  33087=>"101001010",
  33088=>"110001110",
  33089=>"100101110",
  33090=>"100101000",
  33091=>"000101110",
  33092=>"101111111",
  33093=>"101100111",
  33094=>"100001010",
  33095=>"001011001",
  33096=>"001000101",
  33097=>"100010100",
  33098=>"110111100",
  33099=>"011011110",
  33100=>"000100100",
  33101=>"000110010",
  33102=>"100110001",
  33103=>"101000111",
  33104=>"011100110",
  33105=>"100001010",
  33106=>"010010011",
  33107=>"000100110",
  33108=>"100000000",
  33109=>"100011100",
  33110=>"001110000",
  33111=>"000011100",
  33112=>"000110001",
  33113=>"010010010",
  33114=>"100001001",
  33115=>"011110111",
  33116=>"110101101",
  33117=>"011001110",
  33118=>"100001011",
  33119=>"011001011",
  33120=>"110110011",
  33121=>"010000001",
  33122=>"000010011",
  33123=>"111110111",
  33124=>"111011101",
  33125=>"001110000",
  33126=>"101001011",
  33127=>"101100010",
  33128=>"100001001",
  33129=>"000010000",
  33130=>"011110100",
  33131=>"000011110",
  33132=>"111101110",
  33133=>"111010000",
  33134=>"000101111",
  33135=>"010010000",
  33136=>"011010100",
  33137=>"001110011",
  33138=>"101111000",
  33139=>"100111111",
  33140=>"011010001",
  33141=>"010011000",
  33142=>"111101001",
  33143=>"011111110",
  33144=>"101001110",
  33145=>"010000001",
  33146=>"001101001",
  33147=>"010001001",
  33148=>"100100010",
  33149=>"111110111",
  33150=>"101101010",
  33151=>"111111111",
  33152=>"100010001",
  33153=>"000011010",
  33154=>"101101110",
  33155=>"000000111",
  33156=>"111101010",
  33157=>"111100100",
  33158=>"000111101",
  33159=>"111111011",
  33160=>"100001110",
  33161=>"010010010",
  33162=>"000100100",
  33163=>"001001011",
  33164=>"001001110",
  33165=>"010111000",
  33166=>"100101001",
  33167=>"010001010",
  33168=>"110101111",
  33169=>"100110101",
  33170=>"010100010",
  33171=>"100000010",
  33172=>"111101010",
  33173=>"111011110",
  33174=>"110010110",
  33175=>"100111111",
  33176=>"011100010",
  33177=>"011011011",
  33178=>"100001001",
  33179=>"010001110",
  33180=>"001001110",
  33181=>"110111111",
  33182=>"001100001",
  33183=>"110000100",
  33184=>"011111000",
  33185=>"111011000",
  33186=>"110010000",
  33187=>"100000011",
  33188=>"101010101",
  33189=>"110001010",
  33190=>"101011010",
  33191=>"010010111",
  33192=>"110110111",
  33193=>"100100100",
  33194=>"110000001",
  33195=>"011001110",
  33196=>"110011101",
  33197=>"111000000",
  33198=>"010110100",
  33199=>"010101010",
  33200=>"100000001",
  33201=>"001110100",
  33202=>"100001000",
  33203=>"010101011",
  33204=>"111100101",
  33205=>"000000101",
  33206=>"111000011",
  33207=>"110001010",
  33208=>"111001001",
  33209=>"100001011",
  33210=>"011011000",
  33211=>"011001111",
  33212=>"001010001",
  33213=>"001111010",
  33214=>"100100110",
  33215=>"001011101",
  33216=>"010001111",
  33217=>"010001100",
  33218=>"001100110",
  33219=>"000010010",
  33220=>"110011100",
  33221=>"001101000",
  33222=>"111101000",
  33223=>"010111010",
  33224=>"010001011",
  33225=>"010101010",
  33226=>"110001000",
  33227=>"110111100",
  33228=>"101110001",
  33229=>"011000101",
  33230=>"010101100",
  33231=>"100101001",
  33232=>"101000000",
  33233=>"111100110",
  33234=>"111001000",
  33235=>"000011001",
  33236=>"110010100",
  33237=>"110001100",
  33238=>"100100010",
  33239=>"001010011",
  33240=>"011101010",
  33241=>"000000010",
  33242=>"110100110",
  33243=>"110101100",
  33244=>"000101101",
  33245=>"111011000",
  33246=>"010111100",
  33247=>"111000010",
  33248=>"000000011",
  33249=>"111101110",
  33250=>"111011100",
  33251=>"111001100",
  33252=>"001101100",
  33253=>"111101111",
  33254=>"011011000",
  33255=>"111001110",
  33256=>"101110100",
  33257=>"110011000",
  33258=>"000100000",
  33259=>"000010000",
  33260=>"000111101",
  33261=>"001110100",
  33262=>"100000010",
  33263=>"111100110",
  33264=>"110111101",
  33265=>"001100000",
  33266=>"100000010",
  33267=>"010001010",
  33268=>"101110100",
  33269=>"101001100",
  33270=>"101001010",
  33271=>"000110110",
  33272=>"000001000",
  33273=>"010000001",
  33274=>"111111011",
  33275=>"101111011",
  33276=>"010011100",
  33277=>"111101100",
  33278=>"000010110",
  33279=>"111101100",
  33280=>"011110011",
  33281=>"001100110",
  33282=>"001011001",
  33283=>"110001101",
  33284=>"000110111",
  33285=>"000011001",
  33286=>"010110011",
  33287=>"111101111",
  33288=>"010010100",
  33289=>"110100111",
  33290=>"000110110",
  33291=>"000011111",
  33292=>"101101001",
  33293=>"111001111",
  33294=>"000000100",
  33295=>"000001000",
  33296=>"110100000",
  33297=>"000001011",
  33298=>"101011010",
  33299=>"110111011",
  33300=>"000000000",
  33301=>"010011110",
  33302=>"000100100",
  33303=>"001101010",
  33304=>"001000001",
  33305=>"011101111",
  33306=>"000000001",
  33307=>"110100001",
  33308=>"111111100",
  33309=>"011000000",
  33310=>"110001001",
  33311=>"111010001",
  33312=>"011001010",
  33313=>"101010001",
  33314=>"110001000",
  33315=>"011110110",
  33316=>"000011011",
  33317=>"111010011",
  33318=>"011110111",
  33319=>"010101010",
  33320=>"100111010",
  33321=>"110101101",
  33322=>"101110011",
  33323=>"010011100",
  33324=>"110000000",
  33325=>"110001011",
  33326=>"101001000",
  33327=>"111101101",
  33328=>"101100011",
  33329=>"101011001",
  33330=>"010101101",
  33331=>"010100001",
  33332=>"101000011",
  33333=>"101101010",
  33334=>"010010011",
  33335=>"111110101",
  33336=>"000000001",
  33337=>"000010011",
  33338=>"110010110",
  33339=>"000111011",
  33340=>"101000111",
  33341=>"100000100",
  33342=>"001001100",
  33343=>"100011010",
  33344=>"001000100",
  33345=>"001101011",
  33346=>"010111110",
  33347=>"010001001",
  33348=>"100001100",
  33349=>"000011100",
  33350=>"111001001",
  33351=>"111110101",
  33352=>"111100101",
  33353=>"001101111",
  33354=>"100010011",
  33355=>"001101010",
  33356=>"110101000",
  33357=>"100110110",
  33358=>"011100110",
  33359=>"110101010",
  33360=>"111111010",
  33361=>"111111100",
  33362=>"000010111",
  33363=>"100100001",
  33364=>"100101100",
  33365=>"110110100",
  33366=>"001010000",
  33367=>"010011110",
  33368=>"111101111",
  33369=>"010000001",
  33370=>"000110001",
  33371=>"101110100",
  33372=>"110101101",
  33373=>"110101100",
  33374=>"101001101",
  33375=>"101001011",
  33376=>"110100101",
  33377=>"000100011",
  33378=>"001001101",
  33379=>"001000101",
  33380=>"101100100",
  33381=>"010010111",
  33382=>"101110100",
  33383=>"111111111",
  33384=>"101111110",
  33385=>"001100000",
  33386=>"010111001",
  33387=>"010110001",
  33388=>"110011100",
  33389=>"000010001",
  33390=>"010111101",
  33391=>"111001111",
  33392=>"000011110",
  33393=>"101100100",
  33394=>"010010001",
  33395=>"001110001",
  33396=>"111011011",
  33397=>"000011101",
  33398=>"110010001",
  33399=>"011101010",
  33400=>"111100110",
  33401=>"100101110",
  33402=>"111010001",
  33403=>"110010010",
  33404=>"001001110",
  33405=>"001010001",
  33406=>"011110111",
  33407=>"000011000",
  33408=>"011010101",
  33409=>"100101000",
  33410=>"100111110",
  33411=>"100001101",
  33412=>"000111010",
  33413=>"001111101",
  33414=>"111110111",
  33415=>"011111111",
  33416=>"010110000",
  33417=>"100010011",
  33418=>"111111111",
  33419=>"010100101",
  33420=>"000001000",
  33421=>"011000010",
  33422=>"010010101",
  33423=>"011001001",
  33424=>"110000000",
  33425=>"000111001",
  33426=>"001101101",
  33427=>"000101110",
  33428=>"101000000",
  33429=>"001111110",
  33430=>"000000011",
  33431=>"010110010",
  33432=>"011110011",
  33433=>"001110000",
  33434=>"011100010",
  33435=>"110111100",
  33436=>"110001011",
  33437=>"001011011",
  33438=>"001011110",
  33439=>"100110000",
  33440=>"001111100",
  33441=>"000010011",
  33442=>"101000111",
  33443=>"100101100",
  33444=>"110001011",
  33445=>"010010010",
  33446=>"000010111",
  33447=>"001000001",
  33448=>"111100010",
  33449=>"001000011",
  33450=>"011001111",
  33451=>"010010110",
  33452=>"010010110",
  33453=>"011001111",
  33454=>"111011100",
  33455=>"111010101",
  33456=>"010110101",
  33457=>"110101011",
  33458=>"110010010",
  33459=>"000110010",
  33460=>"000001010",
  33461=>"000111000",
  33462=>"100101000",
  33463=>"000101101",
  33464=>"111011001",
  33465=>"110000001",
  33466=>"000111100",
  33467=>"110111011",
  33468=>"110111110",
  33469=>"000000011",
  33470=>"001011100",
  33471=>"000011100",
  33472=>"101100100",
  33473=>"101110100",
  33474=>"010100111",
  33475=>"000110000",
  33476=>"100101111",
  33477=>"101000101",
  33478=>"111101111",
  33479=>"110000110",
  33480=>"111000011",
  33481=>"101100110",
  33482=>"011110010",
  33483=>"000001000",
  33484=>"110010110",
  33485=>"111001001",
  33486=>"111110000",
  33487=>"011101100",
  33488=>"111011010",
  33489=>"010001010",
  33490=>"001100010",
  33491=>"100100101",
  33492=>"111010101",
  33493=>"010110000",
  33494=>"010100001",
  33495=>"011100110",
  33496=>"100010110",
  33497=>"011100001",
  33498=>"001000100",
  33499=>"010000110",
  33500=>"101001100",
  33501=>"010100000",
  33502=>"101001111",
  33503=>"100001100",
  33504=>"110111000",
  33505=>"110101010",
  33506=>"110101001",
  33507=>"001101100",
  33508=>"101101111",
  33509=>"001100110",
  33510=>"000000100",
  33511=>"101011110",
  33512=>"001011011",
  33513=>"111001010",
  33514=>"000000100",
  33515=>"100111010",
  33516=>"100111011",
  33517=>"100000001",
  33518=>"110001110",
  33519=>"010010101",
  33520=>"000001000",
  33521=>"110110100",
  33522=>"010010001",
  33523=>"110101100",
  33524=>"101101000",
  33525=>"011100111",
  33526=>"101111111",
  33527=>"111100101",
  33528=>"100100010",
  33529=>"011001111",
  33530=>"010001100",
  33531=>"000011000",
  33532=>"010011010",
  33533=>"010100001",
  33534=>"000110001",
  33535=>"010011001",
  33536=>"011011010",
  33537=>"000011011",
  33538=>"111010100",
  33539=>"000010111",
  33540=>"001010111",
  33541=>"110100001",
  33542=>"111101001",
  33543=>"001001010",
  33544=>"010111001",
  33545=>"000100111",
  33546=>"001111110",
  33547=>"010111111",
  33548=>"111110010",
  33549=>"110011110",
  33550=>"101011011",
  33551=>"000100010",
  33552=>"000111011",
  33553=>"111110001",
  33554=>"010111010",
  33555=>"110100111",
  33556=>"111110001",
  33557=>"000110010",
  33558=>"011000001",
  33559=>"010010000",
  33560=>"111110011",
  33561=>"010100000",
  33562=>"111010100",
  33563=>"011101101",
  33564=>"100011100",
  33565=>"110111001",
  33566=>"100101010",
  33567=>"100010101",
  33568=>"010011111",
  33569=>"110110101",
  33570=>"111111111",
  33571=>"100110111",
  33572=>"110111100",
  33573=>"011110001",
  33574=>"010111110",
  33575=>"100001110",
  33576=>"010111001",
  33577=>"010100001",
  33578=>"100100111",
  33579=>"100110001",
  33580=>"000111010",
  33581=>"011000010",
  33582=>"111000001",
  33583=>"100001001",
  33584=>"000011011",
  33585=>"011000111",
  33586=>"111001000",
  33587=>"010111111",
  33588=>"110111000",
  33589=>"111101010",
  33590=>"001000100",
  33591=>"001110111",
  33592=>"110011100",
  33593=>"111110001",
  33594=>"111001101",
  33595=>"000001001",
  33596=>"001010100",
  33597=>"110000011",
  33598=>"111010010",
  33599=>"000100000",
  33600=>"101100011",
  33601=>"001111111",
  33602=>"111001011",
  33603=>"110000010",
  33604=>"000000101",
  33605=>"100000100",
  33606=>"110101111",
  33607=>"011101110",
  33608=>"110101101",
  33609=>"000010101",
  33610=>"000010101",
  33611=>"000101010",
  33612=>"101110001",
  33613=>"100011110",
  33614=>"000100010",
  33615=>"000001011",
  33616=>"011000001",
  33617=>"000000110",
  33618=>"000101111",
  33619=>"111000000",
  33620=>"011001111",
  33621=>"111010010",
  33622=>"110101100",
  33623=>"000010010",
  33624=>"110101101",
  33625=>"110011110",
  33626=>"000011101",
  33627=>"101000011",
  33628=>"110110101",
  33629=>"111100001",
  33630=>"001001110",
  33631=>"011101001",
  33632=>"011000100",
  33633=>"001010000",
  33634=>"011010011",
  33635=>"011101000",
  33636=>"000100100",
  33637=>"110100001",
  33638=>"101101111",
  33639=>"000001100",
  33640=>"010010010",
  33641=>"000000011",
  33642=>"100110001",
  33643=>"111011101",
  33644=>"100011001",
  33645=>"001111101",
  33646=>"101001001",
  33647=>"001010101",
  33648=>"001011100",
  33649=>"111110000",
  33650=>"111001100",
  33651=>"101101000",
  33652=>"001111001",
  33653=>"100111000",
  33654=>"001101010",
  33655=>"001101100",
  33656=>"111110111",
  33657=>"000100010",
  33658=>"000111010",
  33659=>"111000011",
  33660=>"000010011",
  33661=>"101001111",
  33662=>"110011000",
  33663=>"100011101",
  33664=>"010100011",
  33665=>"000000100",
  33666=>"110101111",
  33667=>"001100101",
  33668=>"011101000",
  33669=>"110100010",
  33670=>"011100111",
  33671=>"010101111",
  33672=>"001111011",
  33673=>"000100110",
  33674=>"010100000",
  33675=>"101110000",
  33676=>"111101001",
  33677=>"011010111",
  33678=>"010110110",
  33679=>"101100001",
  33680=>"010011101",
  33681=>"011001010",
  33682=>"110100001",
  33683=>"010011010",
  33684=>"011100001",
  33685=>"110000000",
  33686=>"110011101",
  33687=>"101101111",
  33688=>"100001100",
  33689=>"111100110",
  33690=>"110000001",
  33691=>"100101111",
  33692=>"110011001",
  33693=>"111111001",
  33694=>"000001100",
  33695=>"000011011",
  33696=>"101101001",
  33697=>"001110110",
  33698=>"100111010",
  33699=>"010110100",
  33700=>"110011110",
  33701=>"011111101",
  33702=>"000100101",
  33703=>"011010110",
  33704=>"011010001",
  33705=>"000100001",
  33706=>"110010011",
  33707=>"100000001",
  33708=>"111000110",
  33709=>"001011001",
  33710=>"011111011",
  33711=>"011011001",
  33712=>"011111011",
  33713=>"110001010",
  33714=>"101000011",
  33715=>"111001111",
  33716=>"110110110",
  33717=>"000010101",
  33718=>"100110000",
  33719=>"010010101",
  33720=>"111111101",
  33721=>"001110000",
  33722=>"100000011",
  33723=>"011101100",
  33724=>"101001010",
  33725=>"100101100",
  33726=>"100101101",
  33727=>"000110000",
  33728=>"100000010",
  33729=>"101101000",
  33730=>"111111101",
  33731=>"111101011",
  33732=>"110001110",
  33733=>"111101011",
  33734=>"010101100",
  33735=>"000100001",
  33736=>"010000111",
  33737=>"101010011",
  33738=>"100111011",
  33739=>"011001011",
  33740=>"001010000",
  33741=>"001100101",
  33742=>"010000000",
  33743=>"100110000",
  33744=>"000111110",
  33745=>"000111011",
  33746=>"000110100",
  33747=>"011011110",
  33748=>"011110000",
  33749=>"110100011",
  33750=>"010111001",
  33751=>"000011011",
  33752=>"011010110",
  33753=>"010000010",
  33754=>"110011101",
  33755=>"000011101",
  33756=>"010101010",
  33757=>"011011101",
  33758=>"101001001",
  33759=>"111101011",
  33760=>"101100110",
  33761=>"000100110",
  33762=>"001011101",
  33763=>"000001101",
  33764=>"010000010",
  33765=>"001010110",
  33766=>"111100000",
  33767=>"100100000",
  33768=>"000100100",
  33769=>"101010111",
  33770=>"010010101",
  33771=>"001001010",
  33772=>"111101101",
  33773=>"000100011",
  33774=>"011111100",
  33775=>"100101011",
  33776=>"001110100",
  33777=>"100111011",
  33778=>"001100100",
  33779=>"000000101",
  33780=>"100011010",
  33781=>"001100101",
  33782=>"000100101",
  33783=>"111001111",
  33784=>"110001010",
  33785=>"000110000",
  33786=>"100000101",
  33787=>"010010100",
  33788=>"000010000",
  33789=>"111011010",
  33790=>"110000110",
  33791=>"000010111",
  33792=>"000000111",
  33793=>"101110011",
  33794=>"000101010",
  33795=>"100001111",
  33796=>"111101011",
  33797=>"010001010",
  33798=>"011000011",
  33799=>"101100110",
  33800=>"111101101",
  33801=>"011010000",
  33802=>"011010110",
  33803=>"111011110",
  33804=>"100000010",
  33805=>"111100001",
  33806=>"011110110",
  33807=>"111111111",
  33808=>"011010100",
  33809=>"010000100",
  33810=>"010100011",
  33811=>"011111010",
  33812=>"000010001",
  33813=>"010100110",
  33814=>"001111100",
  33815=>"010111011",
  33816=>"101101111",
  33817=>"111011010",
  33818=>"111110101",
  33819=>"110000010",
  33820=>"110111111",
  33821=>"111110011",
  33822=>"010101110",
  33823=>"010111100",
  33824=>"100110010",
  33825=>"011010010",
  33826=>"110010001",
  33827=>"000100000",
  33828=>"101110010",
  33829=>"101000010",
  33830=>"001010000",
  33831=>"111000010",
  33832=>"100010101",
  33833=>"001110101",
  33834=>"000001010",
  33835=>"101100000",
  33836=>"000011000",
  33837=>"001100011",
  33838=>"101010110",
  33839=>"010000011",
  33840=>"100011110",
  33841=>"010110110",
  33842=>"110100000",
  33843=>"111001110",
  33844=>"010010111",
  33845=>"100101000",
  33846=>"000111110",
  33847=>"000100111",
  33848=>"000010011",
  33849=>"001001000",
  33850=>"010001100",
  33851=>"100100100",
  33852=>"001101110",
  33853=>"001110011",
  33854=>"111111100",
  33855=>"010001001",
  33856=>"010001100",
  33857=>"000011010",
  33858=>"110110001",
  33859=>"010111000",
  33860=>"110100110",
  33861=>"010111011",
  33862=>"110110111",
  33863=>"001001011",
  33864=>"100011011",
  33865=>"010001011",
  33866=>"000101110",
  33867=>"000100000",
  33868=>"101010011",
  33869=>"011001110",
  33870=>"001110110",
  33871=>"010011010",
  33872=>"101001111",
  33873=>"101111111",
  33874=>"100010101",
  33875=>"101011000",
  33876=>"101110101",
  33877=>"100011100",
  33878=>"000011100",
  33879=>"101011001",
  33880=>"001101011",
  33881=>"110010110",
  33882=>"010110010",
  33883=>"100010111",
  33884=>"110111101",
  33885=>"110000011",
  33886=>"010000011",
  33887=>"010110000",
  33888=>"001001101",
  33889=>"000101011",
  33890=>"011010111",
  33891=>"000110000",
  33892=>"100001111",
  33893=>"011001000",
  33894=>"101000000",
  33895=>"110100010",
  33896=>"100110010",
  33897=>"100011101",
  33898=>"010000001",
  33899=>"111010001",
  33900=>"011111011",
  33901=>"000001000",
  33902=>"010101101",
  33903=>"110011011",
  33904=>"000100111",
  33905=>"100000101",
  33906=>"010111001",
  33907=>"100101101",
  33908=>"000101111",
  33909=>"011101101",
  33910=>"100101101",
  33911=>"110000110",
  33912=>"011011011",
  33913=>"100001001",
  33914=>"111101111",
  33915=>"110000100",
  33916=>"101100111",
  33917=>"111011100",
  33918=>"100001111",
  33919=>"000010001",
  33920=>"010000100",
  33921=>"111111100",
  33922=>"000001000",
  33923=>"111010111",
  33924=>"110010000",
  33925=>"011001101",
  33926=>"010011110",
  33927=>"011100100",
  33928=>"010111010",
  33929=>"000000001",
  33930=>"101101110",
  33931=>"011010111",
  33932=>"110101011",
  33933=>"010010110",
  33934=>"111111111",
  33935=>"000011101",
  33936=>"100000111",
  33937=>"111101111",
  33938=>"100011010",
  33939=>"100101111",
  33940=>"100001001",
  33941=>"001111100",
  33942=>"000100011",
  33943=>"101000011",
  33944=>"101100010",
  33945=>"010100010",
  33946=>"101010101",
  33947=>"000100000",
  33948=>"100111101",
  33949=>"001011001",
  33950=>"101000101",
  33951=>"001100111",
  33952=>"011110100",
  33953=>"010100001",
  33954=>"011111111",
  33955=>"101001000",
  33956=>"111110000",
  33957=>"001010011",
  33958=>"100100111",
  33959=>"010000001",
  33960=>"001111001",
  33961=>"000100110",
  33962=>"000001011",
  33963=>"111111111",
  33964=>"101101010",
  33965=>"011001100",
  33966=>"001110000",
  33967=>"001011100",
  33968=>"111111001",
  33969=>"011010000",
  33970=>"001011111",
  33971=>"100111110",
  33972=>"010001011",
  33973=>"001101001",
  33974=>"000011011",
  33975=>"100110010",
  33976=>"010100001",
  33977=>"011100100",
  33978=>"101010110",
  33979=>"111101110",
  33980=>"001100110",
  33981=>"110101111",
  33982=>"100110110",
  33983=>"100001110",
  33984=>"001000001",
  33985=>"110010010",
  33986=>"110011111",
  33987=>"010010001",
  33988=>"101101000",
  33989=>"110001000",
  33990=>"100011111",
  33991=>"100001010",
  33992=>"101101110",
  33993=>"111010011",
  33994=>"111011000",
  33995=>"100100010",
  33996=>"010001111",
  33997=>"001010101",
  33998=>"111100110",
  33999=>"000100111",
  34000=>"110011111",
  34001=>"111000000",
  34002=>"111111000",
  34003=>"100001110",
  34004=>"000000110",
  34005=>"001110001",
  34006=>"010101100",
  34007=>"011100000",
  34008=>"000111100",
  34009=>"001010100",
  34010=>"000010010",
  34011=>"001100001",
  34012=>"100101001",
  34013=>"110001011",
  34014=>"100101001",
  34015=>"110010000",
  34016=>"101100101",
  34017=>"100011110",
  34018=>"001011100",
  34019=>"010010110",
  34020=>"010100010",
  34021=>"101001111",
  34022=>"000010001",
  34023=>"111101111",
  34024=>"001000000",
  34025=>"001111011",
  34026=>"010001001",
  34027=>"011000000",
  34028=>"001001000",
  34029=>"000010011",
  34030=>"010100110",
  34031=>"100000111",
  34032=>"100011010",
  34033=>"010010010",
  34034=>"011111111",
  34035=>"011010011",
  34036=>"100011011",
  34037=>"000001000",
  34038=>"011000001",
  34039=>"010111111",
  34040=>"111000100",
  34041=>"111001101",
  34042=>"110111001",
  34043=>"100000100",
  34044=>"101000101",
  34045=>"010011110",
  34046=>"111011010",
  34047=>"010110100",
  34048=>"100010011",
  34049=>"000010101",
  34050=>"100110010",
  34051=>"100010111",
  34052=>"001100011",
  34053=>"010000100",
  34054=>"010011101",
  34055=>"000001100",
  34056=>"101110100",
  34057=>"011011101",
  34058=>"101011001",
  34059=>"111110011",
  34060=>"001111101",
  34061=>"001010100",
  34062=>"111000000",
  34063=>"001000000",
  34064=>"001111100",
  34065=>"011000011",
  34066=>"101111111",
  34067=>"100101001",
  34068=>"111001010",
  34069=>"011000100",
  34070=>"100000101",
  34071=>"000000101",
  34072=>"000010001",
  34073=>"010110000",
  34074=>"011100001",
  34075=>"010000110",
  34076=>"011000000",
  34077=>"100011001",
  34078=>"010001010",
  34079=>"001001100",
  34080=>"010000000",
  34081=>"000011010",
  34082=>"010011010",
  34083=>"101100010",
  34084=>"111100100",
  34085=>"101001110",
  34086=>"110011111",
  34087=>"111001011",
  34088=>"011010011",
  34089=>"010110001",
  34090=>"000010100",
  34091=>"000011000",
  34092=>"000001000",
  34093=>"010011001",
  34094=>"011100111",
  34095=>"111000001",
  34096=>"011000110",
  34097=>"111101111",
  34098=>"111001001",
  34099=>"000111110",
  34100=>"110000100",
  34101=>"011000001",
  34102=>"101110101",
  34103=>"111010000",
  34104=>"000000010",
  34105=>"111010000",
  34106=>"000111011",
  34107=>"000101000",
  34108=>"110110001",
  34109=>"000100110",
  34110=>"110010011",
  34111=>"010101000",
  34112=>"000011001",
  34113=>"100100111",
  34114=>"000000101",
  34115=>"000110010",
  34116=>"001100011",
  34117=>"011101010",
  34118=>"000111010",
  34119=>"000101111",
  34120=>"011011010",
  34121=>"001111011",
  34122=>"010001111",
  34123=>"001010000",
  34124=>"110101000",
  34125=>"001000011",
  34126=>"010101110",
  34127=>"011100001",
  34128=>"011100111",
  34129=>"001100001",
  34130=>"110000001",
  34131=>"111011110",
  34132=>"111110010",
  34133=>"011011001",
  34134=>"000110100",
  34135=>"010011011",
  34136=>"000110011",
  34137=>"000110110",
  34138=>"111000010",
  34139=>"000111101",
  34140=>"100111100",
  34141=>"001001101",
  34142=>"011010101",
  34143=>"001101010",
  34144=>"111000000",
  34145=>"101111111",
  34146=>"101001101",
  34147=>"001001100",
  34148=>"001110000",
  34149=>"100000111",
  34150=>"101000011",
  34151=>"111100111",
  34152=>"110010001",
  34153=>"001010111",
  34154=>"011111001",
  34155=>"000010010",
  34156=>"010100000",
  34157=>"111111001",
  34158=>"110110001",
  34159=>"011111011",
  34160=>"100011010",
  34161=>"110111101",
  34162=>"101110000",
  34163=>"111100101",
  34164=>"000110100",
  34165=>"110011111",
  34166=>"000111110",
  34167=>"100111010",
  34168=>"000111100",
  34169=>"100110000",
  34170=>"010011001",
  34171=>"111111110",
  34172=>"100000101",
  34173=>"100100001",
  34174=>"010001000",
  34175=>"101100010",
  34176=>"000101101",
  34177=>"000111010",
  34178=>"110011000",
  34179=>"110011100",
  34180=>"000001000",
  34181=>"001001111",
  34182=>"001101010",
  34183=>"101101101",
  34184=>"001000111",
  34185=>"010110111",
  34186=>"011111100",
  34187=>"001010001",
  34188=>"101000001",
  34189=>"001000000",
  34190=>"101010110",
  34191=>"111111010",
  34192=>"010011100",
  34193=>"001101000",
  34194=>"000011111",
  34195=>"110110001",
  34196=>"101010011",
  34197=>"000100010",
  34198=>"111111111",
  34199=>"000101110",
  34200=>"101100101",
  34201=>"010001010",
  34202=>"011110011",
  34203=>"100000111",
  34204=>"011110111",
  34205=>"010100000",
  34206=>"001100100",
  34207=>"000101100",
  34208=>"010110000",
  34209=>"101010000",
  34210=>"011011011",
  34211=>"100010011",
  34212=>"100001010",
  34213=>"000100010",
  34214=>"010111010",
  34215=>"001010000",
  34216=>"111011000",
  34217=>"110111001",
  34218=>"101101111",
  34219=>"101100100",
  34220=>"100111111",
  34221=>"100010111",
  34222=>"101001010",
  34223=>"100111011",
  34224=>"011111000",
  34225=>"011010000",
  34226=>"110101000",
  34227=>"000110011",
  34228=>"011011001",
  34229=>"010011000",
  34230=>"110011100",
  34231=>"111010000",
  34232=>"111010111",
  34233=>"000101011",
  34234=>"101001011",
  34235=>"010101000",
  34236=>"100111110",
  34237=>"111011001",
  34238=>"101010101",
  34239=>"010101010",
  34240=>"110111111",
  34241=>"011011110",
  34242=>"101110010",
  34243=>"110010001",
  34244=>"000110111",
  34245=>"001100011",
  34246=>"111010101",
  34247=>"100010010",
  34248=>"001010100",
  34249=>"100100010",
  34250=>"000001000",
  34251=>"000000010",
  34252=>"001100011",
  34253=>"000111100",
  34254=>"010110101",
  34255=>"000011101",
  34256=>"001110101",
  34257=>"010001101",
  34258=>"001101010",
  34259=>"111110101",
  34260=>"011111001",
  34261=>"101101010",
  34262=>"001100011",
  34263=>"011010110",
  34264=>"011011000",
  34265=>"001000010",
  34266=>"101011011",
  34267=>"100010101",
  34268=>"111110101",
  34269=>"101011000",
  34270=>"101010111",
  34271=>"110101101",
  34272=>"010100010",
  34273=>"110001110",
  34274=>"110110001",
  34275=>"100001001",
  34276=>"000101100",
  34277=>"100101010",
  34278=>"011111000",
  34279=>"010100001",
  34280=>"100000000",
  34281=>"000010100",
  34282=>"110110010",
  34283=>"111100110",
  34284=>"100101010",
  34285=>"110101001",
  34286=>"011110111",
  34287=>"011000101",
  34288=>"110101110",
  34289=>"111000000",
  34290=>"010010100",
  34291=>"000011011",
  34292=>"001001110",
  34293=>"111000000",
  34294=>"101100110",
  34295=>"000000000",
  34296=>"100000000",
  34297=>"111010101",
  34298=>"101011100",
  34299=>"101100100",
  34300=>"111010010",
  34301=>"010001110",
  34302=>"000011011",
  34303=>"010010011",
  34304=>"000001100",
  34305=>"111101011",
  34306=>"100101111",
  34307=>"001101011",
  34308=>"110010100",
  34309=>"110000101",
  34310=>"100000111",
  34311=>"011011010",
  34312=>"010110100",
  34313=>"111011011",
  34314=>"111101001",
  34315=>"011001111",
  34316=>"101001100",
  34317=>"010110000",
  34318=>"011110010",
  34319=>"111100000",
  34320=>"010100011",
  34321=>"001001101",
  34322=>"000010000",
  34323=>"010101010",
  34324=>"011111100",
  34325=>"000101100",
  34326=>"111010000",
  34327=>"100111001",
  34328=>"001001101",
  34329=>"010101011",
  34330=>"101010101",
  34331=>"000110101",
  34332=>"000010100",
  34333=>"010100010",
  34334=>"101001100",
  34335=>"111100111",
  34336=>"100001111",
  34337=>"111111110",
  34338=>"010100011",
  34339=>"010010010",
  34340=>"110000101",
  34341=>"111100000",
  34342=>"011010001",
  34343=>"101000101",
  34344=>"101111000",
  34345=>"110000100",
  34346=>"010100001",
  34347=>"111111111",
  34348=>"010101001",
  34349=>"000100101",
  34350=>"010110100",
  34351=>"000010011",
  34352=>"110100110",
  34353=>"000001100",
  34354=>"000001101",
  34355=>"100100110",
  34356=>"011000100",
  34357=>"001100000",
  34358=>"000000000",
  34359=>"100010110",
  34360=>"000110010",
  34361=>"101110010",
  34362=>"101101100",
  34363=>"100101000",
  34364=>"110000001",
  34365=>"010111010",
  34366=>"111001000",
  34367=>"110000010",
  34368=>"001010101",
  34369=>"100100000",
  34370=>"011111010",
  34371=>"010100110",
  34372=>"100111011",
  34373=>"011100111",
  34374=>"110101011",
  34375=>"100101110",
  34376=>"011111001",
  34377=>"011000011",
  34378=>"110111001",
  34379=>"000111111",
  34380=>"001010111",
  34381=>"011110010",
  34382=>"111000010",
  34383=>"101001000",
  34384=>"101010000",
  34385=>"110001001",
  34386=>"011101000",
  34387=>"100011100",
  34388=>"011001110",
  34389=>"111100000",
  34390=>"001001000",
  34391=>"001110110",
  34392=>"111101110",
  34393=>"100101111",
  34394=>"101010000",
  34395=>"100001101",
  34396=>"111100101",
  34397=>"001000111",
  34398=>"100101001",
  34399=>"000010110",
  34400=>"111101010",
  34401=>"010001001",
  34402=>"111111011",
  34403=>"011010001",
  34404=>"010111010",
  34405=>"100100000",
  34406=>"001000010",
  34407=>"101000101",
  34408=>"000101001",
  34409=>"011010010",
  34410=>"110100011",
  34411=>"100010001",
  34412=>"101111111",
  34413=>"100010011",
  34414=>"010100011",
  34415=>"110110101",
  34416=>"001101001",
  34417=>"101000000",
  34418=>"110100101",
  34419=>"010101000",
  34420=>"001101110",
  34421=>"001000011",
  34422=>"010010000",
  34423=>"100000101",
  34424=>"111001011",
  34425=>"110001100",
  34426=>"111011111",
  34427=>"010110100",
  34428=>"001111001",
  34429=>"000100000",
  34430=>"000101001",
  34431=>"011101101",
  34432=>"100010000",
  34433=>"011001010",
  34434=>"011001101",
  34435=>"101000001",
  34436=>"100000110",
  34437=>"100011100",
  34438=>"100011000",
  34439=>"101011100",
  34440=>"110010011",
  34441=>"010101011",
  34442=>"101101011",
  34443=>"000000101",
  34444=>"011100001",
  34445=>"011101100",
  34446=>"101100110",
  34447=>"111110011",
  34448=>"111001001",
  34449=>"111100101",
  34450=>"110010111",
  34451=>"101010001",
  34452=>"000010100",
  34453=>"100000101",
  34454=>"110111000",
  34455=>"100010100",
  34456=>"010010001",
  34457=>"001001010",
  34458=>"011101100",
  34459=>"100100010",
  34460=>"111000011",
  34461=>"101001010",
  34462=>"110000001",
  34463=>"000001000",
  34464=>"011101100",
  34465=>"010010111",
  34466=>"001100100",
  34467=>"111110110",
  34468=>"101010001",
  34469=>"110001010",
  34470=>"000110010",
  34471=>"011110011",
  34472=>"000110010",
  34473=>"011000010",
  34474=>"100110101",
  34475=>"101101100",
  34476=>"010010111",
  34477=>"000111010",
  34478=>"001010111",
  34479=>"000001110",
  34480=>"000111101",
  34481=>"010110110",
  34482=>"100101100",
  34483=>"100100101",
  34484=>"100101101",
  34485=>"001010111",
  34486=>"101001000",
  34487=>"000100010",
  34488=>"011111101",
  34489=>"011110110",
  34490=>"110000011",
  34491=>"101001001",
  34492=>"101100000",
  34493=>"011011111",
  34494=>"010101111",
  34495=>"010110110",
  34496=>"010000100",
  34497=>"010111110",
  34498=>"111001100",
  34499=>"110011011",
  34500=>"110010001",
  34501=>"001010101",
  34502=>"011100001",
  34503=>"011111011",
  34504=>"001001100",
  34505=>"000110010",
  34506=>"011011110",
  34507=>"100001101",
  34508=>"100100010",
  34509=>"010100100",
  34510=>"110000110",
  34511=>"001011111",
  34512=>"111101011",
  34513=>"101001001",
  34514=>"010100001",
  34515=>"101100010",
  34516=>"000001101",
  34517=>"101111111",
  34518=>"011010110",
  34519=>"001000100",
  34520=>"000110110",
  34521=>"111111001",
  34522=>"100100111",
  34523=>"111010010",
  34524=>"101001100",
  34525=>"110101111",
  34526=>"010111111",
  34527=>"100001100",
  34528=>"000100010",
  34529=>"100111000",
  34530=>"100100101",
  34531=>"011100010",
  34532=>"001000011",
  34533=>"010111101",
  34534=>"011001111",
  34535=>"111011111",
  34536=>"011100011",
  34537=>"110100100",
  34538=>"001000000",
  34539=>"001101101",
  34540=>"100110000",
  34541=>"111011000",
  34542=>"101101101",
  34543=>"001010111",
  34544=>"011101011",
  34545=>"011000001",
  34546=>"110010001",
  34547=>"001101111",
  34548=>"000101010",
  34549=>"110001001",
  34550=>"011010010",
  34551=>"010110011",
  34552=>"000011101",
  34553=>"111000100",
  34554=>"111010110",
  34555=>"101011110",
  34556=>"001000100",
  34557=>"001101010",
  34558=>"100100111",
  34559=>"001110111",
  34560=>"100010001",
  34561=>"110000000",
  34562=>"011110000",
  34563=>"110011100",
  34564=>"111100001",
  34565=>"000100101",
  34566=>"010011010",
  34567=>"111011111",
  34568=>"100000101",
  34569=>"101101100",
  34570=>"010101111",
  34571=>"001001000",
  34572=>"100110011",
  34573=>"001000000",
  34574=>"010100011",
  34575=>"101010011",
  34576=>"110000101",
  34577=>"000100100",
  34578=>"001100101",
  34579=>"111110011",
  34580=>"110110101",
  34581=>"001110101",
  34582=>"000010011",
  34583=>"011010000",
  34584=>"100001010",
  34585=>"100011100",
  34586=>"001111110",
  34587=>"110010100",
  34588=>"000011111",
  34589=>"110001100",
  34590=>"011011111",
  34591=>"101001010",
  34592=>"100101001",
  34593=>"100011100",
  34594=>"110110001",
  34595=>"001110110",
  34596=>"101100101",
  34597=>"001111111",
  34598=>"001010101",
  34599=>"111010011",
  34600=>"001010001",
  34601=>"101001000",
  34602=>"001000000",
  34603=>"010111110",
  34604=>"001000101",
  34605=>"100110010",
  34606=>"000110011",
  34607=>"101011111",
  34608=>"100000000",
  34609=>"111000100",
  34610=>"101001000",
  34611=>"011010000",
  34612=>"110100100",
  34613=>"110101101",
  34614=>"011011010",
  34615=>"011110011",
  34616=>"001101000",
  34617=>"001101111",
  34618=>"000110001",
  34619=>"111100100",
  34620=>"001111000",
  34621=>"110000011",
  34622=>"110110000",
  34623=>"101110101",
  34624=>"000100110",
  34625=>"101111100",
  34626=>"111011110",
  34627=>"001000010",
  34628=>"000000010",
  34629=>"110111011",
  34630=>"010010110",
  34631=>"100001010",
  34632=>"110111010",
  34633=>"011111100",
  34634=>"100001100",
  34635=>"110110111",
  34636=>"110011001",
  34637=>"100000101",
  34638=>"001111111",
  34639=>"111011010",
  34640=>"001001001",
  34641=>"110000010",
  34642=>"101011000",
  34643=>"011000111",
  34644=>"111011010",
  34645=>"111010001",
  34646=>"000101111",
  34647=>"110010001",
  34648=>"010000011",
  34649=>"010101100",
  34650=>"010000111",
  34651=>"101100001",
  34652=>"111001011",
  34653=>"100011000",
  34654=>"100100110",
  34655=>"110111101",
  34656=>"100001111",
  34657=>"011100101",
  34658=>"001001111",
  34659=>"011010010",
  34660=>"111111110",
  34661=>"010111101",
  34662=>"011110111",
  34663=>"111110000",
  34664=>"001011011",
  34665=>"101011100",
  34666=>"000010111",
  34667=>"000000000",
  34668=>"011110001",
  34669=>"010100100",
  34670=>"000111010",
  34671=>"111111100",
  34672=>"110100110",
  34673=>"010010111",
  34674=>"001011111",
  34675=>"010001110",
  34676=>"010111001",
  34677=>"111110111",
  34678=>"011010001",
  34679=>"010000101",
  34680=>"011001010",
  34681=>"000010010",
  34682=>"101010111",
  34683=>"101110000",
  34684=>"000011001",
  34685=>"101111011",
  34686=>"000011000",
  34687=>"000101100",
  34688=>"100000000",
  34689=>"001111011",
  34690=>"111000111",
  34691=>"010111000",
  34692=>"000100011",
  34693=>"011111011",
  34694=>"001000101",
  34695=>"000111110",
  34696=>"111101000",
  34697=>"111100001",
  34698=>"010101111",
  34699=>"111101100",
  34700=>"010011001",
  34701=>"111111101",
  34702=>"000101111",
  34703=>"101100111",
  34704=>"000011001",
  34705=>"100000101",
  34706=>"000011010",
  34707=>"110101111",
  34708=>"011011000",
  34709=>"101001111",
  34710=>"011000101",
  34711=>"010101110",
  34712=>"001001100",
  34713=>"111001011",
  34714=>"000011110",
  34715=>"100100001",
  34716=>"001111101",
  34717=>"010110100",
  34718=>"101010100",
  34719=>"100010010",
  34720=>"101110010",
  34721=>"011001100",
  34722=>"010010110",
  34723=>"010000001",
  34724=>"000000100",
  34725=>"111101010",
  34726=>"110111111",
  34727=>"100010111",
  34728=>"110001010",
  34729=>"101000111",
  34730=>"101100000",
  34731=>"110000000",
  34732=>"100000100",
  34733=>"000001011",
  34734=>"000101001",
  34735=>"010110111",
  34736=>"011101101",
  34737=>"011001111",
  34738=>"000000011",
  34739=>"111011001",
  34740=>"111110110",
  34741=>"100100001",
  34742=>"011010001",
  34743=>"101011100",
  34744=>"001000011",
  34745=>"110001100",
  34746=>"100001111",
  34747=>"111110110",
  34748=>"100010010",
  34749=>"000001101",
  34750=>"101010011",
  34751=>"101101111",
  34752=>"011011101",
  34753=>"110101101",
  34754=>"000110001",
  34755=>"000110110",
  34756=>"111100010",
  34757=>"100011101",
  34758=>"011010101",
  34759=>"101000110",
  34760=>"110011010",
  34761=>"001110111",
  34762=>"000010101",
  34763=>"010110111",
  34764=>"001101010",
  34765=>"011111011",
  34766=>"001111000",
  34767=>"010000111",
  34768=>"110110111",
  34769=>"111000001",
  34770=>"001001111",
  34771=>"011110001",
  34772=>"011000111",
  34773=>"101110100",
  34774=>"011010001",
  34775=>"011011101",
  34776=>"011110001",
  34777=>"101010100",
  34778=>"001110010",
  34779=>"000100101",
  34780=>"110001110",
  34781=>"001001000",
  34782=>"010110011",
  34783=>"010101110",
  34784=>"100000111",
  34785=>"110000000",
  34786=>"100111100",
  34787=>"011100111",
  34788=>"111000011",
  34789=>"000110101",
  34790=>"100111000",
  34791=>"010000011",
  34792=>"101111111",
  34793=>"100010001",
  34794=>"000110110",
  34795=>"000000110",
  34796=>"100011000",
  34797=>"000001101",
  34798=>"111001001",
  34799=>"001110001",
  34800=>"001011101",
  34801=>"110001110",
  34802=>"111111000",
  34803=>"110011101",
  34804=>"010011010",
  34805=>"011001100",
  34806=>"011101111",
  34807=>"001011000",
  34808=>"011011000",
  34809=>"000110101",
  34810=>"010101111",
  34811=>"010011001",
  34812=>"110100011",
  34813=>"011111111",
  34814=>"000100010",
  34815=>"010010001",
  34816=>"010101111",
  34817=>"011000101",
  34818=>"111000101",
  34819=>"010100010",
  34820=>"100110010",
  34821=>"101101101",
  34822=>"010001111",
  34823=>"111010011",
  34824=>"011011000",
  34825=>"110000000",
  34826=>"000000011",
  34827=>"000010110",
  34828=>"110010000",
  34829=>"110110111",
  34830=>"100100010",
  34831=>"101101110",
  34832=>"001010101",
  34833=>"101111010",
  34834=>"000101110",
  34835=>"010110000",
  34836=>"111111011",
  34837=>"100001111",
  34838=>"101110000",
  34839=>"111100011",
  34840=>"110111111",
  34841=>"111001110",
  34842=>"001000100",
  34843=>"011010001",
  34844=>"001110010",
  34845=>"010000000",
  34846=>"010111011",
  34847=>"111111100",
  34848=>"110010100",
  34849=>"011010011",
  34850=>"001100111",
  34851=>"000101111",
  34852=>"100101001",
  34853=>"010001101",
  34854=>"110001010",
  34855=>"000011000",
  34856=>"000110011",
  34857=>"100111001",
  34858=>"100111011",
  34859=>"000000101",
  34860=>"000000010",
  34861=>"011011111",
  34862=>"011100000",
  34863=>"110001000",
  34864=>"100111111",
  34865=>"001011111",
  34866=>"111001111",
  34867=>"100100010",
  34868=>"001011110",
  34869=>"011110011",
  34870=>"010011001",
  34871=>"111101001",
  34872=>"000110001",
  34873=>"011010011",
  34874=>"001110110",
  34875=>"101000100",
  34876=>"101011010",
  34877=>"100110010",
  34878=>"000010001",
  34879=>"001100111",
  34880=>"011011111",
  34881=>"011100110",
  34882=>"010001000",
  34883=>"110010101",
  34884=>"100100110",
  34885=>"111101010",
  34886=>"010100110",
  34887=>"100011011",
  34888=>"111101100",
  34889=>"001111000",
  34890=>"111100011",
  34891=>"111100101",
  34892=>"111100010",
  34893=>"000110001",
  34894=>"110110111",
  34895=>"001111101",
  34896=>"001001101",
  34897=>"000001000",
  34898=>"110100000",
  34899=>"001101110",
  34900=>"110011001",
  34901=>"110000000",
  34902=>"111101110",
  34903=>"000001100",
  34904=>"101001101",
  34905=>"010000000",
  34906=>"010011001",
  34907=>"001010110",
  34908=>"110110011",
  34909=>"000110000",
  34910=>"100111100",
  34911=>"010011101",
  34912=>"100011111",
  34913=>"111010110",
  34914=>"010000111",
  34915=>"100101101",
  34916=>"100001101",
  34917=>"011010001",
  34918=>"111001010",
  34919=>"100011111",
  34920=>"111000111",
  34921=>"010001110",
  34922=>"110000110",
  34923=>"000110010",
  34924=>"101111110",
  34925=>"001110101",
  34926=>"001000101",
  34927=>"100000010",
  34928=>"100011110",
  34929=>"010011100",
  34930=>"100001100",
  34931=>"001100100",
  34932=>"010011101",
  34933=>"010010100",
  34934=>"111110111",
  34935=>"000100100",
  34936=>"100100011",
  34937=>"110000000",
  34938=>"000001101",
  34939=>"111010000",
  34940=>"010000010",
  34941=>"001100000",
  34942=>"111011111",
  34943=>"001100001",
  34944=>"001101110",
  34945=>"110110011",
  34946=>"111111111",
  34947=>"010001110",
  34948=>"111111000",
  34949=>"000111011",
  34950=>"011110010",
  34951=>"110000101",
  34952=>"101001101",
  34953=>"000001111",
  34954=>"011100111",
  34955=>"111101011",
  34956=>"011100111",
  34957=>"110011100",
  34958=>"000101111",
  34959=>"001000001",
  34960=>"110110011",
  34961=>"010111110",
  34962=>"000000111",
  34963=>"001011100",
  34964=>"110010001",
  34965=>"111100011",
  34966=>"011011001",
  34967=>"010011100",
  34968=>"001101001",
  34969=>"100011101",
  34970=>"100001011",
  34971=>"000000010",
  34972=>"101111011",
  34973=>"111101100",
  34974=>"111010000",
  34975=>"100101010",
  34976=>"010111010",
  34977=>"000001011",
  34978=>"001111011",
  34979=>"111110100",
  34980=>"001111010",
  34981=>"000111010",
  34982=>"011000100",
  34983=>"010011100",
  34984=>"000000010",
  34985=>"101001110",
  34986=>"011010001",
  34987=>"111010001",
  34988=>"110110101",
  34989=>"011110110",
  34990=>"000101100",
  34991=>"110000001",
  34992=>"101101000",
  34993=>"100101101",
  34994=>"100001100",
  34995=>"010110100",
  34996=>"111101000",
  34997=>"110100000",
  34998=>"000110100",
  34999=>"000100100",
  35000=>"101100101",
  35001=>"111100010",
  35002=>"111101010",
  35003=>"110001100",
  35004=>"010000111",
  35005=>"100000111",
  35006=>"000110011",
  35007=>"011011110",
  35008=>"001100010",
  35009=>"000000100",
  35010=>"011111101",
  35011=>"000011001",
  35012=>"110100000",
  35013=>"001110100",
  35014=>"010110011",
  35015=>"000011010",
  35016=>"111110011",
  35017=>"101101100",
  35018=>"111101100",
  35019=>"100001111",
  35020=>"010100100",
  35021=>"111111111",
  35022=>"011110110",
  35023=>"001010001",
  35024=>"000001000",
  35025=>"110001011",
  35026=>"010101000",
  35027=>"110110001",
  35028=>"100001011",
  35029=>"010100111",
  35030=>"100001001",
  35031=>"100101100",
  35032=>"001111000",
  35033=>"100100011",
  35034=>"111111001",
  35035=>"110111100",
  35036=>"011000000",
  35037=>"011111110",
  35038=>"000101101",
  35039=>"000110100",
  35040=>"001000100",
  35041=>"011110001",
  35042=>"000110101",
  35043=>"001001111",
  35044=>"010100001",
  35045=>"100010001",
  35046=>"110110110",
  35047=>"011001011",
  35048=>"100011011",
  35049=>"000011101",
  35050=>"000100110",
  35051=>"110110110",
  35052=>"011001010",
  35053=>"001100101",
  35054=>"100010001",
  35055=>"110100001",
  35056=>"111000101",
  35057=>"001000000",
  35058=>"011001010",
  35059=>"110010111",
  35060=>"011111000",
  35061=>"011011011",
  35062=>"100010100",
  35063=>"100101110",
  35064=>"001110110",
  35065=>"010010110",
  35066=>"011111110",
  35067=>"011100111",
  35068=>"001011111",
  35069=>"001000000",
  35070=>"101100101",
  35071=>"101100001",
  35072=>"111011101",
  35073=>"110000001",
  35074=>"110110110",
  35075=>"000011101",
  35076=>"000011011",
  35077=>"111001001",
  35078=>"010111111",
  35079=>"111101100",
  35080=>"010000001",
  35081=>"011111001",
  35082=>"000011011",
  35083=>"100000000",
  35084=>"011011111",
  35085=>"110000100",
  35086=>"000101111",
  35087=>"110001110",
  35088=>"010001110",
  35089=>"100011000",
  35090=>"101101101",
  35091=>"000011010",
  35092=>"001001101",
  35093=>"111111100",
  35094=>"110100001",
  35095=>"111011111",
  35096=>"010101110",
  35097=>"101111100",
  35098=>"001000110",
  35099=>"100111111",
  35100=>"111100010",
  35101=>"111000101",
  35102=>"100101110",
  35103=>"110111100",
  35104=>"001101001",
  35105=>"100011111",
  35106=>"011100110",
  35107=>"010100000",
  35108=>"001010011",
  35109=>"010101010",
  35110=>"110101101",
  35111=>"000110010",
  35112=>"000001000",
  35113=>"010001000",
  35114=>"000100001",
  35115=>"001111000",
  35116=>"110111000",
  35117=>"000001000",
  35118=>"100101011",
  35119=>"010010100",
  35120=>"111010101",
  35121=>"101110110",
  35122=>"000000110",
  35123=>"101100001",
  35124=>"110000010",
  35125=>"011101001",
  35126=>"101110011",
  35127=>"100011101",
  35128=>"101101100",
  35129=>"011001111",
  35130=>"101111101",
  35131=>"010000001",
  35132=>"000001001",
  35133=>"001101110",
  35134=>"010000000",
  35135=>"111000111",
  35136=>"010010011",
  35137=>"100011111",
  35138=>"000000110",
  35139=>"000111001",
  35140=>"100011100",
  35141=>"110100010",
  35142=>"010011011",
  35143=>"110000110",
  35144=>"010001000",
  35145=>"001110010",
  35146=>"111011000",
  35147=>"011101010",
  35148=>"010000000",
  35149=>"110000101",
  35150=>"111101101",
  35151=>"000010000",
  35152=>"111000010",
  35153=>"011001111",
  35154=>"000000000",
  35155=>"110101110",
  35156=>"101011011",
  35157=>"110100110",
  35158=>"011000001",
  35159=>"111001011",
  35160=>"110010000",
  35161=>"111011100",
  35162=>"000000000",
  35163=>"000110111",
  35164=>"101011111",
  35165=>"101010110",
  35166=>"111111111",
  35167=>"110011010",
  35168=>"110101111",
  35169=>"100100011",
  35170=>"000111011",
  35171=>"110111110",
  35172=>"101010010",
  35173=>"001101000",
  35174=>"100010000",
  35175=>"001110000",
  35176=>"001100000",
  35177=>"011001110",
  35178=>"011011011",
  35179=>"010000001",
  35180=>"100010101",
  35181=>"001000110",
  35182=>"101111100",
  35183=>"011011010",
  35184=>"010010101",
  35185=>"001111010",
  35186=>"100011011",
  35187=>"101010001",
  35188=>"110100000",
  35189=>"010001100",
  35190=>"000100110",
  35191=>"100110110",
  35192=>"001000111",
  35193=>"101011001",
  35194=>"100111010",
  35195=>"010010001",
  35196=>"001110101",
  35197=>"000000100",
  35198=>"011111001",
  35199=>"001110110",
  35200=>"100011010",
  35201=>"001010011",
  35202=>"010001110",
  35203=>"001010111",
  35204=>"001010000",
  35205=>"001011011",
  35206=>"011111001",
  35207=>"000001110",
  35208=>"111100110",
  35209=>"110011001",
  35210=>"101010011",
  35211=>"001011010",
  35212=>"011011000",
  35213=>"000001011",
  35214=>"110110110",
  35215=>"011000010",
  35216=>"000110001",
  35217=>"000000110",
  35218=>"001110100",
  35219=>"111111011",
  35220=>"111011000",
  35221=>"101100000",
  35222=>"010111110",
  35223=>"101010111",
  35224=>"101111100",
  35225=>"011000100",
  35226=>"111000010",
  35227=>"001010111",
  35228=>"100011111",
  35229=>"001101010",
  35230=>"101110110",
  35231=>"111111111",
  35232=>"111100101",
  35233=>"010000000",
  35234=>"000110111",
  35235=>"001001101",
  35236=>"000111111",
  35237=>"000110010",
  35238=>"001010100",
  35239=>"011000010",
  35240=>"101111001",
  35241=>"001111010",
  35242=>"001101101",
  35243=>"000000000",
  35244=>"011011100",
  35245=>"101000100",
  35246=>"011111110",
  35247=>"011110000",
  35248=>"111010010",
  35249=>"000000010",
  35250=>"111001001",
  35251=>"000101001",
  35252=>"000000101",
  35253=>"111101110",
  35254=>"110100000",
  35255=>"101100010",
  35256=>"101111010",
  35257=>"101001010",
  35258=>"010000001",
  35259=>"000110100",
  35260=>"010010010",
  35261=>"111101011",
  35262=>"011100011",
  35263=>"100011011",
  35264=>"000001000",
  35265=>"000000000",
  35266=>"111101101",
  35267=>"110111101",
  35268=>"101100111",
  35269=>"101000111",
  35270=>"110010100",
  35271=>"000011001",
  35272=>"001111101",
  35273=>"001110111",
  35274=>"110010101",
  35275=>"010011011",
  35276=>"001010100",
  35277=>"100111111",
  35278=>"100111000",
  35279=>"100100010",
  35280=>"101000111",
  35281=>"110100101",
  35282=>"100000011",
  35283=>"100111101",
  35284=>"111110101",
  35285=>"011100000",
  35286=>"010010110",
  35287=>"000010001",
  35288=>"100000010",
  35289=>"010101110",
  35290=>"101011100",
  35291=>"001001011",
  35292=>"111001011",
  35293=>"100011110",
  35294=>"110111101",
  35295=>"110100000",
  35296=>"100101000",
  35297=>"101110010",
  35298=>"100110101",
  35299=>"011111010",
  35300=>"100100111",
  35301=>"110011101",
  35302=>"000100011",
  35303=>"010010111",
  35304=>"100100001",
  35305=>"100100100",
  35306=>"100010001",
  35307=>"010111001",
  35308=>"010010000",
  35309=>"100101111",
  35310=>"001100000",
  35311=>"001110010",
  35312=>"101111101",
  35313=>"100000001",
  35314=>"111110001",
  35315=>"101101011",
  35316=>"011110000",
  35317=>"001010000",
  35318=>"011100000",
  35319=>"110010111",
  35320=>"011001000",
  35321=>"001000001",
  35322=>"100110011",
  35323=>"011010000",
  35324=>"101110111",
  35325=>"010100000",
  35326=>"001000111",
  35327=>"010110010",
  35328=>"111000100",
  35329=>"100101100",
  35330=>"000001011",
  35331=>"000011111",
  35332=>"111001000",
  35333=>"001101100",
  35334=>"101011000",
  35335=>"011111110",
  35336=>"011111001",
  35337=>"010010101",
  35338=>"101011101",
  35339=>"010101110",
  35340=>"011011010",
  35341=>"111100111",
  35342=>"001101000",
  35343=>"011100101",
  35344=>"010010000",
  35345=>"001001000",
  35346=>"010000000",
  35347=>"101001111",
  35348=>"110010111",
  35349=>"100001110",
  35350=>"110001010",
  35351=>"011110110",
  35352=>"111001000",
  35353=>"101101110",
  35354=>"101011100",
  35355=>"000011100",
  35356=>"110110001",
  35357=>"100101100",
  35358=>"110000000",
  35359=>"001011000",
  35360=>"110001101",
  35361=>"110100100",
  35362=>"110010100",
  35363=>"101100011",
  35364=>"111100111",
  35365=>"101100001",
  35366=>"110101111",
  35367=>"101111011",
  35368=>"000101100",
  35369=>"101100100",
  35370=>"011000110",
  35371=>"001000110",
  35372=>"001000010",
  35373=>"010011000",
  35374=>"000010110",
  35375=>"000011000",
  35376=>"001001101",
  35377=>"011011010",
  35378=>"011010101",
  35379=>"010000010",
  35380=>"101010010",
  35381=>"101011011",
  35382=>"000000011",
  35383=>"101111100",
  35384=>"110110111",
  35385=>"110000000",
  35386=>"011101101",
  35387=>"110101100",
  35388=>"101111001",
  35389=>"110010100",
  35390=>"000000001",
  35391=>"111111100",
  35392=>"011111111",
  35393=>"000000011",
  35394=>"000101001",
  35395=>"110000000",
  35396=>"111011011",
  35397=>"011001011",
  35398=>"011110000",
  35399=>"001100000",
  35400=>"000110010",
  35401=>"001101001",
  35402=>"110011001",
  35403=>"010111110",
  35404=>"100100101",
  35405=>"001001011",
  35406=>"110100010",
  35407=>"101000001",
  35408=>"111000101",
  35409=>"111110110",
  35410=>"100101101",
  35411=>"111111011",
  35412=>"110110000",
  35413=>"001100000",
  35414=>"110010111",
  35415=>"011010100",
  35416=>"100001111",
  35417=>"000011011",
  35418=>"111000001",
  35419=>"100101101",
  35420=>"001001000",
  35421=>"010000010",
  35422=>"011001101",
  35423=>"110110100",
  35424=>"101110011",
  35425=>"011001000",
  35426=>"100110110",
  35427=>"000110011",
  35428=>"111100110",
  35429=>"110010110",
  35430=>"111110111",
  35431=>"011011001",
  35432=>"000010001",
  35433=>"000011000",
  35434=>"110000101",
  35435=>"000010100",
  35436=>"101011101",
  35437=>"010000010",
  35438=>"010000101",
  35439=>"011100010",
  35440=>"011000000",
  35441=>"000111101",
  35442=>"010100101",
  35443=>"001010010",
  35444=>"111001011",
  35445=>"111111111",
  35446=>"011110101",
  35447=>"010000000",
  35448=>"010101111",
  35449=>"010011111",
  35450=>"001101110",
  35451=>"111111110",
  35452=>"100001001",
  35453=>"000101101",
  35454=>"010000100",
  35455=>"110011111",
  35456=>"010001100",
  35457=>"101111001",
  35458=>"100100111",
  35459=>"100100001",
  35460=>"100011110",
  35461=>"010100110",
  35462=>"110010010",
  35463=>"111010111",
  35464=>"111000011",
  35465=>"001101001",
  35466=>"001100100",
  35467=>"111110110",
  35468=>"001000110",
  35469=>"111010101",
  35470=>"110110000",
  35471=>"100110111",
  35472=>"100100001",
  35473=>"101111101",
  35474=>"101111100",
  35475=>"011111111",
  35476=>"000100110",
  35477=>"110001100",
  35478=>"111111000",
  35479=>"101001110",
  35480=>"011100100",
  35481=>"100010000",
  35482=>"110010001",
  35483=>"010101011",
  35484=>"010000001",
  35485=>"010000110",
  35486=>"000100000",
  35487=>"100100110",
  35488=>"100101110",
  35489=>"010011001",
  35490=>"010000001",
  35491=>"010011011",
  35492=>"100001010",
  35493=>"000001010",
  35494=>"100010110",
  35495=>"000100000",
  35496=>"110000000",
  35497=>"011001101",
  35498=>"110001101",
  35499=>"101100110",
  35500=>"011100111",
  35501=>"001110001",
  35502=>"110110000",
  35503=>"111001001",
  35504=>"100010100",
  35505=>"010010011",
  35506=>"111111111",
  35507=>"010101000",
  35508=>"001010110",
  35509=>"100010101",
  35510=>"000010000",
  35511=>"110011100",
  35512=>"111001110",
  35513=>"001110011",
  35514=>"101100101",
  35515=>"100011100",
  35516=>"100000111",
  35517=>"100101001",
  35518=>"000000000",
  35519=>"000101001",
  35520=>"011010110",
  35521=>"011011111",
  35522=>"100010100",
  35523=>"011100100",
  35524=>"111001111",
  35525=>"001000000",
  35526=>"110000100",
  35527=>"010000100",
  35528=>"010011101",
  35529=>"001001101",
  35530=>"100010111",
  35531=>"110011000",
  35532=>"101101010",
  35533=>"100000100",
  35534=>"010111111",
  35535=>"101001110",
  35536=>"101110111",
  35537=>"000000001",
  35538=>"001011000",
  35539=>"110010010",
  35540=>"000000010",
  35541=>"101011010",
  35542=>"011111100",
  35543=>"100111001",
  35544=>"111000110",
  35545=>"100010101",
  35546=>"000100101",
  35547=>"010001001",
  35548=>"001110111",
  35549=>"111110100",
  35550=>"101110101",
  35551=>"100010001",
  35552=>"010111001",
  35553=>"011111110",
  35554=>"011101110",
  35555=>"001101101",
  35556=>"011101101",
  35557=>"110010000",
  35558=>"000000101",
  35559=>"110001101",
  35560=>"111000100",
  35561=>"101111111",
  35562=>"111011011",
  35563=>"010111110",
  35564=>"001001010",
  35565=>"100010001",
  35566=>"111111111",
  35567=>"000101001",
  35568=>"110001111",
  35569=>"101100001",
  35570=>"100000111",
  35571=>"001011001",
  35572=>"010111001",
  35573=>"000000001",
  35574=>"101011001",
  35575=>"101000010",
  35576=>"100111101",
  35577=>"010011001",
  35578=>"001110100",
  35579=>"000001011",
  35580=>"011101010",
  35581=>"011111111",
  35582=>"100110011",
  35583=>"001100101",
  35584=>"010110011",
  35585=>"001010011",
  35586=>"001101110",
  35587=>"101111111",
  35588=>"110100110",
  35589=>"100100100",
  35590=>"010010000",
  35591=>"111001101",
  35592=>"111010000",
  35593=>"101111101",
  35594=>"001110010",
  35595=>"101101100",
  35596=>"010010100",
  35597=>"110010110",
  35598=>"011010100",
  35599=>"011001100",
  35600=>"000010100",
  35601=>"100011000",
  35602=>"011100100",
  35603=>"001101111",
  35604=>"000101101",
  35605=>"100110000",
  35606=>"101101000",
  35607=>"011010011",
  35608=>"111000111",
  35609=>"000000100",
  35610=>"100001001",
  35611=>"011100010",
  35612=>"100001101",
  35613=>"001000100",
  35614=>"000111000",
  35615=>"010001101",
  35616=>"000100111",
  35617=>"010001110",
  35618=>"101101011",
  35619=>"110110111",
  35620=>"001100011",
  35621=>"000101100",
  35622=>"010001011",
  35623=>"011110011",
  35624=>"111000101",
  35625=>"000100110",
  35626=>"101011110",
  35627=>"011111011",
  35628=>"011101110",
  35629=>"000000011",
  35630=>"111111110",
  35631=>"011111110",
  35632=>"111001010",
  35633=>"001001001",
  35634=>"010001101",
  35635=>"010010010",
  35636=>"000011001",
  35637=>"100000010",
  35638=>"000000110",
  35639=>"100001110",
  35640=>"010001010",
  35641=>"110100011",
  35642=>"111010001",
  35643=>"110011100",
  35644=>"000100101",
  35645=>"001011000",
  35646=>"011100010",
  35647=>"110010111",
  35648=>"010011001",
  35649=>"101000000",
  35650=>"000001111",
  35651=>"001110010",
  35652=>"101001110",
  35653=>"111001110",
  35654=>"101000101",
  35655=>"001010101",
  35656=>"111110010",
  35657=>"001101111",
  35658=>"100110000",
  35659=>"010101011",
  35660=>"100100010",
  35661=>"101010001",
  35662=>"110111100",
  35663=>"110100101",
  35664=>"011101111",
  35665=>"110111101",
  35666=>"000000000",
  35667=>"111101011",
  35668=>"000011110",
  35669=>"110010011",
  35670=>"111011110",
  35671=>"001101011",
  35672=>"001010000",
  35673=>"110000000",
  35674=>"011001000",
  35675=>"001100000",
  35676=>"110110010",
  35677=>"000100010",
  35678=>"010010011",
  35679=>"000101000",
  35680=>"000010101",
  35681=>"100110010",
  35682=>"000100101",
  35683=>"111000111",
  35684=>"011100011",
  35685=>"101011010",
  35686=>"001001011",
  35687=>"011111000",
  35688=>"110010010",
  35689=>"111000001",
  35690=>"111101010",
  35691=>"011000000",
  35692=>"011011001",
  35693=>"100010110",
  35694=>"000011111",
  35695=>"001011000",
  35696=>"010101000",
  35697=>"111111101",
  35698=>"101011101",
  35699=>"001100000",
  35700=>"111010110",
  35701=>"000000111",
  35702=>"011101111",
  35703=>"010110110",
  35704=>"111111010",
  35705=>"011001001",
  35706=>"011001010",
  35707=>"111100000",
  35708=>"100101010",
  35709=>"000001101",
  35710=>"011100001",
  35711=>"000011100",
  35712=>"100110011",
  35713=>"100111100",
  35714=>"010010100",
  35715=>"010110111",
  35716=>"010111100",
  35717=>"100010001",
  35718=>"010010101",
  35719=>"100101010",
  35720=>"111010101",
  35721=>"110101110",
  35722=>"101101110",
  35723=>"000111111",
  35724=>"000100100",
  35725=>"101000110",
  35726=>"111110100",
  35727=>"110101111",
  35728=>"110001101",
  35729=>"001111111",
  35730=>"010000100",
  35731=>"000101001",
  35732=>"100100010",
  35733=>"001010000",
  35734=>"010101001",
  35735=>"010100001",
  35736=>"010000101",
  35737=>"000000100",
  35738=>"100001100",
  35739=>"100111010",
  35740=>"010010000",
  35741=>"000111001",
  35742=>"110010001",
  35743=>"011010110",
  35744=>"110101011",
  35745=>"101100100",
  35746=>"000010101",
  35747=>"110010110",
  35748=>"010000100",
  35749=>"010011111",
  35750=>"101001111",
  35751=>"100110011",
  35752=>"011111111",
  35753=>"000110100",
  35754=>"100111110",
  35755=>"110001001",
  35756=>"101011111",
  35757=>"000010000",
  35758=>"111111010",
  35759=>"010111110",
  35760=>"111001101",
  35761=>"111101100",
  35762=>"001111000",
  35763=>"100111001",
  35764=>"110111000",
  35765=>"110111111",
  35766=>"101111010",
  35767=>"111101110",
  35768=>"000001100",
  35769=>"110100010",
  35770=>"011010101",
  35771=>"110101110",
  35772=>"110101001",
  35773=>"011010000",
  35774=>"000010000",
  35775=>"011010101",
  35776=>"111101111",
  35777=>"001011100",
  35778=>"111010001",
  35779=>"110011011",
  35780=>"011100100",
  35781=>"010111111",
  35782=>"101100111",
  35783=>"011011111",
  35784=>"100110000",
  35785=>"100011001",
  35786=>"010001001",
  35787=>"101101100",
  35788=>"010100010",
  35789=>"110010001",
  35790=>"100111111",
  35791=>"101000001",
  35792=>"000000100",
  35793=>"000100110",
  35794=>"011100101",
  35795=>"110000100",
  35796=>"000010111",
  35797=>"000010001",
  35798=>"001001111",
  35799=>"110010101",
  35800=>"010011100",
  35801=>"101111001",
  35802=>"100001111",
  35803=>"011000000",
  35804=>"110011110",
  35805=>"000001111",
  35806=>"110010011",
  35807=>"011011111",
  35808=>"011001000",
  35809=>"011010010",
  35810=>"001101100",
  35811=>"010000100",
  35812=>"000100101",
  35813=>"011001111",
  35814=>"011001101",
  35815=>"110111011",
  35816=>"100001010",
  35817=>"110001101",
  35818=>"000011110",
  35819=>"000011111",
  35820=>"010100001",
  35821=>"000000010",
  35822=>"000110111",
  35823=>"000010111",
  35824=>"000110011",
  35825=>"111110111",
  35826=>"011010110",
  35827=>"101001100",
  35828=>"111101111",
  35829=>"110000000",
  35830=>"001000111",
  35831=>"100011101",
  35832=>"011001011",
  35833=>"111110101",
  35834=>"110011010",
  35835=>"010100110",
  35836=>"011000100",
  35837=>"110000110",
  35838=>"001100001",
  35839=>"010111111",
  35840=>"010011100",
  35841=>"000011111",
  35842=>"000110101",
  35843=>"010011100",
  35844=>"010111111",
  35845=>"010011111",
  35846=>"101010000",
  35847=>"111000110",
  35848=>"110001110",
  35849=>"100000100",
  35850=>"110111010",
  35851=>"101111101",
  35852=>"111101001",
  35853=>"000110101",
  35854=>"111101101",
  35855=>"001011111",
  35856=>"110100011",
  35857=>"000000110",
  35858=>"110010000",
  35859=>"111011111",
  35860=>"110100001",
  35861=>"000110101",
  35862=>"001101011",
  35863=>"110101111",
  35864=>"001110001",
  35865=>"001110111",
  35866=>"111010001",
  35867=>"110111010",
  35868=>"111000011",
  35869=>"110100010",
  35870=>"011110000",
  35871=>"110010110",
  35872=>"100101010",
  35873=>"110101000",
  35874=>"001101100",
  35875=>"110110110",
  35876=>"111001001",
  35877=>"011110010",
  35878=>"100000000",
  35879=>"001101000",
  35880=>"011111101",
  35881=>"010011110",
  35882=>"101101100",
  35883=>"111010111",
  35884=>"000000001",
  35885=>"001011110",
  35886=>"010001100",
  35887=>"011000000",
  35888=>"111011011",
  35889=>"010011000",
  35890=>"000000111",
  35891=>"000011000",
  35892=>"000000111",
  35893=>"100100001",
  35894=>"000000010",
  35895=>"100011010",
  35896=>"101001011",
  35897=>"110101000",
  35898=>"101000100",
  35899=>"001010100",
  35900=>"110101110",
  35901=>"010011011",
  35902=>"001001011",
  35903=>"101000001",
  35904=>"000000101",
  35905=>"111100011",
  35906=>"100111001",
  35907=>"110010100",
  35908=>"101111101",
  35909=>"100000110",
  35910=>"000101011",
  35911=>"010101000",
  35912=>"100011101",
  35913=>"010010111",
  35914=>"111100100",
  35915=>"001111001",
  35916=>"100001011",
  35917=>"111101011",
  35918=>"110010110",
  35919=>"111101100",
  35920=>"110111011",
  35921=>"101010110",
  35922=>"111000101",
  35923=>"100011011",
  35924=>"111101010",
  35925=>"101100001",
  35926=>"000100100",
  35927=>"101100101",
  35928=>"110101101",
  35929=>"110100010",
  35930=>"110001110",
  35931=>"010101010",
  35932=>"100000100",
  35933=>"101010111",
  35934=>"110110010",
  35935=>"110100111",
  35936=>"001001111",
  35937=>"001010000",
  35938=>"101101010",
  35939=>"010011100",
  35940=>"011001100",
  35941=>"011011011",
  35942=>"111001000",
  35943=>"000010101",
  35944=>"000000111",
  35945=>"110110010",
  35946=>"000101010",
  35947=>"100011101",
  35948=>"100110101",
  35949=>"000011011",
  35950=>"100011100",
  35951=>"111001000",
  35952=>"000001111",
  35953=>"001101001",
  35954=>"101101000",
  35955=>"110001111",
  35956=>"000001101",
  35957=>"100011010",
  35958=>"110000111",
  35959=>"000010000",
  35960=>"001011100",
  35961=>"001001110",
  35962=>"111110101",
  35963=>"010110011",
  35964=>"100001110",
  35965=>"101100110",
  35966=>"110111100",
  35967=>"001110010",
  35968=>"111110110",
  35969=>"101101100",
  35970=>"101101101",
  35971=>"101001010",
  35972=>"011100011",
  35973=>"111000100",
  35974=>"110001011",
  35975=>"110101111",
  35976=>"000110101",
  35977=>"111100011",
  35978=>"111000101",
  35979=>"000000110",
  35980=>"000100101",
  35981=>"101110011",
  35982=>"100010110",
  35983=>"010110010",
  35984=>"100000110",
  35985=>"100111101",
  35986=>"110100001",
  35987=>"010010101",
  35988=>"011001000",
  35989=>"111010100",
  35990=>"000101010",
  35991=>"111010111",
  35992=>"001101000",
  35993=>"101000001",
  35994=>"111010000",
  35995=>"000000000",
  35996=>"111000101",
  35997=>"111111000",
  35998=>"100100111",
  35999=>"111110011",
  36000=>"100001001",
  36001=>"101011000",
  36002=>"101100111",
  36003=>"110001010",
  36004=>"010111010",
  36005=>"100100111",
  36006=>"101101100",
  36007=>"110000011",
  36008=>"011111110",
  36009=>"101100010",
  36010=>"001000001",
  36011=>"110010000",
  36012=>"011010000",
  36013=>"011010101",
  36014=>"000011001",
  36015=>"111111101",
  36016=>"001101111",
  36017=>"111111001",
  36018=>"100101101",
  36019=>"000100111",
  36020=>"000100110",
  36021=>"110011110",
  36022=>"011001001",
  36023=>"000011001",
  36024=>"101010110",
  36025=>"101011101",
  36026=>"000110001",
  36027=>"100100010",
  36028=>"110011010",
  36029=>"101101001",
  36030=>"000000011",
  36031=>"110110011",
  36032=>"000001110",
  36033=>"000001000",
  36034=>"111100010",
  36035=>"000100000",
  36036=>"110000011",
  36037=>"000001010",
  36038=>"110001011",
  36039=>"101101001",
  36040=>"011111000",
  36041=>"100100100",
  36042=>"010000110",
  36043=>"010001001",
  36044=>"101000010",
  36045=>"001110100",
  36046=>"111101101",
  36047=>"101100010",
  36048=>"111100000",
  36049=>"000111011",
  36050=>"010111101",
  36051=>"111000101",
  36052=>"010100110",
  36053=>"100001100",
  36054=>"001011100",
  36055=>"000001111",
  36056=>"010110100",
  36057=>"011101001",
  36058=>"001001110",
  36059=>"000010101",
  36060=>"111111000",
  36061=>"110001011",
  36062=>"001010001",
  36063=>"111011000",
  36064=>"001001101",
  36065=>"000011011",
  36066=>"001100101",
  36067=>"110100000",
  36068=>"101110011",
  36069=>"101000100",
  36070=>"011000010",
  36071=>"001101010",
  36072=>"000011001",
  36073=>"101001101",
  36074=>"001111100",
  36075=>"110000111",
  36076=>"000000101",
  36077=>"101110010",
  36078=>"001011000",
  36079=>"010000000",
  36080=>"001111100",
  36081=>"001000111",
  36082=>"100011001",
  36083=>"101011111",
  36084=>"111111101",
  36085=>"111110110",
  36086=>"010000000",
  36087=>"001110010",
  36088=>"100101110",
  36089=>"101111100",
  36090=>"000001001",
  36091=>"000001101",
  36092=>"111101111",
  36093=>"111110011",
  36094=>"011101011",
  36095=>"110100000",
  36096=>"010101100",
  36097=>"100000011",
  36098=>"101110110",
  36099=>"110000110",
  36100=>"101011001",
  36101=>"011001111",
  36102=>"100000010",
  36103=>"110000100",
  36104=>"111100010",
  36105=>"000001000",
  36106=>"110001010",
  36107=>"100010111",
  36108=>"110100001",
  36109=>"000001100",
  36110=>"010001101",
  36111=>"000010110",
  36112=>"111001101",
  36113=>"010100011",
  36114=>"100000010",
  36115=>"010101100",
  36116=>"010000100",
  36117=>"101000101",
  36118=>"111000011",
  36119=>"000011100",
  36120=>"100001011",
  36121=>"101101001",
  36122=>"111110001",
  36123=>"100101001",
  36124=>"110101111",
  36125=>"000100101",
  36126=>"101100100",
  36127=>"100000110",
  36128=>"000010101",
  36129=>"011000010",
  36130=>"110100011",
  36131=>"000010001",
  36132=>"110001010",
  36133=>"000111101",
  36134=>"000101001",
  36135=>"111001111",
  36136=>"111101110",
  36137=>"111001011",
  36138=>"000000111",
  36139=>"100010011",
  36140=>"011110010",
  36141=>"100110010",
  36142=>"110000110",
  36143=>"000101010",
  36144=>"110101110",
  36145=>"000110111",
  36146=>"100000000",
  36147=>"101000011",
  36148=>"111111000",
  36149=>"010110101",
  36150=>"000001001",
  36151=>"111100011",
  36152=>"100000011",
  36153=>"110110100",
  36154=>"111110000",
  36155=>"001010000",
  36156=>"001010001",
  36157=>"100010001",
  36158=>"010110010",
  36159=>"100000100",
  36160=>"111101001",
  36161=>"001000010",
  36162=>"110110011",
  36163=>"000101011",
  36164=>"111001011",
  36165=>"100010011",
  36166=>"111000010",
  36167=>"010110101",
  36168=>"000000000",
  36169=>"000011100",
  36170=>"001001000",
  36171=>"000001001",
  36172=>"110000010",
  36173=>"011011011",
  36174=>"101001101",
  36175=>"110101100",
  36176=>"011110101",
  36177=>"100011000",
  36178=>"100110110",
  36179=>"111111001",
  36180=>"001101011",
  36181=>"000000110",
  36182=>"111000010",
  36183=>"100001000",
  36184=>"000110000",
  36185=>"010010011",
  36186=>"110011101",
  36187=>"100101100",
  36188=>"101011000",
  36189=>"111110010",
  36190=>"100001111",
  36191=>"010100010",
  36192=>"000100011",
  36193=>"011000100",
  36194=>"100001100",
  36195=>"010010110",
  36196=>"110100011",
  36197=>"111000011",
  36198=>"000111111",
  36199=>"001100111",
  36200=>"001111011",
  36201=>"101100111",
  36202=>"110101111",
  36203=>"110110010",
  36204=>"101111000",
  36205=>"100000110",
  36206=>"000001011",
  36207=>"110011100",
  36208=>"111001011",
  36209=>"001111101",
  36210=>"101100010",
  36211=>"101100101",
  36212=>"111100010",
  36213=>"110101100",
  36214=>"001010110",
  36215=>"011001111",
  36216=>"011011010",
  36217=>"000001110",
  36218=>"110011001",
  36219=>"111110101",
  36220=>"000010111",
  36221=>"010101011",
  36222=>"111101001",
  36223=>"011010001",
  36224=>"111010011",
  36225=>"001100101",
  36226=>"011100100",
  36227=>"000001101",
  36228=>"111010101",
  36229=>"101101101",
  36230=>"101100010",
  36231=>"001110011",
  36232=>"010010101",
  36233=>"010010011",
  36234=>"010111110",
  36235=>"101110111",
  36236=>"011100100",
  36237=>"011101101",
  36238=>"110111100",
  36239=>"101001001",
  36240=>"100000100",
  36241=>"110100101",
  36242=>"010000001",
  36243=>"010110011",
  36244=>"001010101",
  36245=>"011100101",
  36246=>"010011010",
  36247=>"000111100",
  36248=>"100100110",
  36249=>"011000010",
  36250=>"000100101",
  36251=>"000000100",
  36252=>"110000101",
  36253=>"010010011",
  36254=>"111100111",
  36255=>"001001100",
  36256=>"110011101",
  36257=>"011000100",
  36258=>"001100111",
  36259=>"001011101",
  36260=>"100101000",
  36261=>"000100100",
  36262=>"011100111",
  36263=>"110110111",
  36264=>"010011101",
  36265=>"000000000",
  36266=>"101010110",
  36267=>"001101110",
  36268=>"000001110",
  36269=>"101001111",
  36270=>"010100001",
  36271=>"001111000",
  36272=>"100010101",
  36273=>"101110001",
  36274=>"110001010",
  36275=>"111011001",
  36276=>"101100011",
  36277=>"010010100",
  36278=>"000100100",
  36279=>"011101101",
  36280=>"110100111",
  36281=>"101001001",
  36282=>"110111010",
  36283=>"100000110",
  36284=>"111101110",
  36285=>"110111100",
  36286=>"110101011",
  36287=>"101100101",
  36288=>"010000111",
  36289=>"011100101",
  36290=>"011001100",
  36291=>"010100111",
  36292=>"100000101",
  36293=>"000100001",
  36294=>"001001111",
  36295=>"110011100",
  36296=>"111101110",
  36297=>"001001000",
  36298=>"100011110",
  36299=>"011111000",
  36300=>"110000101",
  36301=>"110100110",
  36302=>"100011000",
  36303=>"000000000",
  36304=>"101010011",
  36305=>"110111100",
  36306=>"001111000",
  36307=>"001101001",
  36308=>"110110011",
  36309=>"101010101",
  36310=>"101110000",
  36311=>"110011100",
  36312=>"000100110",
  36313=>"001011011",
  36314=>"100010000",
  36315=>"011100110",
  36316=>"011010110",
  36317=>"010001000",
  36318=>"000000000",
  36319=>"011010010",
  36320=>"101111100",
  36321=>"000111000",
  36322=>"100010001",
  36323=>"011110010",
  36324=>"000011111",
  36325=>"000101010",
  36326=>"011010011",
  36327=>"010111100",
  36328=>"110000100",
  36329=>"011010100",
  36330=>"001110010",
  36331=>"100000110",
  36332=>"111111101",
  36333=>"101000100",
  36334=>"001100111",
  36335=>"001000110",
  36336=>"110100111",
  36337=>"111000111",
  36338=>"010010001",
  36339=>"011110001",
  36340=>"110001011",
  36341=>"011100100",
  36342=>"111001110",
  36343=>"110000110",
  36344=>"111001011",
  36345=>"110011111",
  36346=>"010000011",
  36347=>"101110100",
  36348=>"000001011",
  36349=>"101110001",
  36350=>"000011110",
  36351=>"101000111",
  36352=>"010111000",
  36353=>"011110010",
  36354=>"101010111",
  36355=>"000110000",
  36356=>"101010000",
  36357=>"111111111",
  36358=>"110011110",
  36359=>"010001010",
  36360=>"101010001",
  36361=>"100011001",
  36362=>"000100011",
  36363=>"010000010",
  36364=>"001111011",
  36365=>"000110001",
  36366=>"010110011",
  36367=>"100101000",
  36368=>"011110111",
  36369=>"000111000",
  36370=>"010100001",
  36371=>"110111110",
  36372=>"110010101",
  36373=>"110111011",
  36374=>"110111101",
  36375=>"001100111",
  36376=>"000110111",
  36377=>"101010001",
  36378=>"010010111",
  36379=>"100101001",
  36380=>"000010110",
  36381=>"010010000",
  36382=>"111011001",
  36383=>"011111101",
  36384=>"011010111",
  36385=>"101001100",
  36386=>"111010110",
  36387=>"110110110",
  36388=>"010110101",
  36389=>"100111111",
  36390=>"110101010",
  36391=>"010011010",
  36392=>"011001001",
  36393=>"001010011",
  36394=>"111101100",
  36395=>"111000101",
  36396=>"100110010",
  36397=>"100010000",
  36398=>"101000100",
  36399=>"101110001",
  36400=>"110100001",
  36401=>"010100001",
  36402=>"101011110",
  36403=>"111010111",
  36404=>"011000010",
  36405=>"111011111",
  36406=>"101101110",
  36407=>"011101001",
  36408=>"110000101",
  36409=>"100101000",
  36410=>"000001010",
  36411=>"111111011",
  36412=>"010010101",
  36413=>"110110100",
  36414=>"101101010",
  36415=>"010001010",
  36416=>"001011011",
  36417=>"011110010",
  36418=>"010011100",
  36419=>"101011001",
  36420=>"101010001",
  36421=>"010000010",
  36422=>"010001100",
  36423=>"100101000",
  36424=>"101000110",
  36425=>"000000010",
  36426=>"010001001",
  36427=>"000111010",
  36428=>"000101011",
  36429=>"011010110",
  36430=>"111001011",
  36431=>"010000111",
  36432=>"001000111",
  36433=>"000010000",
  36434=>"010010000",
  36435=>"110010101",
  36436=>"010101011",
  36437=>"101010010",
  36438=>"100110100",
  36439=>"000100100",
  36440=>"110001011",
  36441=>"100111010",
  36442=>"111111100",
  36443=>"100001010",
  36444=>"011110110",
  36445=>"011100110",
  36446=>"010110011",
  36447=>"101011100",
  36448=>"001011110",
  36449=>"000011000",
  36450=>"011010111",
  36451=>"011110011",
  36452=>"011011011",
  36453=>"010111000",
  36454=>"011001110",
  36455=>"000001111",
  36456=>"000000001",
  36457=>"100010010",
  36458=>"110110111",
  36459=>"110000000",
  36460=>"111100101",
  36461=>"101100110",
  36462=>"000111011",
  36463=>"000100010",
  36464=>"110001101",
  36465=>"000101001",
  36466=>"101100100",
  36467=>"010100011",
  36468=>"011001010",
  36469=>"010010111",
  36470=>"110001000",
  36471=>"100111000",
  36472=>"010010010",
  36473=>"011011000",
  36474=>"010111101",
  36475=>"100111111",
  36476=>"101110110",
  36477=>"000100111",
  36478=>"101111000",
  36479=>"010010110",
  36480=>"001010000",
  36481=>"101111111",
  36482=>"111001000",
  36483=>"001001110",
  36484=>"011101011",
  36485=>"000000010",
  36486=>"110010001",
  36487=>"011001110",
  36488=>"100101110",
  36489=>"111000000",
  36490=>"111111001",
  36491=>"001001101",
  36492=>"001000011",
  36493=>"001010000",
  36494=>"001001011",
  36495=>"111111000",
  36496=>"001111000",
  36497=>"101010111",
  36498=>"001001101",
  36499=>"000011000",
  36500=>"010011011",
  36501=>"011010101",
  36502=>"111010001",
  36503=>"100100011",
  36504=>"101000000",
  36505=>"100011000",
  36506=>"011011110",
  36507=>"110110111",
  36508=>"100011001",
  36509=>"000110011",
  36510=>"010001110",
  36511=>"000100000",
  36512=>"010010001",
  36513=>"001000000",
  36514=>"010111001",
  36515=>"110101000",
  36516=>"111111110",
  36517=>"100000101",
  36518=>"001000001",
  36519=>"001110011",
  36520=>"101011111",
  36521=>"100110010",
  36522=>"000000110",
  36523=>"010110111",
  36524=>"011001010",
  36525=>"100110011",
  36526=>"100010110",
  36527=>"100001010",
  36528=>"110000101",
  36529=>"111000111",
  36530=>"001011100",
  36531=>"001101110",
  36532=>"101110001",
  36533=>"000010101",
  36534=>"110100100",
  36535=>"011111100",
  36536=>"101010101",
  36537=>"101111111",
  36538=>"100011110",
  36539=>"001100011",
  36540=>"100000011",
  36541=>"010011010",
  36542=>"000101001",
  36543=>"100011000",
  36544=>"000010110",
  36545=>"011110001",
  36546=>"111010110",
  36547=>"010100001",
  36548=>"101110001",
  36549=>"000010001",
  36550=>"011010100",
  36551=>"111000111",
  36552=>"111100010",
  36553=>"110100110",
  36554=>"101010000",
  36555=>"110011010",
  36556=>"100110010",
  36557=>"001000111",
  36558=>"011101101",
  36559=>"100011111",
  36560=>"110110100",
  36561=>"101101101",
  36562=>"010011111",
  36563=>"010101011",
  36564=>"010110111",
  36565=>"001101101",
  36566=>"101010110",
  36567=>"000000011",
  36568=>"100101000",
  36569=>"101011100",
  36570=>"111000010",
  36571=>"001010001",
  36572=>"010000010",
  36573=>"000000100",
  36574=>"000010010",
  36575=>"101111110",
  36576=>"001000001",
  36577=>"001010010",
  36578=>"101010011",
  36579=>"001001011",
  36580=>"110001001",
  36581=>"111111001",
  36582=>"100001111",
  36583=>"000000101",
  36584=>"111111110",
  36585=>"000111000",
  36586=>"110100010",
  36587=>"001001101",
  36588=>"001110010",
  36589=>"100110100",
  36590=>"011111110",
  36591=>"011000000",
  36592=>"000001001",
  36593=>"101110100",
  36594=>"000110011",
  36595=>"011100001",
  36596=>"111000011",
  36597=>"110110010",
  36598=>"100101111",
  36599=>"110111100",
  36600=>"000011011",
  36601=>"110100100",
  36602=>"110110000",
  36603=>"010000000",
  36604=>"111001000",
  36605=>"000110010",
  36606=>"011111111",
  36607=>"100111100",
  36608=>"100110010",
  36609=>"011100010",
  36610=>"101100100",
  36611=>"100111000",
  36612=>"011001111",
  36613=>"001001010",
  36614=>"110101100",
  36615=>"001100111",
  36616=>"010111001",
  36617=>"011100010",
  36618=>"111111110",
  36619=>"111000110",
  36620=>"001010010",
  36621=>"111100111",
  36622=>"000000111",
  36623=>"000111011",
  36624=>"000010110",
  36625=>"100100001",
  36626=>"100010000",
  36627=>"101010111",
  36628=>"010010101",
  36629=>"110000000",
  36630=>"110011110",
  36631=>"010011100",
  36632=>"010110100",
  36633=>"011001111",
  36634=>"000011110",
  36635=>"011110110",
  36636=>"111010000",
  36637=>"001110011",
  36638=>"001010110",
  36639=>"011111100",
  36640=>"111101100",
  36641=>"110100000",
  36642=>"111001011",
  36643=>"001000111",
  36644=>"101100010",
  36645=>"101101101",
  36646=>"101111111",
  36647=>"001010010",
  36648=>"110000100",
  36649=>"000110100",
  36650=>"101110010",
  36651=>"110101100",
  36652=>"011001100",
  36653=>"011001010",
  36654=>"011100101",
  36655=>"000000111",
  36656=>"001000100",
  36657=>"011101100",
  36658=>"110011111",
  36659=>"000001100",
  36660=>"011100101",
  36661=>"001001100",
  36662=>"001010010",
  36663=>"110110101",
  36664=>"011100110",
  36665=>"001010000",
  36666=>"101101001",
  36667=>"011110000",
  36668=>"000100010",
  36669=>"101111101",
  36670=>"000011001",
  36671=>"110101111",
  36672=>"001001010",
  36673=>"100111101",
  36674=>"100111010",
  36675=>"110111001",
  36676=>"001100011",
  36677=>"010110100",
  36678=>"111000000",
  36679=>"010111010",
  36680=>"010011011",
  36681=>"000101000",
  36682=>"110111011",
  36683=>"010001001",
  36684=>"000111001",
  36685=>"110001000",
  36686=>"001000011",
  36687=>"011100010",
  36688=>"110110101",
  36689=>"001110011",
  36690=>"110001111",
  36691=>"101111001",
  36692=>"001100100",
  36693=>"111001001",
  36694=>"001001111",
  36695=>"100100101",
  36696=>"001010111",
  36697=>"101100101",
  36698=>"101001110",
  36699=>"011101101",
  36700=>"100101011",
  36701=>"101011001",
  36702=>"111111111",
  36703=>"000100011",
  36704=>"100000110",
  36705=>"110111001",
  36706=>"010101101",
  36707=>"000111100",
  36708=>"110101111",
  36709=>"101101000",
  36710=>"100001101",
  36711=>"111110001",
  36712=>"001000010",
  36713=>"011110111",
  36714=>"111000101",
  36715=>"001000100",
  36716=>"010010011",
  36717=>"001000101",
  36718=>"100110011",
  36719=>"110011101",
  36720=>"010101101",
  36721=>"000111110",
  36722=>"000001011",
  36723=>"100001100",
  36724=>"000000110",
  36725=>"010000000",
  36726=>"010111000",
  36727=>"111101001",
  36728=>"111001011",
  36729=>"110000101",
  36730=>"101101101",
  36731=>"010001010",
  36732=>"110110001",
  36733=>"000010010",
  36734=>"101100100",
  36735=>"010100001",
  36736=>"110011110",
  36737=>"111110011",
  36738=>"000111010",
  36739=>"000001111",
  36740=>"100000010",
  36741=>"011101101",
  36742=>"000100011",
  36743=>"000110001",
  36744=>"100000100",
  36745=>"101111100",
  36746=>"011111011",
  36747=>"111110111",
  36748=>"011111000",
  36749=>"101001001",
  36750=>"100110101",
  36751=>"101001011",
  36752=>"010110111",
  36753=>"011111001",
  36754=>"010000010",
  36755=>"001111010",
  36756=>"001010110",
  36757=>"111001010",
  36758=>"010111111",
  36759=>"000111010",
  36760=>"100111010",
  36761=>"000010100",
  36762=>"010000110",
  36763=>"011010001",
  36764=>"011010001",
  36765=>"001100000",
  36766=>"111011000",
  36767=>"001010000",
  36768=>"001111110",
  36769=>"111000010",
  36770=>"110001101",
  36771=>"010111010",
  36772=>"000011001",
  36773=>"100101011",
  36774=>"010110001",
  36775=>"111011001",
  36776=>"101000110",
  36777=>"010000110",
  36778=>"101110000",
  36779=>"001100110",
  36780=>"000110100",
  36781=>"100000110",
  36782=>"000001011",
  36783=>"100111010",
  36784=>"011001001",
  36785=>"111101010",
  36786=>"100011110",
  36787=>"011011001",
  36788=>"101101001",
  36789=>"001111100",
  36790=>"011101110",
  36791=>"010111100",
  36792=>"010000110",
  36793=>"100000011",
  36794=>"100100001",
  36795=>"000000110",
  36796=>"110001111",
  36797=>"111000101",
  36798=>"100110011",
  36799=>"000100100",
  36800=>"001000110",
  36801=>"100111111",
  36802=>"110100111",
  36803=>"111000010",
  36804=>"011111011",
  36805=>"110110110",
  36806=>"010111010",
  36807=>"011100010",
  36808=>"010010011",
  36809=>"010110101",
  36810=>"111001111",
  36811=>"101011011",
  36812=>"000111001",
  36813=>"011000111",
  36814=>"001000111",
  36815=>"111011111",
  36816=>"110111010",
  36817=>"011110100",
  36818=>"001111100",
  36819=>"111010101",
  36820=>"110010110",
  36821=>"110010000",
  36822=>"100110100",
  36823=>"010100010",
  36824=>"001000101",
  36825=>"010000100",
  36826=>"000110011",
  36827=>"000011000",
  36828=>"001000000",
  36829=>"100000101",
  36830=>"100101111",
  36831=>"110100000",
  36832=>"011001010",
  36833=>"100100111",
  36834=>"110000110",
  36835=>"100010101",
  36836=>"000000000",
  36837=>"000101010",
  36838=>"001100101",
  36839=>"111000110",
  36840=>"010011001",
  36841=>"010011000",
  36842=>"000110100",
  36843=>"000111110",
  36844=>"101110010",
  36845=>"010001101",
  36846=>"100000000",
  36847=>"000111110",
  36848=>"111111110",
  36849=>"000100101",
  36850=>"000110000",
  36851=>"111100001",
  36852=>"010001111",
  36853=>"010001011",
  36854=>"011001001",
  36855=>"010100010",
  36856=>"001011011",
  36857=>"001111111",
  36858=>"010001011",
  36859=>"101111111",
  36860=>"010011110",
  36861=>"001001010",
  36862=>"110100011",
  36863=>"011110010",
  36864=>"111010011",
  36865=>"001001010",
  36866=>"100101001",
  36867=>"111010110",
  36868=>"011010010",
  36869=>"000011001",
  36870=>"100001000",
  36871=>"000001011",
  36872=>"000000110",
  36873=>"111111100",
  36874=>"000101111",
  36875=>"111000010",
  36876=>"110110011",
  36877=>"000100101",
  36878=>"011000001",
  36879=>"010111111",
  36880=>"100100111",
  36881=>"011001110",
  36882=>"000010100",
  36883=>"000110001",
  36884=>"001000011",
  36885=>"101110111",
  36886=>"111011011",
  36887=>"110101011",
  36888=>"010011111",
  36889=>"000000001",
  36890=>"001110001",
  36891=>"000100100",
  36892=>"111000111",
  36893=>"110110010",
  36894=>"001100000",
  36895=>"001111100",
  36896=>"111000100",
  36897=>"001100100",
  36898=>"011000011",
  36899=>"000101010",
  36900=>"110010001",
  36901=>"000100110",
  36902=>"010000011",
  36903=>"000001100",
  36904=>"111111000",
  36905=>"010100111",
  36906=>"001111111",
  36907=>"100011100",
  36908=>"101101100",
  36909=>"111010101",
  36910=>"011000001",
  36911=>"101000100",
  36912=>"110100111",
  36913=>"011111111",
  36914=>"101000011",
  36915=>"101100101",
  36916=>"111100011",
  36917=>"100001010",
  36918=>"111010000",
  36919=>"100000010",
  36920=>"100001100",
  36921=>"111111010",
  36922=>"110101011",
  36923=>"110001010",
  36924=>"011101000",
  36925=>"010000110",
  36926=>"000101000",
  36927=>"010001010",
  36928=>"100001010",
  36929=>"001110001",
  36930=>"000010100",
  36931=>"100000000",
  36932=>"001010010",
  36933=>"111001110",
  36934=>"100001001",
  36935=>"111110100",
  36936=>"111001010",
  36937=>"101110010",
  36938=>"100111101",
  36939=>"100001110",
  36940=>"111101001",
  36941=>"100001010",
  36942=>"011010010",
  36943=>"010100000",
  36944=>"011110010",
  36945=>"100011010",
  36946=>"000101100",
  36947=>"111011010",
  36948=>"001000101",
  36949=>"100010001",
  36950=>"001011101",
  36951=>"000100101",
  36952=>"111011000",
  36953=>"101101110",
  36954=>"011100111",
  36955=>"110001110",
  36956=>"101101010",
  36957=>"100100011",
  36958=>"000100010",
  36959=>"000010110",
  36960=>"100000111",
  36961=>"110010010",
  36962=>"100000010",
  36963=>"101101101",
  36964=>"000100001",
  36965=>"011100100",
  36966=>"010101001",
  36967=>"011001111",
  36968=>"000011010",
  36969=>"011110111",
  36970=>"011001001",
  36971=>"111000101",
  36972=>"011110110",
  36973=>"001111111",
  36974=>"011101011",
  36975=>"000111011",
  36976=>"010010010",
  36977=>"001001100",
  36978=>"011000000",
  36979=>"110101010",
  36980=>"100011011",
  36981=>"111101101",
  36982=>"000010100",
  36983=>"000000000",
  36984=>"010111100",
  36985=>"001100011",
  36986=>"000101100",
  36987=>"011111100",
  36988=>"010101000",
  36989=>"111110111",
  36990=>"000111110",
  36991=>"110011100",
  36992=>"010011000",
  36993=>"000011011",
  36994=>"100001000",
  36995=>"010110100",
  36996=>"101100101",
  36997=>"000101111",
  36998=>"001111110",
  36999=>"010000011",
  37000=>"010001111",
  37001=>"011100111",
  37002=>"010000110",
  37003=>"110111100",
  37004=>"011010111",
  37005=>"011111011",
  37006=>"000100110",
  37007=>"100101001",
  37008=>"011111111",
  37009=>"010010000",
  37010=>"110111011",
  37011=>"000001101",
  37012=>"001101100",
  37013=>"011110101",
  37014=>"011010111",
  37015=>"110010010",
  37016=>"011010100",
  37017=>"001010110",
  37018=>"001111111",
  37019=>"111000000",
  37020=>"101100000",
  37021=>"100110110",
  37022=>"110010111",
  37023=>"110011000",
  37024=>"010111110",
  37025=>"011000001",
  37026=>"110010111",
  37027=>"000100111",
  37028=>"110110000",
  37029=>"010000101",
  37030=>"001111011",
  37031=>"111100010",
  37032=>"000010100",
  37033=>"111011110",
  37034=>"101011001",
  37035=>"111101010",
  37036=>"001010110",
  37037=>"111101111",
  37038=>"000010111",
  37039=>"111001110",
  37040=>"110101100",
  37041=>"100110111",
  37042=>"000100000",
  37043=>"010011111",
  37044=>"000100111",
  37045=>"100100000",
  37046=>"110010001",
  37047=>"010000011",
  37048=>"110001100",
  37049=>"001010000",
  37050=>"111111101",
  37051=>"011000101",
  37052=>"101101011",
  37053=>"100001101",
  37054=>"110111011",
  37055=>"010000101",
  37056=>"110000111",
  37057=>"110000000",
  37058=>"000001000",
  37059=>"100110100",
  37060=>"100001111",
  37061=>"000000000",
  37062=>"110001111",
  37063=>"100010000",
  37064=>"111111010",
  37065=>"001101100",
  37066=>"111010010",
  37067=>"100001000",
  37068=>"001011101",
  37069=>"100111111",
  37070=>"111011011",
  37071=>"010110001",
  37072=>"110110101",
  37073=>"100100001",
  37074=>"001100000",
  37075=>"000000011",
  37076=>"011011111",
  37077=>"100101100",
  37078=>"100011110",
  37079=>"100111010",
  37080=>"000011011",
  37081=>"111100001",
  37082=>"010010101",
  37083=>"110010100",
  37084=>"000100101",
  37085=>"010110001",
  37086=>"010010010",
  37087=>"000000111",
  37088=>"000100101",
  37089=>"100110001",
  37090=>"010101100",
  37091=>"001100011",
  37092=>"111011010",
  37093=>"011000100",
  37094=>"110000110",
  37095=>"001110100",
  37096=>"011101000",
  37097=>"100010010",
  37098=>"110010110",
  37099=>"100010110",
  37100=>"101011001",
  37101=>"000101001",
  37102=>"010111111",
  37103=>"110110011",
  37104=>"100011101",
  37105=>"001001111",
  37106=>"001011000",
  37107=>"000000011",
  37108=>"100101101",
  37109=>"101101000",
  37110=>"111000111",
  37111=>"110111111",
  37112=>"100001101",
  37113=>"110010010",
  37114=>"100000011",
  37115=>"001010000",
  37116=>"001010101",
  37117=>"101011001",
  37118=>"101111001",
  37119=>"001010111",
  37120=>"101110010",
  37121=>"000011100",
  37122=>"101100111",
  37123=>"111010001",
  37124=>"000001111",
  37125=>"001110001",
  37126=>"000100001",
  37127=>"101010001",
  37128=>"010110111",
  37129=>"110111011",
  37130=>"000001111",
  37131=>"010110100",
  37132=>"101100110",
  37133=>"110111101",
  37134=>"100101101",
  37135=>"110010110",
  37136=>"001001010",
  37137=>"011110101",
  37138=>"101001001",
  37139=>"110111100",
  37140=>"111110110",
  37141=>"111001010",
  37142=>"000110010",
  37143=>"100110110",
  37144=>"001100001",
  37145=>"001011111",
  37146=>"100100000",
  37147=>"000111100",
  37148=>"110111110",
  37149=>"101010111",
  37150=>"010000010",
  37151=>"000100100",
  37152=>"011000010",
  37153=>"000001010",
  37154=>"000010001",
  37155=>"010001010",
  37156=>"100011011",
  37157=>"101010000",
  37158=>"101111101",
  37159=>"110000000",
  37160=>"110011010",
  37161=>"111100101",
  37162=>"001110011",
  37163=>"100111100",
  37164=>"001101110",
  37165=>"111011000",
  37166=>"110000100",
  37167=>"110100100",
  37168=>"110101011",
  37169=>"100011100",
  37170=>"000011010",
  37171=>"110011010",
  37172=>"100000010",
  37173=>"101101011",
  37174=>"000011011",
  37175=>"001111111",
  37176=>"010011010",
  37177=>"001111010",
  37178=>"000011100",
  37179=>"100100111",
  37180=>"010110011",
  37181=>"101010111",
  37182=>"110110100",
  37183=>"011101010",
  37184=>"110111000",
  37185=>"100100101",
  37186=>"001100101",
  37187=>"001101000",
  37188=>"101111110",
  37189=>"110010010",
  37190=>"100001101",
  37191=>"001011001",
  37192=>"000000000",
  37193=>"111001000",
  37194=>"001101111",
  37195=>"100101100",
  37196=>"111000100",
  37197=>"111001110",
  37198=>"011000010",
  37199=>"011110111",
  37200=>"101001001",
  37201=>"111100101",
  37202=>"100010101",
  37203=>"110001011",
  37204=>"110111011",
  37205=>"110110011",
  37206=>"111011100",
  37207=>"100110101",
  37208=>"000010010",
  37209=>"100110011",
  37210=>"001000011",
  37211=>"000010100",
  37212=>"110000011",
  37213=>"001110010",
  37214=>"100110110",
  37215=>"001000111",
  37216=>"101110001",
  37217=>"110000010",
  37218=>"101000010",
  37219=>"001001110",
  37220=>"101111000",
  37221=>"100101010",
  37222=>"011100100",
  37223=>"100000010",
  37224=>"000011011",
  37225=>"001011011",
  37226=>"000110111",
  37227=>"001001000",
  37228=>"100100010",
  37229=>"111101111",
  37230=>"001011011",
  37231=>"000101111",
  37232=>"001000110",
  37233=>"101011101",
  37234=>"101111111",
  37235=>"001010111",
  37236=>"111000011",
  37237=>"111110011",
  37238=>"010011100",
  37239=>"010010111",
  37240=>"111110001",
  37241=>"111111111",
  37242=>"011100001",
  37243=>"011110000",
  37244=>"011000011",
  37245=>"011100010",
  37246=>"111010101",
  37247=>"010101011",
  37248=>"101110110",
  37249=>"000101001",
  37250=>"000010110",
  37251=>"010011000",
  37252=>"101100111",
  37253=>"100111000",
  37254=>"010000101",
  37255=>"111100111",
  37256=>"110101101",
  37257=>"001001011",
  37258=>"001011111",
  37259=>"000100011",
  37260=>"011101001",
  37261=>"011001001",
  37262=>"110101001",
  37263=>"010010010",
  37264=>"111101001",
  37265=>"001011100",
  37266=>"000110000",
  37267=>"001001001",
  37268=>"101010001",
  37269=>"110001111",
  37270=>"101111000",
  37271=>"000111101",
  37272=>"111110110",
  37273=>"101111101",
  37274=>"110101111",
  37275=>"010001100",
  37276=>"010100001",
  37277=>"100011011",
  37278=>"011110001",
  37279=>"011111100",
  37280=>"110110110",
  37281=>"101100000",
  37282=>"100101111",
  37283=>"000000111",
  37284=>"011111001",
  37285=>"111110100",
  37286=>"011000100",
  37287=>"100110011",
  37288=>"111101000",
  37289=>"010101010",
  37290=>"100011101",
  37291=>"100000011",
  37292=>"111111010",
  37293=>"001001100",
  37294=>"111101110",
  37295=>"000110110",
  37296=>"000000000",
  37297=>"110110001",
  37298=>"000000010",
  37299=>"100000010",
  37300=>"111001100",
  37301=>"101011111",
  37302=>"000111100",
  37303=>"001100000",
  37304=>"110011100",
  37305=>"010101011",
  37306=>"011011001",
  37307=>"110111011",
  37308=>"011111011",
  37309=>"100000111",
  37310=>"110111110",
  37311=>"110000110",
  37312=>"010100011",
  37313=>"010000110",
  37314=>"110000000",
  37315=>"111011010",
  37316=>"110101011",
  37317=>"101111111",
  37318=>"000010000",
  37319=>"101001010",
  37320=>"111100101",
  37321=>"001000101",
  37322=>"111110011",
  37323=>"010010101",
  37324=>"101100100",
  37325=>"101110100",
  37326=>"011111000",
  37327=>"111010010",
  37328=>"011001100",
  37329=>"101000000",
  37330=>"110100001",
  37331=>"001100111",
  37332=>"011010010",
  37333=>"001000000",
  37334=>"111000001",
  37335=>"001100110",
  37336=>"010100011",
  37337=>"100010001",
  37338=>"110010010",
  37339=>"110110101",
  37340=>"010101010",
  37341=>"011100101",
  37342=>"101000111",
  37343=>"100011100",
  37344=>"001111001",
  37345=>"100111001",
  37346=>"010010101",
  37347=>"110001100",
  37348=>"111000010",
  37349=>"000110000",
  37350=>"010110011",
  37351=>"101000001",
  37352=>"011111100",
  37353=>"011010101",
  37354=>"000101101",
  37355=>"110101011",
  37356=>"110111101",
  37357=>"001011101",
  37358=>"010000001",
  37359=>"000101001",
  37360=>"000010011",
  37361=>"100111111",
  37362=>"001000000",
  37363=>"011010001",
  37364=>"111110111",
  37365=>"111100001",
  37366=>"010110011",
  37367=>"000000111",
  37368=>"110110000",
  37369=>"010000111",
  37370=>"001001110",
  37371=>"111111101",
  37372=>"010000101",
  37373=>"111101010",
  37374=>"000001011",
  37375=>"011101010",
  37376=>"011100001",
  37377=>"000011100",
  37378=>"101000001",
  37379=>"001011110",
  37380=>"000101011",
  37381=>"011110011",
  37382=>"001101110",
  37383=>"000010111",
  37384=>"101110101",
  37385=>"001101100",
  37386=>"110100010",
  37387=>"110100011",
  37388=>"100100111",
  37389=>"101011010",
  37390=>"111110101",
  37391=>"010011010",
  37392=>"111001001",
  37393=>"100101110",
  37394=>"111001101",
  37395=>"000001100",
  37396=>"100001101",
  37397=>"011001011",
  37398=>"001111011",
  37399=>"111110010",
  37400=>"010001110",
  37401=>"010001000",
  37402=>"101001000",
  37403=>"000111100",
  37404=>"101010001",
  37405=>"100010100",
  37406=>"111110110",
  37407=>"110110110",
  37408=>"100100100",
  37409=>"001110110",
  37410=>"001000000",
  37411=>"111110111",
  37412=>"001110000",
  37413=>"111101100",
  37414=>"010011001",
  37415=>"001010011",
  37416=>"000011010",
  37417=>"101010010",
  37418=>"011111110",
  37419=>"110100100",
  37420=>"011110011",
  37421=>"001001001",
  37422=>"110111001",
  37423=>"100110011",
  37424=>"111001110",
  37425=>"010110011",
  37426=>"000101100",
  37427=>"100101010",
  37428=>"000000001",
  37429=>"111000111",
  37430=>"011111000",
  37431=>"111011010",
  37432=>"111101001",
  37433=>"000110111",
  37434=>"111100110",
  37435=>"111101100",
  37436=>"001011110",
  37437=>"101111110",
  37438=>"101110111",
  37439=>"101110011",
  37440=>"001100000",
  37441=>"101100100",
  37442=>"000000010",
  37443=>"101000110",
  37444=>"101100110",
  37445=>"011000100",
  37446=>"011000011",
  37447=>"001110010",
  37448=>"000110100",
  37449=>"011111111",
  37450=>"110100010",
  37451=>"111100011",
  37452=>"011101010",
  37453=>"101011101",
  37454=>"110110110",
  37455=>"110111101",
  37456=>"011000001",
  37457=>"010010111",
  37458=>"100001111",
  37459=>"000011100",
  37460=>"010011011",
  37461=>"100001001",
  37462=>"001000001",
  37463=>"000001000",
  37464=>"010001011",
  37465=>"101100011",
  37466=>"000000010",
  37467=>"001010001",
  37468=>"000000100",
  37469=>"001010001",
  37470=>"000011001",
  37471=>"111010101",
  37472=>"111101111",
  37473=>"001110000",
  37474=>"000111111",
  37475=>"101101001",
  37476=>"011111110",
  37477=>"101101100",
  37478=>"100111101",
  37479=>"000010101",
  37480=>"000110101",
  37481=>"001000010",
  37482=>"000101010",
  37483=>"111110011",
  37484=>"000010010",
  37485=>"000000101",
  37486=>"010011000",
  37487=>"010010000",
  37488=>"100000011",
  37489=>"011010010",
  37490=>"011001000",
  37491=>"110001010",
  37492=>"110001001",
  37493=>"110111000",
  37494=>"010010111",
  37495=>"000111000",
  37496=>"000011011",
  37497=>"011000110",
  37498=>"111101111",
  37499=>"001010110",
  37500=>"111001101",
  37501=>"000001011",
  37502=>"001011100",
  37503=>"001011110",
  37504=>"011001011",
  37505=>"111101101",
  37506=>"100110110",
  37507=>"110001110",
  37508=>"001011100",
  37509=>"110011110",
  37510=>"100100111",
  37511=>"100100111",
  37512=>"001101011",
  37513=>"100010110",
  37514=>"101011010",
  37515=>"101111111",
  37516=>"000111111",
  37517=>"010110010",
  37518=>"101110111",
  37519=>"000001101",
  37520=>"100000011",
  37521=>"101111111",
  37522=>"110110011",
  37523=>"011101000",
  37524=>"010010000",
  37525=>"001100100",
  37526=>"000111110",
  37527=>"011100001",
  37528=>"010101011",
  37529=>"110011010",
  37530=>"100100000",
  37531=>"111111111",
  37532=>"101100100",
  37533=>"101000011",
  37534=>"100011001",
  37535=>"000101111",
  37536=>"110000000",
  37537=>"010001011",
  37538=>"101000100",
  37539=>"010011000",
  37540=>"100000111",
  37541=>"011110100",
  37542=>"000110010",
  37543=>"100110001",
  37544=>"110101100",
  37545=>"101100001",
  37546=>"000000110",
  37547=>"100110000",
  37548=>"111001000",
  37549=>"011100010",
  37550=>"110011000",
  37551=>"111101010",
  37552=>"010110011",
  37553=>"000000101",
  37554=>"010011100",
  37555=>"110111001",
  37556=>"000111011",
  37557=>"010111011",
  37558=>"111001001",
  37559=>"100111010",
  37560=>"010000000",
  37561=>"101101100",
  37562=>"100001010",
  37563=>"110010011",
  37564=>"101110110",
  37565=>"011000111",
  37566=>"000110011",
  37567=>"001000100",
  37568=>"010101000",
  37569=>"001101101",
  37570=>"111101000",
  37571=>"101100111",
  37572=>"010000011",
  37573=>"101011001",
  37574=>"101010111",
  37575=>"000110111",
  37576=>"111000010",
  37577=>"011110110",
  37578=>"101001100",
  37579=>"110011000",
  37580=>"101001000",
  37581=>"111111111",
  37582=>"111101111",
  37583=>"110010111",
  37584=>"000000101",
  37585=>"001111111",
  37586=>"000010000",
  37587=>"110010110",
  37588=>"011011111",
  37589=>"000100000",
  37590=>"110010000",
  37591=>"010100000",
  37592=>"001011000",
  37593=>"111011110",
  37594=>"110000001",
  37595=>"000010100",
  37596=>"001100100",
  37597=>"011111010",
  37598=>"010001001",
  37599=>"101111011",
  37600=>"011101010",
  37601=>"010001000",
  37602=>"010101111",
  37603=>"010100110",
  37604=>"000100010",
  37605=>"111110011",
  37606=>"100000111",
  37607=>"000010100",
  37608=>"000111100",
  37609=>"001101101",
  37610=>"101000111",
  37611=>"000110101",
  37612=>"000000110",
  37613=>"011011000",
  37614=>"011100110",
  37615=>"100100101",
  37616=>"100011100",
  37617=>"101100101",
  37618=>"000010111",
  37619=>"010101000",
  37620=>"111111010",
  37621=>"010110101",
  37622=>"010011001",
  37623=>"010110111",
  37624=>"001110000",
  37625=>"100010110",
  37626=>"000001001",
  37627=>"011000011",
  37628=>"000110000",
  37629=>"011110110",
  37630=>"001010100",
  37631=>"000111100",
  37632=>"001000011",
  37633=>"001100001",
  37634=>"101001000",
  37635=>"111000100",
  37636=>"110111111",
  37637=>"001010110",
  37638=>"000000011",
  37639=>"000101101",
  37640=>"111001011",
  37641=>"000000101",
  37642=>"010111110",
  37643=>"111101111",
  37644=>"010111101",
  37645=>"001100100",
  37646=>"100010011",
  37647=>"100110100",
  37648=>"010111100",
  37649=>"010100110",
  37650=>"010110111",
  37651=>"110111001",
  37652=>"111000011",
  37653=>"010110100",
  37654=>"001010011",
  37655=>"011011111",
  37656=>"100011101",
  37657=>"001101001",
  37658=>"000100110",
  37659=>"000000011",
  37660=>"010010100",
  37661=>"111110011",
  37662=>"000111110",
  37663=>"001011010",
  37664=>"011110100",
  37665=>"111110110",
  37666=>"111110110",
  37667=>"111110101",
  37668=>"010001001",
  37669=>"110111111",
  37670=>"110100111",
  37671=>"001101010",
  37672=>"111101110",
  37673=>"101101100",
  37674=>"010111111",
  37675=>"100000010",
  37676=>"100101100",
  37677=>"000100000",
  37678=>"100110010",
  37679=>"001110011",
  37680=>"100100010",
  37681=>"011111100",
  37682=>"000110010",
  37683=>"111100100",
  37684=>"001011000",
  37685=>"111010000",
  37686=>"001101000",
  37687=>"000111101",
  37688=>"001111001",
  37689=>"111000010",
  37690=>"111101011",
  37691=>"000101011",
  37692=>"111000100",
  37693=>"001101000",
  37694=>"011110000",
  37695=>"110101101",
  37696=>"100010001",
  37697=>"011010001",
  37698=>"000100010",
  37699=>"101100110",
  37700=>"011100101",
  37701=>"101010010",
  37702=>"010111110",
  37703=>"101111001",
  37704=>"011110110",
  37705=>"101111011",
  37706=>"100111010",
  37707=>"001101100",
  37708=>"011010011",
  37709=>"010100101",
  37710=>"010110011",
  37711=>"000010001",
  37712=>"000011011",
  37713=>"101010110",
  37714=>"000101000",
  37715=>"001110011",
  37716=>"000111001",
  37717=>"010101101",
  37718=>"001100101",
  37719=>"101111000",
  37720=>"111111011",
  37721=>"101110010",
  37722=>"101100111",
  37723=>"110111111",
  37724=>"010010011",
  37725=>"111111001",
  37726=>"001011011",
  37727=>"100010111",
  37728=>"111111000",
  37729=>"010001100",
  37730=>"001000011",
  37731=>"001100010",
  37732=>"001000010",
  37733=>"001100100",
  37734=>"100100000",
  37735=>"110010001",
  37736=>"100000000",
  37737=>"010011000",
  37738=>"111011010",
  37739=>"111000111",
  37740=>"101001001",
  37741=>"011111000",
  37742=>"001101111",
  37743=>"000101001",
  37744=>"011111100",
  37745=>"010001001",
  37746=>"110101111",
  37747=>"100001011",
  37748=>"000011101",
  37749=>"010010010",
  37750=>"011110010",
  37751=>"000100010",
  37752=>"100111111",
  37753=>"101000001",
  37754=>"000001101",
  37755=>"010001001",
  37756=>"100100001",
  37757=>"001100010",
  37758=>"101100011",
  37759=>"010010011",
  37760=>"101001001",
  37761=>"010111001",
  37762=>"011000000",
  37763=>"000100111",
  37764=>"111011001",
  37765=>"000000000",
  37766=>"101011001",
  37767=>"100010001",
  37768=>"100101010",
  37769=>"110111110",
  37770=>"100101011",
  37771=>"011010010",
  37772=>"011101001",
  37773=>"101011001",
  37774=>"010010111",
  37775=>"111000100",
  37776=>"001001001",
  37777=>"001110010",
  37778=>"001001101",
  37779=>"111000101",
  37780=>"111110111",
  37781=>"110101100",
  37782=>"010111010",
  37783=>"011110111",
  37784=>"101001011",
  37785=>"010100111",
  37786=>"001110010",
  37787=>"000010000",
  37788=>"111101010",
  37789=>"001011000",
  37790=>"110000010",
  37791=>"000100110",
  37792=>"101100111",
  37793=>"100101101",
  37794=>"000011111",
  37795=>"111111100",
  37796=>"100110011",
  37797=>"000001001",
  37798=>"110111111",
  37799=>"110000100",
  37800=>"011010001",
  37801=>"110010011",
  37802=>"000100001",
  37803=>"110111010",
  37804=>"101011101",
  37805=>"110110010",
  37806=>"010001001",
  37807=>"101111101",
  37808=>"110111000",
  37809=>"011011110",
  37810=>"000010110",
  37811=>"100100111",
  37812=>"011100100",
  37813=>"010100101",
  37814=>"000100110",
  37815=>"000110110",
  37816=>"011111111",
  37817=>"010111000",
  37818=>"101111011",
  37819=>"010010010",
  37820=>"100001000",
  37821=>"010111110",
  37822=>"011110100",
  37823=>"001110101",
  37824=>"110000101",
  37825=>"110100110",
  37826=>"100010011",
  37827=>"010000000",
  37828=>"111111101",
  37829=>"010011101",
  37830=>"100101100",
  37831=>"111101010",
  37832=>"110100100",
  37833=>"110001100",
  37834=>"101001111",
  37835=>"001101010",
  37836=>"010111100",
  37837=>"011110111",
  37838=>"010000101",
  37839=>"100111110",
  37840=>"100010100",
  37841=>"110001100",
  37842=>"001111111",
  37843=>"100000001",
  37844=>"101101111",
  37845=>"100001100",
  37846=>"100011001",
  37847=>"000000001",
  37848=>"100111101",
  37849=>"000110101",
  37850=>"111000001",
  37851=>"101001011",
  37852=>"001110101",
  37853=>"000101110",
  37854=>"010101010",
  37855=>"001010001",
  37856=>"001001000",
  37857=>"001001100",
  37858=>"110111110",
  37859=>"001010011",
  37860=>"010000001",
  37861=>"101001011",
  37862=>"000001100",
  37863=>"101001011",
  37864=>"110010001",
  37865=>"111110010",
  37866=>"100101110",
  37867=>"111001000",
  37868=>"100111010",
  37869=>"000011111",
  37870=>"001010001",
  37871=>"111010100",
  37872=>"100010010",
  37873=>"111100110",
  37874=>"110100100",
  37875=>"010111010",
  37876=>"010100010",
  37877=>"000100010",
  37878=>"110111011",
  37879=>"010101110",
  37880=>"100111111",
  37881=>"111010011",
  37882=>"110011000",
  37883=>"011011110",
  37884=>"010001111",
  37885=>"101101010",
  37886=>"000000101",
  37887=>"011000001",
  37888=>"111101111",
  37889=>"001000101",
  37890=>"010010111",
  37891=>"010011000",
  37892=>"100100110",
  37893=>"100010001",
  37894=>"001001111",
  37895=>"100101100",
  37896=>"010010100",
  37897=>"001111101",
  37898=>"011111100",
  37899=>"000110111",
  37900=>"001101111",
  37901=>"001000110",
  37902=>"010010101",
  37903=>"101100011",
  37904=>"011111100",
  37905=>"011001111",
  37906=>"001100010",
  37907=>"111100010",
  37908=>"111110100",
  37909=>"001000111",
  37910=>"000000010",
  37911=>"001001100",
  37912=>"001111011",
  37913=>"111011110",
  37914=>"110010100",
  37915=>"101100001",
  37916=>"111000001",
  37917=>"110011011",
  37918=>"010100010",
  37919=>"101111001",
  37920=>"000100000",
  37921=>"101110101",
  37922=>"110001111",
  37923=>"011010110",
  37924=>"101110110",
  37925=>"000101000",
  37926=>"001111101",
  37927=>"111011000",
  37928=>"101100011",
  37929=>"100110101",
  37930=>"011011100",
  37931=>"000110010",
  37932=>"111101000",
  37933=>"111001111",
  37934=>"101101011",
  37935=>"100000101",
  37936=>"101111000",
  37937=>"000101101",
  37938=>"011001111",
  37939=>"110010000",
  37940=>"001000001",
  37941=>"000001000",
  37942=>"010001111",
  37943=>"011101010",
  37944=>"011010000",
  37945=>"100001000",
  37946=>"011101111",
  37947=>"111100001",
  37948=>"001000111",
  37949=>"100101100",
  37950=>"011011000",
  37951=>"011000010",
  37952=>"110100111",
  37953=>"001001010",
  37954=>"011010101",
  37955=>"000110111",
  37956=>"001110000",
  37957=>"001111010",
  37958=>"111110111",
  37959=>"000000010",
  37960=>"000111100",
  37961=>"010110001",
  37962=>"010000101",
  37963=>"001001100",
  37964=>"111100110",
  37965=>"100100011",
  37966=>"111001110",
  37967=>"001111011",
  37968=>"111111100",
  37969=>"001111101",
  37970=>"010111011",
  37971=>"010011110",
  37972=>"000101001",
  37973=>"111110100",
  37974=>"001101011",
  37975=>"100011101",
  37976=>"111110100",
  37977=>"101011000",
  37978=>"011110101",
  37979=>"010000100",
  37980=>"011101010",
  37981=>"001000010",
  37982=>"010100001",
  37983=>"101100001",
  37984=>"001111111",
  37985=>"111101011",
  37986=>"001011011",
  37987=>"100111011",
  37988=>"011010110",
  37989=>"110001011",
  37990=>"010100000",
  37991=>"001110010",
  37992=>"011001110",
  37993=>"011110111",
  37994=>"111110000",
  37995=>"011000000",
  37996=>"000000100",
  37997=>"011111111",
  37998=>"010010001",
  37999=>"111100001",
  38000=>"001001000",
  38001=>"100011101",
  38002=>"100001011",
  38003=>"100001110",
  38004=>"101001110",
  38005=>"111001000",
  38006=>"110110011",
  38007=>"111111010",
  38008=>"010011101",
  38009=>"101101110",
  38010=>"011100000",
  38011=>"001000010",
  38012=>"010010100",
  38013=>"000000101",
  38014=>"101100111",
  38015=>"100000011",
  38016=>"100011010",
  38017=>"000111111",
  38018=>"101000000",
  38019=>"100001100",
  38020=>"100110010",
  38021=>"001101000",
  38022=>"110101011",
  38023=>"111000000",
  38024=>"101100010",
  38025=>"000011110",
  38026=>"110011010",
  38027=>"010100001",
  38028=>"000010100",
  38029=>"111101110",
  38030=>"101101110",
  38031=>"000111110",
  38032=>"111001011",
  38033=>"010001000",
  38034=>"011000011",
  38035=>"110000010",
  38036=>"110100110",
  38037=>"100100000",
  38038=>"001001101",
  38039=>"100000010",
  38040=>"100111011",
  38041=>"110001100",
  38042=>"010011111",
  38043=>"100001101",
  38044=>"010000000",
  38045=>"011101100",
  38046=>"100001101",
  38047=>"101000101",
  38048=>"111011000",
  38049=>"101001111",
  38050=>"000110000",
  38051=>"111111000",
  38052=>"100101110",
  38053=>"001000101",
  38054=>"110000101",
  38055=>"111011100",
  38056=>"001111000",
  38057=>"011010011",
  38058=>"101001110",
  38059=>"101111110",
  38060=>"000110011",
  38061=>"010111101",
  38062=>"010110010",
  38063=>"101010001",
  38064=>"101001101",
  38065=>"011001000",
  38066=>"010010011",
  38067=>"001101000",
  38068=>"010000000",
  38069=>"101001000",
  38070=>"100111101",
  38071=>"010100000",
  38072=>"000100010",
  38073=>"000101100",
  38074=>"000100110",
  38075=>"100001011",
  38076=>"100101010",
  38077=>"000001010",
  38078=>"001000100",
  38079=>"110001101",
  38080=>"111100110",
  38081=>"111110101",
  38082=>"001011011",
  38083=>"111111011",
  38084=>"110010111",
  38085=>"110110101",
  38086=>"001011001",
  38087=>"111111110",
  38088=>"111111100",
  38089=>"111101111",
  38090=>"010110101",
  38091=>"010001010",
  38092=>"110100110",
  38093=>"101000100",
  38094=>"001100111",
  38095=>"010011100",
  38096=>"010011011",
  38097=>"110010011",
  38098=>"010000101",
  38099=>"100100011",
  38100=>"001000100",
  38101=>"010101000",
  38102=>"011010011",
  38103=>"011011101",
  38104=>"000000010",
  38105=>"010101000",
  38106=>"110010100",
  38107=>"110000100",
  38108=>"010000110",
  38109=>"001010110",
  38110=>"011011101",
  38111=>"100001100",
  38112=>"000100111",
  38113=>"100001101",
  38114=>"110010011",
  38115=>"010000001",
  38116=>"010011110",
  38117=>"011001001",
  38118=>"111010101",
  38119=>"010101110",
  38120=>"000110111",
  38121=>"100101001",
  38122=>"101101101",
  38123=>"100100010",
  38124=>"010100110",
  38125=>"100010100",
  38126=>"110000010",
  38127=>"001000111",
  38128=>"011001011",
  38129=>"111101001",
  38130=>"101001000",
  38131=>"110111110",
  38132=>"000011111",
  38133=>"110110100",
  38134=>"111100100",
  38135=>"101000001",
  38136=>"101111011",
  38137=>"001000101",
  38138=>"000111110",
  38139=>"100101111",
  38140=>"100000011",
  38141=>"010000111",
  38142=>"111001101",
  38143=>"111001000",
  38144=>"001011011",
  38145=>"011001111",
  38146=>"010001100",
  38147=>"000011000",
  38148=>"011101000",
  38149=>"100110111",
  38150=>"111100010",
  38151=>"001101110",
  38152=>"100111010",
  38153=>"000101101",
  38154=>"100011100",
  38155=>"110100001",
  38156=>"100011000",
  38157=>"000101000",
  38158=>"101011010",
  38159=>"100100111",
  38160=>"110010111",
  38161=>"011111101",
  38162=>"001011001",
  38163=>"000011001",
  38164=>"111011010",
  38165=>"100101001",
  38166=>"100000100",
  38167=>"111010110",
  38168=>"001101011",
  38169=>"010001011",
  38170=>"110100001",
  38171=>"100111101",
  38172=>"100000111",
  38173=>"010111111",
  38174=>"100001110",
  38175=>"000000000",
  38176=>"101110000",
  38177=>"000110001",
  38178=>"111000000",
  38179=>"011101110",
  38180=>"001001101",
  38181=>"010110011",
  38182=>"001000000",
  38183=>"100001111",
  38184=>"100011000",
  38185=>"001001100",
  38186=>"010110011",
  38187=>"010001010",
  38188=>"010000001",
  38189=>"000010100",
  38190=>"110001111",
  38191=>"100111000",
  38192=>"101010101",
  38193=>"000011111",
  38194=>"000110111",
  38195=>"110011100",
  38196=>"100111110",
  38197=>"000011100",
  38198=>"100110110",
  38199=>"110111000",
  38200=>"101010011",
  38201=>"110010100",
  38202=>"101101000",
  38203=>"001001100",
  38204=>"100101100",
  38205=>"111011010",
  38206=>"110010000",
  38207=>"010011101",
  38208=>"000100001",
  38209=>"001000011",
  38210=>"111001000",
  38211=>"001101000",
  38212=>"000111110",
  38213=>"101101100",
  38214=>"000111011",
  38215=>"010011110",
  38216=>"010101011",
  38217=>"001010110",
  38218=>"011001101",
  38219=>"010011000",
  38220=>"010000110",
  38221=>"011001111",
  38222=>"001111010",
  38223=>"011001000",
  38224=>"110000001",
  38225=>"101100001",
  38226=>"111010000",
  38227=>"010110000",
  38228=>"000000101",
  38229=>"000001011",
  38230=>"000100001",
  38231=>"100110011",
  38232=>"000000101",
  38233=>"000010011",
  38234=>"011001011",
  38235=>"100010001",
  38236=>"111000100",
  38237=>"111001001",
  38238=>"011001001",
  38239=>"011111101",
  38240=>"110110010",
  38241=>"101100111",
  38242=>"111001110",
  38243=>"101110111",
  38244=>"110010101",
  38245=>"100010010",
  38246=>"110000110",
  38247=>"110000111",
  38248=>"000100001",
  38249=>"011010001",
  38250=>"111100011",
  38251=>"110010001",
  38252=>"110011101",
  38253=>"111110101",
  38254=>"111110111",
  38255=>"110101110",
  38256=>"101011111",
  38257=>"000101101",
  38258=>"110110101",
  38259=>"000110110",
  38260=>"110111011",
  38261=>"100110101",
  38262=>"000110110",
  38263=>"001001100",
  38264=>"110010010",
  38265=>"011001111",
  38266=>"111001100",
  38267=>"111110110",
  38268=>"000110011",
  38269=>"000100000",
  38270=>"001111011",
  38271=>"111111100",
  38272=>"101000100",
  38273=>"100010010",
  38274=>"101110001",
  38275=>"111011000",
  38276=>"000011101",
  38277=>"000100010",
  38278=>"100000000",
  38279=>"100000010",
  38280=>"011001010",
  38281=>"000010000",
  38282=>"000001000",
  38283=>"110011101",
  38284=>"101100110",
  38285=>"000000101",
  38286=>"100011000",
  38287=>"111101101",
  38288=>"100000111",
  38289=>"110001000",
  38290=>"000100001",
  38291=>"010110111",
  38292=>"010001000",
  38293=>"110010100",
  38294=>"110100111",
  38295=>"011111111",
  38296=>"001111010",
  38297=>"000100000",
  38298=>"111000010",
  38299=>"101001010",
  38300=>"100000101",
  38301=>"101111011",
  38302=>"010011011",
  38303=>"011111011",
  38304=>"111101111",
  38305=>"010100001",
  38306=>"110100101",
  38307=>"000110111",
  38308=>"000110100",
  38309=>"001001000",
  38310=>"010111011",
  38311=>"010100100",
  38312=>"010010011",
  38313=>"101111100",
  38314=>"111011000",
  38315=>"010000010",
  38316=>"110110110",
  38317=>"011101111",
  38318=>"010111110",
  38319=>"100001101",
  38320=>"001011100",
  38321=>"110100100",
  38322=>"000100100",
  38323=>"110010101",
  38324=>"101111000",
  38325=>"100111001",
  38326=>"101111101",
  38327=>"011111011",
  38328=>"011011100",
  38329=>"111001011",
  38330=>"011110111",
  38331=>"010110001",
  38332=>"100010100",
  38333=>"110011001",
  38334=>"100010110",
  38335=>"111111011",
  38336=>"010011010",
  38337=>"001010100",
  38338=>"110010101",
  38339=>"111010010",
  38340=>"001011011",
  38341=>"011000010",
  38342=>"011000110",
  38343=>"000000011",
  38344=>"011100001",
  38345=>"111001100",
  38346=>"011000001",
  38347=>"110110001",
  38348=>"010011001",
  38349=>"000100111",
  38350=>"111010101",
  38351=>"000110111",
  38352=>"101110100",
  38353=>"110010001",
  38354=>"011000011",
  38355=>"110111100",
  38356=>"001111100",
  38357=>"100010011",
  38358=>"000111000",
  38359=>"111001100",
  38360=>"001010101",
  38361=>"010000000",
  38362=>"110100000",
  38363=>"111011000",
  38364=>"000001010",
  38365=>"100011111",
  38366=>"110110000",
  38367=>"100110111",
  38368=>"000101101",
  38369=>"011101001",
  38370=>"000001010",
  38371=>"100010101",
  38372=>"010110010",
  38373=>"010111001",
  38374=>"111001111",
  38375=>"001111011",
  38376=>"001000110",
  38377=>"110011010",
  38378=>"000101100",
  38379=>"000000111",
  38380=>"000010001",
  38381=>"001101101",
  38382=>"010011011",
  38383=>"000001001",
  38384=>"001000110",
  38385=>"110110001",
  38386=>"110001101",
  38387=>"001010001",
  38388=>"000110111",
  38389=>"011100110",
  38390=>"101010010",
  38391=>"110000000",
  38392=>"101101011",
  38393=>"110010100",
  38394=>"100100000",
  38395=>"111110110",
  38396=>"000000101",
  38397=>"001010011",
  38398=>"000111010",
  38399=>"000010101",
  38400=>"011001001",
  38401=>"111101110",
  38402=>"011010000",
  38403=>"001001011",
  38404=>"010111101",
  38405=>"010001011",
  38406=>"100111101",
  38407=>"010110111",
  38408=>"010011110",
  38409=>"001000010",
  38410=>"001111000",
  38411=>"001011001",
  38412=>"100111111",
  38413=>"101011010",
  38414=>"010100001",
  38415=>"011010000",
  38416=>"110111110",
  38417=>"101011100",
  38418=>"111111100",
  38419=>"001001110",
  38420=>"011001101",
  38421=>"111011101",
  38422=>"000101010",
  38423=>"001111011",
  38424=>"111101101",
  38425=>"001110010",
  38426=>"000001011",
  38427=>"111010000",
  38428=>"011111101",
  38429=>"010100001",
  38430=>"111001100",
  38431=>"110000101",
  38432=>"111000000",
  38433=>"100101001",
  38434=>"000010110",
  38435=>"110100010",
  38436=>"100001010",
  38437=>"111110100",
  38438=>"010011101",
  38439=>"111101011",
  38440=>"011110010",
  38441=>"010110111",
  38442=>"010101000",
  38443=>"111110110",
  38444=>"011010001",
  38445=>"101110100",
  38446=>"100000010",
  38447=>"010111010",
  38448=>"000010010",
  38449=>"000011001",
  38450=>"001010110",
  38451=>"101010000",
  38452=>"000101110",
  38453=>"101001111",
  38454=>"000000000",
  38455=>"001011100",
  38456=>"011000100",
  38457=>"100101001",
  38458=>"111010101",
  38459=>"111100111",
  38460=>"110100101",
  38461=>"000000010",
  38462=>"000010011",
  38463=>"110100101",
  38464=>"001011101",
  38465=>"010001101",
  38466=>"100111111",
  38467=>"101011000",
  38468=>"001100100",
  38469=>"100000110",
  38470=>"000001001",
  38471=>"101001111",
  38472=>"010001111",
  38473=>"110001001",
  38474=>"001101010",
  38475=>"100110011",
  38476=>"111010110",
  38477=>"100101111",
  38478=>"100111111",
  38479=>"010100001",
  38480=>"010100000",
  38481=>"100010000",
  38482=>"000111100",
  38483=>"111001111",
  38484=>"111010100",
  38485=>"000001010",
  38486=>"001100000",
  38487=>"101100111",
  38488=>"001001111",
  38489=>"100011101",
  38490=>"011011011",
  38491=>"001011000",
  38492=>"111000101",
  38493=>"000001110",
  38494=>"111100100",
  38495=>"110110001",
  38496=>"111001010",
  38497=>"100010000",
  38498=>"100111100",
  38499=>"011100001",
  38500=>"000101101",
  38501=>"001010111",
  38502=>"100100100",
  38503=>"011011000",
  38504=>"000101111",
  38505=>"000100011",
  38506=>"010111111",
  38507=>"000011110",
  38508=>"110011111",
  38509=>"011101000",
  38510=>"100111011",
  38511=>"100010011",
  38512=>"001101111",
  38513=>"101000001",
  38514=>"101011101",
  38515=>"100101100",
  38516=>"111000011",
  38517=>"010011101",
  38518=>"111001110",
  38519=>"110101000",
  38520=>"100011100",
  38521=>"111011101",
  38522=>"111011100",
  38523=>"011111100",
  38524=>"111010110",
  38525=>"010010011",
  38526=>"100110111",
  38527=>"111011110",
  38528=>"010000101",
  38529=>"011100110",
  38530=>"100100111",
  38531=>"000100010",
  38532=>"011011011",
  38533=>"011111101",
  38534=>"110110111",
  38535=>"011010000",
  38536=>"000011100",
  38537=>"000000100",
  38538=>"011010010",
  38539=>"110010111",
  38540=>"111001101",
  38541=>"010000101",
  38542=>"000000010",
  38543=>"100100101",
  38544=>"001011011",
  38545=>"100111011",
  38546=>"000011111",
  38547=>"110001000",
  38548=>"011010001",
  38549=>"101011111",
  38550=>"111000110",
  38551=>"011001000",
  38552=>"010111011",
  38553=>"011001101",
  38554=>"101000101",
  38555=>"000100101",
  38556=>"011000010",
  38557=>"101100111",
  38558=>"011001110",
  38559=>"111011000",
  38560=>"011100100",
  38561=>"111100000",
  38562=>"010011101",
  38563=>"100111010",
  38564=>"111100110",
  38565=>"010110000",
  38566=>"100101101",
  38567=>"000001101",
  38568=>"001000000",
  38569=>"001101010",
  38570=>"100010100",
  38571=>"001001110",
  38572=>"010100110",
  38573=>"010110000",
  38574=>"011111101",
  38575=>"000101100",
  38576=>"010000111",
  38577=>"011100100",
  38578=>"101011000",
  38579=>"000100100",
  38580=>"111111100",
  38581=>"101001010",
  38582=>"001000011",
  38583=>"011110100",
  38584=>"111011110",
  38585=>"110111111",
  38586=>"111000010",
  38587=>"111000100",
  38588=>"000101011",
  38589=>"101101110",
  38590=>"101001111",
  38591=>"000010001",
  38592=>"001101111",
  38593=>"100101100",
  38594=>"111010101",
  38595=>"110011111",
  38596=>"000100000",
  38597=>"010000010",
  38598=>"000100110",
  38599=>"001101000",
  38600=>"100000111",
  38601=>"010100001",
  38602=>"000100001",
  38603=>"011000011",
  38604=>"110010101",
  38605=>"001111000",
  38606=>"111111101",
  38607=>"111011011",
  38608=>"110011111",
  38609=>"110101001",
  38610=>"110001111",
  38611=>"111011111",
  38612=>"101000011",
  38613=>"010101011",
  38614=>"100110111",
  38615=>"001011001",
  38616=>"011011011",
  38617=>"110110001",
  38618=>"000100000",
  38619=>"011011011",
  38620=>"000100111",
  38621=>"010000100",
  38622=>"100110010",
  38623=>"010100001",
  38624=>"001000101",
  38625=>"111001101",
  38626=>"101100101",
  38627=>"101111000",
  38628=>"010100000",
  38629=>"010111110",
  38630=>"000100101",
  38631=>"011011111",
  38632=>"110011010",
  38633=>"011000000",
  38634=>"111100100",
  38635=>"000001011",
  38636=>"000000111",
  38637=>"001001011",
  38638=>"111001000",
  38639=>"011001100",
  38640=>"100100111",
  38641=>"010011110",
  38642=>"100100101",
  38643=>"100100111",
  38644=>"111110100",
  38645=>"001100000",
  38646=>"010010001",
  38647=>"000101001",
  38648=>"111110110",
  38649=>"111011111",
  38650=>"110001100",
  38651=>"000100011",
  38652=>"101001111",
  38653=>"011111011",
  38654=>"100011011",
  38655=>"111101011",
  38656=>"100100100",
  38657=>"000100100",
  38658=>"010010100",
  38659=>"001010110",
  38660=>"011000010",
  38661=>"110100000",
  38662=>"110101101",
  38663=>"100100110",
  38664=>"110110110",
  38665=>"111000101",
  38666=>"110010001",
  38667=>"010001011",
  38668=>"000101111",
  38669=>"010011000",
  38670=>"101011010",
  38671=>"000110110",
  38672=>"101010011",
  38673=>"011100001",
  38674=>"000011111",
  38675=>"101000111",
  38676=>"100110101",
  38677=>"110111001",
  38678=>"011100101",
  38679=>"100011100",
  38680=>"111001101",
  38681=>"000111100",
  38682=>"000100010",
  38683=>"000100010",
  38684=>"001000000",
  38685=>"000011101",
  38686=>"101011010",
  38687=>"001011011",
  38688=>"000001010",
  38689=>"001000100",
  38690=>"111101010",
  38691=>"100010000",
  38692=>"011011100",
  38693=>"100101111",
  38694=>"000110110",
  38695=>"000001011",
  38696=>"010000000",
  38697=>"100111110",
  38698=>"001010101",
  38699=>"000001010",
  38700=>"000111110",
  38701=>"010001011",
  38702=>"101110010",
  38703=>"101100001",
  38704=>"111011111",
  38705=>"100111010",
  38706=>"000000011",
  38707=>"101110010",
  38708=>"110100001",
  38709=>"101100001",
  38710=>"010100100",
  38711=>"111000001",
  38712=>"001111110",
  38713=>"010101100",
  38714=>"010011000",
  38715=>"110010100",
  38716=>"100011110",
  38717=>"000111100",
  38718=>"101000000",
  38719=>"101000000",
  38720=>"010001010",
  38721=>"010110010",
  38722=>"111110100",
  38723=>"000000100",
  38724=>"110101100",
  38725=>"111101111",
  38726=>"111111010",
  38727=>"101111010",
  38728=>"000111111",
  38729=>"101011111",
  38730=>"110001001",
  38731=>"111100110",
  38732=>"011000001",
  38733=>"101001001",
  38734=>"001101011",
  38735=>"101110100",
  38736=>"101111111",
  38737=>"100100100",
  38738=>"110001101",
  38739=>"010000000",
  38740=>"100101111",
  38741=>"001100001",
  38742=>"101101000",
  38743=>"100001111",
  38744=>"111100010",
  38745=>"111101100",
  38746=>"100111101",
  38747=>"111010000",
  38748=>"000110110",
  38749=>"001111001",
  38750=>"001111010",
  38751=>"010100011",
  38752=>"001001000",
  38753=>"100001000",
  38754=>"010110110",
  38755=>"010000001",
  38756=>"011001100",
  38757=>"010010100",
  38758=>"101101101",
  38759=>"010111001",
  38760=>"001010001",
  38761=>"010100001",
  38762=>"101000100",
  38763=>"011000110",
  38764=>"110110001",
  38765=>"110011101",
  38766=>"110111101",
  38767=>"100101011",
  38768=>"000011011",
  38769=>"011000010",
  38770=>"001101111",
  38771=>"011101001",
  38772=>"001101101",
  38773=>"011111010",
  38774=>"001101101",
  38775=>"101001101",
  38776=>"001011101",
  38777=>"111111111",
  38778=>"001111110",
  38779=>"010101101",
  38780=>"001110011",
  38781=>"100101000",
  38782=>"111101111",
  38783=>"100011110",
  38784=>"011110000",
  38785=>"010100110",
  38786=>"001000101",
  38787=>"000100101",
  38788=>"110100010",
  38789=>"001011001",
  38790=>"100000111",
  38791=>"000011101",
  38792=>"110111001",
  38793=>"010000000",
  38794=>"110110101",
  38795=>"110001101",
  38796=>"001010010",
  38797=>"001100110",
  38798=>"010100001",
  38799=>"101010001",
  38800=>"101110110",
  38801=>"100110010",
  38802=>"101100101",
  38803=>"000110110",
  38804=>"001100101",
  38805=>"110001010",
  38806=>"000011001",
  38807=>"101010001",
  38808=>"101100101",
  38809=>"111101011",
  38810=>"000100101",
  38811=>"110100000",
  38812=>"100101100",
  38813=>"001010110",
  38814=>"101100110",
  38815=>"101000101",
  38816=>"111100111",
  38817=>"111001100",
  38818=>"011001011",
  38819=>"001111101",
  38820=>"101110000",
  38821=>"011000101",
  38822=>"101110110",
  38823=>"001001001",
  38824=>"110010100",
  38825=>"101011011",
  38826=>"110111001",
  38827=>"000111100",
  38828=>"111001000",
  38829=>"000110000",
  38830=>"001001001",
  38831=>"101001001",
  38832=>"100011010",
  38833=>"011101010",
  38834=>"001101111",
  38835=>"011001111",
  38836=>"100100111",
  38837=>"011101111",
  38838=>"110101010",
  38839=>"101100101",
  38840=>"000110000",
  38841=>"000011011",
  38842=>"000000011",
  38843=>"101000001",
  38844=>"001110011",
  38845=>"101100110",
  38846=>"001100000",
  38847=>"101100101",
  38848=>"111001001",
  38849=>"001001000",
  38850=>"010010100",
  38851=>"110101110",
  38852=>"010000000",
  38853=>"111001000",
  38854=>"010111000",
  38855=>"110010000",
  38856=>"001000100",
  38857=>"001010010",
  38858=>"111110110",
  38859=>"000110111",
  38860=>"111111000",
  38861=>"110101001",
  38862=>"000001110",
  38863=>"011010000",
  38864=>"111000011",
  38865=>"100100010",
  38866=>"100100111",
  38867=>"000001000",
  38868=>"101001111",
  38869=>"001110011",
  38870=>"010011011",
  38871=>"110101001",
  38872=>"110101001",
  38873=>"100101101",
  38874=>"010001001",
  38875=>"100010100",
  38876=>"010101101",
  38877=>"110001100",
  38878=>"111001111",
  38879=>"010110001",
  38880=>"001001011",
  38881=>"111001111",
  38882=>"111100100",
  38883=>"001111000",
  38884=>"100001011",
  38885=>"100110101",
  38886=>"111110000",
  38887=>"010110101",
  38888=>"100101000",
  38889=>"000000000",
  38890=>"011000110",
  38891=>"000001111",
  38892=>"011001100",
  38893=>"101000100",
  38894=>"010011001",
  38895=>"010010000",
  38896=>"111111010",
  38897=>"110011001",
  38898=>"000011010",
  38899=>"011001100",
  38900=>"110100100",
  38901=>"110010010",
  38902=>"011111111",
  38903=>"101110000",
  38904=>"001111101",
  38905=>"110100101",
  38906=>"010101100",
  38907=>"010101011",
  38908=>"111101000",
  38909=>"010100000",
  38910=>"111011101",
  38911=>"011100111",
  38912=>"110110010",
  38913=>"101110000",
  38914=>"010001000",
  38915=>"110000100",
  38916=>"110000100",
  38917=>"110010000",
  38918=>"000110001",
  38919=>"010111100",
  38920=>"010011111",
  38921=>"000010101",
  38922=>"110100110",
  38923=>"010010101",
  38924=>"001000011",
  38925=>"000001110",
  38926=>"101010101",
  38927=>"110000011",
  38928=>"000011100",
  38929=>"111110001",
  38930=>"111001101",
  38931=>"011101010",
  38932=>"101111101",
  38933=>"101110100",
  38934=>"011011011",
  38935=>"110010100",
  38936=>"000100110",
  38937=>"010100000",
  38938=>"111110010",
  38939=>"101111110",
  38940=>"001011111",
  38941=>"001000011",
  38942=>"100110010",
  38943=>"011010010",
  38944=>"001111000",
  38945=>"111000100",
  38946=>"111110100",
  38947=>"000011011",
  38948=>"011100011",
  38949=>"001001001",
  38950=>"111101011",
  38951=>"010000101",
  38952=>"010101011",
  38953=>"110111101",
  38954=>"000000001",
  38955=>"100000011",
  38956=>"110110111",
  38957=>"100101001",
  38958=>"110111101",
  38959=>"011101100",
  38960=>"011110110",
  38961=>"111110001",
  38962=>"110110001",
  38963=>"111011001",
  38964=>"010100011",
  38965=>"011011001",
  38966=>"110011010",
  38967=>"001110101",
  38968=>"100110001",
  38969=>"001100111",
  38970=>"111011001",
  38971=>"100001011",
  38972=>"100001101",
  38973=>"100010000",
  38974=>"000110111",
  38975=>"111100001",
  38976=>"011110101",
  38977=>"001010100",
  38978=>"001010110",
  38979=>"011011010",
  38980=>"000111100",
  38981=>"011000110",
  38982=>"011111111",
  38983=>"111111010",
  38984=>"000110111",
  38985=>"100011110",
  38986=>"100011010",
  38987=>"100101000",
  38988=>"011010010",
  38989=>"011100111",
  38990=>"010111011",
  38991=>"110011000",
  38992=>"111101111",
  38993=>"111101100",
  38994=>"101000000",
  38995=>"000011001",
  38996=>"100110000",
  38997=>"010001111",
  38998=>"100100110",
  38999=>"101000011",
  39000=>"001001111",
  39001=>"001101110",
  39002=>"010100001",
  39003=>"101000011",
  39004=>"100100001",
  39005=>"001001110",
  39006=>"010000111",
  39007=>"000100011",
  39008=>"110110001",
  39009=>"101000000",
  39010=>"101000111",
  39011=>"010111001",
  39012=>"000100101",
  39013=>"100100111",
  39014=>"100000000",
  39015=>"000010000",
  39016=>"111000000",
  39017=>"111001101",
  39018=>"011000001",
  39019=>"010101010",
  39020=>"100110001",
  39021=>"010110110",
  39022=>"101000101",
  39023=>"111001000",
  39024=>"011110010",
  39025=>"000100001",
  39026=>"000000011",
  39027=>"001100000",
  39028=>"101111001",
  39029=>"000110011",
  39030=>"000100011",
  39031=>"101110011",
  39032=>"000101001",
  39033=>"000100001",
  39034=>"000011111",
  39035=>"001101000",
  39036=>"100111010",
  39037=>"110000101",
  39038=>"101111001",
  39039=>"000011010",
  39040=>"001101010",
  39041=>"010011100",
  39042=>"011011001",
  39043=>"110001010",
  39044=>"110001001",
  39045=>"100101011",
  39046=>"011011101",
  39047=>"111100100",
  39048=>"101001000",
  39049=>"001011011",
  39050=>"100111000",
  39051=>"101001000",
  39052=>"010101000",
  39053=>"001101011",
  39054=>"100111001",
  39055=>"111101010",
  39056=>"100100000",
  39057=>"000010010",
  39058=>"111011011",
  39059=>"000010001",
  39060=>"101010111",
  39061=>"001010001",
  39062=>"111011000",
  39063=>"101101011",
  39064=>"000000110",
  39065=>"100011001",
  39066=>"111110101",
  39067=>"000111100",
  39068=>"100010010",
  39069=>"010010011",
  39070=>"000111000",
  39071=>"101111000",
  39072=>"001011100",
  39073=>"101101000",
  39074=>"111001101",
  39075=>"001100010",
  39076=>"110010101",
  39077=>"100000111",
  39078=>"111101010",
  39079=>"010011010",
  39080=>"111010111",
  39081=>"010111011",
  39082=>"001111110",
  39083=>"100010101",
  39084=>"111100111",
  39085=>"101001000",
  39086=>"100011111",
  39087=>"111001111",
  39088=>"011111111",
  39089=>"010110111",
  39090=>"001000110",
  39091=>"111110000",
  39092=>"111100101",
  39093=>"100110101",
  39094=>"010010001",
  39095=>"101100110",
  39096=>"011010101",
  39097=>"001101011",
  39098=>"011000000",
  39099=>"001111110",
  39100=>"011011010",
  39101=>"011101000",
  39102=>"010001011",
  39103=>"101010100",
  39104=>"001101011",
  39105=>"100101010",
  39106=>"100100000",
  39107=>"110110000",
  39108=>"000110011",
  39109=>"110011001",
  39110=>"010100110",
  39111=>"000111100",
  39112=>"100101100",
  39113=>"001110010",
  39114=>"000000011",
  39115=>"111010000",
  39116=>"011100010",
  39117=>"111100001",
  39118=>"011010000",
  39119=>"000100100",
  39120=>"100011101",
  39121=>"010100111",
  39122=>"111100010",
  39123=>"100101001",
  39124=>"100101000",
  39125=>"011101101",
  39126=>"101000100",
  39127=>"001001011",
  39128=>"010010011",
  39129=>"101100001",
  39130=>"000111011",
  39131=>"000000010",
  39132=>"110011011",
  39133=>"100111001",
  39134=>"111101001",
  39135=>"111011011",
  39136=>"010110001",
  39137=>"000100010",
  39138=>"011000100",
  39139=>"011001000",
  39140=>"111000110",
  39141=>"101100001",
  39142=>"111110111",
  39143=>"010111111",
  39144=>"101101110",
  39145=>"100010100",
  39146=>"100010110",
  39147=>"001000101",
  39148=>"111101011",
  39149=>"001001101",
  39150=>"010000001",
  39151=>"001010111",
  39152=>"110010010",
  39153=>"111011001",
  39154=>"100010100",
  39155=>"011110001",
  39156=>"101101100",
  39157=>"111011011",
  39158=>"111101000",
  39159=>"100110000",
  39160=>"101011100",
  39161=>"111001011",
  39162=>"101000011",
  39163=>"100000101",
  39164=>"100110101",
  39165=>"011111001",
  39166=>"011101101",
  39167=>"010010010",
  39168=>"100001110",
  39169=>"111110011",
  39170=>"010110011",
  39171=>"010100011",
  39172=>"010000100",
  39173=>"001110110",
  39174=>"000111000",
  39175=>"110010100",
  39176=>"101100101",
  39177=>"010101101",
  39178=>"000111101",
  39179=>"010100101",
  39180=>"101001110",
  39181=>"011010010",
  39182=>"010010010",
  39183=>"101111000",
  39184=>"011000000",
  39185=>"010001000",
  39186=>"110000110",
  39187=>"100101110",
  39188=>"011000011",
  39189=>"001011110",
  39190=>"110100101",
  39191=>"111011101",
  39192=>"010110100",
  39193=>"010101100",
  39194=>"001000101",
  39195=>"100101100",
  39196=>"000110101",
  39197=>"111000100",
  39198=>"101011010",
  39199=>"111100010",
  39200=>"010000000",
  39201=>"001111001",
  39202=>"011000110",
  39203=>"001010001",
  39204=>"100110001",
  39205=>"010111010",
  39206=>"011010001",
  39207=>"110000101",
  39208=>"100101000",
  39209=>"010001011",
  39210=>"000011000",
  39211=>"110110111",
  39212=>"110100001",
  39213=>"100111100",
  39214=>"111010110",
  39215=>"100010110",
  39216=>"110111100",
  39217=>"101101101",
  39218=>"001011101",
  39219=>"101111000",
  39220=>"111000100",
  39221=>"111111001",
  39222=>"010100110",
  39223=>"100010000",
  39224=>"000010011",
  39225=>"111111111",
  39226=>"101101001",
  39227=>"101001010",
  39228=>"110010000",
  39229=>"101101010",
  39230=>"010101000",
  39231=>"010100011",
  39232=>"000010001",
  39233=>"011000010",
  39234=>"001001010",
  39235=>"101001111",
  39236=>"110010100",
  39237=>"111011000",
  39238=>"111101110",
  39239=>"110001001",
  39240=>"100101101",
  39241=>"011011001",
  39242=>"101111101",
  39243=>"000000111",
  39244=>"110111101",
  39245=>"110100010",
  39246=>"110001111",
  39247=>"111110110",
  39248=>"010100111",
  39249=>"010001110",
  39250=>"001000010",
  39251=>"001000100",
  39252=>"010011100",
  39253=>"110101001",
  39254=>"111111000",
  39255=>"101100111",
  39256=>"100011010",
  39257=>"101110010",
  39258=>"001001110",
  39259=>"101100100",
  39260=>"111001101",
  39261=>"011011000",
  39262=>"101010110",
  39263=>"100001100",
  39264=>"101100010",
  39265=>"011011110",
  39266=>"010011000",
  39267=>"000101100",
  39268=>"101111011",
  39269=>"111011000",
  39270=>"101001111",
  39271=>"000010010",
  39272=>"011111111",
  39273=>"000000000",
  39274=>"111110101",
  39275=>"001001101",
  39276=>"111011101",
  39277=>"101110110",
  39278=>"111101101",
  39279=>"100011111",
  39280=>"101011011",
  39281=>"000100011",
  39282=>"110100101",
  39283=>"111100111",
  39284=>"001000101",
  39285=>"000111111",
  39286=>"001110110",
  39287=>"101101110",
  39288=>"100000000",
  39289=>"111110010",
  39290=>"011001111",
  39291=>"110100101",
  39292=>"011110000",
  39293=>"010111011",
  39294=>"111100000",
  39295=>"101010100",
  39296=>"010100110",
  39297=>"000011110",
  39298=>"011001100",
  39299=>"000001110",
  39300=>"001110111",
  39301=>"111010101",
  39302=>"111001010",
  39303=>"011000011",
  39304=>"010000111",
  39305=>"011001010",
  39306=>"001011001",
  39307=>"000011111",
  39308=>"100111110",
  39309=>"000000010",
  39310=>"010100000",
  39311=>"010011101",
  39312=>"111000011",
  39313=>"100111101",
  39314=>"111111100",
  39315=>"111110011",
  39316=>"101000111",
  39317=>"000100010",
  39318=>"010010101",
  39319=>"011100110",
  39320=>"100001010",
  39321=>"101101010",
  39322=>"111101000",
  39323=>"110100001",
  39324=>"111000001",
  39325=>"100011000",
  39326=>"110001011",
  39327=>"111110010",
  39328=>"101011101",
  39329=>"101101101",
  39330=>"010100110",
  39331=>"001010010",
  39332=>"110101111",
  39333=>"100001101",
  39334=>"111111100",
  39335=>"100101000",
  39336=>"101101110",
  39337=>"000000100",
  39338=>"101000001",
  39339=>"001000011",
  39340=>"011000111",
  39341=>"010000001",
  39342=>"111000011",
  39343=>"111010101",
  39344=>"010100110",
  39345=>"011101111",
  39346=>"101111010",
  39347=>"011111011",
  39348=>"010111110",
  39349=>"000000111",
  39350=>"010110110",
  39351=>"000111110",
  39352=>"101000010",
  39353=>"001010111",
  39354=>"000011000",
  39355=>"000100100",
  39356=>"111000101",
  39357=>"011110001",
  39358=>"010111000",
  39359=>"101010001",
  39360=>"011000000",
  39361=>"000001101",
  39362=>"010111010",
  39363=>"101001011",
  39364=>"011100101",
  39365=>"111100011",
  39366=>"001011100",
  39367=>"000111111",
  39368=>"100000010",
  39369=>"010000010",
  39370=>"001111101",
  39371=>"001010000",
  39372=>"111110101",
  39373=>"100110011",
  39374=>"000111111",
  39375=>"001100101",
  39376=>"100010101",
  39377=>"011100001",
  39378=>"101111100",
  39379=>"110110101",
  39380=>"010010110",
  39381=>"010101100",
  39382=>"010000001",
  39383=>"110110111",
  39384=>"010010011",
  39385=>"111010111",
  39386=>"101110100",
  39387=>"100100010",
  39388=>"110011110",
  39389=>"000000110",
  39390=>"010110001",
  39391=>"001001100",
  39392=>"000111011",
  39393=>"111110011",
  39394=>"000001011",
  39395=>"100001010",
  39396=>"010111100",
  39397=>"101111101",
  39398=>"100011101",
  39399=>"001101110",
  39400=>"001110101",
  39401=>"000110110",
  39402=>"101111011",
  39403=>"100000111",
  39404=>"100101111",
  39405=>"010111000",
  39406=>"101100101",
  39407=>"110100000",
  39408=>"011001110",
  39409=>"000000101",
  39410=>"101101101",
  39411=>"000111111",
  39412=>"001000000",
  39413=>"001000110",
  39414=>"010011011",
  39415=>"000001000",
  39416=>"010101111",
  39417=>"111110000",
  39418=>"110000101",
  39419=>"110111000",
  39420=>"111110100",
  39421=>"100000010",
  39422=>"011010010",
  39423=>"011010011",
  39424=>"000000100",
  39425=>"001010010",
  39426=>"100100011",
  39427=>"111101111",
  39428=>"011010001",
  39429=>"101111110",
  39430=>"111111000",
  39431=>"100001010",
  39432=>"001001101",
  39433=>"100100111",
  39434=>"010110101",
  39435=>"110010101",
  39436=>"110000110",
  39437=>"110100010",
  39438=>"010011011",
  39439=>"101111101",
  39440=>"011010110",
  39441=>"010010111",
  39442=>"110010000",
  39443=>"010010100",
  39444=>"001101100",
  39445=>"000110111",
  39446=>"101001011",
  39447=>"100111101",
  39448=>"100100011",
  39449=>"001100101",
  39450=>"011100111",
  39451=>"001100000",
  39452=>"100101111",
  39453=>"101000001",
  39454=>"001000000",
  39455=>"010100111",
  39456=>"000011000",
  39457=>"001011111",
  39458=>"111000000",
  39459=>"110001100",
  39460=>"110101000",
  39461=>"101001001",
  39462=>"110010101",
  39463=>"010001101",
  39464=>"010000010",
  39465=>"001010001",
  39466=>"010111101",
  39467=>"011001111",
  39468=>"111011111",
  39469=>"010011001",
  39470=>"011101101",
  39471=>"010010011",
  39472=>"011000010",
  39473=>"111101100",
  39474=>"001000011",
  39475=>"001001001",
  39476=>"111010001",
  39477=>"110110011",
  39478=>"101010000",
  39479=>"111100011",
  39480=>"111111011",
  39481=>"100111001",
  39482=>"000101110",
  39483=>"100101111",
  39484=>"011101010",
  39485=>"101011001",
  39486=>"000010000",
  39487=>"001000111",
  39488=>"011111011",
  39489=>"100000111",
  39490=>"011011101",
  39491=>"111100010",
  39492=>"000110101",
  39493=>"010101001",
  39494=>"111010001",
  39495=>"101101101",
  39496=>"001101111",
  39497=>"100110101",
  39498=>"000011010",
  39499=>"010111110",
  39500=>"010010101",
  39501=>"101000010",
  39502=>"011011111",
  39503=>"001110101",
  39504=>"110010000",
  39505=>"110111101",
  39506=>"010000100",
  39507=>"001000010",
  39508=>"100011011",
  39509=>"001101110",
  39510=>"010101001",
  39511=>"101001101",
  39512=>"000011100",
  39513=>"110010110",
  39514=>"000000000",
  39515=>"001000110",
  39516=>"110111111",
  39517=>"100011001",
  39518=>"100000010",
  39519=>"101010001",
  39520=>"100100101",
  39521=>"111000110",
  39522=>"010110011",
  39523=>"100101110",
  39524=>"010100110",
  39525=>"000110101",
  39526=>"111111011",
  39527=>"000000100",
  39528=>"101000010",
  39529=>"011001100",
  39530=>"001011110",
  39531=>"000100000",
  39532=>"000011110",
  39533=>"001000001",
  39534=>"001010000",
  39535=>"111000100",
  39536=>"100011101",
  39537=>"100001010",
  39538=>"011100010",
  39539=>"111100100",
  39540=>"101110101",
  39541=>"111110101",
  39542=>"110001010",
  39543=>"011101111",
  39544=>"110100010",
  39545=>"100001011",
  39546=>"011111010",
  39547=>"100101110",
  39548=>"000010111",
  39549=>"000001011",
  39550=>"101000010",
  39551=>"000001010",
  39552=>"100110111",
  39553=>"101101000",
  39554=>"111000001",
  39555=>"000001000",
  39556=>"100101011",
  39557=>"100110110",
  39558=>"000100110",
  39559=>"010111011",
  39560=>"101101000",
  39561=>"000001101",
  39562=>"110001101",
  39563=>"100101111",
  39564=>"000000101",
  39565=>"010011110",
  39566=>"010011011",
  39567=>"111111111",
  39568=>"000111111",
  39569=>"110010001",
  39570=>"100000010",
  39571=>"100101100",
  39572=>"100011111",
  39573=>"001010010",
  39574=>"011110011",
  39575=>"101011001",
  39576=>"011001001",
  39577=>"110000011",
  39578=>"000101110",
  39579=>"101010100",
  39580=>"101000100",
  39581=>"101101000",
  39582=>"100011000",
  39583=>"100011101",
  39584=>"111011000",
  39585=>"101001001",
  39586=>"101110001",
  39587=>"010111111",
  39588=>"101100000",
  39589=>"001010011",
  39590=>"000001010",
  39591=>"100010010",
  39592=>"001011001",
  39593=>"000000000",
  39594=>"101001011",
  39595=>"101000100",
  39596=>"100000100",
  39597=>"011000110",
  39598=>"000101010",
  39599=>"100010111",
  39600=>"100000101",
  39601=>"011110000",
  39602=>"100100011",
  39603=>"001011001",
  39604=>"011001000",
  39605=>"011100100",
  39606=>"001110111",
  39607=>"000010000",
  39608=>"101000101",
  39609=>"001001001",
  39610=>"010001000",
  39611=>"001001110",
  39612=>"001111011",
  39613=>"101001101",
  39614=>"000110001",
  39615=>"000101110",
  39616=>"000101100",
  39617=>"111000010",
  39618=>"111110100",
  39619=>"010010110",
  39620=>"010100010",
  39621=>"010010111",
  39622=>"111001101",
  39623=>"101111001",
  39624=>"110110111",
  39625=>"001100111",
  39626=>"100000100",
  39627=>"001000001",
  39628=>"011001110",
  39629=>"011100100",
  39630=>"001110010",
  39631=>"010100000",
  39632=>"000101101",
  39633=>"110000011",
  39634=>"011110011",
  39635=>"000100111",
  39636=>"101001010",
  39637=>"111110010",
  39638=>"110100111",
  39639=>"011101000",
  39640=>"011111001",
  39641=>"110001011",
  39642=>"111110001",
  39643=>"000101010",
  39644=>"100010010",
  39645=>"111100100",
  39646=>"111011010",
  39647=>"011111001",
  39648=>"000000110",
  39649=>"100101001",
  39650=>"011001010",
  39651=>"000111010",
  39652=>"001101001",
  39653=>"010010000",
  39654=>"001011100",
  39655=>"000110100",
  39656=>"010010011",
  39657=>"001000011",
  39658=>"001110110",
  39659=>"100000111",
  39660=>"110111100",
  39661=>"101001001",
  39662=>"110110001",
  39663=>"000000100",
  39664=>"110111001",
  39665=>"011101001",
  39666=>"111000100",
  39667=>"100110001",
  39668=>"001110001",
  39669=>"011100111",
  39670=>"110000101",
  39671=>"101000000",
  39672=>"011010011",
  39673=>"000000101",
  39674=>"101110001",
  39675=>"100001101",
  39676=>"000101111",
  39677=>"101000010",
  39678=>"100101101",
  39679=>"111010000",
  39680=>"100110000",
  39681=>"101100010",
  39682=>"111101010",
  39683=>"101010010",
  39684=>"110111101",
  39685=>"100010000",
  39686=>"010010010",
  39687=>"001111010",
  39688=>"101101011",
  39689=>"010101001",
  39690=>"000111000",
  39691=>"001100001",
  39692=>"100111110",
  39693=>"011000111",
  39694=>"000111100",
  39695=>"110011000",
  39696=>"011000110",
  39697=>"100110001",
  39698=>"110011110",
  39699=>"000000011",
  39700=>"100110111",
  39701=>"010010011",
  39702=>"111001001",
  39703=>"010100100",
  39704=>"101101001",
  39705=>"011100000",
  39706=>"000010001",
  39707=>"001111111",
  39708=>"110111011",
  39709=>"100101100",
  39710=>"100111000",
  39711=>"100110010",
  39712=>"111001001",
  39713=>"110011100",
  39714=>"011111011",
  39715=>"000011000",
  39716=>"010000010",
  39717=>"101010111",
  39718=>"010101100",
  39719=>"110111000",
  39720=>"110011110",
  39721=>"001101011",
  39722=>"110001011",
  39723=>"000011000",
  39724=>"110011011",
  39725=>"101000011",
  39726=>"001000011",
  39727=>"100111001",
  39728=>"000101100",
  39729=>"010100101",
  39730=>"110000100",
  39731=>"110010011",
  39732=>"011110111",
  39733=>"101010111",
  39734=>"100110000",
  39735=>"110011100",
  39736=>"001111101",
  39737=>"110111011",
  39738=>"111100110",
  39739=>"010100000",
  39740=>"111101000",
  39741=>"111101001",
  39742=>"100110001",
  39743=>"101001000",
  39744=>"101101110",
  39745=>"001100000",
  39746=>"111000011",
  39747=>"110011101",
  39748=>"111001101",
  39749=>"010111010",
  39750=>"000100001",
  39751=>"001111010",
  39752=>"011001010",
  39753=>"000000100",
  39754=>"111011110",
  39755=>"011101001",
  39756=>"111111010",
  39757=>"010101011",
  39758=>"100110100",
  39759=>"011010111",
  39760=>"111101111",
  39761=>"111101100",
  39762=>"011001000",
  39763=>"000000110",
  39764=>"011111000",
  39765=>"000110100",
  39766=>"101111001",
  39767=>"000110001",
  39768=>"010101110",
  39769=>"010101001",
  39770=>"101111100",
  39771=>"001011001",
  39772=>"101110110",
  39773=>"000001110",
  39774=>"010110011",
  39775=>"101111010",
  39776=>"010100001",
  39777=>"110101011",
  39778=>"010001100",
  39779=>"011011111",
  39780=>"111001101",
  39781=>"001011101",
  39782=>"011110000",
  39783=>"101000000",
  39784=>"111100100",
  39785=>"010101111",
  39786=>"100010100",
  39787=>"101000110",
  39788=>"000001101",
  39789=>"110010010",
  39790=>"101000110",
  39791=>"011110000",
  39792=>"111000110",
  39793=>"011110001",
  39794=>"101101100",
  39795=>"001000011",
  39796=>"100110111",
  39797=>"000010110",
  39798=>"010100001",
  39799=>"100111111",
  39800=>"100100110",
  39801=>"001000111",
  39802=>"000000100",
  39803=>"011111010",
  39804=>"111110000",
  39805=>"100111110",
  39806=>"100110101",
  39807=>"011000000",
  39808=>"011101001",
  39809=>"011011111",
  39810=>"101100011",
  39811=>"000011110",
  39812=>"110011100",
  39813=>"101011010",
  39814=>"111000011",
  39815=>"010000010",
  39816=>"101011101",
  39817=>"000000010",
  39818=>"101001101",
  39819=>"111001101",
  39820=>"010100010",
  39821=>"101010110",
  39822=>"001000110",
  39823=>"101011101",
  39824=>"111111010",
  39825=>"110001110",
  39826=>"111101000",
  39827=>"101101010",
  39828=>"001001101",
  39829=>"000101000",
  39830=>"110111111",
  39831=>"001000000",
  39832=>"000110100",
  39833=>"110100000",
  39834=>"111101110",
  39835=>"101001100",
  39836=>"101110011",
  39837=>"001001110",
  39838=>"100000001",
  39839=>"100010010",
  39840=>"100010010",
  39841=>"010001001",
  39842=>"001001010",
  39843=>"110100011",
  39844=>"010011000",
  39845=>"011000111",
  39846=>"100100101",
  39847=>"000001111",
  39848=>"111110101",
  39849=>"010101100",
  39850=>"100001010",
  39851=>"000011110",
  39852=>"111010111",
  39853=>"101111100",
  39854=>"111110110",
  39855=>"001100010",
  39856=>"111001001",
  39857=>"010000011",
  39858=>"101101000",
  39859=>"001010101",
  39860=>"111110110",
  39861=>"100010111",
  39862=>"101100110",
  39863=>"001100010",
  39864=>"000101101",
  39865=>"010111100",
  39866=>"011100011",
  39867=>"010101011",
  39868=>"110110011",
  39869=>"100100100",
  39870=>"111011011",
  39871=>"011000100",
  39872=>"101001101",
  39873=>"010011001",
  39874=>"010000111",
  39875=>"001010000",
  39876=>"000110101",
  39877=>"111111000",
  39878=>"101010001",
  39879=>"000101001",
  39880=>"000110110",
  39881=>"000000011",
  39882=>"001010101",
  39883=>"000000000",
  39884=>"111101110",
  39885=>"000100111",
  39886=>"000110101",
  39887=>"010000011",
  39888=>"000111110",
  39889=>"001011001",
  39890=>"101010110",
  39891=>"101000111",
  39892=>"011001000",
  39893=>"101000111",
  39894=>"110100101",
  39895=>"111111001",
  39896=>"100001101",
  39897=>"111010111",
  39898=>"001000000",
  39899=>"000001000",
  39900=>"000010100",
  39901=>"001110101",
  39902=>"011110000",
  39903=>"001011100",
  39904=>"111011110",
  39905=>"001110100",
  39906=>"110000100",
  39907=>"100000100",
  39908=>"111101100",
  39909=>"011010111",
  39910=>"011011011",
  39911=>"111101111",
  39912=>"111001100",
  39913=>"000000011",
  39914=>"110100011",
  39915=>"000010010",
  39916=>"111000110",
  39917=>"101111011",
  39918=>"101000101",
  39919=>"011011010",
  39920=>"010110000",
  39921=>"011101110",
  39922=>"011010100",
  39923=>"110011110",
  39924=>"110010111",
  39925=>"111000010",
  39926=>"101100100",
  39927=>"110110010",
  39928=>"000001010",
  39929=>"111010110",
  39930=>"011110111",
  39931=>"001010001",
  39932=>"110000101",
  39933=>"001011111",
  39934=>"011011110",
  39935=>"111010001",
  39936=>"100100011",
  39937=>"000000101",
  39938=>"101111011",
  39939=>"101011111",
  39940=>"000100011",
  39941=>"001001110",
  39942=>"011010100",
  39943=>"011001000",
  39944=>"101100000",
  39945=>"000011000",
  39946=>"011001011",
  39947=>"101111110",
  39948=>"001000111",
  39949=>"110010100",
  39950=>"100010011",
  39951=>"001011000",
  39952=>"010001011",
  39953=>"011101101",
  39954=>"101100110",
  39955=>"110100100",
  39956=>"110010000",
  39957=>"000011111",
  39958=>"001111101",
  39959=>"100001010",
  39960=>"001101101",
  39961=>"001000010",
  39962=>"010111011",
  39963=>"101011010",
  39964=>"001110110",
  39965=>"101100000",
  39966=>"100101000",
  39967=>"100000101",
  39968=>"000100001",
  39969=>"101011011",
  39970=>"100011110",
  39971=>"010110001",
  39972=>"111101100",
  39973=>"111100001",
  39974=>"001000101",
  39975=>"001100100",
  39976=>"011001000",
  39977=>"001100111",
  39978=>"111010010",
  39979=>"001110001",
  39980=>"000111001",
  39981=>"001011100",
  39982=>"111000001",
  39983=>"100111110",
  39984=>"001001101",
  39985=>"010001011",
  39986=>"011000000",
  39987=>"010000011",
  39988=>"100001100",
  39989=>"000000000",
  39990=>"111011000",
  39991=>"000001111",
  39992=>"010010001",
  39993=>"100000011",
  39994=>"110011111",
  39995=>"010000010",
  39996=>"100111110",
  39997=>"111111110",
  39998=>"000101011",
  39999=>"001111101",
  40000=>"110111111",
  40001=>"001100000",
  40002=>"100010001",
  40003=>"000110011",
  40004=>"000000001",
  40005=>"000110000",
  40006=>"011011111",
  40007=>"110010000",
  40008=>"110100010",
  40009=>"011000111",
  40010=>"100111000",
  40011=>"001000110",
  40012=>"000110011",
  40013=>"110000001",
  40014=>"001110001",
  40015=>"101111000",
  40016=>"110001011",
  40017=>"000110100",
  40018=>"011101100",
  40019=>"001110110",
  40020=>"101110110",
  40021=>"001000110",
  40022=>"100111001",
  40023=>"110001111",
  40024=>"000110011",
  40025=>"011101101",
  40026=>"011001100",
  40027=>"000000100",
  40028=>"100011100",
  40029=>"100001011",
  40030=>"100011011",
  40031=>"100101010",
  40032=>"110001010",
  40033=>"000000001",
  40034=>"100101100",
  40035=>"000100011",
  40036=>"110001001",
  40037=>"111110001",
  40038=>"001000100",
  40039=>"001101001",
  40040=>"110101110",
  40041=>"000101000",
  40042=>"101101111",
  40043=>"000001010",
  40044=>"010110100",
  40045=>"001111111",
  40046=>"001011011",
  40047=>"010001110",
  40048=>"000011011",
  40049=>"100011100",
  40050=>"001011101",
  40051=>"001111111",
  40052=>"011000011",
  40053=>"111000110",
  40054=>"100110000",
  40055=>"100011111",
  40056=>"000111110",
  40057=>"011011101",
  40058=>"000100101",
  40059=>"011011111",
  40060=>"111101111",
  40061=>"101010000",
  40062=>"000000010",
  40063=>"101011001",
  40064=>"000010011",
  40065=>"010000011",
  40066=>"011011101",
  40067=>"000100011",
  40068=>"010000100",
  40069=>"011011110",
  40070=>"000011010",
  40071=>"011111001",
  40072=>"010000101",
  40073=>"110100101",
  40074=>"000010001",
  40075=>"111011011",
  40076=>"111011101",
  40077=>"110000110",
  40078=>"101001001",
  40079=>"111000001",
  40080=>"001111000",
  40081=>"000100111",
  40082=>"110001110",
  40083=>"011111110",
  40084=>"111000000",
  40085=>"101010001",
  40086=>"010011111",
  40087=>"010110111",
  40088=>"000110010",
  40089=>"100010010",
  40090=>"000010111",
  40091=>"001010001",
  40092=>"101110011",
  40093=>"011111011",
  40094=>"111101000",
  40095=>"100110010",
  40096=>"000110000",
  40097=>"010011001",
  40098=>"110111010",
  40099=>"001110100",
  40100=>"010000001",
  40101=>"100100011",
  40102=>"011101100",
  40103=>"111011111",
  40104=>"101000010",
  40105=>"100010101",
  40106=>"101001100",
  40107=>"010100110",
  40108=>"001100001",
  40109=>"000000100",
  40110=>"011100000",
  40111=>"100110100",
  40112=>"111010100",
  40113=>"100010101",
  40114=>"011100111",
  40115=>"000101111",
  40116=>"001011100",
  40117=>"100010000",
  40118=>"000011010",
  40119=>"100010100",
  40120=>"110010100",
  40121=>"010101000",
  40122=>"000001010",
  40123=>"111101000",
  40124=>"111100011",
  40125=>"010011101",
  40126=>"010011100",
  40127=>"001000000",
  40128=>"100010100",
  40129=>"001011110",
  40130=>"101001111",
  40131=>"101010100",
  40132=>"000110011",
  40133=>"010001110",
  40134=>"000100110",
  40135=>"010001010",
  40136=>"111110101",
  40137=>"010111011",
  40138=>"011110001",
  40139=>"110011101",
  40140=>"010101001",
  40141=>"111100000",
  40142=>"100100011",
  40143=>"000001001",
  40144=>"100000011",
  40145=>"111000000",
  40146=>"001000010",
  40147=>"101101001",
  40148=>"001001001",
  40149=>"010100000",
  40150=>"111100001",
  40151=>"011000110",
  40152=>"101110111",
  40153=>"100011000",
  40154=>"110010001",
  40155=>"001111001",
  40156=>"110001010",
  40157=>"011010110",
  40158=>"110100011",
  40159=>"001011111",
  40160=>"011011100",
  40161=>"011101101",
  40162=>"100001001",
  40163=>"110010000",
  40164=>"110101110",
  40165=>"010001111",
  40166=>"000000010",
  40167=>"010111111",
  40168=>"101110011",
  40169=>"111100000",
  40170=>"001001110",
  40171=>"111010011",
  40172=>"101110110",
  40173=>"110000001",
  40174=>"100001011",
  40175=>"011001111",
  40176=>"000001000",
  40177=>"111001110",
  40178=>"111001101",
  40179=>"011100100",
  40180=>"101100011",
  40181=>"010001011",
  40182=>"111011000",
  40183=>"011100101",
  40184=>"000000111",
  40185=>"011000001",
  40186=>"110001110",
  40187=>"110010000",
  40188=>"011010011",
  40189=>"011011011",
  40190=>"011000010",
  40191=>"010010111",
  40192=>"010111010",
  40193=>"111010001",
  40194=>"011011000",
  40195=>"010010001",
  40196=>"111001001",
  40197=>"001000010",
  40198=>"000010110",
  40199=>"111010111",
  40200=>"111001100",
  40201=>"000000001",
  40202=>"111101000",
  40203=>"100000101",
  40204=>"001100111",
  40205=>"001010110",
  40206=>"001101010",
  40207=>"000010111",
  40208=>"100100110",
  40209=>"010000101",
  40210=>"100111011",
  40211=>"100110111",
  40212=>"110010000",
  40213=>"000001000",
  40214=>"001001110",
  40215=>"110101101",
  40216=>"100011011",
  40217=>"001000110",
  40218=>"111000010",
  40219=>"011110011",
  40220=>"001011100",
  40221=>"111110111",
  40222=>"101101001",
  40223=>"000000111",
  40224=>"101001101",
  40225=>"110110000",
  40226=>"011011000",
  40227=>"001110111",
  40228=>"110001111",
  40229=>"000101011",
  40230=>"110111110",
  40231=>"000100101",
  40232=>"101101111",
  40233=>"111010111",
  40234=>"000111010",
  40235=>"111000000",
  40236=>"100110010",
  40237=>"110001110",
  40238=>"111101111",
  40239=>"001100001",
  40240=>"010110010",
  40241=>"100010100",
  40242=>"101010011",
  40243=>"001100001",
  40244=>"101101110",
  40245=>"001000000",
  40246=>"111111010",
  40247=>"100110111",
  40248=>"010110001",
  40249=>"010001001",
  40250=>"110100100",
  40251=>"011101111",
  40252=>"110000111",
  40253=>"011110100",
  40254=>"011001011",
  40255=>"010110011",
  40256=>"001001001",
  40257=>"010100110",
  40258=>"010110110",
  40259=>"111001000",
  40260=>"010110110",
  40261=>"000000111",
  40262=>"010100100",
  40263=>"100101110",
  40264=>"010110100",
  40265=>"110101010",
  40266=>"010101111",
  40267=>"010100000",
  40268=>"000100110",
  40269=>"100010010",
  40270=>"000100000",
  40271=>"101000100",
  40272=>"100000101",
  40273=>"111000010",
  40274=>"001011011",
  40275=>"000001011",
  40276=>"110100000",
  40277=>"010110000",
  40278=>"000001010",
  40279=>"001010000",
  40280=>"000100001",
  40281=>"111110011",
  40282=>"110110110",
  40283=>"100011110",
  40284=>"100110111",
  40285=>"000011111",
  40286=>"101101001",
  40287=>"101101110",
  40288=>"011001010",
  40289=>"101010010",
  40290=>"011100100",
  40291=>"010001010",
  40292=>"111011011",
  40293=>"000100111",
  40294=>"101010001",
  40295=>"111111111",
  40296=>"101011111",
  40297=>"101010100",
  40298=>"010001100",
  40299=>"110000010",
  40300=>"001101111",
  40301=>"001011111",
  40302=>"001100011",
  40303=>"100001101",
  40304=>"100001001",
  40305=>"111000110",
  40306=>"010000111",
  40307=>"011101110",
  40308=>"010000100",
  40309=>"101011110",
  40310=>"001101101",
  40311=>"110101100",
  40312=>"010011000",
  40313=>"010011010",
  40314=>"101001111",
  40315=>"111111001",
  40316=>"101001111",
  40317=>"010101010",
  40318=>"100100010",
  40319=>"000100100",
  40320=>"001001111",
  40321=>"100001011",
  40322=>"101101101",
  40323=>"010001001",
  40324=>"101010111",
  40325=>"000010101",
  40326=>"101000100",
  40327=>"101011101",
  40328=>"111111000",
  40329=>"000100110",
  40330=>"110000000",
  40331=>"000100111",
  40332=>"000100110",
  40333=>"000101100",
  40334=>"110101000",
  40335=>"110001110",
  40336=>"110000110",
  40337=>"001011010",
  40338=>"110111100",
  40339=>"001101100",
  40340=>"011001010",
  40341=>"110110011",
  40342=>"001000110",
  40343=>"101100111",
  40344=>"001111011",
  40345=>"011110110",
  40346=>"111010110",
  40347=>"000011011",
  40348=>"110110010",
  40349=>"000111011",
  40350=>"100011110",
  40351=>"111011101",
  40352=>"100000000",
  40353=>"110100100",
  40354=>"001011011",
  40355=>"000100000",
  40356=>"110111101",
  40357=>"101110111",
  40358=>"101110000",
  40359=>"101100111",
  40360=>"101001001",
  40361=>"011010100",
  40362=>"100011100",
  40363=>"001101111",
  40364=>"100111001",
  40365=>"011100101",
  40366=>"100111101",
  40367=>"000001011",
  40368=>"011100001",
  40369=>"110110101",
  40370=>"100111101",
  40371=>"010010011",
  40372=>"111110100",
  40373=>"001010001",
  40374=>"001110000",
  40375=>"110111100",
  40376=>"111001001",
  40377=>"111011001",
  40378=>"011001100",
  40379=>"110010100",
  40380=>"000110000",
  40381=>"001110111",
  40382=>"101001101",
  40383=>"001000110",
  40384=>"000000000",
  40385=>"101010001",
  40386=>"001100000",
  40387=>"110110001",
  40388=>"011000111",
  40389=>"100101010",
  40390=>"000011011",
  40391=>"111010010",
  40392=>"011001011",
  40393=>"001010110",
  40394=>"000111101",
  40395=>"100011111",
  40396=>"001001001",
  40397=>"001111100",
  40398=>"010111100",
  40399=>"011001100",
  40400=>"001011100",
  40401=>"001111110",
  40402=>"010000000",
  40403=>"011111010",
  40404=>"000011001",
  40405=>"101010010",
  40406=>"101010101",
  40407=>"100001010",
  40408=>"111111010",
  40409=>"110110111",
  40410=>"111111010",
  40411=>"111001110",
  40412=>"110101000",
  40413=>"110010001",
  40414=>"001000010",
  40415=>"101110001",
  40416=>"010110101",
  40417=>"000101010",
  40418=>"110111011",
  40419=>"010011101",
  40420=>"101000100",
  40421=>"110100001",
  40422=>"000110100",
  40423=>"110011001",
  40424=>"010110000",
  40425=>"001001101",
  40426=>"010001010",
  40427=>"001001010",
  40428=>"000101000",
  40429=>"000000010",
  40430=>"100100011",
  40431=>"100110010",
  40432=>"000011111",
  40433=>"000110111",
  40434=>"110011000",
  40435=>"110100110",
  40436=>"001010101",
  40437=>"001011000",
  40438=>"111011100",
  40439=>"010001111",
  40440=>"010110000",
  40441=>"111000101",
  40442=>"000110010",
  40443=>"110011110",
  40444=>"101001101",
  40445=>"011101000",
  40446=>"000011001",
  40447=>"111101110",
  40448=>"010010110",
  40449=>"111011000",
  40450=>"011000101",
  40451=>"101101000",
  40452=>"110100100",
  40453=>"001100001",
  40454=>"100100101",
  40455=>"000111011",
  40456=>"101110001",
  40457=>"100001011",
  40458=>"101110100",
  40459=>"001000101",
  40460=>"010101011",
  40461=>"110111100",
  40462=>"111110100",
  40463=>"000000000",
  40464=>"101111000",
  40465=>"011010010",
  40466=>"010110010",
  40467=>"000011010",
  40468=>"011101010",
  40469=>"110101111",
  40470=>"011010100",
  40471=>"010111010",
  40472=>"101011101",
  40473=>"000000111",
  40474=>"010101111",
  40475=>"101101110",
  40476=>"101000100",
  40477=>"100101001",
  40478=>"111110110",
  40479=>"001110100",
  40480=>"001100111",
  40481=>"111111010",
  40482=>"101101101",
  40483=>"100010000",
  40484=>"010101111",
  40485=>"100011110",
  40486=>"001011000",
  40487=>"100111100",
  40488=>"110010100",
  40489=>"111101111",
  40490=>"000110101",
  40491=>"000010000",
  40492=>"100110111",
  40493=>"000000001",
  40494=>"110100110",
  40495=>"000100000",
  40496=>"001010001",
  40497=>"101011001",
  40498=>"101110100",
  40499=>"010001000",
  40500=>"011001101",
  40501=>"011000101",
  40502=>"100010000",
  40503=>"011101101",
  40504=>"100000011",
  40505=>"000101111",
  40506=>"111010011",
  40507=>"011101000",
  40508=>"001000111",
  40509=>"011010000",
  40510=>"110011011",
  40511=>"111000010",
  40512=>"001100010",
  40513=>"001011101",
  40514=>"000000000",
  40515=>"000110001",
  40516=>"010011100",
  40517=>"101101011",
  40518=>"010100100",
  40519=>"000110000",
  40520=>"101001000",
  40521=>"101101101",
  40522=>"010000110",
  40523=>"110111110",
  40524=>"010100011",
  40525=>"011011011",
  40526=>"001010010",
  40527=>"101000010",
  40528=>"100001100",
  40529=>"111011101",
  40530=>"001001011",
  40531=>"010011100",
  40532=>"010001011",
  40533=>"000100111",
  40534=>"100100001",
  40535=>"111101000",
  40536=>"010110110",
  40537=>"001101000",
  40538=>"001011011",
  40539=>"111010010",
  40540=>"101101110",
  40541=>"110100000",
  40542=>"000101111",
  40543=>"000101000",
  40544=>"110011110",
  40545=>"000010011",
  40546=>"000010100",
  40547=>"000101100",
  40548=>"110101000",
  40549=>"110001000",
  40550=>"111001111",
  40551=>"001000010",
  40552=>"000000010",
  40553=>"111111011",
  40554=>"101111110",
  40555=>"001011100",
  40556=>"000000011",
  40557=>"111011101",
  40558=>"010001001",
  40559=>"101011101",
  40560=>"100110001",
  40561=>"001001101",
  40562=>"110101010",
  40563=>"100101010",
  40564=>"001000111",
  40565=>"110010101",
  40566=>"111111100",
  40567=>"000010000",
  40568=>"010110010",
  40569=>"010001100",
  40570=>"111111001",
  40571=>"111010011",
  40572=>"101111011",
  40573=>"010001100",
  40574=>"000010010",
  40575=>"100100001",
  40576=>"001001011",
  40577=>"000101010",
  40578=>"010100000",
  40579=>"011010011",
  40580=>"000000011",
  40581=>"100110111",
  40582=>"110001111",
  40583=>"011111111",
  40584=>"001100000",
  40585=>"101011110",
  40586=>"001001110",
  40587=>"001000000",
  40588=>"111111101",
  40589=>"111110110",
  40590=>"010011000",
  40591=>"011101001",
  40592=>"011100000",
  40593=>"001100110",
  40594=>"110000111",
  40595=>"111111010",
  40596=>"101001110",
  40597=>"110111010",
  40598=>"011001010",
  40599=>"100011001",
  40600=>"010111100",
  40601=>"000011010",
  40602=>"010110000",
  40603=>"100011111",
  40604=>"000111101",
  40605=>"111100110",
  40606=>"000000011",
  40607=>"001000101",
  40608=>"100100010",
  40609=>"010110011",
  40610=>"110001000",
  40611=>"111000110",
  40612=>"110001010",
  40613=>"101000111",
  40614=>"001010101",
  40615=>"011000011",
  40616=>"011100000",
  40617=>"100110111",
  40618=>"011010010",
  40619=>"100110000",
  40620=>"001101101",
  40621=>"001000011",
  40622=>"101000010",
  40623=>"001111010",
  40624=>"111010100",
  40625=>"100100100",
  40626=>"110011110",
  40627=>"011101100",
  40628=>"100011011",
  40629=>"101001101",
  40630=>"001011000",
  40631=>"101011011",
  40632=>"100010000",
  40633=>"111011000",
  40634=>"011111011",
  40635=>"110010000",
  40636=>"110001011",
  40637=>"101001011",
  40638=>"110110011",
  40639=>"001100011",
  40640=>"010111111",
  40641=>"000000110",
  40642=>"010000100",
  40643=>"000111101",
  40644=>"000101110",
  40645=>"111001100",
  40646=>"011110100",
  40647=>"011111010",
  40648=>"110100111",
  40649=>"100011100",
  40650=>"101001000",
  40651=>"001100111",
  40652=>"110111111",
  40653=>"001101010",
  40654=>"010101111",
  40655=>"000110011",
  40656=>"001100000",
  40657=>"011001111",
  40658=>"010110000",
  40659=>"011110101",
  40660=>"010001001",
  40661=>"101000100",
  40662=>"000100110",
  40663=>"111001001",
  40664=>"010100011",
  40665=>"111000110",
  40666=>"000001000",
  40667=>"011110110",
  40668=>"010000110",
  40669=>"000100100",
  40670=>"110111011",
  40671=>"001111000",
  40672=>"010101111",
  40673=>"000100100",
  40674=>"101110110",
  40675=>"010110010",
  40676=>"101101100",
  40677=>"000011100",
  40678=>"011000110",
  40679=>"111010111",
  40680=>"111101011",
  40681=>"110011101",
  40682=>"110110011",
  40683=>"011110111",
  40684=>"110011110",
  40685=>"110001111",
  40686=>"000011111",
  40687=>"000010001",
  40688=>"011000110",
  40689=>"000011010",
  40690=>"011100000",
  40691=>"011110000",
  40692=>"110111011",
  40693=>"001100000",
  40694=>"101101010",
  40695=>"001011110",
  40696=>"111010100",
  40697=>"010101101",
  40698=>"001001001",
  40699=>"010000100",
  40700=>"101000101",
  40701=>"010111001",
  40702=>"001010101",
  40703=>"101010000",
  40704=>"001010000",
  40705=>"111011001",
  40706=>"100100010",
  40707=>"000011101",
  40708=>"000000001",
  40709=>"110111101",
  40710=>"000011001",
  40711=>"001000011",
  40712=>"100000111",
  40713=>"101110111",
  40714=>"100011110",
  40715=>"101010110",
  40716=>"101010001",
  40717=>"100111100",
  40718=>"010010100",
  40719=>"000101001",
  40720=>"110011000",
  40721=>"001011000",
  40722=>"100111111",
  40723=>"000011011",
  40724=>"111011011",
  40725=>"110000101",
  40726=>"010000001",
  40727=>"011111110",
  40728=>"010011010",
  40729=>"001010111",
  40730=>"100111111",
  40731=>"001010011",
  40732=>"011001000",
  40733=>"110011110",
  40734=>"001110111",
  40735=>"111111011",
  40736=>"110000011",
  40737=>"101100110",
  40738=>"101111001",
  40739=>"100101001",
  40740=>"000010110",
  40741=>"101000011",
  40742=>"100000101",
  40743=>"001000101",
  40744=>"101111110",
  40745=>"110110101",
  40746=>"000011110",
  40747=>"110101000",
  40748=>"010010101",
  40749=>"100110111",
  40750=>"111110001",
  40751=>"101111000",
  40752=>"011010001",
  40753=>"101111010",
  40754=>"111101101",
  40755=>"001100110",
  40756=>"110010001",
  40757=>"100100010",
  40758=>"000111001",
  40759=>"110100111",
  40760=>"101110010",
  40761=>"100010110",
  40762=>"010110001",
  40763=>"001101101",
  40764=>"111000001",
  40765=>"100100000",
  40766=>"111011110",
  40767=>"110100111",
  40768=>"100110011",
  40769=>"100111001",
  40770=>"101010111",
  40771=>"100000110",
  40772=>"100110100",
  40773=>"000001111",
  40774=>"100010001",
  40775=>"111001001",
  40776=>"001111111",
  40777=>"010110110",
  40778=>"000100111",
  40779=>"000100110",
  40780=>"000101010",
  40781=>"010100001",
  40782=>"010100111",
  40783=>"010010010",
  40784=>"010010111",
  40785=>"100100100",
  40786=>"010101111",
  40787=>"000100011",
  40788=>"101111000",
  40789=>"000100110",
  40790=>"010110010",
  40791=>"111101001",
  40792=>"010110100",
  40793=>"110000000",
  40794=>"001101010",
  40795=>"000110111",
  40796=>"111011111",
  40797=>"111101010",
  40798=>"101101000",
  40799=>"000001000",
  40800=>"110001100",
  40801=>"111110111",
  40802=>"111010000",
  40803=>"011101110",
  40804=>"111111111",
  40805=>"100010001",
  40806=>"000001000",
  40807=>"110001110",
  40808=>"111000010",
  40809=>"010101011",
  40810=>"110011111",
  40811=>"001110111",
  40812=>"110000000",
  40813=>"101101100",
  40814=>"011000000",
  40815=>"010010010",
  40816=>"000010000",
  40817=>"100111110",
  40818=>"000011010",
  40819=>"100110000",
  40820=>"111100111",
  40821=>"111111111",
  40822=>"111001000",
  40823=>"111010110",
  40824=>"101101000",
  40825=>"100011011",
  40826=>"101000101",
  40827=>"101000010",
  40828=>"001100011",
  40829=>"101100101",
  40830=>"000100001",
  40831=>"101011011",
  40832=>"010010000",
  40833=>"111011000",
  40834=>"100001011",
  40835=>"100010111",
  40836=>"001111000",
  40837=>"010000001",
  40838=>"110101111",
  40839=>"010110111",
  40840=>"011111011",
  40841=>"001000110",
  40842=>"010111111",
  40843=>"010010011",
  40844=>"111000010",
  40845=>"101110000",
  40846=>"000101011",
  40847=>"010000000",
  40848=>"000001000",
  40849=>"100000001",
  40850=>"110001010",
  40851=>"100111111",
  40852=>"100100001",
  40853=>"000110001",
  40854=>"111011000",
  40855=>"001010000",
  40856=>"100111111",
  40857=>"010010111",
  40858=>"101000111",
  40859=>"110010000",
  40860=>"101001100",
  40861=>"101111110",
  40862=>"111011010",
  40863=>"110011101",
  40864=>"100100110",
  40865=>"111101010",
  40866=>"000100001",
  40867=>"101011011",
  40868=>"111100000",
  40869=>"011101011",
  40870=>"111001010",
  40871=>"100111001",
  40872=>"110001000",
  40873=>"111000110",
  40874=>"011010011",
  40875=>"110100100",
  40876=>"111100010",
  40877=>"000111111",
  40878=>"101001110",
  40879=>"111001000",
  40880=>"001100110",
  40881=>"100001000",
  40882=>"100111100",
  40883=>"000000000",
  40884=>"101100010",
  40885=>"111111000",
  40886=>"100001010",
  40887=>"101111011",
  40888=>"010010001",
  40889=>"111000110",
  40890=>"000010100",
  40891=>"111101010",
  40892=>"011000111",
  40893=>"100000010",
  40894=>"010111101",
  40895=>"000110010",
  40896=>"110101110",
  40897=>"011001110",
  40898=>"100000111",
  40899=>"100100110",
  40900=>"000010000",
  40901=>"011000000",
  40902=>"100100011",
  40903=>"000100011",
  40904=>"000100110",
  40905=>"101110011",
  40906=>"010000111",
  40907=>"111110111",
  40908=>"010100100",
  40909=>"111000101",
  40910=>"001011101",
  40911=>"001000001",
  40912=>"111010110",
  40913=>"111011001",
  40914=>"110101110",
  40915=>"000100000",
  40916=>"000011101",
  40917=>"101011011",
  40918=>"100001101",
  40919=>"111011100",
  40920=>"100011011",
  40921=>"100101111",
  40922=>"001000111",
  40923=>"100000111",
  40924=>"011001111",
  40925=>"110001100",
  40926=>"101111111",
  40927=>"111100011",
  40928=>"000000100",
  40929=>"010010000",
  40930=>"000101110",
  40931=>"111010110",
  40932=>"100010100",
  40933=>"001000000",
  40934=>"011111101",
  40935=>"010011111",
  40936=>"111100111",
  40937=>"100110111",
  40938=>"001000110",
  40939=>"010011110",
  40940=>"101000101",
  40941=>"110000001",
  40942=>"100011111",
  40943=>"110001111",
  40944=>"011101010",
  40945=>"011011010",
  40946=>"100001000",
  40947=>"100101001",
  40948=>"000110001",
  40949=>"101111001",
  40950=>"000000000",
  40951=>"011010101",
  40952=>"011100100",
  40953=>"100001110",
  40954=>"101001111",
  40955=>"100100100",
  40956=>"010000010",
  40957=>"000000101",
  40958=>"100101100",
  40959=>"100000001",
  40960=>"111010000",
  40961=>"101011110",
  40962=>"000000101",
  40963=>"010111001",
  40964=>"100100010",
  40965=>"000001110",
  40966=>"000111101",
  40967=>"111011001",
  40968=>"000000011",
  40969=>"000011100",
  40970=>"111001000",
  40971=>"000111110",
  40972=>"110010001",
  40973=>"101111101",
  40974=>"000001000",
  40975=>"010001001",
  40976=>"111100001",
  40977=>"001010010",
  40978=>"100000110",
  40979=>"001011000",
  40980=>"001011110",
  40981=>"110011100",
  40982=>"010000010",
  40983=>"111010100",
  40984=>"111011000",
  40985=>"100001011",
  40986=>"110010100",
  40987=>"110110010",
  40988=>"111011101",
  40989=>"011000100",
  40990=>"100010001",
  40991=>"111101001",
  40992=>"101100000",
  40993=>"000000100",
  40994=>"110101010",
  40995=>"101001111",
  40996=>"110100010",
  40997=>"101110000",
  40998=>"110001101",
  40999=>"010000000",
  41000=>"101000111",
  41001=>"110011001",
  41002=>"111001010",
  41003=>"100010101",
  41004=>"011011011",
  41005=>"010101110",
  41006=>"001001101",
  41007=>"101101100",
  41008=>"110011001",
  41009=>"101110110",
  41010=>"111111110",
  41011=>"000011101",
  41012=>"110000100",
  41013=>"110101010",
  41014=>"111111111",
  41015=>"000000000",
  41016=>"001010011",
  41017=>"001011010",
  41018=>"000110001",
  41019=>"000110010",
  41020=>"000000100",
  41021=>"011010001",
  41022=>"000011000",
  41023=>"000110101",
  41024=>"010001000",
  41025=>"001000000",
  41026=>"011000110",
  41027=>"010101100",
  41028=>"111011000",
  41029=>"111010100",
  41030=>"111000011",
  41031=>"010001101",
  41032=>"111100101",
  41033=>"111111011",
  41034=>"001100101",
  41035=>"101011111",
  41036=>"001000010",
  41037=>"110100000",
  41038=>"111011010",
  41039=>"110001101",
  41040=>"101100001",
  41041=>"001101100",
  41042=>"010101001",
  41043=>"100111011",
  41044=>"010000101",
  41045=>"010101101",
  41046=>"101100111",
  41047=>"110100000",
  41048=>"101100101",
  41049=>"101100111",
  41050=>"110000011",
  41051=>"000100000",
  41052=>"100001011",
  41053=>"101010101",
  41054=>"100010000",
  41055=>"100111000",
  41056=>"010011111",
  41057=>"100111101",
  41058=>"010110110",
  41059=>"001001100",
  41060=>"000101011",
  41061=>"101111100",
  41062=>"000100111",
  41063=>"010100111",
  41064=>"100001110",
  41065=>"111100010",
  41066=>"011011001",
  41067=>"100001001",
  41068=>"000001110",
  41069=>"101000010",
  41070=>"101010101",
  41071=>"000010101",
  41072=>"010010010",
  41073=>"111011011",
  41074=>"111001000",
  41075=>"100000110",
  41076=>"000100000",
  41077=>"100011000",
  41078=>"101101010",
  41079=>"011101011",
  41080=>"110111101",
  41081=>"100000010",
  41082=>"001100010",
  41083=>"100101000",
  41084=>"000101001",
  41085=>"011011001",
  41086=>"000000011",
  41087=>"101000110",
  41088=>"011110000",
  41089=>"001000100",
  41090=>"010100001",
  41091=>"100010100",
  41092=>"000010010",
  41093=>"011110111",
  41094=>"001011111",
  41095=>"111011100",
  41096=>"010110110",
  41097=>"001101101",
  41098=>"100100101",
  41099=>"111101001",
  41100=>"010010011",
  41101=>"100100000",
  41102=>"010100110",
  41103=>"010000010",
  41104=>"011100100",
  41105=>"000010110",
  41106=>"101001011",
  41107=>"110111110",
  41108=>"110111000",
  41109=>"000111111",
  41110=>"100111101",
  41111=>"011100000",
  41112=>"111101011",
  41113=>"100111000",
  41114=>"011101100",
  41115=>"110110010",
  41116=>"011011100",
  41117=>"110111010",
  41118=>"000001101",
  41119=>"110111101",
  41120=>"000000101",
  41121=>"111100001",
  41122=>"111110111",
  41123=>"000010101",
  41124=>"111111110",
  41125=>"110010111",
  41126=>"010001010",
  41127=>"000110100",
  41128=>"100111000",
  41129=>"010001100",
  41130=>"001010110",
  41131=>"111001111",
  41132=>"111101001",
  41133=>"001011010",
  41134=>"101110100",
  41135=>"011101111",
  41136=>"010110000",
  41137=>"000001000",
  41138=>"011011010",
  41139=>"101110100",
  41140=>"110011001",
  41141=>"001110100",
  41142=>"000001110",
  41143=>"000011000",
  41144=>"011101111",
  41145=>"000101111",
  41146=>"000010010",
  41147=>"001001001",
  41148=>"111001110",
  41149=>"101111110",
  41150=>"000100001",
  41151=>"001111100",
  41152=>"101110100",
  41153=>"100111100",
  41154=>"000000000",
  41155=>"010000110",
  41156=>"100010110",
  41157=>"111101101",
  41158=>"111011111",
  41159=>"010010110",
  41160=>"110111101",
  41161=>"111011100",
  41162=>"110111000",
  41163=>"101110100",
  41164=>"000000110",
  41165=>"100011011",
  41166=>"101011101",
  41167=>"001011100",
  41168=>"000011011",
  41169=>"000100100",
  41170=>"010101000",
  41171=>"000101100",
  41172=>"010010000",
  41173=>"001001001",
  41174=>"000011101",
  41175=>"000110010",
  41176=>"101101010",
  41177=>"101101000",
  41178=>"101100000",
  41179=>"011110001",
  41180=>"011011001",
  41181=>"001001000",
  41182=>"011100110",
  41183=>"100101110",
  41184=>"010111000",
  41185=>"111000101",
  41186=>"001001101",
  41187=>"000000001",
  41188=>"100000001",
  41189=>"001000110",
  41190=>"000011110",
  41191=>"000000111",
  41192=>"000101010",
  41193=>"001110001",
  41194=>"011100111",
  41195=>"001000011",
  41196=>"001000000",
  41197=>"000010101",
  41198=>"111001000",
  41199=>"010110101",
  41200=>"101111110",
  41201=>"100010111",
  41202=>"011001000",
  41203=>"110010011",
  41204=>"111001110",
  41205=>"101000011",
  41206=>"110110111",
  41207=>"001110001",
  41208=>"110111101",
  41209=>"001111000",
  41210=>"000100100",
  41211=>"010101000",
  41212=>"101101000",
  41213=>"101000000",
  41214=>"010110110",
  41215=>"100101111",
  41216=>"001100101",
  41217=>"101000100",
  41218=>"110000000",
  41219=>"110001001",
  41220=>"010010110",
  41221=>"000101000",
  41222=>"001000000",
  41223=>"111001100",
  41224=>"100010001",
  41225=>"001010010",
  41226=>"101010101",
  41227=>"001000010",
  41228=>"111000110",
  41229=>"010001100",
  41230=>"101000011",
  41231=>"000100010",
  41232=>"111111011",
  41233=>"000000001",
  41234=>"010000110",
  41235=>"011101100",
  41236=>"001010110",
  41237=>"101001011",
  41238=>"001000000",
  41239=>"101100111",
  41240=>"011000011",
  41241=>"010100110",
  41242=>"111010011",
  41243=>"011001010",
  41244=>"001101001",
  41245=>"010010111",
  41246=>"100101010",
  41247=>"110000111",
  41248=>"011000100",
  41249=>"101000110",
  41250=>"010111111",
  41251=>"111001011",
  41252=>"001110100",
  41253=>"110001011",
  41254=>"000011000",
  41255=>"100000001",
  41256=>"010100110",
  41257=>"100011011",
  41258=>"101111110",
  41259=>"011000101",
  41260=>"101011000",
  41261=>"000000010",
  41262=>"001000000",
  41263=>"111101011",
  41264=>"011001111",
  41265=>"001101101",
  41266=>"111100011",
  41267=>"100100110",
  41268=>"010101100",
  41269=>"010100000",
  41270=>"000100110",
  41271=>"011010111",
  41272=>"101011110",
  41273=>"110000011",
  41274=>"110010000",
  41275=>"110011010",
  41276=>"111111011",
  41277=>"111111101",
  41278=>"100001000",
  41279=>"110101100",
  41280=>"101000011",
  41281=>"101101100",
  41282=>"001111010",
  41283=>"100001101",
  41284=>"011010100",
  41285=>"110101010",
  41286=>"011010001",
  41287=>"110101110",
  41288=>"100111010",
  41289=>"111001010",
  41290=>"011011001",
  41291=>"111101001",
  41292=>"010000110",
  41293=>"111111011",
  41294=>"100011010",
  41295=>"101101101",
  41296=>"001111100",
  41297=>"110000110",
  41298=>"110010100",
  41299=>"001000100",
  41300=>"111100110",
  41301=>"011001000",
  41302=>"100110011",
  41303=>"101101000",
  41304=>"000100001",
  41305=>"010000001",
  41306=>"100010010",
  41307=>"100010011",
  41308=>"100100100",
  41309=>"011011110",
  41310=>"100100000",
  41311=>"000010001",
  41312=>"000110011",
  41313=>"110101101",
  41314=>"001011011",
  41315=>"010100011",
  41316=>"110011100",
  41317=>"110001110",
  41318=>"101001101",
  41319=>"110101000",
  41320=>"001101111",
  41321=>"010010001",
  41322=>"010011111",
  41323=>"100011110",
  41324=>"001111100",
  41325=>"000111010",
  41326=>"100101101",
  41327=>"110110010",
  41328=>"011011011",
  41329=>"011111110",
  41330=>"110000010",
  41331=>"101000111",
  41332=>"101101110",
  41333=>"111111011",
  41334=>"010011010",
  41335=>"011000111",
  41336=>"111100101",
  41337=>"110011001",
  41338=>"111110011",
  41339=>"010101110",
  41340=>"011111110",
  41341=>"111011110",
  41342=>"110001111",
  41343=>"111010110",
  41344=>"001010011",
  41345=>"111011001",
  41346=>"001010110",
  41347=>"000011000",
  41348=>"100000111",
  41349=>"100000011",
  41350=>"001101010",
  41351=>"111000010",
  41352=>"000000010",
  41353=>"011010100",
  41354=>"010101000",
  41355=>"111001001",
  41356=>"000111111",
  41357=>"111001011",
  41358=>"000111011",
  41359=>"001100111",
  41360=>"000110100",
  41361=>"001001101",
  41362=>"011011101",
  41363=>"001101101",
  41364=>"111000101",
  41365=>"111111010",
  41366=>"000100000",
  41367=>"100100001",
  41368=>"000000011",
  41369=>"000000011",
  41370=>"110100111",
  41371=>"011100100",
  41372=>"011001010",
  41373=>"001010000",
  41374=>"101011000",
  41375=>"001000001",
  41376=>"010010010",
  41377=>"100010011",
  41378=>"101001010",
  41379=>"111001000",
  41380=>"011000111",
  41381=>"111001100",
  41382=>"111101011",
  41383=>"100100110",
  41384=>"111111110",
  41385=>"001100011",
  41386=>"000111011",
  41387=>"101010101",
  41388=>"000000011",
  41389=>"101001000",
  41390=>"000110111",
  41391=>"010000110",
  41392=>"100000110",
  41393=>"100000000",
  41394=>"010010110",
  41395=>"110000001",
  41396=>"100011000",
  41397=>"101011101",
  41398=>"110011010",
  41399=>"010101001",
  41400=>"011011001",
  41401=>"111010010",
  41402=>"101001101",
  41403=>"100000010",
  41404=>"100100000",
  41405=>"111111110",
  41406=>"010001110",
  41407=>"101110000",
  41408=>"110111011",
  41409=>"001001101",
  41410=>"011001001",
  41411=>"000001111",
  41412=>"001001110",
  41413=>"100101000",
  41414=>"110001111",
  41415=>"000000101",
  41416=>"011011100",
  41417=>"010110000",
  41418=>"011011100",
  41419=>"000000110",
  41420=>"111000100",
  41421=>"100001111",
  41422=>"000011100",
  41423=>"000001000",
  41424=>"110111010",
  41425=>"011000001",
  41426=>"001001110",
  41427=>"111100000",
  41428=>"001100001",
  41429=>"000101001",
  41430=>"001110111",
  41431=>"010000001",
  41432=>"100100011",
  41433=>"001011101",
  41434=>"010000011",
  41435=>"111010100",
  41436=>"100100111",
  41437=>"111111110",
  41438=>"001111111",
  41439=>"011101100",
  41440=>"110101110",
  41441=>"111101100",
  41442=>"010110101",
  41443=>"011111110",
  41444=>"010011000",
  41445=>"000010001",
  41446=>"110110000",
  41447=>"001011101",
  41448=>"111111111",
  41449=>"101100110",
  41450=>"001010010",
  41451=>"110001100",
  41452=>"100001111",
  41453=>"111011111",
  41454=>"110100100",
  41455=>"101001001",
  41456=>"011010111",
  41457=>"101000010",
  41458=>"111001111",
  41459=>"000000100",
  41460=>"001010100",
  41461=>"010011100",
  41462=>"100101110",
  41463=>"001001011",
  41464=>"110111110",
  41465=>"011001000",
  41466=>"111100011",
  41467=>"111011000",
  41468=>"001101010",
  41469=>"110000101",
  41470=>"011000111",
  41471=>"010000011",
  41472=>"001001100",
  41473=>"100100011",
  41474=>"100100110",
  41475=>"000001001",
  41476=>"111111010",
  41477=>"101110100",
  41478=>"110000011",
  41479=>"111101001",
  41480=>"010011010",
  41481=>"000100001",
  41482=>"010111100",
  41483=>"000000100",
  41484=>"001010010",
  41485=>"111001010",
  41486=>"010001110",
  41487=>"011000001",
  41488=>"001101101",
  41489=>"011111001",
  41490=>"111001110",
  41491=>"111101100",
  41492=>"011000100",
  41493=>"000000010",
  41494=>"011000100",
  41495=>"010000100",
  41496=>"011000110",
  41497=>"111011101",
  41498=>"110101111",
  41499=>"100001110",
  41500=>"001000000",
  41501=>"100100010",
  41502=>"011010011",
  41503=>"110001110",
  41504=>"101000000",
  41505=>"000110111",
  41506=>"110010111",
  41507=>"101001000",
  41508=>"111001110",
  41509=>"001001111",
  41510=>"010011111",
  41511=>"010000100",
  41512=>"110101111",
  41513=>"011110001",
  41514=>"110110011",
  41515=>"111001010",
  41516=>"011110110",
  41517=>"110111100",
  41518=>"101101100",
  41519=>"010011110",
  41520=>"001011011",
  41521=>"101010011",
  41522=>"101101110",
  41523=>"000100100",
  41524=>"001101101",
  41525=>"010100000",
  41526=>"101110111",
  41527=>"001101010",
  41528=>"111010011",
  41529=>"111101100",
  41530=>"110000010",
  41531=>"110101001",
  41532=>"110000100",
  41533=>"110010011",
  41534=>"000101101",
  41535=>"100000101",
  41536=>"001111001",
  41537=>"011000010",
  41538=>"010011001",
  41539=>"100100110",
  41540=>"010001000",
  41541=>"000000110",
  41542=>"000010000",
  41543=>"111100100",
  41544=>"101111000",
  41545=>"001010001",
  41546=>"000101111",
  41547=>"100001110",
  41548=>"001011010",
  41549=>"010001011",
  41550=>"111101001",
  41551=>"101000111",
  41552=>"110111010",
  41553=>"110111111",
  41554=>"111100010",
  41555=>"010101111",
  41556=>"110010011",
  41557=>"110010000",
  41558=>"011101101",
  41559=>"000100000",
  41560=>"001011111",
  41561=>"000001000",
  41562=>"010100000",
  41563=>"001000011",
  41564=>"110001000",
  41565=>"100100010",
  41566=>"100111000",
  41567=>"100011110",
  41568=>"111111000",
  41569=>"010100111",
  41570=>"101111110",
  41571=>"110001001",
  41572=>"000011000",
  41573=>"001011010",
  41574=>"100011010",
  41575=>"110011000",
  41576=>"001000000",
  41577=>"011110110",
  41578=>"101111000",
  41579=>"110001000",
  41580=>"101111110",
  41581=>"110001111",
  41582=>"011011100",
  41583=>"010110111",
  41584=>"101100000",
  41585=>"111001111",
  41586=>"101011011",
  41587=>"100010010",
  41588=>"110010111",
  41589=>"010111110",
  41590=>"111000011",
  41591=>"000110101",
  41592=>"011100101",
  41593=>"110011011",
  41594=>"110101111",
  41595=>"111100001",
  41596=>"001001000",
  41597=>"000010100",
  41598=>"011110000",
  41599=>"110000111",
  41600=>"101010000",
  41601=>"010111111",
  41602=>"111101010",
  41603=>"001000101",
  41604=>"111111011",
  41605=>"011111110",
  41606=>"001011011",
  41607=>"011010000",
  41608=>"111010010",
  41609=>"000000001",
  41610=>"100100001",
  41611=>"001100110",
  41612=>"010000000",
  41613=>"100000000",
  41614=>"000011100",
  41615=>"001010100",
  41616=>"110001111",
  41617=>"111100001",
  41618=>"100000101",
  41619=>"000111111",
  41620=>"000011110",
  41621=>"011111010",
  41622=>"000001001",
  41623=>"000101000",
  41624=>"101000001",
  41625=>"111111110",
  41626=>"001001001",
  41627=>"100001000",
  41628=>"011100110",
  41629=>"101110101",
  41630=>"100111010",
  41631=>"010110011",
  41632=>"010011001",
  41633=>"110011110",
  41634=>"111101010",
  41635=>"110100011",
  41636=>"010011010",
  41637=>"100101101",
  41638=>"100010111",
  41639=>"101101101",
  41640=>"100001011",
  41641=>"110101001",
  41642=>"010100111",
  41643=>"110001001",
  41644=>"101100101",
  41645=>"010000100",
  41646=>"011010010",
  41647=>"000101110",
  41648=>"100111111",
  41649=>"100011110",
  41650=>"111011111",
  41651=>"000010001",
  41652=>"111111100",
  41653=>"011111111",
  41654=>"100100110",
  41655=>"100110000",
  41656=>"000011001",
  41657=>"100100111",
  41658=>"100001011",
  41659=>"101110110",
  41660=>"101011001",
  41661=>"000000100",
  41662=>"000100001",
  41663=>"101111011",
  41664=>"100110000",
  41665=>"100001111",
  41666=>"011001100",
  41667=>"000001001",
  41668=>"001000110",
  41669=>"100110111",
  41670=>"001101100",
  41671=>"000011000",
  41672=>"001111101",
  41673=>"100001001",
  41674=>"100010110",
  41675=>"000110010",
  41676=>"011111010",
  41677=>"010010101",
  41678=>"111011000",
  41679=>"101010110",
  41680=>"000000001",
  41681=>"010010111",
  41682=>"101011110",
  41683=>"010111101",
  41684=>"100100100",
  41685=>"001111111",
  41686=>"011100000",
  41687=>"110011101",
  41688=>"100100100",
  41689=>"110100011",
  41690=>"111101110",
  41691=>"001111110",
  41692=>"000101101",
  41693=>"000100110",
  41694=>"010100000",
  41695=>"001000001",
  41696=>"000001101",
  41697=>"011101101",
  41698=>"100110100",
  41699=>"011001001",
  41700=>"001101000",
  41701=>"001000000",
  41702=>"000100010",
  41703=>"111001000",
  41704=>"011110010",
  41705=>"001001110",
  41706=>"000010101",
  41707=>"111011001",
  41708=>"000110001",
  41709=>"011111110",
  41710=>"010101110",
  41711=>"111101111",
  41712=>"100010100",
  41713=>"011010011",
  41714=>"000011111",
  41715=>"001010101",
  41716=>"111101111",
  41717=>"100101100",
  41718=>"100100011",
  41719=>"010011010",
  41720=>"101101110",
  41721=>"000101101",
  41722=>"000100101",
  41723=>"100100010",
  41724=>"000011101",
  41725=>"011010011",
  41726=>"011010011",
  41727=>"000101000",
  41728=>"001011011",
  41729=>"101011010",
  41730=>"001010100",
  41731=>"111110101",
  41732=>"101111011",
  41733=>"110101111",
  41734=>"111011001",
  41735=>"001001101",
  41736=>"111000101",
  41737=>"000000001",
  41738=>"101010100",
  41739=>"101010001",
  41740=>"100110000",
  41741=>"100101101",
  41742=>"001100010",
  41743=>"101111111",
  41744=>"000011001",
  41745=>"000111101",
  41746=>"111111011",
  41747=>"000000100",
  41748=>"101001100",
  41749=>"101010110",
  41750=>"101101110",
  41751=>"010100001",
  41752=>"011111001",
  41753=>"111100010",
  41754=>"010111010",
  41755=>"111100010",
  41756=>"000011110",
  41757=>"100010000",
  41758=>"011111011",
  41759=>"011001001",
  41760=>"001100000",
  41761=>"000010101",
  41762=>"110110001",
  41763=>"101111100",
  41764=>"111111101",
  41765=>"101110110",
  41766=>"110011000",
  41767=>"000011011",
  41768=>"001011000",
  41769=>"100110011",
  41770=>"111111101",
  41771=>"000111101",
  41772=>"011011010",
  41773=>"000000000",
  41774=>"110001101",
  41775=>"000110100",
  41776=>"000100000",
  41777=>"100000111",
  41778=>"001000101",
  41779=>"101101111",
  41780=>"001010110",
  41781=>"000111000",
  41782=>"001100100",
  41783=>"011010000",
  41784=>"010110100",
  41785=>"000010001",
  41786=>"001110110",
  41787=>"010100110",
  41788=>"010111000",
  41789=>"000011000",
  41790=>"010001110",
  41791=>"111101011",
  41792=>"000011000",
  41793=>"101000111",
  41794=>"000000010",
  41795=>"101100111",
  41796=>"000100110",
  41797=>"111001100",
  41798=>"111100110",
  41799=>"000010110",
  41800=>"100000110",
  41801=>"100100110",
  41802=>"110011111",
  41803=>"101001111",
  41804=>"101101101",
  41805=>"111101011",
  41806=>"000000111",
  41807=>"110101000",
  41808=>"110001000",
  41809=>"111000000",
  41810=>"100111001",
  41811=>"110011110",
  41812=>"100110100",
  41813=>"111001000",
  41814=>"100101100",
  41815=>"110110010",
  41816=>"000001100",
  41817=>"010101101",
  41818=>"001101110",
  41819=>"101101010",
  41820=>"100111010",
  41821=>"101110000",
  41822=>"000011011",
  41823=>"010000000",
  41824=>"011111111",
  41825=>"000100110",
  41826=>"010000000",
  41827=>"010000010",
  41828=>"001011001",
  41829=>"001011001",
  41830=>"110110000",
  41831=>"110010111",
  41832=>"111000001",
  41833=>"110101111",
  41834=>"100110101",
  41835=>"011011111",
  41836=>"100110000",
  41837=>"001010110",
  41838=>"000001110",
  41839=>"100110101",
  41840=>"110010000",
  41841=>"001000001",
  41842=>"000010100",
  41843=>"100100100",
  41844=>"000011010",
  41845=>"111111100",
  41846=>"101001110",
  41847=>"111001010",
  41848=>"001011111",
  41849=>"001100010",
  41850=>"000000101",
  41851=>"110010000",
  41852=>"000111001",
  41853=>"010101011",
  41854=>"001110000",
  41855=>"111111101",
  41856=>"001011110",
  41857=>"011110001",
  41858=>"010000111",
  41859=>"101000011",
  41860=>"000001001",
  41861=>"110110100",
  41862=>"100111101",
  41863=>"010010001",
  41864=>"011000100",
  41865=>"010010000",
  41866=>"111001110",
  41867=>"111100101",
  41868=>"011001101",
  41869=>"000000001",
  41870=>"000001100",
  41871=>"111010111",
  41872=>"101010101",
  41873=>"000001000",
  41874=>"010111100",
  41875=>"000111100",
  41876=>"011111011",
  41877=>"000011010",
  41878=>"110000010",
  41879=>"111000110",
  41880=>"001000001",
  41881=>"011000100",
  41882=>"110111011",
  41883=>"101100110",
  41884=>"111001100",
  41885=>"010111100",
  41886=>"111111100",
  41887=>"101001101",
  41888=>"010010101",
  41889=>"100110101",
  41890=>"111001000",
  41891=>"111100011",
  41892=>"010100000",
  41893=>"001111111",
  41894=>"001000111",
  41895=>"010001010",
  41896=>"101101010",
  41897=>"010111001",
  41898=>"001101011",
  41899=>"011101011",
  41900=>"101001001",
  41901=>"011001100",
  41902=>"001111101",
  41903=>"011011000",
  41904=>"100110000",
  41905=>"110001100",
  41906=>"011001100",
  41907=>"111011111",
  41908=>"010010110",
  41909=>"010110010",
  41910=>"111010111",
  41911=>"100011101",
  41912=>"110011111",
  41913=>"110000101",
  41914=>"010010100",
  41915=>"100010100",
  41916=>"010010001",
  41917=>"010000010",
  41918=>"111100100",
  41919=>"000010000",
  41920=>"000110010",
  41921=>"001010000",
  41922=>"100000110",
  41923=>"101010011",
  41924=>"001000010",
  41925=>"101010011",
  41926=>"000100111",
  41927=>"010001011",
  41928=>"010100010",
  41929=>"001100111",
  41930=>"000111001",
  41931=>"000110111",
  41932=>"111110110",
  41933=>"010110110",
  41934=>"100101110",
  41935=>"011000100",
  41936=>"101001010",
  41937=>"110110100",
  41938=>"000001101",
  41939=>"010000000",
  41940=>"100000001",
  41941=>"110000001",
  41942=>"100101110",
  41943=>"011000101",
  41944=>"101011011",
  41945=>"000000011",
  41946=>"011000001",
  41947=>"100000001",
  41948=>"001010000",
  41949=>"101101010",
  41950=>"010110001",
  41951=>"001010010",
  41952=>"100111011",
  41953=>"110000001",
  41954=>"001010000",
  41955=>"001111001",
  41956=>"110100011",
  41957=>"100111010",
  41958=>"110111101",
  41959=>"001000010",
  41960=>"001111000",
  41961=>"111000111",
  41962=>"100011111",
  41963=>"011110011",
  41964=>"001100101",
  41965=>"101110011",
  41966=>"111100111",
  41967=>"011001010",
  41968=>"101101001",
  41969=>"001011011",
  41970=>"000010110",
  41971=>"110111100",
  41972=>"110110010",
  41973=>"110100110",
  41974=>"001000100",
  41975=>"111101101",
  41976=>"001101111",
  41977=>"010001010",
  41978=>"100100010",
  41979=>"010100000",
  41980=>"111101011",
  41981=>"010001101",
  41982=>"011001101",
  41983=>"011011000",
  41984=>"011010001",
  41985=>"010000001",
  41986=>"111101110",
  41987=>"101110001",
  41988=>"111101001",
  41989=>"110000101",
  41990=>"110101100",
  41991=>"110101111",
  41992=>"000011110",
  41993=>"100011111",
  41994=>"001001110",
  41995=>"010000000",
  41996=>"010001011",
  41997=>"000101001",
  41998=>"011001101",
  41999=>"100000111",
  42000=>"000110000",
  42001=>"100110101",
  42002=>"001010101",
  42003=>"110000111",
  42004=>"010011111",
  42005=>"110010100",
  42006=>"000110001",
  42007=>"000000110",
  42008=>"000010001",
  42009=>"111101110",
  42010=>"010110011",
  42011=>"101110110",
  42012=>"110000110",
  42013=>"110000011",
  42014=>"001111101",
  42015=>"010011110",
  42016=>"011010110",
  42017=>"100011100",
  42018=>"000000000",
  42019=>"100001111",
  42020=>"001011101",
  42021=>"001011110",
  42022=>"011011011",
  42023=>"010100000",
  42024=>"010000010",
  42025=>"001001101",
  42026=>"111011111",
  42027=>"010000100",
  42028=>"011000000",
  42029=>"110111001",
  42030=>"111010100",
  42031=>"110001101",
  42032=>"111101101",
  42033=>"001001110",
  42034=>"001000001",
  42035=>"101100001",
  42036=>"101000110",
  42037=>"011110000",
  42038=>"101010110",
  42039=>"011011110",
  42040=>"010001101",
  42041=>"001001001",
  42042=>"001001011",
  42043=>"001000111",
  42044=>"011110010",
  42045=>"000001100",
  42046=>"111110000",
  42047=>"110110110",
  42048=>"110110010",
  42049=>"101100101",
  42050=>"000001001",
  42051=>"111001001",
  42052=>"000000000",
  42053=>"110001000",
  42054=>"110101001",
  42055=>"111110000",
  42056=>"001110110",
  42057=>"101110111",
  42058=>"110100100",
  42059=>"100000000",
  42060=>"001110111",
  42061=>"100100111",
  42062=>"001000011",
  42063=>"011011011",
  42064=>"000001111",
  42065=>"100101011",
  42066=>"001001101",
  42067=>"110010111",
  42068=>"010001110",
  42069=>"111101100",
  42070=>"001110100",
  42071=>"010101000",
  42072=>"011001101",
  42073=>"110101110",
  42074=>"111110110",
  42075=>"000000000",
  42076=>"001010010",
  42077=>"100001111",
  42078=>"110001111",
  42079=>"000100000",
  42080=>"110000101",
  42081=>"011111101",
  42082=>"011101110",
  42083=>"010010010",
  42084=>"100110001",
  42085=>"110111011",
  42086=>"001001110",
  42087=>"100010001",
  42088=>"010000110",
  42089=>"001000001",
  42090=>"010101010",
  42091=>"001010001",
  42092=>"101110111",
  42093=>"111110011",
  42094=>"101000100",
  42095=>"011101001",
  42096=>"110010101",
  42097=>"111000000",
  42098=>"101010111",
  42099=>"010111101",
  42100=>"001000011",
  42101=>"101010010",
  42102=>"111111110",
  42103=>"000110011",
  42104=>"101101111",
  42105=>"010000101",
  42106=>"010100011",
  42107=>"100111000",
  42108=>"101110110",
  42109=>"110100000",
  42110=>"010000000",
  42111=>"001100011",
  42112=>"110010010",
  42113=>"101110111",
  42114=>"111110100",
  42115=>"110100111",
  42116=>"111111000",
  42117=>"000011111",
  42118=>"101001011",
  42119=>"100111011",
  42120=>"100010010",
  42121=>"110101111",
  42122=>"001111001",
  42123=>"110001001",
  42124=>"111010101",
  42125=>"010111011",
  42126=>"010010101",
  42127=>"110000011",
  42128=>"100000101",
  42129=>"111110101",
  42130=>"111000100",
  42131=>"101111000",
  42132=>"000111001",
  42133=>"110111001",
  42134=>"111111001",
  42135=>"001010110",
  42136=>"001010001",
  42137=>"011010100",
  42138=>"100010001",
  42139=>"010001000",
  42140=>"011100101",
  42141=>"101110001",
  42142=>"111001111",
  42143=>"010100101",
  42144=>"010100010",
  42145=>"100010010",
  42146=>"011001011",
  42147=>"001100000",
  42148=>"111101011",
  42149=>"101110010",
  42150=>"000101000",
  42151=>"100011110",
  42152=>"110001110",
  42153=>"001000010",
  42154=>"100101001",
  42155=>"001010100",
  42156=>"111010110",
  42157=>"000011110",
  42158=>"110110010",
  42159=>"000000000",
  42160=>"110100011",
  42161=>"010001101",
  42162=>"000001110",
  42163=>"001110111",
  42164=>"111111000",
  42165=>"110010001",
  42166=>"111001010",
  42167=>"000101011",
  42168=>"010011100",
  42169=>"101101111",
  42170=>"111010000",
  42171=>"010110111",
  42172=>"100001101",
  42173=>"000010111",
  42174=>"000000100",
  42175=>"000010111",
  42176=>"010010100",
  42177=>"000000111",
  42178=>"101011111",
  42179=>"010001111",
  42180=>"001000111",
  42181=>"100000101",
  42182=>"000100110",
  42183=>"101110011",
  42184=>"000111101",
  42185=>"011010001",
  42186=>"001011011",
  42187=>"101001001",
  42188=>"001101100",
  42189=>"000110000",
  42190=>"000110011",
  42191=>"101100101",
  42192=>"100111000",
  42193=>"110111110",
  42194=>"010110101",
  42195=>"100111110",
  42196=>"011010001",
  42197=>"100000000",
  42198=>"011011100",
  42199=>"011011110",
  42200=>"101100000",
  42201=>"000100001",
  42202=>"101011010",
  42203=>"110000100",
  42204=>"111000110",
  42205=>"111011000",
  42206=>"101100101",
  42207=>"011010011",
  42208=>"001011100",
  42209=>"101011110",
  42210=>"110010001",
  42211=>"101101011",
  42212=>"101000100",
  42213=>"111110110",
  42214=>"000111010",
  42215=>"011100100",
  42216=>"101010100",
  42217=>"001000010",
  42218=>"001000001",
  42219=>"001101100",
  42220=>"110011000",
  42221=>"000010101",
  42222=>"011100110",
  42223=>"000100100",
  42224=>"110111110",
  42225=>"011101111",
  42226=>"101010011",
  42227=>"000101101",
  42228=>"111101011",
  42229=>"010011010",
  42230=>"000011100",
  42231=>"100011110",
  42232=>"001101000",
  42233=>"111100101",
  42234=>"000010010",
  42235=>"011001010",
  42236=>"101001011",
  42237=>"001101101",
  42238=>"011010110",
  42239=>"110110110",
  42240=>"010111010",
  42241=>"010011111",
  42242=>"010011010",
  42243=>"100000100",
  42244=>"001000010",
  42245=>"010010001",
  42246=>"010001110",
  42247=>"000001011",
  42248=>"101001011",
  42249=>"100001111",
  42250=>"111111110",
  42251=>"111110111",
  42252=>"011001011",
  42253=>"001110100",
  42254=>"100110101",
  42255=>"110100000",
  42256=>"010010110",
  42257=>"101111111",
  42258=>"111111111",
  42259=>"010111111",
  42260=>"000000111",
  42261=>"011111101",
  42262=>"000000000",
  42263=>"111001101",
  42264=>"101110010",
  42265=>"100111111",
  42266=>"111101101",
  42267=>"010111111",
  42268=>"110111000",
  42269=>"111011111",
  42270=>"000001110",
  42271=>"001010111",
  42272=>"011001000",
  42273=>"011110001",
  42274=>"100110110",
  42275=>"100111001",
  42276=>"100001101",
  42277=>"011100111",
  42278=>"101010001",
  42279=>"011110111",
  42280=>"011110101",
  42281=>"101100101",
  42282=>"100100111",
  42283=>"100000000",
  42284=>"011111101",
  42285=>"110110100",
  42286=>"000001110",
  42287=>"000000100",
  42288=>"011010000",
  42289=>"000101011",
  42290=>"110111011",
  42291=>"100111000",
  42292=>"101111010",
  42293=>"111101100",
  42294=>"000011111",
  42295=>"011101111",
  42296=>"100001011",
  42297=>"101000111",
  42298=>"000010100",
  42299=>"000101011",
  42300=>"000101011",
  42301=>"001011110",
  42302=>"101111010",
  42303=>"110101111",
  42304=>"111001101",
  42305=>"110101001",
  42306=>"010111101",
  42307=>"010000100",
  42308=>"100011000",
  42309=>"010100011",
  42310=>"111001101",
  42311=>"100110110",
  42312=>"101111011",
  42313=>"001011101",
  42314=>"110010000",
  42315=>"101010111",
  42316=>"100110010",
  42317=>"110111100",
  42318=>"000001001",
  42319=>"000010000",
  42320=>"111000000",
  42321=>"001011110",
  42322=>"010101101",
  42323=>"111101101",
  42324=>"101110111",
  42325=>"111101001",
  42326=>"110101010",
  42327=>"101000010",
  42328=>"010001101",
  42329=>"100100100",
  42330=>"110011011",
  42331=>"000100011",
  42332=>"011111001",
  42333=>"010110011",
  42334=>"000101000",
  42335=>"001111000",
  42336=>"000010010",
  42337=>"011000101",
  42338=>"001011000",
  42339=>"111010111",
  42340=>"001011001",
  42341=>"011011000",
  42342=>"001000011",
  42343=>"001000000",
  42344=>"100010001",
  42345=>"000000001",
  42346=>"000011001",
  42347=>"110101010",
  42348=>"010111000",
  42349=>"000000010",
  42350=>"011101101",
  42351=>"001101101",
  42352=>"001000111",
  42353=>"100001110",
  42354=>"110100010",
  42355=>"110100111",
  42356=>"000001101",
  42357=>"110100101",
  42358=>"001010101",
  42359=>"011111001",
  42360=>"110011101",
  42361=>"000001111",
  42362=>"110011100",
  42363=>"011000011",
  42364=>"110011001",
  42365=>"111100100",
  42366=>"001110001",
  42367=>"111110100",
  42368=>"101011111",
  42369=>"100100000",
  42370=>"100101001",
  42371=>"111000111",
  42372=>"100011010",
  42373=>"010110000",
  42374=>"010100111",
  42375=>"101110010",
  42376=>"001011000",
  42377=>"001001100",
  42378=>"000100111",
  42379=>"101011000",
  42380=>"101000111",
  42381=>"111000000",
  42382=>"000100110",
  42383=>"010111111",
  42384=>"111001011",
  42385=>"011110011",
  42386=>"010010111",
  42387=>"111010011",
  42388=>"100001010",
  42389=>"110000011",
  42390=>"110011100",
  42391=>"001101111",
  42392=>"001111010",
  42393=>"101011001",
  42394=>"101000010",
  42395=>"101101101",
  42396=>"000000000",
  42397=>"110101011",
  42398=>"100111110",
  42399=>"010100111",
  42400=>"111111100",
  42401=>"110000010",
  42402=>"000011001",
  42403=>"110110100",
  42404=>"101110110",
  42405=>"000000001",
  42406=>"011101100",
  42407=>"001011100",
  42408=>"100100100",
  42409=>"011000110",
  42410=>"010010001",
  42411=>"110010011",
  42412=>"110110100",
  42413=>"111011101",
  42414=>"101101000",
  42415=>"111011010",
  42416=>"011110011",
  42417=>"100000111",
  42418=>"101110111",
  42419=>"101000111",
  42420=>"111111110",
  42421=>"010110011",
  42422=>"001011100",
  42423=>"111001111",
  42424=>"100111101",
  42425=>"110111101",
  42426=>"000000000",
  42427=>"111010110",
  42428=>"100000100",
  42429=>"100001111",
  42430=>"001101010",
  42431=>"101100111",
  42432=>"011110101",
  42433=>"000001000",
  42434=>"111101100",
  42435=>"111011001",
  42436=>"000110111",
  42437=>"111100000",
  42438=>"000010001",
  42439=>"000110100",
  42440=>"010100010",
  42441=>"001101111",
  42442=>"001000001",
  42443=>"100000011",
  42444=>"000100101",
  42445=>"000010111",
  42446=>"010000011",
  42447=>"101010111",
  42448=>"000111110",
  42449=>"011100001",
  42450=>"011101001",
  42451=>"100101110",
  42452=>"111101011",
  42453=>"101100001",
  42454=>"010110001",
  42455=>"111111100",
  42456=>"111000100",
  42457=>"001111100",
  42458=>"011100001",
  42459=>"101010001",
  42460=>"011100011",
  42461=>"110101010",
  42462=>"000001100",
  42463=>"010111111",
  42464=>"110000100",
  42465=>"010100011",
  42466=>"111011011",
  42467=>"101111000",
  42468=>"111100111",
  42469=>"110111111",
  42470=>"101101111",
  42471=>"001111000",
  42472=>"011011001",
  42473=>"011111001",
  42474=>"000101111",
  42475=>"101111011",
  42476=>"011101000",
  42477=>"000101000",
  42478=>"110000111",
  42479=>"100100001",
  42480=>"001001100",
  42481=>"010101100",
  42482=>"111110010",
  42483=>"101011011",
  42484=>"111001110",
  42485=>"011010001",
  42486=>"011100011",
  42487=>"111010111",
  42488=>"100101110",
  42489=>"001100111",
  42490=>"111011100",
  42491=>"011100001",
  42492=>"110010111",
  42493=>"001111001",
  42494=>"000100001",
  42495=>"101000000",
  42496=>"100000000",
  42497=>"100000111",
  42498=>"001110111",
  42499=>"000111100",
  42500=>"010011001",
  42501=>"110010010",
  42502=>"010000010",
  42503=>"111110010",
  42504=>"000010010",
  42505=>"111101111",
  42506=>"011110000",
  42507=>"100100011",
  42508=>"001001000",
  42509=>"101100111",
  42510=>"111000000",
  42511=>"111111001",
  42512=>"010010101",
  42513=>"110010001",
  42514=>"101100110",
  42515=>"101101000",
  42516=>"101000010",
  42517=>"000110111",
  42518=>"011101110",
  42519=>"001111000",
  42520=>"111101101",
  42521=>"110011100",
  42522=>"011000010",
  42523=>"000011010",
  42524=>"000111011",
  42525=>"001000000",
  42526=>"000011110",
  42527=>"101100111",
  42528=>"010011100",
  42529=>"100011100",
  42530=>"001001001",
  42531=>"011001100",
  42532=>"011010101",
  42533=>"011011011",
  42534=>"001011111",
  42535=>"111011001",
  42536=>"000100110",
  42537=>"010010101",
  42538=>"111100011",
  42539=>"010010010",
  42540=>"110110110",
  42541=>"000000111",
  42542=>"110110100",
  42543=>"001110111",
  42544=>"011010100",
  42545=>"110011111",
  42546=>"111100101",
  42547=>"000000000",
  42548=>"110000010",
  42549=>"001110111",
  42550=>"100100101",
  42551=>"110010011",
  42552=>"110110010",
  42553=>"111110110",
  42554=>"001101100",
  42555=>"110111101",
  42556=>"100000111",
  42557=>"010010111",
  42558=>"001100111",
  42559=>"000000100",
  42560=>"100001111",
  42561=>"010111000",
  42562=>"111100100",
  42563=>"000111001",
  42564=>"110110000",
  42565=>"111110101",
  42566=>"000100000",
  42567=>"000110000",
  42568=>"000110011",
  42569=>"111101110",
  42570=>"001000101",
  42571=>"111101001",
  42572=>"010011101",
  42573=>"101000111",
  42574=>"111110100",
  42575=>"111010101",
  42576=>"100111111",
  42577=>"111010001",
  42578=>"111110101",
  42579=>"110110101",
  42580=>"001001000",
  42581=>"000000110",
  42582=>"100100101",
  42583=>"101100111",
  42584=>"000101000",
  42585=>"110111100",
  42586=>"110110001",
  42587=>"010100111",
  42588=>"110100011",
  42589=>"111000110",
  42590=>"010000111",
  42591=>"011110110",
  42592=>"100111000",
  42593=>"100111010",
  42594=>"000001001",
  42595=>"111011000",
  42596=>"010111110",
  42597=>"101000000",
  42598=>"110000110",
  42599=>"011101010",
  42600=>"111011011",
  42601=>"010111110",
  42602=>"011110001",
  42603=>"011110111",
  42604=>"110100011",
  42605=>"010000010",
  42606=>"101001110",
  42607=>"001111110",
  42608=>"001101001",
  42609=>"111101000",
  42610=>"011001001",
  42611=>"111101111",
  42612=>"000010110",
  42613=>"111100011",
  42614=>"011011101",
  42615=>"000011101",
  42616=>"110011010",
  42617=>"101000101",
  42618=>"100011010",
  42619=>"000100011",
  42620=>"110001010",
  42621=>"111000001",
  42622=>"110111010",
  42623=>"011000101",
  42624=>"001100101",
  42625=>"001100000",
  42626=>"011001101",
  42627=>"011000100",
  42628=>"001100001",
  42629=>"101001000",
  42630=>"101000011",
  42631=>"011000110",
  42632=>"100001010",
  42633=>"111011010",
  42634=>"110100110",
  42635=>"000101010",
  42636=>"101011000",
  42637=>"000110100",
  42638=>"111011110",
  42639=>"000000000",
  42640=>"100011000",
  42641=>"011110000",
  42642=>"011110111",
  42643=>"001000101",
  42644=>"001011111",
  42645=>"011000110",
  42646=>"010010100",
  42647=>"001111110",
  42648=>"111111011",
  42649=>"010010010",
  42650=>"110110110",
  42651=>"111010101",
  42652=>"010010100",
  42653=>"100100010",
  42654=>"011100100",
  42655=>"101111011",
  42656=>"101100110",
  42657=>"011000010",
  42658=>"111011101",
  42659=>"100001011",
  42660=>"011110001",
  42661=>"000111110",
  42662=>"010001111",
  42663=>"011001101",
  42664=>"011001111",
  42665=>"001000101",
  42666=>"101101010",
  42667=>"011010100",
  42668=>"111001010",
  42669=>"101111100",
  42670=>"100111010",
  42671=>"111100010",
  42672=>"011001011",
  42673=>"001100101",
  42674=>"011100111",
  42675=>"110011100",
  42676=>"100000111",
  42677=>"000001111",
  42678=>"100001000",
  42679=>"000001111",
  42680=>"010001001",
  42681=>"110001100",
  42682=>"000110001",
  42683=>"111101001",
  42684=>"101101001",
  42685=>"110001010",
  42686=>"110110100",
  42687=>"000000011",
  42688=>"111111110",
  42689=>"000111011",
  42690=>"001100110",
  42691=>"011101111",
  42692=>"000111101",
  42693=>"000010111",
  42694=>"111010101",
  42695=>"111001101",
  42696=>"111000111",
  42697=>"111111011",
  42698=>"011010111",
  42699=>"111000000",
  42700=>"111001110",
  42701=>"110001000",
  42702=>"101000001",
  42703=>"110100101",
  42704=>"000111101",
  42705=>"101111001",
  42706=>"000011111",
  42707=>"100010001",
  42708=>"011100001",
  42709=>"100000010",
  42710=>"000111000",
  42711=>"010110110",
  42712=>"100101010",
  42713=>"000100000",
  42714=>"110110001",
  42715=>"111101001",
  42716=>"110101100",
  42717=>"011000101",
  42718=>"111100110",
  42719=>"111101001",
  42720=>"100011110",
  42721=>"011010100",
  42722=>"100010100",
  42723=>"101011010",
  42724=>"010111101",
  42725=>"010000101",
  42726=>"101011101",
  42727=>"010000010",
  42728=>"100100011",
  42729=>"010111100",
  42730=>"011100010",
  42731=>"100110011",
  42732=>"111011110",
  42733=>"000100000",
  42734=>"100010010",
  42735=>"101110000",
  42736=>"011111010",
  42737=>"010100110",
  42738=>"000101101",
  42739=>"111010100",
  42740=>"101111100",
  42741=>"000110001",
  42742=>"111010010",
  42743=>"001101010",
  42744=>"010100100",
  42745=>"101100011",
  42746=>"101101110",
  42747=>"000010000",
  42748=>"111010100",
  42749=>"010000101",
  42750=>"111101100",
  42751=>"010011000",
  42752=>"000101110",
  42753=>"000110000",
  42754=>"000001011",
  42755=>"110101010",
  42756=>"011111111",
  42757=>"111011000",
  42758=>"011101001",
  42759=>"000010001",
  42760=>"111011001",
  42761=>"011011011",
  42762=>"110111001",
  42763=>"001011111",
  42764=>"001100001",
  42765=>"011100000",
  42766=>"101000011",
  42767=>"101111001",
  42768=>"000000111",
  42769=>"111101110",
  42770=>"111111100",
  42771=>"000011111",
  42772=>"110001100",
  42773=>"111110101",
  42774=>"110110011",
  42775=>"001110010",
  42776=>"011111000",
  42777=>"010000001",
  42778=>"000000100",
  42779=>"110001010",
  42780=>"011000011",
  42781=>"011110101",
  42782=>"000000000",
  42783=>"010110010",
  42784=>"111111111",
  42785=>"101100111",
  42786=>"001110100",
  42787=>"110000010",
  42788=>"001111010",
  42789=>"001100011",
  42790=>"011010011",
  42791=>"110110000",
  42792=>"011010011",
  42793=>"011100111",
  42794=>"111000100",
  42795=>"101110110",
  42796=>"001011110",
  42797=>"001000111",
  42798=>"000001000",
  42799=>"110101110",
  42800=>"001000110",
  42801=>"000000001",
  42802=>"101010001",
  42803=>"001000011",
  42804=>"101101100",
  42805=>"010111111",
  42806=>"010010111",
  42807=>"010100111",
  42808=>"001111010",
  42809=>"100011100",
  42810=>"010101110",
  42811=>"001110100",
  42812=>"101101010",
  42813=>"011110000",
  42814=>"110111110",
  42815=>"111111110",
  42816=>"000001010",
  42817=>"000011111",
  42818=>"010000000",
  42819=>"000000001",
  42820=>"001101111",
  42821=>"100010011",
  42822=>"000100101",
  42823=>"010101011",
  42824=>"011000000",
  42825=>"000110001",
  42826=>"001111001",
  42827=>"111100000",
  42828=>"001110011",
  42829=>"010101110",
  42830=>"001010110",
  42831=>"101010111",
  42832=>"100100000",
  42833=>"110010100",
  42834=>"010110011",
  42835=>"111010101",
  42836=>"000101100",
  42837=>"000100101",
  42838=>"111000010",
  42839=>"111010011",
  42840=>"101101100",
  42841=>"010010101",
  42842=>"100110010",
  42843=>"111011010",
  42844=>"111011100",
  42845=>"110101110",
  42846=>"000010011",
  42847=>"000001001",
  42848=>"111011010",
  42849=>"111010001",
  42850=>"001000111",
  42851=>"011011111",
  42852=>"000000000",
  42853=>"101111010",
  42854=>"101001111",
  42855=>"011011101",
  42856=>"000100010",
  42857=>"010100011",
  42858=>"010011111",
  42859=>"110001000",
  42860=>"110011000",
  42861=>"111000110",
  42862=>"100010000",
  42863=>"010110110",
  42864=>"111001111",
  42865=>"011101101",
  42866=>"011011101",
  42867=>"101100000",
  42868=>"100000001",
  42869=>"101101001",
  42870=>"100101001",
  42871=>"010100101",
  42872=>"011111101",
  42873=>"100001000",
  42874=>"001010010",
  42875=>"100010011",
  42876=>"011000110",
  42877=>"001100010",
  42878=>"111100110",
  42879=>"011110100",
  42880=>"001010110",
  42881=>"011011011",
  42882=>"110010001",
  42883=>"111100110",
  42884=>"110011101",
  42885=>"000011011",
  42886=>"110001001",
  42887=>"100000001",
  42888=>"101010011",
  42889=>"100110110",
  42890=>"100010100",
  42891=>"111100111",
  42892=>"101011010",
  42893=>"110000011",
  42894=>"100000111",
  42895=>"000110100",
  42896=>"011100111",
  42897=>"001100000",
  42898=>"001000000",
  42899=>"010100111",
  42900=>"010011111",
  42901=>"111100100",
  42902=>"100100010",
  42903=>"001110010",
  42904=>"110001000",
  42905=>"010110010",
  42906=>"011000100",
  42907=>"000000011",
  42908=>"001011111",
  42909=>"100010010",
  42910=>"111110101",
  42911=>"010010000",
  42912=>"101011111",
  42913=>"111011110",
  42914=>"101010111",
  42915=>"111010001",
  42916=>"011111000",
  42917=>"011000011",
  42918=>"000100100",
  42919=>"011110110",
  42920=>"101000001",
  42921=>"000101001",
  42922=>"100100001",
  42923=>"101110101",
  42924=>"011010101",
  42925=>"011000101",
  42926=>"111111001",
  42927=>"010000000",
  42928=>"110100111",
  42929=>"001100011",
  42930=>"000010010",
  42931=>"100111010",
  42932=>"011101000",
  42933=>"001111110",
  42934=>"100000011",
  42935=>"000001100",
  42936=>"110111110",
  42937=>"010110110",
  42938=>"010100101",
  42939=>"011011101",
  42940=>"100101110",
  42941=>"110010111",
  42942=>"000000010",
  42943=>"100011101",
  42944=>"101011101",
  42945=>"110100000",
  42946=>"000101010",
  42947=>"101111100",
  42948=>"011100101",
  42949=>"101010001",
  42950=>"111011101",
  42951=>"011101111",
  42952=>"101000000",
  42953=>"100110011",
  42954=>"111111101",
  42955=>"111011000",
  42956=>"001101011",
  42957=>"010110111",
  42958=>"100010110",
  42959=>"111101111",
  42960=>"111001110",
  42961=>"111000111",
  42962=>"111001101",
  42963=>"010000100",
  42964=>"000010000",
  42965=>"100101000",
  42966=>"010000100",
  42967=>"001001111",
  42968=>"101000010",
  42969=>"100101001",
  42970=>"000000011",
  42971=>"100000000",
  42972=>"000101101",
  42973=>"000011110",
  42974=>"000111111",
  42975=>"010101101",
  42976=>"110111000",
  42977=>"101100100",
  42978=>"101111101",
  42979=>"000000111",
  42980=>"111001100",
  42981=>"011001111",
  42982=>"001000010",
  42983=>"001001000",
  42984=>"001000000",
  42985=>"011110000",
  42986=>"000100010",
  42987=>"011111111",
  42988=>"110110010",
  42989=>"000011000",
  42990=>"110001101",
  42991=>"000000110",
  42992=>"101111111",
  42993=>"001111010",
  42994=>"010000110",
  42995=>"000010100",
  42996=>"100110110",
  42997=>"110111101",
  42998=>"110100100",
  42999=>"111110101",
  43000=>"101011011",
  43001=>"100111010",
  43002=>"110001110",
  43003=>"101110011",
  43004=>"000101101",
  43005=>"101100000",
  43006=>"000111010",
  43007=>"011001010",
  43008=>"010111010",
  43009=>"111010101",
  43010=>"111010000",
  43011=>"100100000",
  43012=>"001001011",
  43013=>"001000010",
  43014=>"111101101",
  43015=>"111110101",
  43016=>"000000011",
  43017=>"110000111",
  43018=>"110001000",
  43019=>"111011001",
  43020=>"010110010",
  43021=>"011110001",
  43022=>"001110010",
  43023=>"000101000",
  43024=>"000010100",
  43025=>"010011101",
  43026=>"010011111",
  43027=>"101010101",
  43028=>"100001000",
  43029=>"001100010",
  43030=>"100101100",
  43031=>"111111111",
  43032=>"000010101",
  43033=>"000000000",
  43034=>"010110001",
  43035=>"110111100",
  43036=>"110111000",
  43037=>"010010111",
  43038=>"111010100",
  43039=>"110110001",
  43040=>"010010110",
  43041=>"111000111",
  43042=>"010001011",
  43043=>"001000001",
  43044=>"100110100",
  43045=>"111110101",
  43046=>"100001111",
  43047=>"100010110",
  43048=>"100000000",
  43049=>"111011110",
  43050=>"001010000",
  43051=>"111010110",
  43052=>"000110111",
  43053=>"000001001",
  43054=>"011011011",
  43055=>"001101000",
  43056=>"010001110",
  43057=>"010100010",
  43058=>"001111000",
  43059=>"000010010",
  43060=>"100100000",
  43061=>"000010001",
  43062=>"011101110",
  43063=>"001010111",
  43064=>"100000001",
  43065=>"101000000",
  43066=>"001100111",
  43067=>"000001001",
  43068=>"111101111",
  43069=>"100000001",
  43070=>"011010100",
  43071=>"100101010",
  43072=>"100000000",
  43073=>"100100000",
  43074=>"000001011",
  43075=>"010010010",
  43076=>"100100010",
  43077=>"001010111",
  43078=>"011001011",
  43079=>"110101101",
  43080=>"011111010",
  43081=>"101111011",
  43082=>"100111010",
  43083=>"010111001",
  43084=>"010011000",
  43085=>"011101001",
  43086=>"001001100",
  43087=>"110110101",
  43088=>"110011111",
  43089=>"010110101",
  43090=>"000000110",
  43091=>"000011011",
  43092=>"111110101",
  43093=>"000000011",
  43094=>"010010110",
  43095=>"110010100",
  43096=>"101011111",
  43097=>"111000011",
  43098=>"100100100",
  43099=>"000001010",
  43100=>"000100111",
  43101=>"000000111",
  43102=>"011011000",
  43103=>"100011010",
  43104=>"100010110",
  43105=>"011010110",
  43106=>"110011111",
  43107=>"001000010",
  43108=>"100011010",
  43109=>"011110001",
  43110=>"010101100",
  43111=>"001100101",
  43112=>"011011100",
  43113=>"110110111",
  43114=>"101100000",
  43115=>"111000000",
  43116=>"110010101",
  43117=>"110100111",
  43118=>"001111001",
  43119=>"000100111",
  43120=>"010100100",
  43121=>"000110000",
  43122=>"110101000",
  43123=>"001000001",
  43124=>"001000010",
  43125=>"101101101",
  43126=>"100101001",
  43127=>"110010010",
  43128=>"010100110",
  43129=>"010001011",
  43130=>"000000001",
  43131=>"000100111",
  43132=>"101011111",
  43133=>"000111101",
  43134=>"010101011",
  43135=>"101100011",
  43136=>"011100111",
  43137=>"000010110",
  43138=>"001010010",
  43139=>"000001101",
  43140=>"110101010",
  43141=>"001110000",
  43142=>"000011010",
  43143=>"110110111",
  43144=>"010010101",
  43145=>"110001101",
  43146=>"101000010",
  43147=>"101010100",
  43148=>"100111001",
  43149=>"100000100",
  43150=>"000111111",
  43151=>"101100110",
  43152=>"000100100",
  43153=>"001010101",
  43154=>"111000010",
  43155=>"010110110",
  43156=>"000001100",
  43157=>"101001101",
  43158=>"101111100",
  43159=>"001011100",
  43160=>"101110010",
  43161=>"110111011",
  43162=>"010011000",
  43163=>"010011101",
  43164=>"011000111",
  43165=>"101000011",
  43166=>"000100011",
  43167=>"101000110",
  43168=>"101010110",
  43169=>"110110001",
  43170=>"010101001",
  43171=>"000010100",
  43172=>"110111010",
  43173=>"111011110",
  43174=>"100110100",
  43175=>"000000001",
  43176=>"011001001",
  43177=>"010000100",
  43178=>"110001000",
  43179=>"010010001",
  43180=>"110111011",
  43181=>"101100001",
  43182=>"000010001",
  43183=>"000101010",
  43184=>"011001001",
  43185=>"110110100",
  43186=>"110111111",
  43187=>"101100110",
  43188=>"010010000",
  43189=>"000010111",
  43190=>"011001101",
  43191=>"101110000",
  43192=>"111111001",
  43193=>"000010001",
  43194=>"000010101",
  43195=>"010000001",
  43196=>"010100110",
  43197=>"100000001",
  43198=>"100101100",
  43199=>"000100000",
  43200=>"110110111",
  43201=>"011000011",
  43202=>"111111010",
  43203=>"100011010",
  43204=>"010100111",
  43205=>"111100000",
  43206=>"010000100",
  43207=>"110010010",
  43208=>"001000101",
  43209=>"110111101",
  43210=>"001011111",
  43211=>"000011011",
  43212=>"110000110",
  43213=>"010010000",
  43214=>"000100111",
  43215=>"001010000",
  43216=>"110001001",
  43217=>"100000011",
  43218=>"011001010",
  43219=>"101101100",
  43220=>"100000111",
  43221=>"111000101",
  43222=>"111011001",
  43223=>"101110001",
  43224=>"110101010",
  43225=>"111100010",
  43226=>"011101101",
  43227=>"010011110",
  43228=>"110110011",
  43229=>"010111010",
  43230=>"001111001",
  43231=>"110000111",
  43232=>"111011000",
  43233=>"010010011",
  43234=>"110111111",
  43235=>"111100001",
  43236=>"100011111",
  43237=>"110110100",
  43238=>"110111111",
  43239=>"000010100",
  43240=>"100000111",
  43241=>"010111100",
  43242=>"000000011",
  43243=>"111011000",
  43244=>"001010000",
  43245=>"010000001",
  43246=>"011010111",
  43247=>"000100010",
  43248=>"100000011",
  43249=>"000011001",
  43250=>"101111010",
  43251=>"100110011",
  43252=>"101110100",
  43253=>"011010111",
  43254=>"100011010",
  43255=>"100101100",
  43256=>"110000100",
  43257=>"100101111",
  43258=>"110011111",
  43259=>"001001001",
  43260=>"000101111",
  43261=>"001111111",
  43262=>"110111111",
  43263=>"010011111",
  43264=>"011010001",
  43265=>"101010111",
  43266=>"011000110",
  43267=>"001010000",
  43268=>"001101111",
  43269=>"000101011",
  43270=>"000011001",
  43271=>"101101001",
  43272=>"111011110",
  43273=>"001000100",
  43274=>"100111101",
  43275=>"001000110",
  43276=>"000001000",
  43277=>"001000110",
  43278=>"000010101",
  43279=>"010000100",
  43280=>"001110111",
  43281=>"011000001",
  43282=>"011001100",
  43283=>"101011101",
  43284=>"001100111",
  43285=>"101011010",
  43286=>"000000101",
  43287=>"100000100",
  43288=>"000111100",
  43289=>"010111100",
  43290=>"001001111",
  43291=>"010100100",
  43292=>"011110100",
  43293=>"111110101",
  43294=>"110001010",
  43295=>"100001000",
  43296=>"100010100",
  43297=>"111110110",
  43298=>"100100100",
  43299=>"100001011",
  43300=>"100001110",
  43301=>"111000000",
  43302=>"010101010",
  43303=>"111010011",
  43304=>"000000000",
  43305=>"011000000",
  43306=>"111101111",
  43307=>"000001111",
  43308=>"110111001",
  43309=>"110000001",
  43310=>"111100101",
  43311=>"010010110",
  43312=>"010110010",
  43313=>"111011001",
  43314=>"011001111",
  43315=>"101100001",
  43316=>"000011001",
  43317=>"001001001",
  43318=>"001101001",
  43319=>"001010100",
  43320=>"000110111",
  43321=>"100101111",
  43322=>"000010010",
  43323=>"101100101",
  43324=>"011100000",
  43325=>"100111100",
  43326=>"111001000",
  43327=>"101000001",
  43328=>"010100100",
  43329=>"011001110",
  43330=>"110010111",
  43331=>"000011000",
  43332=>"000100101",
  43333=>"100100001",
  43334=>"010000000",
  43335=>"100011001",
  43336=>"100001011",
  43337=>"010111011",
  43338=>"010000010",
  43339=>"100101101",
  43340=>"111001110",
  43341=>"001110100",
  43342=>"101100110",
  43343=>"011010000",
  43344=>"110000101",
  43345=>"000110010",
  43346=>"101110010",
  43347=>"111011011",
  43348=>"011101011",
  43349=>"000110111",
  43350=>"001110010",
  43351=>"001011101",
  43352=>"000111011",
  43353=>"111011001",
  43354=>"111110111",
  43355=>"000001111",
  43356=>"111110011",
  43357=>"000111011",
  43358=>"111000000",
  43359=>"000000011",
  43360=>"011101111",
  43361=>"000011000",
  43362=>"010100000",
  43363=>"000011111",
  43364=>"110101010",
  43365=>"011001101",
  43366=>"000010011",
  43367=>"010111000",
  43368=>"001101000",
  43369=>"010011110",
  43370=>"000001101",
  43371=>"111010011",
  43372=>"101011010",
  43373=>"101000011",
  43374=>"001000001",
  43375=>"101001100",
  43376=>"000101100",
  43377=>"010111101",
  43378=>"011110010",
  43379=>"010101011",
  43380=>"010001101",
  43381=>"111011000",
  43382=>"000011001",
  43383=>"011100010",
  43384=>"001110100",
  43385=>"000100111",
  43386=>"100000101",
  43387=>"000100110",
  43388=>"001111010",
  43389=>"100000100",
  43390=>"001111110",
  43391=>"001010110",
  43392=>"100001011",
  43393=>"110110000",
  43394=>"001001011",
  43395=>"001100110",
  43396=>"011001011",
  43397=>"110101001",
  43398=>"011001110",
  43399=>"001101100",
  43400=>"111001010",
  43401=>"001100000",
  43402=>"100011011",
  43403=>"110001010",
  43404=>"000010110",
  43405=>"011010101",
  43406=>"001001001",
  43407=>"111011001",
  43408=>"010110100",
  43409=>"110101001",
  43410=>"000001001",
  43411=>"000011011",
  43412=>"101101001",
  43413=>"011000000",
  43414=>"111000101",
  43415=>"000111110",
  43416=>"010100000",
  43417=>"101000101",
  43418=>"011110000",
  43419=>"001000100",
  43420=>"011111010",
  43421=>"100010010",
  43422=>"101101110",
  43423=>"101000001",
  43424=>"110111000",
  43425=>"000110100",
  43426=>"110111100",
  43427=>"000000101",
  43428=>"101010000",
  43429=>"111001010",
  43430=>"001000001",
  43431=>"000010010",
  43432=>"000001111",
  43433=>"000100111",
  43434=>"111110100",
  43435=>"101100111",
  43436=>"111101001",
  43437=>"010011011",
  43438=>"000000011",
  43439=>"011000101",
  43440=>"010000110",
  43441=>"011000011",
  43442=>"110110011",
  43443=>"110100011",
  43444=>"000010000",
  43445=>"110010101",
  43446=>"010110001",
  43447=>"100010100",
  43448=>"101101010",
  43449=>"101000111",
  43450=>"110011000",
  43451=>"101010010",
  43452=>"100010100",
  43453=>"011011111",
  43454=>"001001100",
  43455=>"010010010",
  43456=>"011010101",
  43457=>"011101111",
  43458=>"001101010",
  43459=>"101100101",
  43460=>"000101000",
  43461=>"001101101",
  43462=>"000000001",
  43463=>"001000010",
  43464=>"100010101",
  43465=>"011001110",
  43466=>"011111101",
  43467=>"110111100",
  43468=>"011100000",
  43469=>"011001111",
  43470=>"011111101",
  43471=>"100000010",
  43472=>"101111111",
  43473=>"010110111",
  43474=>"001111110",
  43475=>"000010111",
  43476=>"111101000",
  43477=>"010100010",
  43478=>"010110100",
  43479=>"000000100",
  43480=>"100100111",
  43481=>"000010000",
  43482=>"001011110",
  43483=>"110101011",
  43484=>"111000101",
  43485=>"110111000",
  43486=>"000010110",
  43487=>"000110010",
  43488=>"100010110",
  43489=>"111001001",
  43490=>"010110111",
  43491=>"101111000",
  43492=>"100000100",
  43493=>"110010011",
  43494=>"101100011",
  43495=>"000011011",
  43496=>"111101111",
  43497=>"110110101",
  43498=>"111111001",
  43499=>"111000001",
  43500=>"111011010",
  43501=>"111000000",
  43502=>"101011100",
  43503=>"010110010",
  43504=>"100011101",
  43505=>"011000000",
  43506=>"101001110",
  43507=>"101100000",
  43508=>"100001010",
  43509=>"101101100",
  43510=>"111000011",
  43511=>"001001110",
  43512=>"001110010",
  43513=>"001001001",
  43514=>"001101010",
  43515=>"011001111",
  43516=>"110010110",
  43517=>"010001110",
  43518=>"101100111",
  43519=>"000101010",
  43520=>"100000101",
  43521=>"011001000",
  43522=>"001110011",
  43523=>"111000100",
  43524=>"000000100",
  43525=>"100111110",
  43526=>"010011000",
  43527=>"101110001",
  43528=>"001110010",
  43529=>"011101111",
  43530=>"101011010",
  43531=>"011001011",
  43532=>"011011010",
  43533=>"001100100",
  43534=>"001111111",
  43535=>"111001111",
  43536=>"100000101",
  43537=>"010011001",
  43538=>"100110001",
  43539=>"110001101",
  43540=>"000111110",
  43541=>"101011010",
  43542=>"101101110",
  43543=>"011000010",
  43544=>"110100000",
  43545=>"011111001",
  43546=>"100100010",
  43547=>"100011010",
  43548=>"000010011",
  43549=>"000010111",
  43550=>"001100010",
  43551=>"010001010",
  43552=>"100100100",
  43553=>"110101101",
  43554=>"101000001",
  43555=>"110011000",
  43556=>"000100111",
  43557=>"100001001",
  43558=>"110010101",
  43559=>"010011101",
  43560=>"101000000",
  43561=>"011100010",
  43562=>"000011001",
  43563=>"011110111",
  43564=>"000111000",
  43565=>"001000011",
  43566=>"001001100",
  43567=>"010010111",
  43568=>"010000010",
  43569=>"001010111",
  43570=>"111011101",
  43571=>"110000111",
  43572=>"100101101",
  43573=>"100001101",
  43574=>"101111010",
  43575=>"100001011",
  43576=>"000101101",
  43577=>"101111011",
  43578=>"011001111",
  43579=>"001100011",
  43580=>"110110101",
  43581=>"000000000",
  43582=>"110110010",
  43583=>"110010011",
  43584=>"110001100",
  43585=>"101101110",
  43586=>"101001111",
  43587=>"110100111",
  43588=>"000001111",
  43589=>"111000100",
  43590=>"111011100",
  43591=>"000011010",
  43592=>"101101110",
  43593=>"110011101",
  43594=>"111010011",
  43595=>"101100100",
  43596=>"111100101",
  43597=>"101011011",
  43598=>"000011010",
  43599=>"110101111",
  43600=>"011011101",
  43601=>"111001111",
  43602=>"001010011",
  43603=>"111010010",
  43604=>"010101011",
  43605=>"011010110",
  43606=>"000001100",
  43607=>"011010011",
  43608=>"000101010",
  43609=>"000010111",
  43610=>"110011010",
  43611=>"001100001",
  43612=>"000100101",
  43613=>"111110110",
  43614=>"111110011",
  43615=>"101101000",
  43616=>"010010110",
  43617=>"000001000",
  43618=>"001001100",
  43619=>"000010110",
  43620=>"110111001",
  43621=>"000101011",
  43622=>"001010101",
  43623=>"011000000",
  43624=>"000100001",
  43625=>"111111101",
  43626=>"111101011",
  43627=>"000100100",
  43628=>"011000100",
  43629=>"100010110",
  43630=>"010000000",
  43631=>"110000100",
  43632=>"011011111",
  43633=>"110010101",
  43634=>"000100000",
  43635=>"011111000",
  43636=>"110111101",
  43637=>"011100000",
  43638=>"111011110",
  43639=>"000000011",
  43640=>"011010101",
  43641=>"011010010",
  43642=>"100011000",
  43643=>"111101001",
  43644=>"100000011",
  43645=>"100111010",
  43646=>"101001011",
  43647=>"111010100",
  43648=>"110111100",
  43649=>"000101001",
  43650=>"100101110",
  43651=>"001001010",
  43652=>"000101000",
  43653=>"111110001",
  43654=>"110001001",
  43655=>"101101011",
  43656=>"111011111",
  43657=>"011111101",
  43658=>"100010001",
  43659=>"100010010",
  43660=>"111001000",
  43661=>"101111001",
  43662=>"101000000",
  43663=>"111110101",
  43664=>"110000100",
  43665=>"110011001",
  43666=>"100101010",
  43667=>"111100101",
  43668=>"001010111",
  43669=>"110100100",
  43670=>"100000110",
  43671=>"110011100",
  43672=>"001000001",
  43673=>"111100011",
  43674=>"010000110",
  43675=>"000011000",
  43676=>"100100110",
  43677=>"001001010",
  43678=>"111101110",
  43679=>"010000110",
  43680=>"000000001",
  43681=>"111000110",
  43682=>"000011000",
  43683=>"010101111",
  43684=>"110111011",
  43685=>"111111101",
  43686=>"101011101",
  43687=>"010001001",
  43688=>"101011010",
  43689=>"000100000",
  43690=>"111101100",
  43691=>"111001100",
  43692=>"010011011",
  43693=>"010111110",
  43694=>"000111001",
  43695=>"011101011",
  43696=>"110010010",
  43697=>"011000111",
  43698=>"001011110",
  43699=>"011101111",
  43700=>"101000010",
  43701=>"010111100",
  43702=>"100100110",
  43703=>"111111001",
  43704=>"101100000",
  43705=>"101011111",
  43706=>"011101111",
  43707=>"101111011",
  43708=>"111011111",
  43709=>"010011000",
  43710=>"001011101",
  43711=>"111011011",
  43712=>"010100001",
  43713=>"111011001",
  43714=>"000000000",
  43715=>"000100000",
  43716=>"000000110",
  43717=>"111111001",
  43718=>"010111010",
  43719=>"010001110",
  43720=>"111100001",
  43721=>"101100101",
  43722=>"100100010",
  43723=>"100111000",
  43724=>"100010011",
  43725=>"101101000",
  43726=>"011100011",
  43727=>"101100010",
  43728=>"111111000",
  43729=>"101010110",
  43730=>"110101101",
  43731=>"101000000",
  43732=>"001100011",
  43733=>"000101110",
  43734=>"001101000",
  43735=>"100010001",
  43736=>"110100000",
  43737=>"010000010",
  43738=>"001000110",
  43739=>"001011000",
  43740=>"011100110",
  43741=>"010111100",
  43742=>"010000101",
  43743=>"010011110",
  43744=>"110011011",
  43745=>"100010010",
  43746=>"011000010",
  43747=>"101000001",
  43748=>"010101100",
  43749=>"000011011",
  43750=>"000000000",
  43751=>"111111110",
  43752=>"111011000",
  43753=>"110010000",
  43754=>"101110100",
  43755=>"000101001",
  43756=>"001111100",
  43757=>"000001000",
  43758=>"111100100",
  43759=>"111111000",
  43760=>"110111010",
  43761=>"110000001",
  43762=>"001010111",
  43763=>"111011101",
  43764=>"100001111",
  43765=>"011101001",
  43766=>"110011111",
  43767=>"000001011",
  43768=>"111110110",
  43769=>"110000110",
  43770=>"011001100",
  43771=>"010011001",
  43772=>"100101010",
  43773=>"110101010",
  43774=>"001000110",
  43775=>"010100000",
  43776=>"111010100",
  43777=>"111110101",
  43778=>"000010001",
  43779=>"000011111",
  43780=>"011000000",
  43781=>"111011010",
  43782=>"011110011",
  43783=>"110010001",
  43784=>"110000000",
  43785=>"010111011",
  43786=>"110010001",
  43787=>"110000110",
  43788=>"001110000",
  43789=>"100010000",
  43790=>"100110100",
  43791=>"111000100",
  43792=>"000001000",
  43793=>"110100010",
  43794=>"001000011",
  43795=>"100111001",
  43796=>"111101101",
  43797=>"001100001",
  43798=>"010011001",
  43799=>"111000000",
  43800=>"100110000",
  43801=>"110011110",
  43802=>"101011000",
  43803=>"001101111",
  43804=>"101100111",
  43805=>"001101111",
  43806=>"011110100",
  43807=>"000100011",
  43808=>"001010111",
  43809=>"001010011",
  43810=>"011011011",
  43811=>"111010011",
  43812=>"110001100",
  43813=>"110111110",
  43814=>"000011110",
  43815=>"111100001",
  43816=>"100011010",
  43817=>"100110111",
  43818=>"110000000",
  43819=>"101111111",
  43820=>"000101000",
  43821=>"011010111",
  43822=>"101011010",
  43823=>"100111001",
  43824=>"000101110",
  43825=>"101101011",
  43826=>"100110011",
  43827=>"110001010",
  43828=>"000000111",
  43829=>"100000111",
  43830=>"100100110",
  43831=>"000100101",
  43832=>"001101011",
  43833=>"010101000",
  43834=>"111100101",
  43835=>"010101111",
  43836=>"000000000",
  43837=>"101110100",
  43838=>"000000000",
  43839=>"010100000",
  43840=>"000110110",
  43841=>"001011100",
  43842=>"010100111",
  43843=>"101001100",
  43844=>"110100000",
  43845=>"001010100",
  43846=>"100010011",
  43847=>"111010110",
  43848=>"101101001",
  43849=>"100110001",
  43850=>"111001111",
  43851=>"101010110",
  43852=>"101011111",
  43853=>"110111100",
  43854=>"000110110",
  43855=>"110010100",
  43856=>"110010010",
  43857=>"000110111",
  43858=>"100110000",
  43859=>"011110011",
  43860=>"111010100",
  43861=>"111100001",
  43862=>"001111010",
  43863=>"100011010",
  43864=>"000110001",
  43865=>"011010010",
  43866=>"010000111",
  43867=>"010000100",
  43868=>"100100110",
  43869=>"110100101",
  43870=>"000101011",
  43871=>"110110000",
  43872=>"110111000",
  43873=>"001101100",
  43874=>"100001101",
  43875=>"111000011",
  43876=>"000000001",
  43877=>"111000000",
  43878=>"001111100",
  43879=>"111010001",
  43880=>"100111101",
  43881=>"100000010",
  43882=>"100010110",
  43883=>"100000010",
  43884=>"110001011",
  43885=>"100101111",
  43886=>"001011101",
  43887=>"101110111",
  43888=>"010001101",
  43889=>"101111011",
  43890=>"001111111",
  43891=>"110010111",
  43892=>"011111000",
  43893=>"100100100",
  43894=>"110011101",
  43895=>"111000000",
  43896=>"000000111",
  43897=>"011111101",
  43898=>"111011111",
  43899=>"101101111",
  43900=>"000010101",
  43901=>"110110101",
  43902=>"001011101",
  43903=>"011000101",
  43904=>"100101011",
  43905=>"001100001",
  43906=>"001011111",
  43907=>"010000100",
  43908=>"000100000",
  43909=>"110001000",
  43910=>"100100111",
  43911=>"001100101",
  43912=>"111011111",
  43913=>"111010000",
  43914=>"111010011",
  43915=>"000100111",
  43916=>"000010001",
  43917=>"000011010",
  43918=>"011100011",
  43919=>"011100100",
  43920=>"100111110",
  43921=>"000101100",
  43922=>"110010001",
  43923=>"001011010",
  43924=>"101001010",
  43925=>"000000001",
  43926=>"100110010",
  43927=>"001000000",
  43928=>"100001111",
  43929=>"110111000",
  43930=>"000011001",
  43931=>"101001000",
  43932=>"001000011",
  43933=>"000101010",
  43934=>"100111010",
  43935=>"000111011",
  43936=>"110100101",
  43937=>"001101111",
  43938=>"101111100",
  43939=>"011001100",
  43940=>"010001011",
  43941=>"011111101",
  43942=>"111100011",
  43943=>"011001000",
  43944=>"010101110",
  43945=>"100010100",
  43946=>"011011101",
  43947=>"101111011",
  43948=>"101010101",
  43949=>"010101001",
  43950=>"100011010",
  43951=>"010111110",
  43952=>"011010001",
  43953=>"011000011",
  43954=>"111000000",
  43955=>"010101000",
  43956=>"101010011",
  43957=>"011011111",
  43958=>"011001011",
  43959=>"101000001",
  43960=>"111010111",
  43961=>"000100000",
  43962=>"110000000",
  43963=>"110001100",
  43964=>"001111000",
  43965=>"011010000",
  43966=>"010001001",
  43967=>"000100000",
  43968=>"100010111",
  43969=>"100011111",
  43970=>"000000001",
  43971=>"001000000",
  43972=>"100001111",
  43973=>"110010011",
  43974=>"110101111",
  43975=>"010001111",
  43976=>"000001110",
  43977=>"010010000",
  43978=>"111101110",
  43979=>"000110011",
  43980=>"010100111",
  43981=>"111010001",
  43982=>"010000000",
  43983=>"111010101",
  43984=>"100101011",
  43985=>"111011001",
  43986=>"110011111",
  43987=>"000100010",
  43988=>"010100110",
  43989=>"010100100",
  43990=>"010110011",
  43991=>"110110010",
  43992=>"101101010",
  43993=>"011100010",
  43994=>"010011111",
  43995=>"101101101",
  43996=>"000010001",
  43997=>"101101101",
  43998=>"110100001",
  43999=>"111001000",
  44000=>"000101001",
  44001=>"100011111",
  44002=>"011101011",
  44003=>"001110101",
  44004=>"111110011",
  44005=>"000110101",
  44006=>"010111100",
  44007=>"001011010",
  44008=>"000000000",
  44009=>"101110011",
  44010=>"110010101",
  44011=>"001010001",
  44012=>"110110111",
  44013=>"111000000",
  44014=>"000001001",
  44015=>"001111011",
  44016=>"011001100",
  44017=>"010000010",
  44018=>"010000000",
  44019=>"101111111",
  44020=>"010011110",
  44021=>"101110001",
  44022=>"101111010",
  44023=>"110010011",
  44024=>"111110000",
  44025=>"010100111",
  44026=>"111011001",
  44027=>"000000010",
  44028=>"000110011",
  44029=>"001101100",
  44030=>"010001000",
  44031=>"110101111",
  44032=>"110001101",
  44033=>"011100001",
  44034=>"011010110",
  44035=>"110010010",
  44036=>"110000001",
  44037=>"110011101",
  44038=>"000110011",
  44039=>"011100001",
  44040=>"010001001",
  44041=>"101101000",
  44042=>"001010100",
  44043=>"011011110",
  44044=>"010101101",
  44045=>"110010011",
  44046=>"110111101",
  44047=>"111111010",
  44048=>"111110000",
  44049=>"011110011",
  44050=>"001110000",
  44051=>"100100110",
  44052=>"010010011",
  44053=>"000101100",
  44054=>"010111111",
  44055=>"010000100",
  44056=>"001110000",
  44057=>"101001110",
  44058=>"011101010",
  44059=>"111111110",
  44060=>"111011000",
  44061=>"010000010",
  44062=>"100101111",
  44063=>"010100000",
  44064=>"000111110",
  44065=>"011110110",
  44066=>"100111000",
  44067=>"010001110",
  44068=>"110111100",
  44069=>"111010101",
  44070=>"001101111",
  44071=>"110100111",
  44072=>"100000010",
  44073=>"001101110",
  44074=>"110011111",
  44075=>"111100001",
  44076=>"000110100",
  44077=>"000101001",
  44078=>"101110100",
  44079=>"100011110",
  44080=>"000111011",
  44081=>"010111010",
  44082=>"111110001",
  44083=>"111000011",
  44084=>"001101111",
  44085=>"101010001",
  44086=>"011001111",
  44087=>"101101001",
  44088=>"001100111",
  44089=>"110011010",
  44090=>"000001001",
  44091=>"100100001",
  44092=>"010010101",
  44093=>"101010111",
  44094=>"011010010",
  44095=>"101000110",
  44096=>"110001010",
  44097=>"100000010",
  44098=>"101111110",
  44099=>"100101000",
  44100=>"110101100",
  44101=>"001001101",
  44102=>"010111110",
  44103=>"000101000",
  44104=>"100101100",
  44105=>"001100001",
  44106=>"001010111",
  44107=>"010000101",
  44108=>"010100100",
  44109=>"011010100",
  44110=>"011111111",
  44111=>"011001011",
  44112=>"111010010",
  44113=>"100100111",
  44114=>"000100110",
  44115=>"001000100",
  44116=>"011010010",
  44117=>"101001001",
  44118=>"011101100",
  44119=>"001011101",
  44120=>"111011000",
  44121=>"100101110",
  44122=>"000101001",
  44123=>"111101010",
  44124=>"010111101",
  44125=>"111110001",
  44126=>"010100111",
  44127=>"001101000",
  44128=>"000000101",
  44129=>"001111100",
  44130=>"101000001",
  44131=>"000000010",
  44132=>"011010000",
  44133=>"001100111",
  44134=>"110110011",
  44135=>"111011100",
  44136=>"110001011",
  44137=>"100110101",
  44138=>"000001101",
  44139=>"111000010",
  44140=>"100100101",
  44141=>"110111100",
  44142=>"001110011",
  44143=>"111001010",
  44144=>"101001010",
  44145=>"011111110",
  44146=>"000011111",
  44147=>"100001011",
  44148=>"101010111",
  44149=>"000011010",
  44150=>"110111010",
  44151=>"111000110",
  44152=>"100101110",
  44153=>"110000101",
  44154=>"001010001",
  44155=>"110111011",
  44156=>"000100000",
  44157=>"001011111",
  44158=>"011101011",
  44159=>"110101001",
  44160=>"010111001",
  44161=>"111111100",
  44162=>"001100011",
  44163=>"010101000",
  44164=>"000110000",
  44165=>"110101110",
  44166=>"000010000",
  44167=>"001100110",
  44168=>"011010000",
  44169=>"000001010",
  44170=>"101100101",
  44171=>"110010101",
  44172=>"011100000",
  44173=>"111000101",
  44174=>"011111010",
  44175=>"111110000",
  44176=>"000101100",
  44177=>"100000001",
  44178=>"101000001",
  44179=>"100111101",
  44180=>"101010100",
  44181=>"110010101",
  44182=>"100001011",
  44183=>"011110111",
  44184=>"100010101",
  44185=>"010011001",
  44186=>"000100110",
  44187=>"101100001",
  44188=>"000000001",
  44189=>"100101010",
  44190=>"010011010",
  44191=>"010001011",
  44192=>"010010101",
  44193=>"001111000",
  44194=>"001001001",
  44195=>"110000010",
  44196=>"001101010",
  44197=>"000101100",
  44198=>"101111101",
  44199=>"010010100",
  44200=>"000111000",
  44201=>"010001010",
  44202=>"100101110",
  44203=>"011111010",
  44204=>"111101011",
  44205=>"101100011",
  44206=>"111011111",
  44207=>"010101000",
  44208=>"001000100",
  44209=>"100001111",
  44210=>"000011000",
  44211=>"010011011",
  44212=>"111100000",
  44213=>"111110101",
  44214=>"110101101",
  44215=>"111000010",
  44216=>"010110110",
  44217=>"101101101",
  44218=>"011000101",
  44219=>"000010110",
  44220=>"011100010",
  44221=>"100000001",
  44222=>"101010100",
  44223=>"000001000",
  44224=>"001001100",
  44225=>"001000100",
  44226=>"010001110",
  44227=>"010011001",
  44228=>"000101000",
  44229=>"010010111",
  44230=>"100110000",
  44231=>"111000011",
  44232=>"000100000",
  44233=>"110001110",
  44234=>"111111101",
  44235=>"011011101",
  44236=>"001010000",
  44237=>"110100000",
  44238=>"000001111",
  44239=>"010101001",
  44240=>"101100111",
  44241=>"011011000",
  44242=>"001101100",
  44243=>"111111101",
  44244=>"111110000",
  44245=>"110110101",
  44246=>"101111000",
  44247=>"000001011",
  44248=>"101000111",
  44249=>"001011010",
  44250=>"001000010",
  44251=>"001000101",
  44252=>"000111111",
  44253=>"011101110",
  44254=>"110110001",
  44255=>"010111100",
  44256=>"111001100",
  44257=>"110010010",
  44258=>"110001001",
  44259=>"010110110",
  44260=>"111101110",
  44261=>"110101111",
  44262=>"111001100",
  44263=>"011100101",
  44264=>"001111110",
  44265=>"011010000",
  44266=>"001111000",
  44267=>"010000011",
  44268=>"100110100",
  44269=>"100001110",
  44270=>"001000001",
  44271=>"000000000",
  44272=>"001011101",
  44273=>"101011100",
  44274=>"000101111",
  44275=>"101011011",
  44276=>"111101000",
  44277=>"000101100",
  44278=>"011110010",
  44279=>"000100011",
  44280=>"001001010",
  44281=>"011001000",
  44282=>"000111110",
  44283=>"000010011",
  44284=>"011111001",
  44285=>"101000001",
  44286=>"111000010",
  44287=>"111111001",
  44288=>"111010100",
  44289=>"101101100",
  44290=>"101111001",
  44291=>"001110100",
  44292=>"000000100",
  44293=>"010101000",
  44294=>"111111101",
  44295=>"010000101",
  44296=>"100110010",
  44297=>"101110111",
  44298=>"101101111",
  44299=>"010100110",
  44300=>"001101010",
  44301=>"011101100",
  44302=>"100100100",
  44303=>"011011111",
  44304=>"001110011",
  44305=>"111000011",
  44306=>"110101110",
  44307=>"011110000",
  44308=>"001011111",
  44309=>"111001101",
  44310=>"011010011",
  44311=>"100111010",
  44312=>"110101110",
  44313=>"001100100",
  44314=>"100010100",
  44315=>"101000011",
  44316=>"000001010",
  44317=>"110110001",
  44318=>"010000010",
  44319=>"011010101",
  44320=>"101011010",
  44321=>"110000110",
  44322=>"111000000",
  44323=>"010110110",
  44324=>"011011000",
  44325=>"101001100",
  44326=>"011010111",
  44327=>"101100110",
  44328=>"000001001",
  44329=>"001010100",
  44330=>"111011110",
  44331=>"111110011",
  44332=>"100001001",
  44333=>"110000110",
  44334=>"101000010",
  44335=>"001111000",
  44336=>"001010101",
  44337=>"111110110",
  44338=>"010001000",
  44339=>"100010100",
  44340=>"110111000",
  44341=>"000000010",
  44342=>"010101100",
  44343=>"100100110",
  44344=>"100011110",
  44345=>"000000110",
  44346=>"101000100",
  44347=>"000000000",
  44348=>"110111000",
  44349=>"100000011",
  44350=>"000000110",
  44351=>"000011100",
  44352=>"010001110",
  44353=>"011000011",
  44354=>"000101010",
  44355=>"100011000",
  44356=>"110011110",
  44357=>"011101000",
  44358=>"100001000",
  44359=>"011111010",
  44360=>"010010011",
  44361=>"001000011",
  44362=>"000110100",
  44363=>"001101110",
  44364=>"111010001",
  44365=>"111000111",
  44366=>"101100010",
  44367=>"100111001",
  44368=>"101010000",
  44369=>"001110000",
  44370=>"110110011",
  44371=>"010101011",
  44372=>"011001010",
  44373=>"001011000",
  44374=>"001111111",
  44375=>"111111111",
  44376=>"001101000",
  44377=>"000111011",
  44378=>"110101100",
  44379=>"100000011",
  44380=>"000101111",
  44381=>"001101000",
  44382=>"111000010",
  44383=>"001000111",
  44384=>"000111111",
  44385=>"111011010",
  44386=>"001001110",
  44387=>"001100000",
  44388=>"000010101",
  44389=>"100111101",
  44390=>"111111110",
  44391=>"000100000",
  44392=>"001100011",
  44393=>"111100001",
  44394=>"111101000",
  44395=>"100101101",
  44396=>"101100101",
  44397=>"111100110",
  44398=>"011011100",
  44399=>"011011100",
  44400=>"101000011",
  44401=>"101010100",
  44402=>"111101000",
  44403=>"001000111",
  44404=>"001010111",
  44405=>"011111010",
  44406=>"101001010",
  44407=>"001010001",
  44408=>"010000110",
  44409=>"111011101",
  44410=>"110011001",
  44411=>"001011110",
  44412=>"111101100",
  44413=>"111110110",
  44414=>"110101000",
  44415=>"001011010",
  44416=>"111000011",
  44417=>"011000100",
  44418=>"111001101",
  44419=>"000100010",
  44420=>"000011100",
  44421=>"000110110",
  44422=>"111110000",
  44423=>"001110100",
  44424=>"000001101",
  44425=>"111011100",
  44426=>"000111110",
  44427=>"100000101",
  44428=>"111111000",
  44429=>"101101111",
  44430=>"001000101",
  44431=>"101011100",
  44432=>"101001111",
  44433=>"011000011",
  44434=>"000111010",
  44435=>"011111110",
  44436=>"001001100",
  44437=>"101001101",
  44438=>"001110010",
  44439=>"000001001",
  44440=>"000001000",
  44441=>"010100101",
  44442=>"100010001",
  44443=>"100111001",
  44444=>"101101000",
  44445=>"100001111",
  44446=>"111010111",
  44447=>"010110111",
  44448=>"101100111",
  44449=>"000000010",
  44450=>"001001000",
  44451=>"111011000",
  44452=>"100011100",
  44453=>"000000000",
  44454=>"101011101",
  44455=>"111011001",
  44456=>"000000010",
  44457=>"011110110",
  44458=>"000001111",
  44459=>"100110110",
  44460=>"001000001",
  44461=>"010110101",
  44462=>"101001111",
  44463=>"110100111",
  44464=>"000101011",
  44465=>"110100110",
  44466=>"000011110",
  44467=>"001111111",
  44468=>"010000010",
  44469=>"110110110",
  44470=>"101000111",
  44471=>"100000110",
  44472=>"100000001",
  44473=>"101100100",
  44474=>"000011001",
  44475=>"010000000",
  44476=>"000001111",
  44477=>"011010110",
  44478=>"111000101",
  44479=>"110101000",
  44480=>"000001100",
  44481=>"000010000",
  44482=>"000011011",
  44483=>"000101001",
  44484=>"000001000",
  44485=>"011001101",
  44486=>"010001111",
  44487=>"000100000",
  44488=>"000000010",
  44489=>"001010101",
  44490=>"111000010",
  44491=>"001010100",
  44492=>"111101010",
  44493=>"001111111",
  44494=>"001000001",
  44495=>"010111100",
  44496=>"001111111",
  44497=>"001110011",
  44498=>"111101100",
  44499=>"100010000",
  44500=>"000001101",
  44501=>"011010001",
  44502=>"101000101",
  44503=>"000010101",
  44504=>"110011100",
  44505=>"001111000",
  44506=>"110111001",
  44507=>"111001000",
  44508=>"000100100",
  44509=>"110111001",
  44510=>"101011101",
  44511=>"011001011",
  44512=>"010001100",
  44513=>"001010000",
  44514=>"100110010",
  44515=>"110101110",
  44516=>"100110001",
  44517=>"001101001",
  44518=>"000100111",
  44519=>"000001111",
  44520=>"011101110",
  44521=>"110000111",
  44522=>"101110000",
  44523=>"100000101",
  44524=>"010000000",
  44525=>"010010001",
  44526=>"000100010",
  44527=>"001111000",
  44528=>"010000011",
  44529=>"100101101",
  44530=>"011010111",
  44531=>"000100011",
  44532=>"100000110",
  44533=>"010001000",
  44534=>"011001000",
  44535=>"011100010",
  44536=>"000100000",
  44537=>"110110111",
  44538=>"000111011",
  44539=>"110010100",
  44540=>"001101011",
  44541=>"000001011",
  44542=>"110110001",
  44543=>"001110111",
  44544=>"010000101",
  44545=>"111011101",
  44546=>"111100100",
  44547=>"000000000",
  44548=>"001111000",
  44549=>"001001010",
  44550=>"100000001",
  44551=>"011110111",
  44552=>"001011010",
  44553=>"000011010",
  44554=>"000110100",
  44555=>"101101101",
  44556=>"110001001",
  44557=>"000010000",
  44558=>"100111100",
  44559=>"010110000",
  44560=>"100000010",
  44561=>"000011110",
  44562=>"010011010",
  44563=>"001011110",
  44564=>"100101010",
  44565=>"100000010",
  44566=>"110010100",
  44567=>"111010111",
  44568=>"100100100",
  44569=>"100000010",
  44570=>"010000011",
  44571=>"111001001",
  44572=>"011000110",
  44573=>"011101000",
  44574=>"110001101",
  44575=>"101010001",
  44576=>"011111110",
  44577=>"010000010",
  44578=>"000000110",
  44579=>"000010101",
  44580=>"010010011",
  44581=>"110000001",
  44582=>"101101100",
  44583=>"101000111",
  44584=>"001101010",
  44585=>"001011100",
  44586=>"000100011",
  44587=>"011011101",
  44588=>"101011110",
  44589=>"101111001",
  44590=>"101111110",
  44591=>"000101000",
  44592=>"100100001",
  44593=>"010000111",
  44594=>"110111010",
  44595=>"110000010",
  44596=>"100100101",
  44597=>"000111000",
  44598=>"011000111",
  44599=>"011000010",
  44600=>"010110010",
  44601=>"011100100",
  44602=>"000111010",
  44603=>"100101111",
  44604=>"000110000",
  44605=>"111011011",
  44606=>"010000101",
  44607=>"101001100",
  44608=>"000011010",
  44609=>"000001100",
  44610=>"001110000",
  44611=>"010111101",
  44612=>"001101110",
  44613=>"110011110",
  44614=>"100010101",
  44615=>"110111011",
  44616=>"001000110",
  44617=>"000100011",
  44618=>"101111100",
  44619=>"001110101",
  44620=>"010101101",
  44621=>"100101101",
  44622=>"100101101",
  44623=>"001111010",
  44624=>"010011111",
  44625=>"100001001",
  44626=>"010111101",
  44627=>"010000111",
  44628=>"111101010",
  44629=>"111101101",
  44630=>"110101011",
  44631=>"010000110",
  44632=>"101111111",
  44633=>"111000100",
  44634=>"000011111",
  44635=>"001101100",
  44636=>"010000100",
  44637=>"111100001",
  44638=>"101000001",
  44639=>"110011100",
  44640=>"111000101",
  44641=>"100111001",
  44642=>"100001101",
  44643=>"001100001",
  44644=>"011010000",
  44645=>"000000000",
  44646=>"001111100",
  44647=>"010101111",
  44648=>"011000001",
  44649=>"011011110",
  44650=>"000100101",
  44651=>"001101110",
  44652=>"001011101",
  44653=>"110111011",
  44654=>"111010110",
  44655=>"010111101",
  44656=>"000010000",
  44657=>"000010010",
  44658=>"110001011",
  44659=>"000010000",
  44660=>"001000000",
  44661=>"010110010",
  44662=>"101110011",
  44663=>"100011101",
  44664=>"000001100",
  44665=>"100101100",
  44666=>"001010000",
  44667=>"110101110",
  44668=>"111001100",
  44669=>"010001001",
  44670=>"101110000",
  44671=>"100000101",
  44672=>"101101101",
  44673=>"001100011",
  44674=>"101001001",
  44675=>"010000000",
  44676=>"000010100",
  44677=>"010001000",
  44678=>"011110100",
  44679=>"011010001",
  44680=>"000100001",
  44681=>"111010111",
  44682=>"010111100",
  44683=>"100110101",
  44684=>"010111011",
  44685=>"111100101",
  44686=>"111110100",
  44687=>"000100000",
  44688=>"010000110",
  44689=>"111100010",
  44690=>"111101000",
  44691=>"001000001",
  44692=>"010010101",
  44693=>"010011100",
  44694=>"000011101",
  44695=>"110100001",
  44696=>"001100111",
  44697=>"110101001",
  44698=>"110011100",
  44699=>"111000111",
  44700=>"111011011",
  44701=>"011101111",
  44702=>"110100110",
  44703=>"000111011",
  44704=>"110110111",
  44705=>"111000100",
  44706=>"101101100",
  44707=>"101001011",
  44708=>"111000101",
  44709=>"101010000",
  44710=>"000100110",
  44711=>"000011111",
  44712=>"010010010",
  44713=>"000100000",
  44714=>"111000101",
  44715=>"001000111",
  44716=>"110111010",
  44717=>"010010001",
  44718=>"110101000",
  44719=>"101011101",
  44720=>"000000111",
  44721=>"101101101",
  44722=>"101111000",
  44723=>"110000001",
  44724=>"010101100",
  44725=>"110001011",
  44726=>"101011111",
  44727=>"000001100",
  44728=>"110111000",
  44729=>"101000001",
  44730=>"101111100",
  44731=>"110001101",
  44732=>"001111001",
  44733=>"000010010",
  44734=>"000000000",
  44735=>"010101010",
  44736=>"010101011",
  44737=>"110111110",
  44738=>"011110011",
  44739=>"100000101",
  44740=>"000111100",
  44741=>"110011101",
  44742=>"011101011",
  44743=>"110011000",
  44744=>"010111100",
  44745=>"101100101",
  44746=>"100111001",
  44747=>"000010011",
  44748=>"001010000",
  44749=>"110110110",
  44750=>"111000000",
  44751=>"011011000",
  44752=>"011111101",
  44753=>"101000111",
  44754=>"110111101",
  44755=>"000111111",
  44756=>"001001001",
  44757=>"111010000",
  44758=>"000111111",
  44759=>"100011100",
  44760=>"000110111",
  44761=>"100111011",
  44762=>"100111110",
  44763=>"111110011",
  44764=>"010001000",
  44765=>"000000010",
  44766=>"010110101",
  44767=>"010001000",
  44768=>"000010010",
  44769=>"100000001",
  44770=>"000000110",
  44771=>"111011111",
  44772=>"000101111",
  44773=>"111101101",
  44774=>"101011100",
  44775=>"000000101",
  44776=>"010001010",
  44777=>"001001000",
  44778=>"101010100",
  44779=>"011101110",
  44780=>"001000010",
  44781=>"101111101",
  44782=>"010110001",
  44783=>"010000010",
  44784=>"000110110",
  44785=>"110011001",
  44786=>"110011100",
  44787=>"101010001",
  44788=>"010001010",
  44789=>"001110010",
  44790=>"001011111",
  44791=>"001101010",
  44792=>"001101001",
  44793=>"110010110",
  44794=>"100010011",
  44795=>"110100111",
  44796=>"010100011",
  44797=>"010111101",
  44798=>"100001000",
  44799=>"010001111",
  44800=>"111011100",
  44801=>"010001000",
  44802=>"010000001",
  44803=>"000111100",
  44804=>"001111000",
  44805=>"110101010",
  44806=>"101001101",
  44807=>"111001011",
  44808=>"001101101",
  44809=>"110100000",
  44810=>"101010000",
  44811=>"000101110",
  44812=>"111011100",
  44813=>"000000110",
  44814=>"011100110",
  44815=>"111001101",
  44816=>"111111000",
  44817=>"011001111",
  44818=>"001001001",
  44819=>"100100000",
  44820=>"100100110",
  44821=>"100000111",
  44822=>"110010010",
  44823=>"000100100",
  44824=>"011001000",
  44825=>"100111001",
  44826=>"000000101",
  44827=>"101101000",
  44828=>"011110100",
  44829=>"000010100",
  44830=>"000110100",
  44831=>"111111000",
  44832=>"100111101",
  44833=>"101010111",
  44834=>"000000101",
  44835=>"001011100",
  44836=>"010010010",
  44837=>"011101001",
  44838=>"001010100",
  44839=>"011000111",
  44840=>"000010011",
  44841=>"101110011",
  44842=>"101101000",
  44843=>"101000111",
  44844=>"011101100",
  44845=>"000010010",
  44846=>"000011000",
  44847=>"001101100",
  44848=>"011011011",
  44849=>"100101011",
  44850=>"010010000",
  44851=>"100000000",
  44852=>"010110011",
  44853=>"011101101",
  44854=>"110110111",
  44855=>"110000011",
  44856=>"100000010",
  44857=>"000000010",
  44858=>"000000110",
  44859=>"010100010",
  44860=>"011110011",
  44861=>"001101110",
  44862=>"101011000",
  44863=>"010011100",
  44864=>"100000000",
  44865=>"010001010",
  44866=>"110101001",
  44867=>"100011111",
  44868=>"101110001",
  44869=>"110001101",
  44870=>"101001100",
  44871=>"011000001",
  44872=>"110011110",
  44873=>"000111001",
  44874=>"110000001",
  44875=>"010001000",
  44876=>"011010110",
  44877=>"000011011",
  44878=>"011101101",
  44879=>"110101101",
  44880=>"101100001",
  44881=>"111101110",
  44882=>"011001001",
  44883=>"010010011",
  44884=>"000010110",
  44885=>"100110101",
  44886=>"001101110",
  44887=>"111111010",
  44888=>"110000000",
  44889=>"100001011",
  44890=>"011010010",
  44891=>"010111101",
  44892=>"010000110",
  44893=>"010010101",
  44894=>"011011001",
  44895=>"000100101",
  44896=>"011111100",
  44897=>"101100001",
  44898=>"100001101",
  44899=>"111011101",
  44900=>"000100011",
  44901=>"000000010",
  44902=>"000110100",
  44903=>"011001010",
  44904=>"000110101",
  44905=>"110111010",
  44906=>"000110000",
  44907=>"010111110",
  44908=>"100011100",
  44909=>"010000000",
  44910=>"110101101",
  44911=>"011010110",
  44912=>"010100110",
  44913=>"011001011",
  44914=>"010110101",
  44915=>"001000100",
  44916=>"101010001",
  44917=>"110110100",
  44918=>"100001000",
  44919=>"000100100",
  44920=>"000000100",
  44921=>"001001011",
  44922=>"100010000",
  44923=>"111101000",
  44924=>"010110001",
  44925=>"101110110",
  44926=>"111101100",
  44927=>"000010100",
  44928=>"000000010",
  44929=>"010101101",
  44930=>"001101010",
  44931=>"001011110",
  44932=>"000001100",
  44933=>"111111011",
  44934=>"011000010",
  44935=>"000010000",
  44936=>"000100001",
  44937=>"100100000",
  44938=>"000001010",
  44939=>"100111100",
  44940=>"000101010",
  44941=>"111101110",
  44942=>"001000101",
  44943=>"100000001",
  44944=>"110100000",
  44945=>"000001011",
  44946=>"100000001",
  44947=>"100110011",
  44948=>"101001010",
  44949=>"001100001",
  44950=>"010010011",
  44951=>"111011111",
  44952=>"101111111",
  44953=>"100100101",
  44954=>"011001100",
  44955=>"000010000",
  44956=>"111010010",
  44957=>"011010111",
  44958=>"101101110",
  44959=>"001011111",
  44960=>"000001100",
  44961=>"010101000",
  44962=>"010110101",
  44963=>"000001010",
  44964=>"000011100",
  44965=>"010010000",
  44966=>"010100000",
  44967=>"000001010",
  44968=>"001000111",
  44969=>"100100001",
  44970=>"110100001",
  44971=>"111100011",
  44972=>"011000011",
  44973=>"010100000",
  44974=>"100100110",
  44975=>"111000100",
  44976=>"011000001",
  44977=>"111100000",
  44978=>"000101100",
  44979=>"001000000",
  44980=>"001010010",
  44981=>"000111001",
  44982=>"000001011",
  44983=>"010100110",
  44984=>"011001100",
  44985=>"101100011",
  44986=>"110101110",
  44987=>"100111100",
  44988=>"101101001",
  44989=>"010001000",
  44990=>"111110110",
  44991=>"100001101",
  44992=>"110111001",
  44993=>"010010001",
  44994=>"010110010",
  44995=>"101101000",
  44996=>"100001100",
  44997=>"111101100",
  44998=>"101000010",
  44999=>"000100100",
  45000=>"100010001",
  45001=>"100101101",
  45002=>"111011111",
  45003=>"101111111",
  45004=>"100001101",
  45005=>"110010011",
  45006=>"100111010",
  45007=>"000000101",
  45008=>"100110110",
  45009=>"101001101",
  45010=>"010001101",
  45011=>"000010101",
  45012=>"101111101",
  45013=>"011000111",
  45014=>"010100101",
  45015=>"010010001",
  45016=>"111101111",
  45017=>"110110111",
  45018=>"010010111",
  45019=>"010110110",
  45020=>"101100100",
  45021=>"011100110",
  45022=>"110100110",
  45023=>"101010011",
  45024=>"000010000",
  45025=>"001001101",
  45026=>"001101101",
  45027=>"000011000",
  45028=>"000001001",
  45029=>"000101111",
  45030=>"000101111",
  45031=>"110111001",
  45032=>"011010110",
  45033=>"001000101",
  45034=>"100011111",
  45035=>"010011101",
  45036=>"101110100",
  45037=>"111010011",
  45038=>"001000110",
  45039=>"010011011",
  45040=>"001100001",
  45041=>"011011001",
  45042=>"111111011",
  45043=>"110000011",
  45044=>"100101011",
  45045=>"010100111",
  45046=>"111010000",
  45047=>"100010001",
  45048=>"000100101",
  45049=>"100000101",
  45050=>"110010000",
  45051=>"101010001",
  45052=>"000100001",
  45053=>"000011101",
  45054=>"000010101",
  45055=>"110000110",
  45056=>"101001111",
  45057=>"001000110",
  45058=>"100001011",
  45059=>"111001110",
  45060=>"100110011",
  45061=>"100100100",
  45062=>"100010000",
  45063=>"110110101",
  45064=>"011001101",
  45065=>"110011110",
  45066=>"111010001",
  45067=>"000010101",
  45068=>"101101100",
  45069=>"011111111",
  45070=>"010001011",
  45071=>"111101110",
  45072=>"010010001",
  45073=>"001101110",
  45074=>"001011111",
  45075=>"101110100",
  45076=>"111101010",
  45077=>"110100101",
  45078=>"000001100",
  45079=>"111100100",
  45080=>"000101100",
  45081=>"111101000",
  45082=>"100101000",
  45083=>"000111001",
  45084=>"000110010",
  45085=>"111011001",
  45086=>"001011110",
  45087=>"111011100",
  45088=>"100101101",
  45089=>"011000000",
  45090=>"101011101",
  45091=>"110110011",
  45092=>"100111101",
  45093=>"100001011",
  45094=>"100010100",
  45095=>"000100100",
  45096=>"110001100",
  45097=>"111101001",
  45098=>"100101010",
  45099=>"110001010",
  45100=>"000000100",
  45101=>"100000110",
  45102=>"100101100",
  45103=>"011111000",
  45104=>"001001010",
  45105=>"101000011",
  45106=>"011001111",
  45107=>"101010110",
  45108=>"111101110",
  45109=>"110100000",
  45110=>"000101110",
  45111=>"101011111",
  45112=>"100000010",
  45113=>"011100111",
  45114=>"011100110",
  45115=>"111000100",
  45116=>"101101001",
  45117=>"101000111",
  45118=>"011011000",
  45119=>"010001001",
  45120=>"011110110",
  45121=>"011111000",
  45122=>"010010100",
  45123=>"111111011",
  45124=>"000001000",
  45125=>"011100010",
  45126=>"001000010",
  45127=>"000101110",
  45128=>"101101111",
  45129=>"000001011",
  45130=>"111011010",
  45131=>"001010010",
  45132=>"110010001",
  45133=>"000100000",
  45134=>"011010001",
  45135=>"001111111",
  45136=>"101000100",
  45137=>"000010010",
  45138=>"010010100",
  45139=>"110000111",
  45140=>"010101010",
  45141=>"100111001",
  45142=>"110100001",
  45143=>"010000001",
  45144=>"011000010",
  45145=>"010000000",
  45146=>"000100010",
  45147=>"101101001",
  45148=>"000110001",
  45149=>"000010111",
  45150=>"101110101",
  45151=>"000101001",
  45152=>"001010001",
  45153=>"101101001",
  45154=>"010001010",
  45155=>"010101001",
  45156=>"101101000",
  45157=>"001011101",
  45158=>"100100100",
  45159=>"110011100",
  45160=>"111001101",
  45161=>"011111100",
  45162=>"111000100",
  45163=>"101100100",
  45164=>"001000101",
  45165=>"100000100",
  45166=>"011000100",
  45167=>"010001000",
  45168=>"110100010",
  45169=>"001011011",
  45170=>"001001001",
  45171=>"110100001",
  45172=>"000010101",
  45173=>"000100111",
  45174=>"111111110",
  45175=>"011001111",
  45176=>"100010101",
  45177=>"000110001",
  45178=>"111101111",
  45179=>"101101110",
  45180=>"101010100",
  45181=>"000011110",
  45182=>"011000010",
  45183=>"011000010",
  45184=>"011010111",
  45185=>"110111110",
  45186=>"100011010",
  45187=>"100100000",
  45188=>"000001100",
  45189=>"110111001",
  45190=>"111001101",
  45191=>"111000011",
  45192=>"101001101",
  45193=>"001101001",
  45194=>"100100000",
  45195=>"000000111",
  45196=>"000001001",
  45197=>"110111101",
  45198=>"110001000",
  45199=>"011000111",
  45200=>"110011000",
  45201=>"101000000",
  45202=>"010001000",
  45203=>"001001010",
  45204=>"000010100",
  45205=>"101011100",
  45206=>"001101010",
  45207=>"101100010",
  45208=>"110000011",
  45209=>"100100110",
  45210=>"000010010",
  45211=>"100011001",
  45212=>"001011011",
  45213=>"100110110",
  45214=>"010110110",
  45215=>"000010110",
  45216=>"000110001",
  45217=>"101001010",
  45218=>"000110111",
  45219=>"010011011",
  45220=>"100100000",
  45221=>"100011001",
  45222=>"000000100",
  45223=>"010100110",
  45224=>"010011001",
  45225=>"100100000",
  45226=>"011100000",
  45227=>"000000110",
  45228=>"101100100",
  45229=>"111011101",
  45230=>"001101110",
  45231=>"111000111",
  45232=>"101100001",
  45233=>"100010001",
  45234=>"101101101",
  45235=>"000000000",
  45236=>"011010001",
  45237=>"111111101",
  45238=>"010111100",
  45239=>"100000100",
  45240=>"111001011",
  45241=>"010001001",
  45242=>"010000000",
  45243=>"100000101",
  45244=>"010010000",
  45245=>"010110000",
  45246=>"101101101",
  45247=>"110100010",
  45248=>"000101000",
  45249=>"010101000",
  45250=>"110110111",
  45251=>"010001110",
  45252=>"101010000",
  45253=>"010000111",
  45254=>"110001101",
  45255=>"000000010",
  45256=>"101011100",
  45257=>"100000100",
  45258=>"001110010",
  45259=>"100011011",
  45260=>"000100010",
  45261=>"101100111",
  45262=>"000111110",
  45263=>"011100100",
  45264=>"000010010",
  45265=>"010100110",
  45266=>"001001010",
  45267=>"010111100",
  45268=>"100111100",
  45269=>"011101011",
  45270=>"001000101",
  45271=>"011110101",
  45272=>"111101010",
  45273=>"101110010",
  45274=>"100110101",
  45275=>"111001101",
  45276=>"000101100",
  45277=>"110001001",
  45278=>"111000101",
  45279=>"001010111",
  45280=>"101011001",
  45281=>"001110001",
  45282=>"100110000",
  45283=>"101010000",
  45284=>"100001001",
  45285=>"101001101",
  45286=>"011001011",
  45287=>"101111001",
  45288=>"010010000",
  45289=>"000100111",
  45290=>"111111101",
  45291=>"000100111",
  45292=>"110110001",
  45293=>"100000011",
  45294=>"000100011",
  45295=>"001000000",
  45296=>"001110000",
  45297=>"001011011",
  45298=>"101100100",
  45299=>"011010110",
  45300=>"010001110",
  45301=>"111100000",
  45302=>"010011001",
  45303=>"001001001",
  45304=>"000111001",
  45305=>"011111111",
  45306=>"101100011",
  45307=>"101001001",
  45308=>"000101000",
  45309=>"000100111",
  45310=>"100011100",
  45311=>"100101100",
  45312=>"110100010",
  45313=>"110000100",
  45314=>"001001110",
  45315=>"111000000",
  45316=>"000111011",
  45317=>"000011001",
  45318=>"001110000",
  45319=>"101111011",
  45320=>"111100010",
  45321=>"010001010",
  45322=>"001110000",
  45323=>"001001101",
  45324=>"001000111",
  45325=>"000101010",
  45326=>"001110011",
  45327=>"010111011",
  45328=>"110010101",
  45329=>"001010000",
  45330=>"001001100",
  45331=>"011001001",
  45332=>"100110001",
  45333=>"100101111",
  45334=>"011001101",
  45335=>"110000101",
  45336=>"111100111",
  45337=>"100010001",
  45338=>"101010101",
  45339=>"110111001",
  45340=>"100001000",
  45341=>"101010100",
  45342=>"011010000",
  45343=>"100011110",
  45344=>"110001101",
  45345=>"001001111",
  45346=>"010010110",
  45347=>"110111011",
  45348=>"101000011",
  45349=>"000111010",
  45350=>"110100101",
  45351=>"001101101",
  45352=>"100011101",
  45353=>"000100011",
  45354=>"111110010",
  45355=>"110101010",
  45356=>"001100000",
  45357=>"100001111",
  45358=>"110100000",
  45359=>"010100110",
  45360=>"001110110",
  45361=>"111111010",
  45362=>"011101011",
  45363=>"101101001",
  45364=>"000010001",
  45365=>"100110101",
  45366=>"001100011",
  45367=>"011100011",
  45368=>"111001000",
  45369=>"011110000",
  45370=>"111011010",
  45371=>"001010111",
  45372=>"011100010",
  45373=>"101110101",
  45374=>"111111100",
  45375=>"111111111",
  45376=>"011001001",
  45377=>"100010110",
  45378=>"101001011",
  45379=>"101100001",
  45380=>"010100100",
  45381=>"110100011",
  45382=>"000000111",
  45383=>"100101000",
  45384=>"101011010",
  45385=>"100011010",
  45386=>"100000011",
  45387=>"000110101",
  45388=>"000011100",
  45389=>"101100010",
  45390=>"100010010",
  45391=>"010001111",
  45392=>"001001000",
  45393=>"001100110",
  45394=>"001000110",
  45395=>"110100011",
  45396=>"101001001",
  45397=>"000011000",
  45398=>"000001001",
  45399=>"010001010",
  45400=>"010101000",
  45401=>"100010001",
  45402=>"100110000",
  45403=>"101010001",
  45404=>"110001001",
  45405=>"011111001",
  45406=>"000101000",
  45407=>"011110011",
  45408=>"100011110",
  45409=>"010001011",
  45410=>"111110001",
  45411=>"101010111",
  45412=>"100011001",
  45413=>"000010011",
  45414=>"000011101",
  45415=>"100111111",
  45416=>"001000001",
  45417=>"111100100",
  45418=>"101101010",
  45419=>"100111011",
  45420=>"010010110",
  45421=>"000111011",
  45422=>"000100010",
  45423=>"101111011",
  45424=>"000111101",
  45425=>"100010010",
  45426=>"110110101",
  45427=>"000111000",
  45428=>"101000101",
  45429=>"111011010",
  45430=>"111111111",
  45431=>"111001110",
  45432=>"111101000",
  45433=>"011000101",
  45434=>"100011110",
  45435=>"001100001",
  45436=>"011010010",
  45437=>"111001100",
  45438=>"010001010",
  45439=>"100101010",
  45440=>"100010100",
  45441=>"111111001",
  45442=>"111100010",
  45443=>"101011000",
  45444=>"111000001",
  45445=>"000001000",
  45446=>"000101001",
  45447=>"111011101",
  45448=>"101111100",
  45449=>"100011000",
  45450=>"000010011",
  45451=>"111111011",
  45452=>"000111100",
  45453=>"110111001",
  45454=>"000011011",
  45455=>"010111101",
  45456=>"011110111",
  45457=>"011100111",
  45458=>"001011100",
  45459=>"010010110",
  45460=>"101111111",
  45461=>"101000111",
  45462=>"110111011",
  45463=>"111110001",
  45464=>"000000101",
  45465=>"101110100",
  45466=>"011101100",
  45467=>"101011010",
  45468=>"000001110",
  45469=>"101111100",
  45470=>"000100001",
  45471=>"001110101",
  45472=>"011110110",
  45473=>"111000011",
  45474=>"001101011",
  45475=>"111100100",
  45476=>"000011111",
  45477=>"001000010",
  45478=>"000110110",
  45479=>"111011001",
  45480=>"100101011",
  45481=>"111011110",
  45482=>"110100000",
  45483=>"011101111",
  45484=>"101001111",
  45485=>"000110111",
  45486=>"000101010",
  45487=>"000011101",
  45488=>"101111101",
  45489=>"100110111",
  45490=>"100001001",
  45491=>"001101001",
  45492=>"111010000",
  45493=>"101011100",
  45494=>"001001100",
  45495=>"110010010",
  45496=>"000111001",
  45497=>"011110111",
  45498=>"010000001",
  45499=>"011001100",
  45500=>"111110010",
  45501=>"100110100",
  45502=>"000111100",
  45503=>"000111101",
  45504=>"010001110",
  45505=>"110111010",
  45506=>"001111111",
  45507=>"101111111",
  45508=>"000001000",
  45509=>"010111000",
  45510=>"111000001",
  45511=>"100111110",
  45512=>"101010110",
  45513=>"111010010",
  45514=>"011101000",
  45515=>"001110011",
  45516=>"100100010",
  45517=>"111111011",
  45518=>"010010001",
  45519=>"011010000",
  45520=>"110111101",
  45521=>"101110001",
  45522=>"100010011",
  45523=>"000110111",
  45524=>"110001010",
  45525=>"000011110",
  45526=>"000100000",
  45527=>"100111100",
  45528=>"001111111",
  45529=>"001101001",
  45530=>"010100101",
  45531=>"111010111",
  45532=>"100111010",
  45533=>"111101110",
  45534=>"010111111",
  45535=>"110000100",
  45536=>"101001011",
  45537=>"010010111",
  45538=>"111110101",
  45539=>"001101101",
  45540=>"011010100",
  45541=>"000111000",
  45542=>"101010100",
  45543=>"011000100",
  45544=>"010110110",
  45545=>"001001000",
  45546=>"000010010",
  45547=>"111100000",
  45548=>"110110111",
  45549=>"011111000",
  45550=>"110010111",
  45551=>"011000001",
  45552=>"111001010",
  45553=>"110000111",
  45554=>"110010100",
  45555=>"011010000",
  45556=>"000110000",
  45557=>"011100010",
  45558=>"011100011",
  45559=>"111000011",
  45560=>"100101101",
  45561=>"001110001",
  45562=>"010011001",
  45563=>"111011000",
  45564=>"010011110",
  45565=>"011101110",
  45566=>"001111101",
  45567=>"111100100",
  45568=>"001001001",
  45569=>"111001001",
  45570=>"010100000",
  45571=>"011001111",
  45572=>"011011101",
  45573=>"101100110",
  45574=>"111000001",
  45575=>"101010010",
  45576=>"100000011",
  45577=>"100100111",
  45578=>"011010101",
  45579=>"100000010",
  45580=>"010001001",
  45581=>"101000010",
  45582=>"100101001",
  45583=>"000110011",
  45584=>"100000011",
  45585=>"010001000",
  45586=>"110101111",
  45587=>"111111010",
  45588=>"011001100",
  45589=>"011110100",
  45590=>"110000000",
  45591=>"001011011",
  45592=>"100011000",
  45593=>"001000001",
  45594=>"001001110",
  45595=>"010010010",
  45596=>"011000100",
  45597=>"011100111",
  45598=>"110100100",
  45599=>"010111111",
  45600=>"110000101",
  45601=>"010101101",
  45602=>"110111111",
  45603=>"111101001",
  45604=>"011111110",
  45605=>"111100101",
  45606=>"111010001",
  45607=>"100111101",
  45608=>"010001010",
  45609=>"110000011",
  45610=>"110001110",
  45611=>"000111100",
  45612=>"110001110",
  45613=>"110100011",
  45614=>"100101101",
  45615=>"101000001",
  45616=>"011111110",
  45617=>"111001110",
  45618=>"111010011",
  45619=>"101111000",
  45620=>"101100001",
  45621=>"001101000",
  45622=>"111000011",
  45623=>"101110010",
  45624=>"001000100",
  45625=>"010001110",
  45626=>"111010101",
  45627=>"101111010",
  45628=>"000001100",
  45629=>"000100001",
  45630=>"101111011",
  45631=>"101111100",
  45632=>"111101101",
  45633=>"001111100",
  45634=>"101010111",
  45635=>"111101010",
  45636=>"111111010",
  45637=>"011001011",
  45638=>"001110000",
  45639=>"000000001",
  45640=>"111000111",
  45641=>"100110010",
  45642=>"001011100",
  45643=>"100101000",
  45644=>"100101110",
  45645=>"010110000",
  45646=>"000010111",
  45647=>"001110100",
  45648=>"100111001",
  45649=>"110110100",
  45650=>"011101011",
  45651=>"110001000",
  45652=>"001111000",
  45653=>"000000010",
  45654=>"110000100",
  45655=>"101100100",
  45656=>"000111000",
  45657=>"010101000",
  45658=>"111101111",
  45659=>"000011100",
  45660=>"100110110",
  45661=>"100100010",
  45662=>"110000110",
  45663=>"110101001",
  45664=>"001111001",
  45665=>"011000101",
  45666=>"011010111",
  45667=>"011000111",
  45668=>"100010101",
  45669=>"101000111",
  45670=>"000110100",
  45671=>"000100011",
  45672=>"010000011",
  45673=>"111000010",
  45674=>"110000011",
  45675=>"111101110",
  45676=>"010001111",
  45677=>"001000001",
  45678=>"000000010",
  45679=>"100001011",
  45680=>"101101100",
  45681=>"110001110",
  45682=>"111010110",
  45683=>"111110011",
  45684=>"110000011",
  45685=>"010000011",
  45686=>"001101111",
  45687=>"010111111",
  45688=>"101101110",
  45689=>"111100010",
  45690=>"011111100",
  45691=>"001000110",
  45692=>"000001000",
  45693=>"111111100",
  45694=>"011100101",
  45695=>"100111101",
  45696=>"111100101",
  45697=>"100010110",
  45698=>"001001010",
  45699=>"011110111",
  45700=>"110100101",
  45701=>"101000110",
  45702=>"100001101",
  45703=>"010010001",
  45704=>"100000111",
  45705=>"100101110",
  45706=>"100000100",
  45707=>"011101100",
  45708=>"110001100",
  45709=>"000001100",
  45710=>"101100000",
  45711=>"011011100",
  45712=>"111111101",
  45713=>"111101100",
  45714=>"010101000",
  45715=>"101110111",
  45716=>"011010010",
  45717=>"001000011",
  45718=>"001101001",
  45719=>"011010110",
  45720=>"001110110",
  45721=>"000101110",
  45722=>"100100001",
  45723=>"001100011",
  45724=>"010101001",
  45725=>"001001100",
  45726=>"100110100",
  45727=>"110100000",
  45728=>"100110101",
  45729=>"111110011",
  45730=>"100001010",
  45731=>"010110010",
  45732=>"000010111",
  45733=>"111111110",
  45734=>"111101011",
  45735=>"100000000",
  45736=>"001001010",
  45737=>"110011010",
  45738=>"000110000",
  45739=>"001100100",
  45740=>"000101100",
  45741=>"001100110",
  45742=>"111001001",
  45743=>"011101011",
  45744=>"101010010",
  45745=>"100010111",
  45746=>"111011111",
  45747=>"110011011",
  45748=>"000011100",
  45749=>"000011101",
  45750=>"000110011",
  45751=>"111000101",
  45752=>"011001101",
  45753=>"000110001",
  45754=>"001001001",
  45755=>"010011000",
  45756=>"001111011",
  45757=>"011000110",
  45758=>"101111110",
  45759=>"111111010",
  45760=>"010100101",
  45761=>"001111001",
  45762=>"010000011",
  45763=>"000100001",
  45764=>"101110010",
  45765=>"101100001",
  45766=>"001010101",
  45767=>"010101101",
  45768=>"011001100",
  45769=>"101011010",
  45770=>"001110000",
  45771=>"100101101",
  45772=>"111010101",
  45773=>"000111100",
  45774=>"001001110",
  45775=>"001000000",
  45776=>"000001011",
  45777=>"101000110",
  45778=>"100100110",
  45779=>"011001000",
  45780=>"100001010",
  45781=>"111000101",
  45782=>"100001100",
  45783=>"110101010",
  45784=>"101000101",
  45785=>"001110110",
  45786=>"111100011",
  45787=>"111111010",
  45788=>"010100110",
  45789=>"101101000",
  45790=>"101101001",
  45791=>"100001011",
  45792=>"010101000",
  45793=>"011011000",
  45794=>"110000111",
  45795=>"010100111",
  45796=>"101000111",
  45797=>"010101011",
  45798=>"100010100",
  45799=>"110000101",
  45800=>"011000000",
  45801=>"101000110",
  45802=>"011000010",
  45803=>"111011000",
  45804=>"100101110",
  45805=>"000011100",
  45806=>"111011010",
  45807=>"010011011",
  45808=>"000111111",
  45809=>"000000010",
  45810=>"110010010",
  45811=>"001110011",
  45812=>"011111000",
  45813=>"011111001",
  45814=>"011011011",
  45815=>"000110000",
  45816=>"001011010",
  45817=>"010110100",
  45818=>"001100001",
  45819=>"010111100",
  45820=>"011110010",
  45821=>"000000001",
  45822=>"000001011",
  45823=>"110111111",
  45824=>"010110010",
  45825=>"111101110",
  45826=>"110101101",
  45827=>"110001010",
  45828=>"100110011",
  45829=>"010101100",
  45830=>"000111000",
  45831=>"110110111",
  45832=>"011100011",
  45833=>"101101001",
  45834=>"011010001",
  45835=>"110001101",
  45836=>"100101000",
  45837=>"000110111",
  45838=>"111101111",
  45839=>"000011111",
  45840=>"000101000",
  45841=>"011111100",
  45842=>"010001010",
  45843=>"100100010",
  45844=>"111000001",
  45845=>"010100000",
  45846=>"000000000",
  45847=>"000100010",
  45848=>"111010001",
  45849=>"111010010",
  45850=>"101010111",
  45851=>"110011101",
  45852=>"011110000",
  45853=>"010110110",
  45854=>"111001100",
  45855=>"100000000",
  45856=>"111010011",
  45857=>"101000101",
  45858=>"100110011",
  45859=>"010111011",
  45860=>"101100100",
  45861=>"000000010",
  45862=>"001011000",
  45863=>"110000110",
  45864=>"110000101",
  45865=>"010100001",
  45866=>"010111111",
  45867=>"111110011",
  45868=>"011110001",
  45869=>"000001010",
  45870=>"010101110",
  45871=>"101101010",
  45872=>"011000010",
  45873=>"000100000",
  45874=>"100110101",
  45875=>"101001100",
  45876=>"011000101",
  45877=>"100010110",
  45878=>"000101111",
  45879=>"010110010",
  45880=>"100010000",
  45881=>"110000110",
  45882=>"111110111",
  45883=>"101011111",
  45884=>"101000011",
  45885=>"010101101",
  45886=>"000000100",
  45887=>"111110111",
  45888=>"101011110",
  45889=>"110011001",
  45890=>"010000001",
  45891=>"011101111",
  45892=>"100001001",
  45893=>"011011001",
  45894=>"001001000",
  45895=>"110111111",
  45896=>"100110011",
  45897=>"000110101",
  45898=>"000100110",
  45899=>"001000001",
  45900=>"010010010",
  45901=>"110100000",
  45902=>"111100000",
  45903=>"100111001",
  45904=>"000000000",
  45905=>"101010101",
  45906=>"011110100",
  45907=>"100111000",
  45908=>"000100000",
  45909=>"100010001",
  45910=>"010011100",
  45911=>"100010000",
  45912=>"110110001",
  45913=>"011011111",
  45914=>"011111110",
  45915=>"001001100",
  45916=>"000011000",
  45917=>"110010110",
  45918=>"100000111",
  45919=>"000000011",
  45920=>"011110010",
  45921=>"111110110",
  45922=>"010001010",
  45923=>"011001100",
  45924=>"010101011",
  45925=>"000111001",
  45926=>"100000111",
  45927=>"010101111",
  45928=>"001010111",
  45929=>"011110001",
  45930=>"101111110",
  45931=>"011110101",
  45932=>"110011001",
  45933=>"001111000",
  45934=>"010011011",
  45935=>"001100010",
  45936=>"001101101",
  45937=>"111111100",
  45938=>"000010111",
  45939=>"011111110",
  45940=>"101010000",
  45941=>"000011101",
  45942=>"000001101",
  45943=>"011011100",
  45944=>"011010100",
  45945=>"010110101",
  45946=>"110000111",
  45947=>"010110010",
  45948=>"111100100",
  45949=>"000011000",
  45950=>"001010010",
  45951=>"100001010",
  45952=>"111101001",
  45953=>"110110110",
  45954=>"110111110",
  45955=>"000111010",
  45956=>"010011010",
  45957=>"000110001",
  45958=>"100101110",
  45959=>"101110010",
  45960=>"101011011",
  45961=>"011000100",
  45962=>"001000101",
  45963=>"000001000",
  45964=>"011101110",
  45965=>"101111011",
  45966=>"010101111",
  45967=>"100101110",
  45968=>"111001111",
  45969=>"111100110",
  45970=>"011101100",
  45971=>"111000110",
  45972=>"110000110",
  45973=>"110111111",
  45974=>"101101100",
  45975=>"101010100",
  45976=>"110111000",
  45977=>"010100101",
  45978=>"111111111",
  45979=>"101010011",
  45980=>"011011110",
  45981=>"010011000",
  45982=>"011101001",
  45983=>"010110110",
  45984=>"001101010",
  45985=>"000101010",
  45986=>"111010111",
  45987=>"010101000",
  45988=>"001000100",
  45989=>"100101101",
  45990=>"001101011",
  45991=>"111101101",
  45992=>"111011111",
  45993=>"111111111",
  45994=>"010110010",
  45995=>"001101010",
  45996=>"001000111",
  45997=>"011110001",
  45998=>"111011110",
  45999=>"111111101",
  46000=>"101101001",
  46001=>"001001100",
  46002=>"011000001",
  46003=>"101110010",
  46004=>"110010010",
  46005=>"110110001",
  46006=>"101011001",
  46007=>"010000011",
  46008=>"111100110",
  46009=>"101110000",
  46010=>"011010101",
  46011=>"110100101",
  46012=>"001001011",
  46013=>"110101111",
  46014=>"100000000",
  46015=>"111111001",
  46016=>"100100111",
  46017=>"100111010",
  46018=>"101100010",
  46019=>"110111000",
  46020=>"100101011",
  46021=>"010101111",
  46022=>"010111101",
  46023=>"111010101",
  46024=>"000000010",
  46025=>"010101000",
  46026=>"100011000",
  46027=>"111100011",
  46028=>"101000000",
  46029=>"101000010",
  46030=>"111100101",
  46031=>"100000100",
  46032=>"010111111",
  46033=>"100001001",
  46034=>"101110100",
  46035=>"110000010",
  46036=>"000000100",
  46037=>"111000011",
  46038=>"101101011",
  46039=>"101100100",
  46040=>"001111100",
  46041=>"000001010",
  46042=>"101111010",
  46043=>"000000100",
  46044=>"110100001",
  46045=>"111011101",
  46046=>"110000000",
  46047=>"001000001",
  46048=>"100111010",
  46049=>"000100101",
  46050=>"010011101",
  46051=>"011000000",
  46052=>"101100000",
  46053=>"110001101",
  46054=>"100110000",
  46055=>"100010110",
  46056=>"001011000",
  46057=>"011101111",
  46058=>"001000101",
  46059=>"011001101",
  46060=>"001010011",
  46061=>"111000010",
  46062=>"111110001",
  46063=>"100011000",
  46064=>"100000110",
  46065=>"101000010",
  46066=>"010110110",
  46067=>"100011110",
  46068=>"111001100",
  46069=>"000000101",
  46070=>"011010101",
  46071=>"101010011",
  46072=>"010101010",
  46073=>"010010001",
  46074=>"000010101",
  46075=>"011011110",
  46076=>"001011001",
  46077=>"101010111",
  46078=>"101110000",
  46079=>"000000011",
  46080=>"110001111",
  46081=>"000001010",
  46082=>"010010001",
  46083=>"011010001",
  46084=>"100100001",
  46085=>"001010100",
  46086=>"110110110",
  46087=>"111010000",
  46088=>"011101111",
  46089=>"001100100",
  46090=>"010110000",
  46091=>"111111001",
  46092=>"011000010",
  46093=>"111101110",
  46094=>"010001000",
  46095=>"111101010",
  46096=>"010100010",
  46097=>"011011010",
  46098=>"001111100",
  46099=>"111011011",
  46100=>"000110100",
  46101=>"110100111",
  46102=>"000011100",
  46103=>"011100000",
  46104=>"011000101",
  46105=>"000001111",
  46106=>"011111010",
  46107=>"111001111",
  46108=>"101010000",
  46109=>"011111100",
  46110=>"011101101",
  46111=>"010010000",
  46112=>"110111111",
  46113=>"001011011",
  46114=>"100001101",
  46115=>"001010000",
  46116=>"011110100",
  46117=>"011110110",
  46118=>"111110011",
  46119=>"110010010",
  46120=>"100110111",
  46121=>"101000111",
  46122=>"111100010",
  46123=>"010000101",
  46124=>"000111011",
  46125=>"011010111",
  46126=>"010100111",
  46127=>"010110010",
  46128=>"110001001",
  46129=>"000000000",
  46130=>"010001011",
  46131=>"100111100",
  46132=>"111001001",
  46133=>"111101000",
  46134=>"111001010",
  46135=>"001101000",
  46136=>"011000000",
  46137=>"101000101",
  46138=>"000111100",
  46139=>"100101010",
  46140=>"000110100",
  46141=>"100010111",
  46142=>"111101110",
  46143=>"110000011",
  46144=>"100000001",
  46145=>"101010000",
  46146=>"001001001",
  46147=>"111000110",
  46148=>"001011000",
  46149=>"111110100",
  46150=>"000010111",
  46151=>"100100000",
  46152=>"011110110",
  46153=>"100011111",
  46154=>"110010000",
  46155=>"001101000",
  46156=>"110110010",
  46157=>"111001111",
  46158=>"110000011",
  46159=>"111001001",
  46160=>"101010000",
  46161=>"111000010",
  46162=>"110011100",
  46163=>"110011111",
  46164=>"011111001",
  46165=>"101101000",
  46166=>"111100001",
  46167=>"111010000",
  46168=>"111100010",
  46169=>"100111000",
  46170=>"111001100",
  46171=>"011100010",
  46172=>"000010010",
  46173=>"101100111",
  46174=>"110101110",
  46175=>"110100000",
  46176=>"011001100",
  46177=>"010000000",
  46178=>"011111101",
  46179=>"100111110",
  46180=>"010100100",
  46181=>"111110101",
  46182=>"110101110",
  46183=>"100111000",
  46184=>"111011111",
  46185=>"001100011",
  46186=>"010111100",
  46187=>"111110001",
  46188=>"010101101",
  46189=>"101000101",
  46190=>"110010101",
  46191=>"110101010",
  46192=>"000000111",
  46193=>"011011010",
  46194=>"101101101",
  46195=>"111010011",
  46196=>"110010001",
  46197=>"101000010",
  46198=>"111110000",
  46199=>"111011010",
  46200=>"111111011",
  46201=>"010111111",
  46202=>"110100111",
  46203=>"010110011",
  46204=>"001011111",
  46205=>"100001001",
  46206=>"000000101",
  46207=>"111111001",
  46208=>"111000111",
  46209=>"111011110",
  46210=>"101110010",
  46211=>"110011000",
  46212=>"111001110",
  46213=>"001101011",
  46214=>"110111100",
  46215=>"111101110",
  46216=>"101111111",
  46217=>"111001010",
  46218=>"001100001",
  46219=>"010001001",
  46220=>"110101010",
  46221=>"100001001",
  46222=>"010001110",
  46223=>"111001000",
  46224=>"000011010",
  46225=>"010100110",
  46226=>"100011110",
  46227=>"010010001",
  46228=>"100011011",
  46229=>"111001000",
  46230=>"000010010",
  46231=>"111010111",
  46232=>"000001100",
  46233=>"111011111",
  46234=>"100010101",
  46235=>"010101101",
  46236=>"100111101",
  46237=>"111111010",
  46238=>"011011100",
  46239=>"111000011",
  46240=>"000111110",
  46241=>"000011101",
  46242=>"110100011",
  46243=>"001000010",
  46244=>"001010001",
  46245=>"001101010",
  46246=>"110001010",
  46247=>"001001010",
  46248=>"111000000",
  46249=>"001101000",
  46250=>"101011101",
  46251=>"000110100",
  46252=>"111110110",
  46253=>"111100011",
  46254=>"111000110",
  46255=>"110011011",
  46256=>"011000011",
  46257=>"001010111",
  46258=>"001011001",
  46259=>"000100001",
  46260=>"001001010",
  46261=>"111010010",
  46262=>"110011110",
  46263=>"100011100",
  46264=>"010001100",
  46265=>"011010100",
  46266=>"001110101",
  46267=>"010000011",
  46268=>"010110010",
  46269=>"000011000",
  46270=>"100100101",
  46271=>"000111011",
  46272=>"011000110",
  46273=>"010101010",
  46274=>"010011000",
  46275=>"110010101",
  46276=>"011000110",
  46277=>"011100000",
  46278=>"100011111",
  46279=>"011100111",
  46280=>"101111101",
  46281=>"110100001",
  46282=>"001100111",
  46283=>"001110001",
  46284=>"000011011",
  46285=>"010000100",
  46286=>"111010101",
  46287=>"101001001",
  46288=>"100110111",
  46289=>"101100101",
  46290=>"100001011",
  46291=>"111110000",
  46292=>"011000100",
  46293=>"001100010",
  46294=>"100001001",
  46295=>"101100110",
  46296=>"010111011",
  46297=>"010101111",
  46298=>"101000011",
  46299=>"011111100",
  46300=>"010100000",
  46301=>"101111101",
  46302=>"101100000",
  46303=>"100000011",
  46304=>"001101100",
  46305=>"011010101",
  46306=>"100000001",
  46307=>"000011010",
  46308=>"100000000",
  46309=>"001011000",
  46310=>"000101011",
  46311=>"110011010",
  46312=>"010000000",
  46313=>"111110110",
  46314=>"111110101",
  46315=>"110100011",
  46316=>"101010100",
  46317=>"100010101",
  46318=>"101111110",
  46319=>"000110000",
  46320=>"100111010",
  46321=>"101101111",
  46322=>"111111111",
  46323=>"111111011",
  46324=>"100011111",
  46325=>"101110001",
  46326=>"100000000",
  46327=>"111101111",
  46328=>"001001111",
  46329=>"111101010",
  46330=>"110111110",
  46331=>"001010100",
  46332=>"111010010",
  46333=>"110100010",
  46334=>"111010101",
  46335=>"010010110",
  46336=>"111011110",
  46337=>"010010110",
  46338=>"110110001",
  46339=>"010010001",
  46340=>"111110100",
  46341=>"010110110",
  46342=>"010110101",
  46343=>"001001111",
  46344=>"011001111",
  46345=>"110110001",
  46346=>"000111111",
  46347=>"111011000",
  46348=>"010111011",
  46349=>"011010010",
  46350=>"110000010",
  46351=>"110011110",
  46352=>"011110110",
  46353=>"100010100",
  46354=>"010001001",
  46355=>"111000011",
  46356=>"100000110",
  46357=>"101000001",
  46358=>"011111010",
  46359=>"110001011",
  46360=>"100010110",
  46361=>"011110110",
  46362=>"101111000",
  46363=>"101011110",
  46364=>"111110010",
  46365=>"001100110",
  46366=>"000100010",
  46367=>"000000111",
  46368=>"111101110",
  46369=>"011010011",
  46370=>"100010110",
  46371=>"101101000",
  46372=>"001000001",
  46373=>"011111010",
  46374=>"000110100",
  46375=>"101001001",
  46376=>"000011100",
  46377=>"010110110",
  46378=>"000110010",
  46379=>"101100110",
  46380=>"111000010",
  46381=>"111111001",
  46382=>"000000011",
  46383=>"011000100",
  46384=>"010001000",
  46385=>"010100001",
  46386=>"101110001",
  46387=>"111001000",
  46388=>"001100100",
  46389=>"001011001",
  46390=>"111001011",
  46391=>"111010011",
  46392=>"101000101",
  46393=>"110101010",
  46394=>"111010000",
  46395=>"001010010",
  46396=>"011010001",
  46397=>"001011100",
  46398=>"101110111",
  46399=>"111001100",
  46400=>"011011101",
  46401=>"011010111",
  46402=>"101100101",
  46403=>"011001100",
  46404=>"101011010",
  46405=>"000100010",
  46406=>"100000010",
  46407=>"110010011",
  46408=>"100001001",
  46409=>"101100101",
  46410=>"011101010",
  46411=>"010110001",
  46412=>"001000110",
  46413=>"000110101",
  46414=>"010101111",
  46415=>"001100000",
  46416=>"100001100",
  46417=>"100010100",
  46418=>"010110011",
  46419=>"111011011",
  46420=>"100100010",
  46421=>"100110010",
  46422=>"001000101",
  46423=>"100000001",
  46424=>"101101000",
  46425=>"010000010",
  46426=>"100101101",
  46427=>"010000100",
  46428=>"111110000",
  46429=>"000101011",
  46430=>"101110111",
  46431=>"000111010",
  46432=>"011000011",
  46433=>"001111111",
  46434=>"010001011",
  46435=>"011001000",
  46436=>"110010111",
  46437=>"101000011",
  46438=>"001000011",
  46439=>"101110000",
  46440=>"001011110",
  46441=>"001101010",
  46442=>"011010010",
  46443=>"110111110",
  46444=>"110110101",
  46445=>"111101100",
  46446=>"100110011",
  46447=>"001000100",
  46448=>"111100110",
  46449=>"000111110",
  46450=>"100101110",
  46451=>"000101001",
  46452=>"111101011",
  46453=>"001000001",
  46454=>"101010001",
  46455=>"010000100",
  46456=>"110011110",
  46457=>"011100111",
  46458=>"110101100",
  46459=>"111110110",
  46460=>"111110110",
  46461=>"100100110",
  46462=>"100100101",
  46463=>"100011101",
  46464=>"100100110",
  46465=>"100100011",
  46466=>"101001110",
  46467=>"100001111",
  46468=>"010101101",
  46469=>"000100101",
  46470=>"011000011",
  46471=>"100010101",
  46472=>"001010111",
  46473=>"000000011",
  46474=>"000001110",
  46475=>"111110111",
  46476=>"010001000",
  46477=>"110111100",
  46478=>"001101101",
  46479=>"110000100",
  46480=>"001100100",
  46481=>"100100000",
  46482=>"011100010",
  46483=>"000110010",
  46484=>"101101010",
  46485=>"000110010",
  46486=>"101000100",
  46487=>"111001101",
  46488=>"101111010",
  46489=>"000100101",
  46490=>"011010001",
  46491=>"101111110",
  46492=>"110000010",
  46493=>"011111110",
  46494=>"011001011",
  46495=>"010100100",
  46496=>"001110011",
  46497=>"111010100",
  46498=>"000011101",
  46499=>"111010000",
  46500=>"010000001",
  46501=>"001110111",
  46502=>"010111101",
  46503=>"000110010",
  46504=>"011101110",
  46505=>"011011011",
  46506=>"100110111",
  46507=>"000110111",
  46508=>"111110010",
  46509=>"011110111",
  46510=>"100011111",
  46511=>"000111111",
  46512=>"110101001",
  46513=>"010000111",
  46514=>"010110110",
  46515=>"111100001",
  46516=>"101010000",
  46517=>"111111100",
  46518=>"001011110",
  46519=>"010111101",
  46520=>"011000000",
  46521=>"111001101",
  46522=>"100000101",
  46523=>"110101010",
  46524=>"000011110",
  46525=>"110010111",
  46526=>"001001010",
  46527=>"100100010",
  46528=>"010000101",
  46529=>"001101111",
  46530=>"110111011",
  46531=>"010010111",
  46532=>"000000101",
  46533=>"110000010",
  46534=>"111100000",
  46535=>"100010000",
  46536=>"100110100",
  46537=>"001000110",
  46538=>"000010100",
  46539=>"101101000",
  46540=>"001111010",
  46541=>"110010011",
  46542=>"101100010",
  46543=>"011100111",
  46544=>"110111111",
  46545=>"010000000",
  46546=>"001001010",
  46547=>"111011111",
  46548=>"000100001",
  46549=>"011000010",
  46550=>"000101110",
  46551=>"100101100",
  46552=>"111100111",
  46553=>"000011000",
  46554=>"011100101",
  46555=>"010101010",
  46556=>"101010011",
  46557=>"010010011",
  46558=>"000010000",
  46559=>"100011110",
  46560=>"001101010",
  46561=>"000010001",
  46562=>"111110110",
  46563=>"010110111",
  46564=>"010110111",
  46565=>"000100111",
  46566=>"011010000",
  46567=>"111011110",
  46568=>"101100100",
  46569=>"101100011",
  46570=>"100111001",
  46571=>"110001111",
  46572=>"110010101",
  46573=>"110101100",
  46574=>"100101010",
  46575=>"110011111",
  46576=>"100000011",
  46577=>"101000101",
  46578=>"000110101",
  46579=>"111101101",
  46580=>"111010001",
  46581=>"011001110",
  46582=>"110011000",
  46583=>"011111110",
  46584=>"101000111",
  46585=>"111111110",
  46586=>"000100001",
  46587=>"111001010",
  46588=>"111000100",
  46589=>"001011100",
  46590=>"111110001",
  46591=>"110001110",
  46592=>"000111001",
  46593=>"010101000",
  46594=>"001101100",
  46595=>"101100001",
  46596=>"101011110",
  46597=>"110111011",
  46598=>"000000000",
  46599=>"000001111",
  46600=>"110100110",
  46601=>"001000110",
  46602=>"010011011",
  46603=>"111010000",
  46604=>"001001010",
  46605=>"001111110",
  46606=>"110010111",
  46607=>"101101110",
  46608=>"110001110",
  46609=>"010100101",
  46610=>"111010010",
  46611=>"011101011",
  46612=>"001110010",
  46613=>"011101110",
  46614=>"100101100",
  46615=>"101110001",
  46616=>"000010111",
  46617=>"000110111",
  46618=>"111001011",
  46619=>"000110000",
  46620=>"111000110",
  46621=>"010101010",
  46622=>"110000000",
  46623=>"110001110",
  46624=>"011001010",
  46625=>"001010000",
  46626=>"000100101",
  46627=>"111100101",
  46628=>"010011011",
  46629=>"111010100",
  46630=>"100100010",
  46631=>"110000000",
  46632=>"010000101",
  46633=>"000000110",
  46634=>"100011111",
  46635=>"100000100",
  46636=>"111110101",
  46637=>"110100011",
  46638=>"100101000",
  46639=>"111110101",
  46640=>"011110110",
  46641=>"011010100",
  46642=>"011000001",
  46643=>"000100011",
  46644=>"100101110",
  46645=>"000011101",
  46646=>"010010000",
  46647=>"000111011",
  46648=>"110011111",
  46649=>"001010110",
  46650=>"101011001",
  46651=>"001100101",
  46652=>"111011011",
  46653=>"000111100",
  46654=>"001010101",
  46655=>"110101001",
  46656=>"010100010",
  46657=>"110011010",
  46658=>"100000101",
  46659=>"000000000",
  46660=>"110111111",
  46661=>"110101000",
  46662=>"110000101",
  46663=>"111000000",
  46664=>"110010101",
  46665=>"011011101",
  46666=>"110111010",
  46667=>"100110100",
  46668=>"111010001",
  46669=>"110000101",
  46670=>"011111001",
  46671=>"011111101",
  46672=>"101110101",
  46673=>"010000101",
  46674=>"101111100",
  46675=>"000111001",
  46676=>"100100100",
  46677=>"100100010",
  46678=>"000111010",
  46679=>"100111010",
  46680=>"011111111",
  46681=>"110100011",
  46682=>"110011010",
  46683=>"110010111",
  46684=>"000100010",
  46685=>"100010001",
  46686=>"111110110",
  46687=>"100001101",
  46688=>"111011001",
  46689=>"100001111",
  46690=>"011000111",
  46691=>"000001011",
  46692=>"001000111",
  46693=>"001100111",
  46694=>"001110001",
  46695=>"001011101",
  46696=>"111010111",
  46697=>"000100100",
  46698=>"100111011",
  46699=>"101010011",
  46700=>"100111000",
  46701=>"010001100",
  46702=>"111010111",
  46703=>"111101100",
  46704=>"011111100",
  46705=>"100110111",
  46706=>"111011001",
  46707=>"000111101",
  46708=>"000000111",
  46709=>"011100100",
  46710=>"011000001",
  46711=>"010010001",
  46712=>"001010110",
  46713=>"011100101",
  46714=>"011101001",
  46715=>"101010111",
  46716=>"110000100",
  46717=>"001000000",
  46718=>"111010011",
  46719=>"111011111",
  46720=>"100011100",
  46721=>"000100011",
  46722=>"100111000",
  46723=>"010111011",
  46724=>"101010111",
  46725=>"100110101",
  46726=>"101011000",
  46727=>"010111110",
  46728=>"000000011",
  46729=>"110100010",
  46730=>"000110100",
  46731=>"001000110",
  46732=>"101100101",
  46733=>"001101110",
  46734=>"111101001",
  46735=>"010011011",
  46736=>"110000011",
  46737=>"110001111",
  46738=>"010110001",
  46739=>"011110000",
  46740=>"001001001",
  46741=>"001000001",
  46742=>"010111001",
  46743=>"011100001",
  46744=>"100111101",
  46745=>"100101000",
  46746=>"111001001",
  46747=>"101110000",
  46748=>"100101101",
  46749=>"101010001",
  46750=>"111000011",
  46751=>"010100000",
  46752=>"001001100",
  46753=>"001100100",
  46754=>"101111010",
  46755=>"111001101",
  46756=>"010111111",
  46757=>"101000001",
  46758=>"100010100",
  46759=>"110100100",
  46760=>"010110111",
  46761=>"111100001",
  46762=>"000101011",
  46763=>"101111100",
  46764=>"101110111",
  46765=>"110101110",
  46766=>"001010011",
  46767=>"110001100",
  46768=>"010011001",
  46769=>"001011111",
  46770=>"001100000",
  46771=>"100010011",
  46772=>"111101000",
  46773=>"000000000",
  46774=>"111100001",
  46775=>"010110100",
  46776=>"110111110",
  46777=>"001100100",
  46778=>"101000001",
  46779=>"010101100",
  46780=>"000111101",
  46781=>"110011010",
  46782=>"111101111",
  46783=>"100000011",
  46784=>"111001111",
  46785=>"111001101",
  46786=>"011010101",
  46787=>"101000000",
  46788=>"010111010",
  46789=>"010110110",
  46790=>"000011100",
  46791=>"010110001",
  46792=>"011010111",
  46793=>"111110100",
  46794=>"100100010",
  46795=>"000000101",
  46796=>"000010010",
  46797=>"111111001",
  46798=>"101101011",
  46799=>"010010000",
  46800=>"000111010",
  46801=>"100011110",
  46802=>"111111001",
  46803=>"011100100",
  46804=>"111101011",
  46805=>"110000001",
  46806=>"100111010",
  46807=>"110101000",
  46808=>"000000001",
  46809=>"110101110",
  46810=>"101110100",
  46811=>"101110111",
  46812=>"010001000",
  46813=>"110000010",
  46814=>"111011000",
  46815=>"000000001",
  46816=>"010000000",
  46817=>"110000100",
  46818=>"110001001",
  46819=>"110001100",
  46820=>"100001000",
  46821=>"001110111",
  46822=>"101011101",
  46823=>"010110110",
  46824=>"101111101",
  46825=>"001011001",
  46826=>"111111111",
  46827=>"100011111",
  46828=>"110011111",
  46829=>"111011001",
  46830=>"110010100",
  46831=>"100011100",
  46832=>"011110111",
  46833=>"000011001",
  46834=>"010000111",
  46835=>"001101000",
  46836=>"111001000",
  46837=>"011001010",
  46838=>"111111010",
  46839=>"010110011",
  46840=>"100110011",
  46841=>"100111101",
  46842=>"000010111",
  46843=>"111111101",
  46844=>"101011010",
  46845=>"000001111",
  46846=>"000100011",
  46847=>"100110110",
  46848=>"001001111",
  46849=>"101101001",
  46850=>"000000010",
  46851=>"100000011",
  46852=>"111101000",
  46853=>"000000110",
  46854=>"000111100",
  46855=>"011111000",
  46856=>"010111110",
  46857=>"100010100",
  46858=>"000101100",
  46859=>"000100101",
  46860=>"111100011",
  46861=>"100110110",
  46862=>"010000000",
  46863=>"010101000",
  46864=>"101011101",
  46865=>"111001111",
  46866=>"010110110",
  46867=>"000011000",
  46868=>"110001000",
  46869=>"011111010",
  46870=>"101110001",
  46871=>"101001010",
  46872=>"001101000",
  46873=>"100000000",
  46874=>"011100000",
  46875=>"110100110",
  46876=>"001010000",
  46877=>"000001011",
  46878=>"010100101",
  46879=>"011101111",
  46880=>"101001011",
  46881=>"001101111",
  46882=>"101000001",
  46883=>"011111100",
  46884=>"001011110",
  46885=>"000011000",
  46886=>"110111101",
  46887=>"010000001",
  46888=>"001111101",
  46889=>"100110101",
  46890=>"010110010",
  46891=>"001010000",
  46892=>"100010110",
  46893=>"110000001",
  46894=>"111101111",
  46895=>"010000101",
  46896=>"111101100",
  46897=>"010111010",
  46898=>"100111100",
  46899=>"100100001",
  46900=>"000101110",
  46901=>"011110101",
  46902=>"110110101",
  46903=>"111011110",
  46904=>"001011010",
  46905=>"001000001",
  46906=>"110011001",
  46907=>"010010000",
  46908=>"110111101",
  46909=>"011110110",
  46910=>"000010001",
  46911=>"110001111",
  46912=>"001010001",
  46913=>"111100001",
  46914=>"011010011",
  46915=>"110101111",
  46916=>"111011001",
  46917=>"010010010",
  46918=>"100001011",
  46919=>"010110101",
  46920=>"000111011",
  46921=>"010000101",
  46922=>"011111110",
  46923=>"000101000",
  46924=>"000110000",
  46925=>"111110000",
  46926=>"101101100",
  46927=>"100001001",
  46928=>"100000111",
  46929=>"000011101",
  46930=>"101110010",
  46931=>"011101000",
  46932=>"010000001",
  46933=>"000100100",
  46934=>"001111001",
  46935=>"011110100",
  46936=>"011010110",
  46937=>"110111110",
  46938=>"010101011",
  46939=>"110111000",
  46940=>"010101001",
  46941=>"010101111",
  46942=>"101110100",
  46943=>"000001010",
  46944=>"011111101",
  46945=>"110111011",
  46946=>"101100001",
  46947=>"000001100",
  46948=>"000000110",
  46949=>"001000100",
  46950=>"001101010",
  46951=>"011000100",
  46952=>"000000011",
  46953=>"000110011",
  46954=>"111110000",
  46955=>"001101110",
  46956=>"011000001",
  46957=>"010000110",
  46958=>"101011100",
  46959=>"011101110",
  46960=>"011101011",
  46961=>"101010110",
  46962=>"101011001",
  46963=>"110000110",
  46964=>"111110011",
  46965=>"000101111",
  46966=>"010011110",
  46967=>"011111100",
  46968=>"111010111",
  46969=>"101010000",
  46970=>"011010010",
  46971=>"101100110",
  46972=>"011000111",
  46973=>"010000101",
  46974=>"011001100",
  46975=>"011001001",
  46976=>"010010010",
  46977=>"111110100",
  46978=>"010010100",
  46979=>"100110011",
  46980=>"011100000",
  46981=>"110110000",
  46982=>"010000101",
  46983=>"100110100",
  46984=>"110000010",
  46985=>"110111010",
  46986=>"111010101",
  46987=>"110011001",
  46988=>"111000001",
  46989=>"001111010",
  46990=>"001001111",
  46991=>"010110011",
  46992=>"001001100",
  46993=>"000010001",
  46994=>"000001000",
  46995=>"010010011",
  46996=>"111000000",
  46997=>"010111111",
  46998=>"100011111",
  46999=>"011111111",
  47000=>"011100111",
  47001=>"010111001",
  47002=>"100111000",
  47003=>"011011001",
  47004=>"000011011",
  47005=>"010011001",
  47006=>"100001000",
  47007=>"111100000",
  47008=>"011011000",
  47009=>"101000100",
  47010=>"101100011",
  47011=>"101100101",
  47012=>"001100110",
  47013=>"111000110",
  47014=>"010110100",
  47015=>"101011001",
  47016=>"001100001",
  47017=>"000011000",
  47018=>"111111010",
  47019=>"111100010",
  47020=>"010111101",
  47021=>"010110110",
  47022=>"010110000",
  47023=>"111111111",
  47024=>"001011101",
  47025=>"110000111",
  47026=>"100010110",
  47027=>"100011001",
  47028=>"010001100",
  47029=>"111110110",
  47030=>"011001111",
  47031=>"011010001",
  47032=>"000001001",
  47033=>"100100000",
  47034=>"001101001",
  47035=>"000000101",
  47036=>"101110100",
  47037=>"111000101",
  47038=>"110010100",
  47039=>"100011001",
  47040=>"010111110",
  47041=>"010000011",
  47042=>"100011000",
  47043=>"101010111",
  47044=>"001111110",
  47045=>"100110010",
  47046=>"100001111",
  47047=>"111001110",
  47048=>"101001001",
  47049=>"111111011",
  47050=>"010100010",
  47051=>"100001101",
  47052=>"101010000",
  47053=>"001001101",
  47054=>"110011111",
  47055=>"101000001",
  47056=>"100111110",
  47057=>"001000111",
  47058=>"001110100",
  47059=>"100111000",
  47060=>"110001101",
  47061=>"000111111",
  47062=>"000100000",
  47063=>"001100100",
  47064=>"100001101",
  47065=>"000110010",
  47066=>"111001010",
  47067=>"001100000",
  47068=>"101010010",
  47069=>"100010000",
  47070=>"101010110",
  47071=>"111010001",
  47072=>"011101111",
  47073=>"011010100",
  47074=>"011110000",
  47075=>"000001100",
  47076=>"000001001",
  47077=>"001001101",
  47078=>"101111110",
  47079=>"110110001",
  47080=>"101100010",
  47081=>"101011111",
  47082=>"110110011",
  47083=>"001000101",
  47084=>"101111001",
  47085=>"001110010",
  47086=>"010001000",
  47087=>"101001111",
  47088=>"111100111",
  47089=>"111101011",
  47090=>"001110110",
  47091=>"110010100",
  47092=>"111111011",
  47093=>"111011010",
  47094=>"000011001",
  47095=>"110110110",
  47096=>"101010110",
  47097=>"011110100",
  47098=>"100110111",
  47099=>"111101100",
  47100=>"101101101",
  47101=>"111111001",
  47102=>"111000000",
  47103=>"101001100",
  47104=>"110110101",
  47105=>"110101010",
  47106=>"111111011",
  47107=>"011001100",
  47108=>"010001000",
  47109=>"101001011",
  47110=>"111111101",
  47111=>"010110111",
  47112=>"101000000",
  47113=>"100101001",
  47114=>"010001111",
  47115=>"111010010",
  47116=>"000001110",
  47117=>"000110100",
  47118=>"111000011",
  47119=>"010011100",
  47120=>"101110001",
  47121=>"011001000",
  47122=>"111001111",
  47123=>"100100001",
  47124=>"101111101",
  47125=>"000001000",
  47126=>"101110110",
  47127=>"100110100",
  47128=>"010110001",
  47129=>"001001111",
  47130=>"100010010",
  47131=>"100100100",
  47132=>"000101101",
  47133=>"100011101",
  47134=>"001001100",
  47135=>"100110010",
  47136=>"111001011",
  47137=>"101000010",
  47138=>"001000001",
  47139=>"000100010",
  47140=>"000111010",
  47141=>"011110100",
  47142=>"100001110",
  47143=>"000010001",
  47144=>"011001000",
  47145=>"011110010",
  47146=>"000011010",
  47147=>"001100001",
  47148=>"111110011",
  47149=>"011110111",
  47150=>"011111010",
  47151=>"100100011",
  47152=>"110100011",
  47153=>"001000110",
  47154=>"100011101",
  47155=>"110100010",
  47156=>"001101010",
  47157=>"001100110",
  47158=>"000100111",
  47159=>"001001001",
  47160=>"000011010",
  47161=>"011010000",
  47162=>"000100010",
  47163=>"101101101",
  47164=>"101110100",
  47165=>"111011111",
  47166=>"100001110",
  47167=>"110101001",
  47168=>"100101001",
  47169=>"011111001",
  47170=>"000010110",
  47171=>"111110100",
  47172=>"001001110",
  47173=>"001101011",
  47174=>"010100110",
  47175=>"101001100",
  47176=>"000000101",
  47177=>"010100011",
  47178=>"011110011",
  47179=>"111100100",
  47180=>"001100000",
  47181=>"101110001",
  47182=>"010100111",
  47183=>"101011010",
  47184=>"101011100",
  47185=>"111000000",
  47186=>"010111101",
  47187=>"010100010",
  47188=>"011111101",
  47189=>"000110000",
  47190=>"011100100",
  47191=>"001100110",
  47192=>"011100010",
  47193=>"100000011",
  47194=>"111100101",
  47195=>"010100000",
  47196=>"110100000",
  47197=>"000000110",
  47198=>"000100000",
  47199=>"000001010",
  47200=>"111000111",
  47201=>"100110100",
  47202=>"100000010",
  47203=>"000000100",
  47204=>"010100101",
  47205=>"000000000",
  47206=>"111011101",
  47207=>"011111110",
  47208=>"101011101",
  47209=>"011001011",
  47210=>"100010010",
  47211=>"000000010",
  47212=>"100010000",
  47213=>"000001000",
  47214=>"100000010",
  47215=>"110111001",
  47216=>"011111000",
  47217=>"100000000",
  47218=>"101011110",
  47219=>"000000101",
  47220=>"101110000",
  47221=>"100101101",
  47222=>"000011111",
  47223=>"110110100",
  47224=>"100011010",
  47225=>"001011101",
  47226=>"010010001",
  47227=>"101101001",
  47228=>"010001101",
  47229=>"101111100",
  47230=>"110001000",
  47231=>"011101011",
  47232=>"010100000",
  47233=>"101111000",
  47234=>"101001101",
  47235=>"000001100",
  47236=>"100010110",
  47237=>"010011111",
  47238=>"111000110",
  47239=>"100100000",
  47240=>"111110000",
  47241=>"101011000",
  47242=>"000100011",
  47243=>"100100001",
  47244=>"100100111",
  47245=>"010100110",
  47246=>"000101011",
  47247=>"001010010",
  47248=>"000110100",
  47249=>"100001001",
  47250=>"110111001",
  47251=>"000010100",
  47252=>"110001000",
  47253=>"010010100",
  47254=>"010101111",
  47255=>"011010101",
  47256=>"010010110",
  47257=>"001010000",
  47258=>"000100111",
  47259=>"001110000",
  47260=>"101101111",
  47261=>"101010101",
  47262=>"110011010",
  47263=>"101011110",
  47264=>"001110111",
  47265=>"111111100",
  47266=>"000100000",
  47267=>"000111110",
  47268=>"110101110",
  47269=>"010101111",
  47270=>"101010001",
  47271=>"111110111",
  47272=>"110110000",
  47273=>"000000000",
  47274=>"101100000",
  47275=>"000111111",
  47276=>"110100100",
  47277=>"101010000",
  47278=>"011001001",
  47279=>"010100100",
  47280=>"111001100",
  47281=>"110110100",
  47282=>"111111001",
  47283=>"001101000",
  47284=>"101010100",
  47285=>"100000111",
  47286=>"110000010",
  47287=>"001101011",
  47288=>"101110010",
  47289=>"010000011",
  47290=>"000010110",
  47291=>"011010011",
  47292=>"111100101",
  47293=>"101010011",
  47294=>"110000000",
  47295=>"011011111",
  47296=>"101100000",
  47297=>"010011010",
  47298=>"111100000",
  47299=>"011111110",
  47300=>"011001101",
  47301=>"010000001",
  47302=>"011011011",
  47303=>"010001111",
  47304=>"000011100",
  47305=>"100001011",
  47306=>"100100100",
  47307=>"000011010",
  47308=>"011001110",
  47309=>"110010011",
  47310=>"101000111",
  47311=>"000100001",
  47312=>"000100100",
  47313=>"001101100",
  47314=>"001110000",
  47315=>"100011111",
  47316=>"011100100",
  47317=>"001101101",
  47318=>"101000011",
  47319=>"111111011",
  47320=>"010101001",
  47321=>"110111111",
  47322=>"000111001",
  47323=>"100001010",
  47324=>"101110111",
  47325=>"001011100",
  47326=>"001100110",
  47327=>"100011010",
  47328=>"110100000",
  47329=>"010011010",
  47330=>"100000000",
  47331=>"110010001",
  47332=>"011011101",
  47333=>"110101000",
  47334=>"110110011",
  47335=>"100101101",
  47336=>"111100001",
  47337=>"110001000",
  47338=>"010010010",
  47339=>"111011000",
  47340=>"100001000",
  47341=>"011001101",
  47342=>"101000110",
  47343=>"010101111",
  47344=>"100001110",
  47345=>"100111100",
  47346=>"001011100",
  47347=>"001001101",
  47348=>"101111011",
  47349=>"111011101",
  47350=>"111100011",
  47351=>"000000110",
  47352=>"001001100",
  47353=>"110100101",
  47354=>"100011011",
  47355=>"101111000",
  47356=>"110110001",
  47357=>"111010000",
  47358=>"111000010",
  47359=>"000010110",
  47360=>"110000110",
  47361=>"000011010",
  47362=>"001101110",
  47363=>"011011111",
  47364=>"110111000",
  47365=>"001010000",
  47366=>"101001010",
  47367=>"110111011",
  47368=>"110100100",
  47369=>"111001110",
  47370=>"100000010",
  47371=>"001111110",
  47372=>"000011101",
  47373=>"000011101",
  47374=>"001011000",
  47375=>"001000110",
  47376=>"010000111",
  47377=>"001000101",
  47378=>"001111101",
  47379=>"110110110",
  47380=>"111111100",
  47381=>"010001101",
  47382=>"011110010",
  47383=>"001000100",
  47384=>"100010010",
  47385=>"000110010",
  47386=>"011100101",
  47387=>"000010110",
  47388=>"101010110",
  47389=>"111101001",
  47390=>"110010100",
  47391=>"000011000",
  47392=>"100101100",
  47393=>"111101111",
  47394=>"100010101",
  47395=>"001100101",
  47396=>"111000110",
  47397=>"100000110",
  47398=>"000001001",
  47399=>"011111110",
  47400=>"100001000",
  47401=>"111110000",
  47402=>"111101010",
  47403=>"011101011",
  47404=>"110001100",
  47405=>"111000000",
  47406=>"110101000",
  47407=>"001011010",
  47408=>"011010001",
  47409=>"011111011",
  47410=>"101010101",
  47411=>"001101011",
  47412=>"110001000",
  47413=>"000110100",
  47414=>"100110101",
  47415=>"111001111",
  47416=>"011111111",
  47417=>"010100101",
  47418=>"100111110",
  47419=>"101111110",
  47420=>"110001000",
  47421=>"101110111",
  47422=>"101110000",
  47423=>"100011001",
  47424=>"110001010",
  47425=>"110100110",
  47426=>"001010001",
  47427=>"000000001",
  47428=>"000000110",
  47429=>"110010101",
  47430=>"011011000",
  47431=>"110111100",
  47432=>"110010010",
  47433=>"011110010",
  47434=>"000010010",
  47435=>"000010011",
  47436=>"101000010",
  47437=>"010110000",
  47438=>"101111110",
  47439=>"010110101",
  47440=>"001011101",
  47441=>"011000111",
  47442=>"010110110",
  47443=>"111111111",
  47444=>"110011010",
  47445=>"011110010",
  47446=>"100100100",
  47447=>"000011000",
  47448=>"100111111",
  47449=>"000011011",
  47450=>"100110010",
  47451=>"111010011",
  47452=>"111111110",
  47453=>"110110011",
  47454=>"111001100",
  47455=>"100111001",
  47456=>"100001011",
  47457=>"100010110",
  47458=>"001101000",
  47459=>"000100110",
  47460=>"110100111",
  47461=>"111101000",
  47462=>"100101001",
  47463=>"010110000",
  47464=>"100100010",
  47465=>"110010011",
  47466=>"100100011",
  47467=>"010000000",
  47468=>"001001110",
  47469=>"100011111",
  47470=>"011101110",
  47471=>"100101010",
  47472=>"101010101",
  47473=>"011000111",
  47474=>"001011111",
  47475=>"110011000",
  47476=>"011000011",
  47477=>"101011101",
  47478=>"100010001",
  47479=>"100110000",
  47480=>"101110011",
  47481=>"010010000",
  47482=>"100101101",
  47483=>"111011001",
  47484=>"011011010",
  47485=>"000101011",
  47486=>"110110111",
  47487=>"000001110",
  47488=>"000001101",
  47489=>"100000011",
  47490=>"100011010",
  47491=>"001101110",
  47492=>"111001100",
  47493=>"010000110",
  47494=>"010111001",
  47495=>"010001000",
  47496=>"101000011",
  47497=>"101010011",
  47498=>"001101010",
  47499=>"011011110",
  47500=>"001000001",
  47501=>"011011010",
  47502=>"101100010",
  47503=>"110111111",
  47504=>"100100010",
  47505=>"110110000",
  47506=>"110011010",
  47507=>"000000001",
  47508=>"111000011",
  47509=>"010110101",
  47510=>"111010111",
  47511=>"101111011",
  47512=>"100100000",
  47513=>"000011111",
  47514=>"000100110",
  47515=>"000010110",
  47516=>"110001000",
  47517=>"000111101",
  47518=>"001001111",
  47519=>"101100101",
  47520=>"010011100",
  47521=>"111001000",
  47522=>"011110000",
  47523=>"010111101",
  47524=>"101011110",
  47525=>"111011010",
  47526=>"011010110",
  47527=>"101101001",
  47528=>"100000001",
  47529=>"010010001",
  47530=>"010100111",
  47531=>"001110000",
  47532=>"011110000",
  47533=>"000111101",
  47534=>"111101100",
  47535=>"011111110",
  47536=>"111111111",
  47537=>"010011111",
  47538=>"110101111",
  47539=>"110111001",
  47540=>"000110010",
  47541=>"111111111",
  47542=>"110000111",
  47543=>"100010011",
  47544=>"011000000",
  47545=>"100011101",
  47546=>"011011001",
  47547=>"100001011",
  47548=>"001101010",
  47549=>"011011110",
  47550=>"101011101",
  47551=>"100111111",
  47552=>"000110111",
  47553=>"001101011",
  47554=>"111100001",
  47555=>"101110011",
  47556=>"111110010",
  47557=>"000101111",
  47558=>"101100010",
  47559=>"000111010",
  47560=>"110100000",
  47561=>"110111111",
  47562=>"100001000",
  47563=>"101001110",
  47564=>"100000111",
  47565=>"001111001",
  47566=>"100101101",
  47567=>"100001001",
  47568=>"101001011",
  47569=>"111110100",
  47570=>"000100100",
  47571=>"011001101",
  47572=>"001101110",
  47573=>"111000000",
  47574=>"110101100",
  47575=>"010001000",
  47576=>"000011000",
  47577=>"010010100",
  47578=>"100101010",
  47579=>"000001001",
  47580=>"001011010",
  47581=>"111101100",
  47582=>"101100100",
  47583=>"111111011",
  47584=>"100110000",
  47585=>"100011110",
  47586=>"100000111",
  47587=>"101001101",
  47588=>"101001101",
  47589=>"111110011",
  47590=>"001111101",
  47591=>"010100100",
  47592=>"101100010",
  47593=>"101000000",
  47594=>"111100010",
  47595=>"111100000",
  47596=>"000101111",
  47597=>"011011101",
  47598=>"100000001",
  47599=>"001110000",
  47600=>"101000011",
  47601=>"000010100",
  47602=>"100111101",
  47603=>"101000101",
  47604=>"000001100",
  47605=>"111111000",
  47606=>"100011011",
  47607=>"100011001",
  47608=>"111001101",
  47609=>"010000100",
  47610=>"011110110",
  47611=>"000001100",
  47612=>"111101100",
  47613=>"100001101",
  47614=>"000111111",
  47615=>"111101010",
  47616=>"000000101",
  47617=>"101001110",
  47618=>"010101101",
  47619=>"110101000",
  47620=>"100111010",
  47621=>"000111110",
  47622=>"110000100",
  47623=>"111101000",
  47624=>"110111111",
  47625=>"010101000",
  47626=>"000011000",
  47627=>"100000110",
  47628=>"011101010",
  47629=>"111111001",
  47630=>"001000000",
  47631=>"000011011",
  47632=>"111010011",
  47633=>"010111101",
  47634=>"010010101",
  47635=>"001000101",
  47636=>"100101101",
  47637=>"010111001",
  47638=>"011000110",
  47639=>"000101010",
  47640=>"110000011",
  47641=>"000100110",
  47642=>"110011100",
  47643=>"100101011",
  47644=>"011011010",
  47645=>"110111010",
  47646=>"001000001",
  47647=>"011110010",
  47648=>"001110111",
  47649=>"010101100",
  47650=>"010111010",
  47651=>"100111100",
  47652=>"101011111",
  47653=>"100101001",
  47654=>"010100001",
  47655=>"111010001",
  47656=>"110110111",
  47657=>"101001011",
  47658=>"000011001",
  47659=>"001101010",
  47660=>"110100000",
  47661=>"000000000",
  47662=>"000111111",
  47663=>"010101111",
  47664=>"101100001",
  47665=>"010011010",
  47666=>"110001000",
  47667=>"110110111",
  47668=>"100011110",
  47669=>"100000000",
  47670=>"001001001",
  47671=>"111011110",
  47672=>"011101111",
  47673=>"111010100",
  47674=>"001010011",
  47675=>"001110011",
  47676=>"100100100",
  47677=>"000000100",
  47678=>"110000000",
  47679=>"100001110",
  47680=>"101001001",
  47681=>"100100110",
  47682=>"011001111",
  47683=>"101100001",
  47684=>"010100010",
  47685=>"011111100",
  47686=>"011100100",
  47687=>"011100100",
  47688=>"000011011",
  47689=>"001000011",
  47690=>"001010101",
  47691=>"000101100",
  47692=>"111010101",
  47693=>"010001000",
  47694=>"001011110",
  47695=>"011000001",
  47696=>"101000111",
  47697=>"110000101",
  47698=>"110000100",
  47699=>"001101110",
  47700=>"011100111",
  47701=>"010110010",
  47702=>"011010110",
  47703=>"100111101",
  47704=>"000101010",
  47705=>"010001101",
  47706=>"100000011",
  47707=>"010110011",
  47708=>"111001111",
  47709=>"010001111",
  47710=>"101000100",
  47711=>"100100010",
  47712=>"001110010",
  47713=>"100000010",
  47714=>"001101011",
  47715=>"000000001",
  47716=>"001110111",
  47717=>"110001111",
  47718=>"011101110",
  47719=>"000111111",
  47720=>"100001101",
  47721=>"111101001",
  47722=>"000001100",
  47723=>"111010000",
  47724=>"110100010",
  47725=>"110010001",
  47726=>"001111010",
  47727=>"101100011",
  47728=>"000110000",
  47729=>"100011000",
  47730=>"100000101",
  47731=>"000110010",
  47732=>"010111000",
  47733=>"100000110",
  47734=>"000111000",
  47735=>"001110010",
  47736=>"010011100",
  47737=>"111010001",
  47738=>"111000110",
  47739=>"011111101",
  47740=>"101101011",
  47741=>"010111111",
  47742=>"101010100",
  47743=>"101011000",
  47744=>"000110000",
  47745=>"101100000",
  47746=>"101011101",
  47747=>"110101000",
  47748=>"111111000",
  47749=>"110110011",
  47750=>"110001100",
  47751=>"011011110",
  47752=>"110111000",
  47753=>"010001011",
  47754=>"000001000",
  47755=>"000100110",
  47756=>"001100110",
  47757=>"110000000",
  47758=>"111010010",
  47759=>"100110111",
  47760=>"110000100",
  47761=>"110010010",
  47762=>"001001001",
  47763=>"000100111",
  47764=>"100101000",
  47765=>"010110000",
  47766=>"010001100",
  47767=>"010111110",
  47768=>"101111100",
  47769=>"011010010",
  47770=>"100000100",
  47771=>"011100001",
  47772=>"110001110",
  47773=>"110011100",
  47774=>"110001000",
  47775=>"000000000",
  47776=>"100011101",
  47777=>"011111110",
  47778=>"101101001",
  47779=>"000110110",
  47780=>"110000011",
  47781=>"010100001",
  47782=>"100100100",
  47783=>"100110000",
  47784=>"111110010",
  47785=>"111101010",
  47786=>"110110010",
  47787=>"010110010",
  47788=>"110000000",
  47789=>"011000001",
  47790=>"010100111",
  47791=>"111010111",
  47792=>"100000000",
  47793=>"011001111",
  47794=>"110111010",
  47795=>"101100110",
  47796=>"111001000",
  47797=>"111011110",
  47798=>"010110101",
  47799=>"101010001",
  47800=>"101101111",
  47801=>"010000100",
  47802=>"010111011",
  47803=>"110010001",
  47804=>"000010100",
  47805=>"011000110",
  47806=>"111101010",
  47807=>"000010100",
  47808=>"110110000",
  47809=>"110111100",
  47810=>"110010000",
  47811=>"010010001",
  47812=>"111001110",
  47813=>"000011001",
  47814=>"111011001",
  47815=>"110011011",
  47816=>"000101110",
  47817=>"101001101",
  47818=>"111010011",
  47819=>"101101100",
  47820=>"101000000",
  47821=>"101010101",
  47822=>"011001110",
  47823=>"011000011",
  47824=>"111110110",
  47825=>"010011110",
  47826=>"110110100",
  47827=>"000101101",
  47828=>"110001101",
  47829=>"101011011",
  47830=>"110101011",
  47831=>"000000010",
  47832=>"101111111",
  47833=>"001010010",
  47834=>"110011100",
  47835=>"111000111",
  47836=>"011100011",
  47837=>"111101100",
  47838=>"010010001",
  47839=>"010001011",
  47840=>"000001100",
  47841=>"010101001",
  47842=>"111001111",
  47843=>"001011110",
  47844=>"011000011",
  47845=>"010000000",
  47846=>"100000101",
  47847=>"101011111",
  47848=>"000100010",
  47849=>"011101110",
  47850=>"011001000",
  47851=>"001001100",
  47852=>"001000101",
  47853=>"000100011",
  47854=>"011010011",
  47855=>"101001000",
  47856=>"111101000",
  47857=>"011111101",
  47858=>"101001101",
  47859=>"110011100",
  47860=>"100010110",
  47861=>"000000111",
  47862=>"110101111",
  47863=>"111110011",
  47864=>"100111000",
  47865=>"101000111",
  47866=>"010110001",
  47867=>"000011111",
  47868=>"011110010",
  47869=>"000100001",
  47870=>"110000100",
  47871=>"101001010",
  47872=>"111101010",
  47873=>"000111101",
  47874=>"010010011",
  47875=>"101111001",
  47876=>"100001000",
  47877=>"000000111",
  47878=>"111001000",
  47879=>"001000011",
  47880=>"010000001",
  47881=>"011010100",
  47882=>"111001100",
  47883=>"111111101",
  47884=>"000011011",
  47885=>"010001111",
  47886=>"101100001",
  47887=>"111100101",
  47888=>"010000011",
  47889=>"100111101",
  47890=>"101101110",
  47891=>"101010110",
  47892=>"001101110",
  47893=>"001000001",
  47894=>"000011101",
  47895=>"101001011",
  47896=>"111000101",
  47897=>"010100011",
  47898=>"001101011",
  47899=>"001001011",
  47900=>"101010101",
  47901=>"010001000",
  47902=>"100110110",
  47903=>"001010101",
  47904=>"010110000",
  47905=>"000001101",
  47906=>"111001010",
  47907=>"000010011",
  47908=>"010010001",
  47909=>"011011100",
  47910=>"101010010",
  47911=>"101111111",
  47912=>"000000001",
  47913=>"101010101",
  47914=>"000101010",
  47915=>"010000101",
  47916=>"100100000",
  47917=>"000001100",
  47918=>"110010000",
  47919=>"110011101",
  47920=>"110000001",
  47921=>"011000100",
  47922=>"101101010",
  47923=>"000010011",
  47924=>"000011011",
  47925=>"111001001",
  47926=>"101001111",
  47927=>"010101100",
  47928=>"110111110",
  47929=>"000111111",
  47930=>"010110000",
  47931=>"101001111",
  47932=>"000001000",
  47933=>"011011011",
  47934=>"010110001",
  47935=>"011111000",
  47936=>"110100000",
  47937=>"001111111",
  47938=>"001000100",
  47939=>"100101110",
  47940=>"011010011",
  47941=>"111001010",
  47942=>"000111101",
  47943=>"111111010",
  47944=>"010011111",
  47945=>"110101010",
  47946=>"111100011",
  47947=>"101010001",
  47948=>"001011010",
  47949=>"111010000",
  47950=>"111101101",
  47951=>"111110111",
  47952=>"101101110",
  47953=>"010111010",
  47954=>"011100110",
  47955=>"101110100",
  47956=>"000001111",
  47957=>"101110000",
  47958=>"001000000",
  47959=>"111011001",
  47960=>"011010101",
  47961=>"110000011",
  47962=>"011110010",
  47963=>"111100101",
  47964=>"110011001",
  47965=>"100010001",
  47966=>"100110010",
  47967=>"100110010",
  47968=>"000110001",
  47969=>"101010011",
  47970=>"000110010",
  47971=>"110110110",
  47972=>"100011010",
  47973=>"000010100",
  47974=>"111100100",
  47975=>"011111110",
  47976=>"100111110",
  47977=>"011001111",
  47978=>"010011100",
  47979=>"100111100",
  47980=>"000100100",
  47981=>"100110110",
  47982=>"101011110",
  47983=>"011110011",
  47984=>"101101010",
  47985=>"001100000",
  47986=>"010101110",
  47987=>"110101001",
  47988=>"010100110",
  47989=>"000000111",
  47990=>"000000101",
  47991=>"011111101",
  47992=>"001100011",
  47993=>"111011000",
  47994=>"110001011",
  47995=>"110110101",
  47996=>"111000101",
  47997=>"101100001",
  47998=>"011110011",
  47999=>"000000010",
  48000=>"000101100",
  48001=>"010110110",
  48002=>"111100110",
  48003=>"110001101",
  48004=>"010001110",
  48005=>"000011001",
  48006=>"001000011",
  48007=>"001011011",
  48008=>"011101111",
  48009=>"000011101",
  48010=>"110100101",
  48011=>"001101101",
  48012=>"010000000",
  48013=>"000100000",
  48014=>"111101010",
  48015=>"111111110",
  48016=>"101100001",
  48017=>"001110100",
  48018=>"110000010",
  48019=>"010000001",
  48020=>"001110001",
  48021=>"100000011",
  48022=>"111111000",
  48023=>"000001010",
  48024=>"011010000",
  48025=>"101011001",
  48026=>"101110010",
  48027=>"110000101",
  48028=>"110000111",
  48029=>"010011010",
  48030=>"010110111",
  48031=>"110000001",
  48032=>"101111111",
  48033=>"000100011",
  48034=>"100000000",
  48035=>"000111100",
  48036=>"010100000",
  48037=>"011001110",
  48038=>"001101001",
  48039=>"010110110",
  48040=>"110001101",
  48041=>"010100000",
  48042=>"010001011",
  48043=>"011100100",
  48044=>"011000001",
  48045=>"011101101",
  48046=>"110110110",
  48047=>"100010110",
  48048=>"101000000",
  48049=>"001010010",
  48050=>"001101000",
  48051=>"000100111",
  48052=>"101101001",
  48053=>"111101110",
  48054=>"000101101",
  48055=>"010110100",
  48056=>"000000001",
  48057=>"100011100",
  48058=>"000110100",
  48059=>"001110010",
  48060=>"100011110",
  48061=>"110111000",
  48062=>"000010001",
  48063=>"001101101",
  48064=>"001000011",
  48065=>"110101010",
  48066=>"100001001",
  48067=>"011000010",
  48068=>"001010111",
  48069=>"011001110",
  48070=>"001011011",
  48071=>"000000010",
  48072=>"111110000",
  48073=>"100111010",
  48074=>"010100001",
  48075=>"101100000",
  48076=>"110000110",
  48077=>"101101011",
  48078=>"100001111",
  48079=>"101001101",
  48080=>"000010011",
  48081=>"111101001",
  48082=>"101100100",
  48083=>"011111011",
  48084=>"011010110",
  48085=>"101010011",
  48086=>"101100000",
  48087=>"001010110",
  48088=>"010000110",
  48089=>"001010101",
  48090=>"010111111",
  48091=>"110001100",
  48092=>"001011011",
  48093=>"101111111",
  48094=>"000101111",
  48095=>"100111101",
  48096=>"110011000",
  48097=>"100100111",
  48098=>"000001100",
  48099=>"111001010",
  48100=>"001001001",
  48101=>"011110111",
  48102=>"000000101",
  48103=>"011111011",
  48104=>"100111100",
  48105=>"110001101",
  48106=>"011011100",
  48107=>"010010011",
  48108=>"011101111",
  48109=>"000001001",
  48110=>"001101010",
  48111=>"010101111",
  48112=>"111000101",
  48113=>"010101000",
  48114=>"000011111",
  48115=>"010100110",
  48116=>"101101110",
  48117=>"000010010",
  48118=>"001000100",
  48119=>"011111110",
  48120=>"001000010",
  48121=>"110111101",
  48122=>"110100111",
  48123=>"010101010",
  48124=>"100111110",
  48125=>"001101101",
  48126=>"110100110",
  48127=>"101111111",
  48128=>"001110101",
  48129=>"011110000",
  48130=>"010110111",
  48131=>"000011101",
  48132=>"001001100",
  48133=>"000000111",
  48134=>"100110011",
  48135=>"010111111",
  48136=>"101001010",
  48137=>"101100111",
  48138=>"100100000",
  48139=>"110101011",
  48140=>"010001011",
  48141=>"001000101",
  48142=>"101101010",
  48143=>"100111000",
  48144=>"110101101",
  48145=>"011110101",
  48146=>"011110101",
  48147=>"000101101",
  48148=>"001001011",
  48149=>"101011000",
  48150=>"100101100",
  48151=>"001011111",
  48152=>"101000011",
  48153=>"100110011",
  48154=>"011010010",
  48155=>"111000010",
  48156=>"010000000",
  48157=>"101111111",
  48158=>"010110001",
  48159=>"100010010",
  48160=>"101110001",
  48161=>"000110011",
  48162=>"001010111",
  48163=>"010101111",
  48164=>"101000010",
  48165=>"101011000",
  48166=>"000000111",
  48167=>"011101011",
  48168=>"101111001",
  48169=>"001100100",
  48170=>"001101010",
  48171=>"101011001",
  48172=>"011101110",
  48173=>"011001110",
  48174=>"111100111",
  48175=>"000000101",
  48176=>"101000111",
  48177=>"100110111",
  48178=>"101111111",
  48179=>"011100000",
  48180=>"101101111",
  48181=>"111001111",
  48182=>"111010011",
  48183=>"011010100",
  48184=>"000101111",
  48185=>"001110000",
  48186=>"001111111",
  48187=>"111010010",
  48188=>"000011100",
  48189=>"010011010",
  48190=>"110010111",
  48191=>"100001100",
  48192=>"010001101",
  48193=>"000100001",
  48194=>"011000110",
  48195=>"011011111",
  48196=>"011100001",
  48197=>"011111010",
  48198=>"110111010",
  48199=>"000100101",
  48200=>"010011111",
  48201=>"001110001",
  48202=>"001011110",
  48203=>"111111111",
  48204=>"110110110",
  48205=>"001111111",
  48206=>"110111100",
  48207=>"111010000",
  48208=>"011000111",
  48209=>"011100111",
  48210=>"110000111",
  48211=>"110100110",
  48212=>"000101001",
  48213=>"001011000",
  48214=>"111110110",
  48215=>"111011000",
  48216=>"111011101",
  48217=>"111111101",
  48218=>"000101000",
  48219=>"001110100",
  48220=>"000011110",
  48221=>"010001010",
  48222=>"010110010",
  48223=>"000010011",
  48224=>"000010111",
  48225=>"100100011",
  48226=>"000111000",
  48227=>"101110110",
  48228=>"111010110",
  48229=>"001001110",
  48230=>"101100101",
  48231=>"111101100",
  48232=>"100001011",
  48233=>"101000111",
  48234=>"110000000",
  48235=>"111110110",
  48236=>"101010010",
  48237=>"110111000",
  48238=>"100000000",
  48239=>"010100111",
  48240=>"111100001",
  48241=>"111110001",
  48242=>"100111010",
  48243=>"010001100",
  48244=>"101111111",
  48245=>"111101100",
  48246=>"110011011",
  48247=>"010110001",
  48248=>"011111100",
  48249=>"011110000",
  48250=>"011111000",
  48251=>"000000100",
  48252=>"011101000",
  48253=>"101100000",
  48254=>"010111110",
  48255=>"111100110",
  48256=>"000001101",
  48257=>"111110111",
  48258=>"010110000",
  48259=>"001111110",
  48260=>"001100101",
  48261=>"001011100",
  48262=>"111001000",
  48263=>"010110011",
  48264=>"011001110",
  48265=>"011110011",
  48266=>"011010010",
  48267=>"101011010",
  48268=>"000011000",
  48269=>"100001011",
  48270=>"100010110",
  48271=>"111010001",
  48272=>"110100011",
  48273=>"010100100",
  48274=>"010111011",
  48275=>"110001110",
  48276=>"001000010",
  48277=>"111000000",
  48278=>"010101011",
  48279=>"101101101",
  48280=>"011010100",
  48281=>"110111110",
  48282=>"110111100",
  48283=>"111100000",
  48284=>"100000011",
  48285=>"011001000",
  48286=>"011001101",
  48287=>"000110000",
  48288=>"001000101",
  48289=>"101111110",
  48290=>"110000010",
  48291=>"110111110",
  48292=>"011101101",
  48293=>"101111001",
  48294=>"100000100",
  48295=>"111001111",
  48296=>"110100011",
  48297=>"110111111",
  48298=>"000011000",
  48299=>"111101001",
  48300=>"101001110",
  48301=>"011110001",
  48302=>"101001001",
  48303=>"100011000",
  48304=>"111010010",
  48305=>"010010001",
  48306=>"001010101",
  48307=>"100101101",
  48308=>"101111001",
  48309=>"001101111",
  48310=>"111010011",
  48311=>"101000000",
  48312=>"000001101",
  48313=>"101011000",
  48314=>"101001010",
  48315=>"110100001",
  48316=>"110110101",
  48317=>"010001000",
  48318=>"011001111",
  48319=>"101111111",
  48320=>"001010101",
  48321=>"001000010",
  48322=>"100100010",
  48323=>"111000101",
  48324=>"011101111",
  48325=>"100000110",
  48326=>"100111000",
  48327=>"101010111",
  48328=>"101011001",
  48329=>"010111111",
  48330=>"111101111",
  48331=>"101001011",
  48332=>"101010110",
  48333=>"001001000",
  48334=>"011100010",
  48335=>"011100110",
  48336=>"101100100",
  48337=>"011010101",
  48338=>"010011010",
  48339=>"111001111",
  48340=>"010101111",
  48341=>"111011001",
  48342=>"010001110",
  48343=>"111010111",
  48344=>"000110111",
  48345=>"000001100",
  48346=>"100111001",
  48347=>"110100000",
  48348=>"100010010",
  48349=>"111000001",
  48350=>"000101000",
  48351=>"100110111",
  48352=>"011010001",
  48353=>"001010001",
  48354=>"001000111",
  48355=>"110110110",
  48356=>"110001000",
  48357=>"011100000",
  48358=>"110011111",
  48359=>"100000001",
  48360=>"010011101",
  48361=>"111011011",
  48362=>"000100000",
  48363=>"101100110",
  48364=>"010110111",
  48365=>"101100100",
  48366=>"011100011",
  48367=>"100010111",
  48368=>"111101111",
  48369=>"110010101",
  48370=>"110010100",
  48371=>"000001001",
  48372=>"101101111",
  48373=>"001101011",
  48374=>"011110001",
  48375=>"101110110",
  48376=>"010101111",
  48377=>"100011111",
  48378=>"010001110",
  48379=>"000000000",
  48380=>"110010001",
  48381=>"100000111",
  48382=>"111011110",
  48383=>"101110110",
  48384=>"010010101",
  48385=>"100111111",
  48386=>"100000110",
  48387=>"111101100",
  48388=>"010111100",
  48389=>"100011100",
  48390=>"010000011",
  48391=>"011010000",
  48392=>"111101111",
  48393=>"101010101",
  48394=>"001011000",
  48395=>"001011111",
  48396=>"010000100",
  48397=>"010011100",
  48398=>"010111101",
  48399=>"000010110",
  48400=>"010010101",
  48401=>"111100001",
  48402=>"110000101",
  48403=>"110110000",
  48404=>"010000111",
  48405=>"110101101",
  48406=>"100111001",
  48407=>"011011101",
  48408=>"110111100",
  48409=>"111111100",
  48410=>"110111101",
  48411=>"011101000",
  48412=>"010010000",
  48413=>"101101110",
  48414=>"001110111",
  48415=>"010111100",
  48416=>"000101010",
  48417=>"101100000",
  48418=>"101101111",
  48419=>"011001011",
  48420=>"001011000",
  48421=>"011111110",
  48422=>"000110000",
  48423=>"010010110",
  48424=>"101011000",
  48425=>"110001010",
  48426=>"101010101",
  48427=>"001011001",
  48428=>"101001110",
  48429=>"010010100",
  48430=>"010000100",
  48431=>"111011000",
  48432=>"011011010",
  48433=>"110000100",
  48434=>"011111000",
  48435=>"000011110",
  48436=>"000000000",
  48437=>"010010001",
  48438=>"011000101",
  48439=>"001100010",
  48440=>"001110000",
  48441=>"011011011",
  48442=>"011011011",
  48443=>"000110100",
  48444=>"010111100",
  48445=>"000001000",
  48446=>"010000100",
  48447=>"011110100",
  48448=>"111001000",
  48449=>"110101110",
  48450=>"000111001",
  48451=>"100000000",
  48452=>"010000010",
  48453=>"000010001",
  48454=>"010010000",
  48455=>"011111110",
  48456=>"101010011",
  48457=>"100001000",
  48458=>"110001111",
  48459=>"001101110",
  48460=>"101110101",
  48461=>"110100000",
  48462=>"111110000",
  48463=>"010000011",
  48464=>"001000001",
  48465=>"100110111",
  48466=>"111010011",
  48467=>"000000111",
  48468=>"011000001",
  48469=>"111000101",
  48470=>"001010110",
  48471=>"011101100",
  48472=>"100101001",
  48473=>"000000010",
  48474=>"110111101",
  48475=>"000001011",
  48476=>"110110100",
  48477=>"100111100",
  48478=>"011000000",
  48479=>"011100100",
  48480=>"001011100",
  48481=>"001100010",
  48482=>"001000001",
  48483=>"000000110",
  48484=>"000100001",
  48485=>"000010001",
  48486=>"011001010",
  48487=>"101110111",
  48488=>"010100011",
  48489=>"100000001",
  48490=>"110100011",
  48491=>"010011111",
  48492=>"101101010",
  48493=>"001000001",
  48494=>"010001101",
  48495=>"001011111",
  48496=>"011011010",
  48497=>"101010111",
  48498=>"111011100",
  48499=>"110101010",
  48500=>"000110000",
  48501=>"011100111",
  48502=>"110000000",
  48503=>"100010001",
  48504=>"101111110",
  48505=>"000111010",
  48506=>"000000101",
  48507=>"011110110",
  48508=>"111101111",
  48509=>"101111011",
  48510=>"000000101",
  48511=>"011000101",
  48512=>"110000100",
  48513=>"101110111",
  48514=>"111111101",
  48515=>"000110101",
  48516=>"101100110",
  48517=>"110101101",
  48518=>"001110000",
  48519=>"000011101",
  48520=>"010111100",
  48521=>"110111001",
  48522=>"110101000",
  48523=>"000100110",
  48524=>"010110101",
  48525=>"110000110",
  48526=>"000101111",
  48527=>"001010101",
  48528=>"101100001",
  48529=>"110000110",
  48530=>"111011100",
  48531=>"011110110",
  48532=>"000110000",
  48533=>"001100010",
  48534=>"101000000",
  48535=>"010000010",
  48536=>"110100101",
  48537=>"000101111",
  48538=>"001001110",
  48539=>"101111010",
  48540=>"110001110",
  48541=>"010010000",
  48542=>"010010001",
  48543=>"101100011",
  48544=>"001011000",
  48545=>"110110010",
  48546=>"001110010",
  48547=>"001001001",
  48548=>"111000100",
  48549=>"100000001",
  48550=>"011011000",
  48551=>"011110101",
  48552=>"010010001",
  48553=>"000001011",
  48554=>"010011011",
  48555=>"111111101",
  48556=>"001000001",
  48557=>"111110110",
  48558=>"100001111",
  48559=>"101011011",
  48560=>"010100101",
  48561=>"110010001",
  48562=>"010001100",
  48563=>"101110010",
  48564=>"000100001",
  48565=>"111111001",
  48566=>"001000001",
  48567=>"001011110",
  48568=>"100110110",
  48569=>"011110000",
  48570=>"000011101",
  48571=>"110110000",
  48572=>"110001011",
  48573=>"010010111",
  48574=>"111001100",
  48575=>"001111101",
  48576=>"101001111",
  48577=>"111100010",
  48578=>"001111101",
  48579=>"011000110",
  48580=>"000011110",
  48581=>"001000101",
  48582=>"111001001",
  48583=>"110100000",
  48584=>"110010011",
  48585=>"000000011",
  48586=>"110000100",
  48587=>"001100100",
  48588=>"001011101",
  48589=>"100010101",
  48590=>"001010111",
  48591=>"001100010",
  48592=>"101011111",
  48593=>"110000001",
  48594=>"010101111",
  48595=>"000001010",
  48596=>"010111001",
  48597=>"000011100",
  48598=>"011010111",
  48599=>"010110111",
  48600=>"111100101",
  48601=>"001101101",
  48602=>"110000111",
  48603=>"111100000",
  48604=>"111001010",
  48605=>"010000000",
  48606=>"100100011",
  48607=>"001100100",
  48608=>"000111011",
  48609=>"000110001",
  48610=>"001110100",
  48611=>"110000001",
  48612=>"101101101",
  48613=>"001010110",
  48614=>"101010010",
  48615=>"100000011",
  48616=>"010111101",
  48617=>"110011010",
  48618=>"100110110",
  48619=>"010101101",
  48620=>"111011000",
  48621=>"100011000",
  48622=>"000101100",
  48623=>"100010011",
  48624=>"101011011",
  48625=>"100001000",
  48626=>"000011101",
  48627=>"100001000",
  48628=>"010001011",
  48629=>"110101000",
  48630=>"010111101",
  48631=>"100101000",
  48632=>"111111111",
  48633=>"000000111",
  48634=>"001101100",
  48635=>"001111011",
  48636=>"100110100",
  48637=>"110001101",
  48638=>"101010000",
  48639=>"111011101",
  48640=>"111000001",
  48641=>"100100100",
  48642=>"111100011",
  48643=>"000111010",
  48644=>"111010100",
  48645=>"001010000",
  48646=>"110000011",
  48647=>"001000010",
  48648=>"010100110",
  48649=>"101010010",
  48650=>"000001010",
  48651=>"111001001",
  48652=>"011010001",
  48653=>"111001000",
  48654=>"011000001",
  48655=>"111101111",
  48656=>"101010111",
  48657=>"100101110",
  48658=>"010000001",
  48659=>"010100110",
  48660=>"100101101",
  48661=>"110100011",
  48662=>"111011110",
  48663=>"001001111",
  48664=>"100000111",
  48665=>"000111011",
  48666=>"010010000",
  48667=>"110111000",
  48668=>"000100010",
  48669=>"100111011",
  48670=>"101101100",
  48671=>"000000000",
  48672=>"110111101",
  48673=>"101011111",
  48674=>"000001100",
  48675=>"001110111",
  48676=>"001010111",
  48677=>"001011101",
  48678=>"110010100",
  48679=>"001110111",
  48680=>"100011110",
  48681=>"110100101",
  48682=>"000000010",
  48683=>"001000010",
  48684=>"000001111",
  48685=>"100010100",
  48686=>"000000001",
  48687=>"010100100",
  48688=>"000011001",
  48689=>"001101100",
  48690=>"110010110",
  48691=>"111111101",
  48692=>"101110110",
  48693=>"100011010",
  48694=>"000001111",
  48695=>"100001011",
  48696=>"001101100",
  48697=>"101111101",
  48698=>"000110101",
  48699=>"000111111",
  48700=>"010001000",
  48701=>"011001101",
  48702=>"100010000",
  48703=>"011000001",
  48704=>"111010100",
  48705=>"111000111",
  48706=>"100100000",
  48707=>"011111010",
  48708=>"110010101",
  48709=>"001001110",
  48710=>"101000000",
  48711=>"111001110",
  48712=>"111110010",
  48713=>"000000111",
  48714=>"111100001",
  48715=>"000100111",
  48716=>"001100010",
  48717=>"010111101",
  48718=>"010000111",
  48719=>"000011111",
  48720=>"100011001",
  48721=>"000101110",
  48722=>"011010110",
  48723=>"000101010",
  48724=>"010001011",
  48725=>"010110111",
  48726=>"000011110",
  48727=>"000110001",
  48728=>"110011011",
  48729=>"011100110",
  48730=>"101110111",
  48731=>"111000000",
  48732=>"000100110",
  48733=>"111011000",
  48734=>"001001001",
  48735=>"101001101",
  48736=>"111010111",
  48737=>"111101101",
  48738=>"000110000",
  48739=>"110111011",
  48740=>"100000010",
  48741=>"110110110",
  48742=>"111010101",
  48743=>"000001011",
  48744=>"101110110",
  48745=>"001001001",
  48746=>"010101011",
  48747=>"111101101",
  48748=>"010001000",
  48749=>"010011011",
  48750=>"111110111",
  48751=>"101001010",
  48752=>"001101101",
  48753=>"010110011",
  48754=>"000011001",
  48755=>"001001110",
  48756=>"011011000",
  48757=>"000000011",
  48758=>"001001101",
  48759=>"101011000",
  48760=>"100000001",
  48761=>"111011101",
  48762=>"000011000",
  48763=>"111101001",
  48764=>"010000010",
  48765=>"110100010",
  48766=>"110001101",
  48767=>"100100011",
  48768=>"000000000",
  48769=>"111000011",
  48770=>"011101000",
  48771=>"001010010",
  48772=>"110010111",
  48773=>"011000110",
  48774=>"101111111",
  48775=>"010001000",
  48776=>"101011010",
  48777=>"110111000",
  48778=>"110000101",
  48779=>"011110101",
  48780=>"100110101",
  48781=>"001001110",
  48782=>"000100100",
  48783=>"100100010",
  48784=>"111010001",
  48785=>"010000101",
  48786=>"010011111",
  48787=>"111000100",
  48788=>"000100001",
  48789=>"101101110",
  48790=>"001000101",
  48791=>"001111010",
  48792=>"111001111",
  48793=>"111101111",
  48794=>"110011111",
  48795=>"111100000",
  48796=>"100111110",
  48797=>"001000000",
  48798=>"011000101",
  48799=>"110010010",
  48800=>"001011011",
  48801=>"100001001",
  48802=>"111110111",
  48803=>"100000000",
  48804=>"110110110",
  48805=>"010110100",
  48806=>"111011010",
  48807=>"010010001",
  48808=>"010100000",
  48809=>"110101010",
  48810=>"000011010",
  48811=>"000001000",
  48812=>"100101010",
  48813=>"101001011",
  48814=>"010000100",
  48815=>"110111010",
  48816=>"101001111",
  48817=>"101000111",
  48818=>"011001100",
  48819=>"101100101",
  48820=>"100010001",
  48821=>"100001111",
  48822=>"010000000",
  48823=>"011010010",
  48824=>"100111111",
  48825=>"010010100",
  48826=>"110110111",
  48827=>"100101111",
  48828=>"000010100",
  48829=>"110111000",
  48830=>"111001011",
  48831=>"110001101",
  48832=>"100110010",
  48833=>"001110001",
  48834=>"101111000",
  48835=>"010101000",
  48836=>"000100001",
  48837=>"000000100",
  48838=>"101100001",
  48839=>"001010001",
  48840=>"001110110",
  48841=>"011001011",
  48842=>"010100010",
  48843=>"110011111",
  48844=>"010100011",
  48845=>"111110110",
  48846=>"101010000",
  48847=>"000100010",
  48848=>"111010100",
  48849=>"011010110",
  48850=>"000110000",
  48851=>"110001110",
  48852=>"100100101",
  48853=>"110100100",
  48854=>"000100110",
  48855=>"000100110",
  48856=>"100101101",
  48857=>"101100111",
  48858=>"100011001",
  48859=>"100101100",
  48860=>"000110100",
  48861=>"000000011",
  48862=>"000110010",
  48863=>"001100100",
  48864=>"010001100",
  48865=>"011011011",
  48866=>"010100011",
  48867=>"111011101",
  48868=>"111110111",
  48869=>"101010001",
  48870=>"110000011",
  48871=>"111101011",
  48872=>"010101100",
  48873=>"111000111",
  48874=>"101011000",
  48875=>"010111001",
  48876=>"100011000",
  48877=>"100110010",
  48878=>"010011010",
  48879=>"111110110",
  48880=>"101100010",
  48881=>"001000011",
  48882=>"010010111",
  48883=>"001111111",
  48884=>"110100110",
  48885=>"001001111",
  48886=>"110111010",
  48887=>"100000011",
  48888=>"100000010",
  48889=>"100100110",
  48890=>"000101001",
  48891=>"011100110",
  48892=>"001000110",
  48893=>"000111001",
  48894=>"001111110",
  48895=>"100111111",
  48896=>"000011100",
  48897=>"011110101",
  48898=>"110101110",
  48899=>"110111111",
  48900=>"001001000",
  48901=>"000010001",
  48902=>"101001001",
  48903=>"110000011",
  48904=>"101101000",
  48905=>"001000100",
  48906=>"001011011",
  48907=>"111111111",
  48908=>"111001001",
  48909=>"011101111",
  48910=>"011011010",
  48911=>"111111101",
  48912=>"101011100",
  48913=>"111000110",
  48914=>"010000011",
  48915=>"011101111",
  48916=>"101111100",
  48917=>"010000110",
  48918=>"111100001",
  48919=>"011101101",
  48920=>"000000110",
  48921=>"100101100",
  48922=>"000011110",
  48923=>"100101001",
  48924=>"101101000",
  48925=>"111011001",
  48926=>"010001010",
  48927=>"101111011",
  48928=>"010011110",
  48929=>"111000101",
  48930=>"111111011",
  48931=>"000100011",
  48932=>"001101011",
  48933=>"110101000",
  48934=>"000000100",
  48935=>"111110101",
  48936=>"011010001",
  48937=>"111100011",
  48938=>"001100010",
  48939=>"111000000",
  48940=>"111011001",
  48941=>"100010010",
  48942=>"000000110",
  48943=>"011000111",
  48944=>"000001011",
  48945=>"110001111",
  48946=>"011110101",
  48947=>"010100000",
  48948=>"111001110",
  48949=>"001011101",
  48950=>"001101001",
  48951=>"110100100",
  48952=>"100110101",
  48953=>"010011010",
  48954=>"101110010",
  48955=>"000101011",
  48956=>"101101001",
  48957=>"100010110",
  48958=>"011110100",
  48959=>"000011101",
  48960=>"001100000",
  48961=>"101111111",
  48962=>"010110111",
  48963=>"110001000",
  48964=>"000101001",
  48965=>"111001001",
  48966=>"111010001",
  48967=>"000011101",
  48968=>"000000010",
  48969=>"100110010",
  48970=>"000101010",
  48971=>"101110101",
  48972=>"101011110",
  48973=>"000000001",
  48974=>"101001001",
  48975=>"001011100",
  48976=>"010110001",
  48977=>"111100000",
  48978=>"010110101",
  48979=>"011101101",
  48980=>"111100010",
  48981=>"111111111",
  48982=>"001111101",
  48983=>"011000111",
  48984=>"100011110",
  48985=>"001010001",
  48986=>"111010001",
  48987=>"111010101",
  48988=>"010100101",
  48989=>"001100110",
  48990=>"100010000",
  48991=>"010000101",
  48992=>"101000011",
  48993=>"000010100",
  48994=>"000010011",
  48995=>"010110110",
  48996=>"001101001",
  48997=>"111000100",
  48998=>"110011111",
  48999=>"110111001",
  49000=>"111101101",
  49001=>"000101111",
  49002=>"000101000",
  49003=>"101010010",
  49004=>"111111111",
  49005=>"111111100",
  49006=>"100011100",
  49007=>"101011100",
  49008=>"101111000",
  49009=>"110011011",
  49010=>"111111111",
  49011=>"000100001",
  49012=>"000001001",
  49013=>"010100011",
  49014=>"000001101",
  49015=>"111110111",
  49016=>"110011100",
  49017=>"010111000",
  49018=>"000011011",
  49019=>"000010001",
  49020=>"000111101",
  49021=>"111011101",
  49022=>"000111111",
  49023=>"001000111",
  49024=>"111001001",
  49025=>"011101000",
  49026=>"110010000",
  49027=>"011100100",
  49028=>"001101101",
  49029=>"101100110",
  49030=>"110010110",
  49031=>"000111101",
  49032=>"001110110",
  49033=>"111010010",
  49034=>"010101000",
  49035=>"111010110",
  49036=>"111011110",
  49037=>"010000000",
  49038=>"101110110",
  49039=>"110111110",
  49040=>"011111101",
  49041=>"000100011",
  49042=>"000010111",
  49043=>"001100000",
  49044=>"100100100",
  49045=>"100110100",
  49046=>"010101000",
  49047=>"110110000",
  49048=>"000011010",
  49049=>"111110000",
  49050=>"110010001",
  49051=>"111001001",
  49052=>"010001111",
  49053=>"001001101",
  49054=>"101110111",
  49055=>"111010011",
  49056=>"000101101",
  49057=>"101100110",
  49058=>"101000100",
  49059=>"010101100",
  49060=>"001101110",
  49061=>"001001010",
  49062=>"001101100",
  49063=>"111101101",
  49064=>"110111000",
  49065=>"101111100",
  49066=>"001110010",
  49067=>"100000110",
  49068=>"100111000",
  49069=>"100001111",
  49070=>"010111000",
  49071=>"101111000",
  49072=>"011011110",
  49073=>"010110101",
  49074=>"001011011",
  49075=>"100101011",
  49076=>"000001001",
  49077=>"001000100",
  49078=>"110111101",
  49079=>"000110111",
  49080=>"001111010",
  49081=>"111011011",
  49082=>"101000011",
  49083=>"001011001",
  49084=>"110001011",
  49085=>"010001000",
  49086=>"111010001",
  49087=>"101001110",
  49088=>"111111000",
  49089=>"111010100",
  49090=>"000101101",
  49091=>"111100100",
  49092=>"001101010",
  49093=>"101011100",
  49094=>"101000001",
  49095=>"110001010",
  49096=>"101000101",
  49097=>"100000011",
  49098=>"110110101",
  49099=>"001001001",
  49100=>"001100001",
  49101=>"000001100",
  49102=>"111111001",
  49103=>"010010010",
  49104=>"111000101",
  49105=>"011111000",
  49106=>"111100100",
  49107=>"001101001",
  49108=>"011001011",
  49109=>"100100010",
  49110=>"110100110",
  49111=>"001110101",
  49112=>"111001111",
  49113=>"101110001",
  49114=>"101111000",
  49115=>"101010100",
  49116=>"100010010",
  49117=>"101111100",
  49118=>"000101000",
  49119=>"001011001",
  49120=>"001001010",
  49121=>"111100001",
  49122=>"111000001",
  49123=>"110101010",
  49124=>"000000011",
  49125=>"100000101",
  49126=>"001001001",
  49127=>"011010110",
  49128=>"010000000",
  49129=>"100001010",
  49130=>"110101100",
  49131=>"110011000",
  49132=>"011110011",
  49133=>"110010110",
  49134=>"001001000",
  49135=>"101110101",
  49136=>"101101000",
  49137=>"011110100",
  49138=>"010101000",
  49139=>"110111011",
  49140=>"111001000",
  49141=>"000100001",
  49142=>"101001111",
  49143=>"000101000",
  49144=>"111011100",
  49145=>"000001110",
  49146=>"101110101",
  49147=>"110011110",
  49148=>"010111111",
  49149=>"111110101",
  49150=>"010101111",
  49151=>"001110100",
  49152=>"001101011",
  49153=>"010100011",
  49154=>"110111011",
  49155=>"000010000",
  49156=>"011110011",
  49157=>"110011001",
  49158=>"100111101",
  49159=>"001111000",
  49160=>"101011010",
  49161=>"000001010",
  49162=>"010101100",
  49163=>"010100000",
  49164=>"110010000",
  49165=>"000000100",
  49166=>"001110101",
  49167=>"000001011",
  49168=>"101000101",
  49169=>"011110101",
  49170=>"100111101",
  49171=>"010010101",
  49172=>"011101000",
  49173=>"111110101",
  49174=>"110101100",
  49175=>"000000100",
  49176=>"111000100",
  49177=>"011011010",
  49178=>"111001101",
  49179=>"011110110",
  49180=>"001110110",
  49181=>"010011110",
  49182=>"110010001",
  49183=>"100001001",
  49184=>"010001100",
  49185=>"110111011",
  49186=>"010010111",
  49187=>"111011010",
  49188=>"010101111",
  49189=>"100111111",
  49190=>"110001001",
  49191=>"110101111",
  49192=>"111001000",
  49193=>"101010100",
  49194=>"110000010",
  49195=>"111000010",
  49196=>"100100110",
  49197=>"010101100",
  49198=>"101001011",
  49199=>"000011011",
  49200=>"010011110",
  49201=>"110111110",
  49202=>"010000100",
  49203=>"011011001",
  49204=>"000011110",
  49205=>"001110101",
  49206=>"110001101",
  49207=>"101111001",
  49208=>"000001001",
  49209=>"101101100",
  49210=>"001000110",
  49211=>"100001100",
  49212=>"100110000",
  49213=>"001111010",
  49214=>"011010101",
  49215=>"000010000",
  49216=>"100011000",
  49217=>"100101100",
  49218=>"001101111",
  49219=>"000101110",
  49220=>"110010000",
  49221=>"101000111",
  49222=>"110010101",
  49223=>"000011010",
  49224=>"011111101",
  49225=>"101010000",
  49226=>"010010010",
  49227=>"101001101",
  49228=>"110110011",
  49229=>"001011110",
  49230=>"000000001",
  49231=>"000010001",
  49232=>"001001011",
  49233=>"101011001",
  49234=>"100110110",
  49235=>"100000010",
  49236=>"011110101",
  49237=>"111001101",
  49238=>"110011111",
  49239=>"101101101",
  49240=>"111110000",
  49241=>"010110111",
  49242=>"101001001",
  49243=>"110001000",
  49244=>"000000010",
  49245=>"100000011",
  49246=>"101111101",
  49247=>"101011100",
  49248=>"011011001",
  49249=>"111101001",
  49250=>"001100010",
  49251=>"010010000",
  49252=>"100100010",
  49253=>"000100100",
  49254=>"001011100",
  49255=>"110001001",
  49256=>"000101000",
  49257=>"011000010",
  49258=>"100001000",
  49259=>"010000100",
  49260=>"110010010",
  49261=>"010110010",
  49262=>"001000101",
  49263=>"000000100",
  49264=>"000111111",
  49265=>"010000000",
  49266=>"011010100",
  49267=>"111100110",
  49268=>"000001001",
  49269=>"001010111",
  49270=>"110101110",
  49271=>"011100100",
  49272=>"000011010",
  49273=>"001101101",
  49274=>"111100110",
  49275=>"111000001",
  49276=>"000111110",
  49277=>"110110110",
  49278=>"101110110",
  49279=>"001010110",
  49280=>"001111110",
  49281=>"101111110",
  49282=>"011000000",
  49283=>"100010000",
  49284=>"001101001",
  49285=>"101101110",
  49286=>"001001001",
  49287=>"100111000",
  49288=>"011101110",
  49289=>"111110000",
  49290=>"011011101",
  49291=>"110001111",
  49292=>"011101101",
  49293=>"110011101",
  49294=>"111111011",
  49295=>"111111111",
  49296=>"001110100",
  49297=>"100010011",
  49298=>"011001001",
  49299=>"110101001",
  49300=>"011011000",
  49301=>"010011100",
  49302=>"000010100",
  49303=>"001110000",
  49304=>"111100100",
  49305=>"000000110",
  49306=>"011010011",
  49307=>"110111011",
  49308=>"000000111",
  49309=>"110100100",
  49310=>"101111111",
  49311=>"110000000",
  49312=>"110110001",
  49313=>"101100110",
  49314=>"011111111",
  49315=>"001101011",
  49316=>"000110100",
  49317=>"010010010",
  49318=>"010110111",
  49319=>"011011000",
  49320=>"111011101",
  49321=>"000010000",
  49322=>"111000110",
  49323=>"100001001",
  49324=>"111110011",
  49325=>"111101010",
  49326=>"101001001",
  49327=>"010110001",
  49328=>"010000101",
  49329=>"010111010",
  49330=>"001000010",
  49331=>"101010101",
  49332=>"011110101",
  49333=>"111101001",
  49334=>"010001010",
  49335=>"111110000",
  49336=>"101100001",
  49337=>"100011000",
  49338=>"110101010",
  49339=>"100001111",
  49340=>"000011001",
  49341=>"110101100",
  49342=>"011110100",
  49343=>"000010001",
  49344=>"010111000",
  49345=>"110100110",
  49346=>"010001001",
  49347=>"111011110",
  49348=>"111110010",
  49349=>"000101010",
  49350=>"010100101",
  49351=>"001010101",
  49352=>"000001100",
  49353=>"111111010",
  49354=>"001001111",
  49355=>"101110101",
  49356=>"010111101",
  49357=>"100101110",
  49358=>"001100101",
  49359=>"110111110",
  49360=>"101011010",
  49361=>"101111110",
  49362=>"000011000",
  49363=>"010000110",
  49364=>"110100100",
  49365=>"110000101",
  49366=>"011111000",
  49367=>"010111101",
  49368=>"000110000",
  49369=>"101100101",
  49370=>"001011000",
  49371=>"001010010",
  49372=>"000001101",
  49373=>"010101110",
  49374=>"001010010",
  49375=>"111101010",
  49376=>"111110000",
  49377=>"110001110",
  49378=>"010000100",
  49379=>"111110001",
  49380=>"010101011",
  49381=>"101100011",
  49382=>"001001000",
  49383=>"111010111",
  49384=>"010001000",
  49385=>"000111100",
  49386=>"000011001",
  49387=>"101111000",
  49388=>"101000001",
  49389=>"111100000",
  49390=>"010001110",
  49391=>"111111001",
  49392=>"000001000",
  49393=>"111111110",
  49394=>"011011001",
  49395=>"001010011",
  49396=>"001010000",
  49397=>"100110111",
  49398=>"101100011",
  49399=>"111011100",
  49400=>"001001011",
  49401=>"010100011",
  49402=>"000011010",
  49403=>"010101001",
  49404=>"010100001",
  49405=>"111001011",
  49406=>"110000110",
  49407=>"101110010",
  49408=>"110010100",
  49409=>"100000010",
  49410=>"110110111",
  49411=>"001001111",
  49412=>"101010101",
  49413=>"100011000",
  49414=>"000001101",
  49415=>"100100110",
  49416=>"000001001",
  49417=>"110100111",
  49418=>"111010101",
  49419=>"111000101",
  49420=>"110110101",
  49421=>"001010101",
  49422=>"110110001",
  49423=>"100010101",
  49424=>"100001000",
  49425=>"001001111",
  49426=>"101011001",
  49427=>"110111100",
  49428=>"001110100",
  49429=>"011001111",
  49430=>"111101011",
  49431=>"001010011",
  49432=>"011101101",
  49433=>"000000111",
  49434=>"100001011",
  49435=>"001000000",
  49436=>"100111001",
  49437=>"111010110",
  49438=>"100100011",
  49439=>"011110000",
  49440=>"010010001",
  49441=>"001111010",
  49442=>"011001111",
  49443=>"100110101",
  49444=>"111101011",
  49445=>"000000010",
  49446=>"011110100",
  49447=>"111110001",
  49448=>"001101010",
  49449=>"111111000",
  49450=>"101001100",
  49451=>"000101100",
  49452=>"000011010",
  49453=>"000000010",
  49454=>"000001110",
  49455=>"111110001",
  49456=>"100001011",
  49457=>"010110000",
  49458=>"000111010",
  49459=>"010001110",
  49460=>"101100010",
  49461=>"000010000",
  49462=>"111000100",
  49463=>"110110011",
  49464=>"000101010",
  49465=>"010010010",
  49466=>"010111101",
  49467=>"000010111",
  49468=>"100000110",
  49469=>"010011101",
  49470=>"101100010",
  49471=>"110111110",
  49472=>"100100010",
  49473=>"111111000",
  49474=>"000001110",
  49475=>"010011110",
  49476=>"011011100",
  49477=>"101000010",
  49478=>"001101110",
  49479=>"001011000",
  49480=>"000010001",
  49481=>"100100001",
  49482=>"011000001",
  49483=>"010010001",
  49484=>"110101010",
  49485=>"000000110",
  49486=>"111100110",
  49487=>"111110001",
  49488=>"100111000",
  49489=>"001100001",
  49490=>"111110010",
  49491=>"111101001",
  49492=>"000110100",
  49493=>"011100000",
  49494=>"111111001",
  49495=>"001110011",
  49496=>"000100001",
  49497=>"001110100",
  49498=>"011111111",
  49499=>"011101110",
  49500=>"000010010",
  49501=>"100000000",
  49502=>"100001101",
  49503=>"011101101",
  49504=>"110100001",
  49505=>"001111110",
  49506=>"110100010",
  49507=>"011101110",
  49508=>"001101000",
  49509=>"000011011",
  49510=>"011111001",
  49511=>"001011100",
  49512=>"000100100",
  49513=>"011000110",
  49514=>"101000001",
  49515=>"101110011",
  49516=>"100000010",
  49517=>"101010001",
  49518=>"110101000",
  49519=>"111000111",
  49520=>"100110101",
  49521=>"101110001",
  49522=>"111000001",
  49523=>"011101101",
  49524=>"001101101",
  49525=>"100111011",
  49526=>"110100111",
  49527=>"011101101",
  49528=>"011010001",
  49529=>"111111101",
  49530=>"101000001",
  49531=>"110001011",
  49532=>"010001001",
  49533=>"110010000",
  49534=>"100000110",
  49535=>"111100111",
  49536=>"110001111",
  49537=>"001100000",
  49538=>"010110111",
  49539=>"111110111",
  49540=>"101000000",
  49541=>"000110100",
  49542=>"110000001",
  49543=>"111111000",
  49544=>"100111000",
  49545=>"101101001",
  49546=>"111101101",
  49547=>"011100001",
  49548=>"100101001",
  49549=>"101110001",
  49550=>"011100110",
  49551=>"110011110",
  49552=>"110000000",
  49553=>"011010100",
  49554=>"000110111",
  49555=>"110101110",
  49556=>"100010101",
  49557=>"110010100",
  49558=>"100110101",
  49559=>"111011111",
  49560=>"101100010",
  49561=>"001001010",
  49562=>"010110110",
  49563=>"000001010",
  49564=>"010101111",
  49565=>"011110010",
  49566=>"101110111",
  49567=>"000011000",
  49568=>"000011100",
  49569=>"010010000",
  49570=>"010101111",
  49571=>"100000101",
  49572=>"100110101",
  49573=>"000000001",
  49574=>"011101100",
  49575=>"001010011",
  49576=>"111001110",
  49577=>"000000101",
  49578=>"110001000",
  49579=>"010000000",
  49580=>"000000111",
  49581=>"111011101",
  49582=>"101011111",
  49583=>"100000011",
  49584=>"000010010",
  49585=>"100011000",
  49586=>"011011000",
  49587=>"001000000",
  49588=>"100000000",
  49589=>"101111110",
  49590=>"101111101",
  49591=>"110001101",
  49592=>"111000001",
  49593=>"001010111",
  49594=>"000101101",
  49595=>"011010101",
  49596=>"001010001",
  49597=>"010000010",
  49598=>"001111111",
  49599=>"010111111",
  49600=>"111100100",
  49601=>"010100110",
  49602=>"111010100",
  49603=>"110110101",
  49604=>"001001101",
  49605=>"011010100",
  49606=>"110111100",
  49607=>"101001110",
  49608=>"001000110",
  49609=>"000011101",
  49610=>"101001000",
  49611=>"101010100",
  49612=>"101100000",
  49613=>"001111101",
  49614=>"110110110",
  49615=>"100101100",
  49616=>"000011111",
  49617=>"101000111",
  49618=>"100001111",
  49619=>"111110001",
  49620=>"100011111",
  49621=>"001101001",
  49622=>"111101101",
  49623=>"101100100",
  49624=>"000101001",
  49625=>"000000010",
  49626=>"101010000",
  49627=>"111100010",
  49628=>"101111111",
  49629=>"101001011",
  49630=>"000110110",
  49631=>"010011100",
  49632=>"111101111",
  49633=>"000011000",
  49634=>"010111100",
  49635=>"001100110",
  49636=>"001010011",
  49637=>"010100110",
  49638=>"110111111",
  49639=>"100111010",
  49640=>"100101100",
  49641=>"001110110",
  49642=>"101010011",
  49643=>"011011000",
  49644=>"001001010",
  49645=>"111001000",
  49646=>"010101011",
  49647=>"001111000",
  49648=>"000000011",
  49649=>"110010010",
  49650=>"111111000",
  49651=>"010011100",
  49652=>"110000101",
  49653=>"101101010",
  49654=>"101101010",
  49655=>"001001111",
  49656=>"100111101",
  49657=>"001001000",
  49658=>"100011100",
  49659=>"101100100",
  49660=>"001000000",
  49661=>"001001100",
  49662=>"001010000",
  49663=>"101111110",
  49664=>"100000001",
  49665=>"100101101",
  49666=>"111000111",
  49667=>"111100010",
  49668=>"111011100",
  49669=>"000011001",
  49670=>"101010011",
  49671=>"000110001",
  49672=>"110001001",
  49673=>"001110100",
  49674=>"010100001",
  49675=>"100100010",
  49676=>"111011111",
  49677=>"110110111",
  49678=>"000000010",
  49679=>"100100010",
  49680=>"000001001",
  49681=>"000001101",
  49682=>"111001010",
  49683=>"101110100",
  49684=>"000011101",
  49685=>"100101000",
  49686=>"010001010",
  49687=>"110001101",
  49688=>"101011001",
  49689=>"010001001",
  49690=>"110000100",
  49691=>"101110111",
  49692=>"000100100",
  49693=>"011010101",
  49694=>"110010101",
  49695=>"111111010",
  49696=>"001101001",
  49697=>"010010010",
  49698=>"111100100",
  49699=>"000011001",
  49700=>"000000111",
  49701=>"001110101",
  49702=>"011001101",
  49703=>"111001000",
  49704=>"000010101",
  49705=>"110101011",
  49706=>"000111000",
  49707=>"001111110",
  49708=>"100000100",
  49709=>"100101000",
  49710=>"001000101",
  49711=>"001000111",
  49712=>"010100001",
  49713=>"100001011",
  49714=>"101110001",
  49715=>"010011110",
  49716=>"101100000",
  49717=>"110010100",
  49718=>"000101101",
  49719=>"100011110",
  49720=>"110010100",
  49721=>"101000110",
  49722=>"111001111",
  49723=>"001001010",
  49724=>"110011100",
  49725=>"111001111",
  49726=>"100001101",
  49727=>"011000000",
  49728=>"000000001",
  49729=>"011000110",
  49730=>"110011110",
  49731=>"111011010",
  49732=>"110110001",
  49733=>"010011011",
  49734=>"000001000",
  49735=>"001010001",
  49736=>"111001100",
  49737=>"110011001",
  49738=>"001101101",
  49739=>"010000111",
  49740=>"101011000",
  49741=>"000110000",
  49742=>"111110111",
  49743=>"110010010",
  49744=>"110001010",
  49745=>"000111101",
  49746=>"101111101",
  49747=>"100000010",
  49748=>"100110000",
  49749=>"101100110",
  49750=>"000101000",
  49751=>"010001111",
  49752=>"100111101",
  49753=>"111011100",
  49754=>"011100001",
  49755=>"110001100",
  49756=>"000010101",
  49757=>"000011111",
  49758=>"010010111",
  49759=>"001111111",
  49760=>"101110110",
  49761=>"111111110",
  49762=>"001110010",
  49763=>"010100111",
  49764=>"110101111",
  49765=>"010111100",
  49766=>"111110011",
  49767=>"001001101",
  49768=>"010000111",
  49769=>"000101001",
  49770=>"101111111",
  49771=>"001001101",
  49772=>"011000101",
  49773=>"000010110",
  49774=>"000001011",
  49775=>"010000101",
  49776=>"011100001",
  49777=>"011100001",
  49778=>"111101111",
  49779=>"010110000",
  49780=>"011100111",
  49781=>"000111111",
  49782=>"011010010",
  49783=>"011110010",
  49784=>"000100000",
  49785=>"010001001",
  49786=>"110101011",
  49787=>"101000000",
  49788=>"101011000",
  49789=>"010100000",
  49790=>"110111011",
  49791=>"001101101",
  49792=>"110111001",
  49793=>"111101001",
  49794=>"010111111",
  49795=>"000011000",
  49796=>"110101100",
  49797=>"100100110",
  49798=>"101000010",
  49799=>"001111101",
  49800=>"111101010",
  49801=>"111101010",
  49802=>"100010001",
  49803=>"101111110",
  49804=>"000100001",
  49805=>"111110101",
  49806=>"000100000",
  49807=>"011110001",
  49808=>"011001101",
  49809=>"111000011",
  49810=>"100010011",
  49811=>"011101101",
  49812=>"101011001",
  49813=>"111110110",
  49814=>"101001001",
  49815=>"110110110",
  49816=>"100010011",
  49817=>"101001010",
  49818=>"110100101",
  49819=>"111001001",
  49820=>"000010001",
  49821=>"000011100",
  49822=>"000001001",
  49823=>"100101110",
  49824=>"000101011",
  49825=>"110000001",
  49826=>"011000001",
  49827=>"111001101",
  49828=>"001011001",
  49829=>"000010011",
  49830=>"110001100",
  49831=>"000010000",
  49832=>"110111110",
  49833=>"010000011",
  49834=>"010001010",
  49835=>"111001110",
  49836=>"001111110",
  49837=>"000001110",
  49838=>"101110111",
  49839=>"000100100",
  49840=>"001100011",
  49841=>"010001000",
  49842=>"000010111",
  49843=>"000000001",
  49844=>"001000111",
  49845=>"001100100",
  49846=>"001000001",
  49847=>"101011110",
  49848=>"101100100",
  49849=>"111101101",
  49850=>"011110101",
  49851=>"010011001",
  49852=>"101111010",
  49853=>"100111001",
  49854=>"001001101",
  49855=>"010000010",
  49856=>"001010100",
  49857=>"010011100",
  49858=>"100001010",
  49859=>"101101111",
  49860=>"110000101",
  49861=>"000000111",
  49862=>"001001000",
  49863=>"110110111",
  49864=>"000010000",
  49865=>"110111011",
  49866=>"111110010",
  49867=>"111110111",
  49868=>"001110100",
  49869=>"000101001",
  49870=>"110110001",
  49871=>"100001000",
  49872=>"100100100",
  49873=>"111011000",
  49874=>"001010101",
  49875=>"001000001",
  49876=>"000100001",
  49877=>"001111011",
  49878=>"100001000",
  49879=>"001011000",
  49880=>"010011000",
  49881=>"101100001",
  49882=>"101010101",
  49883=>"001010101",
  49884=>"001110110",
  49885=>"111011001",
  49886=>"010101100",
  49887=>"110100110",
  49888=>"000011001",
  49889=>"001110011",
  49890=>"101001001",
  49891=>"111111000",
  49892=>"101000010",
  49893=>"011011111",
  49894=>"111111010",
  49895=>"011110100",
  49896=>"110110111",
  49897=>"110010101",
  49898=>"000100001",
  49899=>"011101101",
  49900=>"000010010",
  49901=>"110101110",
  49902=>"110000011",
  49903=>"010101110",
  49904=>"000101101",
  49905=>"000100001",
  49906=>"010110010",
  49907=>"111111111",
  49908=>"101111011",
  49909=>"110100000",
  49910=>"001010011",
  49911=>"100101101",
  49912=>"100100111",
  49913=>"011011001",
  49914=>"100001111",
  49915=>"101110010",
  49916=>"111011001",
  49917=>"101110100",
  49918=>"110010101",
  49919=>"111001010",
  49920=>"111010001",
  49921=>"000101111",
  49922=>"110011110",
  49923=>"101011000",
  49924=>"010001001",
  49925=>"001100111",
  49926=>"111101000",
  49927=>"111111000",
  49928=>"010010111",
  49929=>"100100001",
  49930=>"000101101",
  49931=>"011010100",
  49932=>"001011101",
  49933=>"000111111",
  49934=>"111000111",
  49935=>"111111111",
  49936=>"111110110",
  49937=>"010000000",
  49938=>"100001110",
  49939=>"000101100",
  49940=>"000001111",
  49941=>"110000010",
  49942=>"010000011",
  49943=>"101011000",
  49944=>"010111010",
  49945=>"101001111",
  49946=>"101000000",
  49947=>"010110110",
  49948=>"111110101",
  49949=>"000100111",
  49950=>"111101010",
  49951=>"000110000",
  49952=>"100010100",
  49953=>"110001001",
  49954=>"111001001",
  49955=>"010111100",
  49956=>"011111101",
  49957=>"100000110",
  49958=>"101111010",
  49959=>"010111010",
  49960=>"001111101",
  49961=>"100001010",
  49962=>"010010000",
  49963=>"011110010",
  49964=>"101101011",
  49965=>"000000010",
  49966=>"111110010",
  49967=>"111111110",
  49968=>"101000000",
  49969=>"000111011",
  49970=>"000010111",
  49971=>"110111101",
  49972=>"100111110",
  49973=>"110010010",
  49974=>"001011010",
  49975=>"101101010",
  49976=>"111001101",
  49977=>"100011011",
  49978=>"111111010",
  49979=>"111011110",
  49980=>"001001000",
  49981=>"000001101",
  49982=>"000100111",
  49983=>"000101000",
  49984=>"101000001",
  49985=>"011100011",
  49986=>"000101110",
  49987=>"001111000",
  49988=>"000100101",
  49989=>"000111010",
  49990=>"100010000",
  49991=>"110110000",
  49992=>"000000101",
  49993=>"111101100",
  49994=>"100100100",
  49995=>"011100101",
  49996=>"111101000",
  49997=>"100011110",
  49998=>"000111100",
  49999=>"110100010",
  50000=>"011011001",
  50001=>"100111101",
  50002=>"111110001",
  50003=>"000010010",
  50004=>"011111011",
  50005=>"101001111",
  50006=>"011000100",
  50007=>"001011100",
  50008=>"101000110",
  50009=>"110010010",
  50010=>"000101111",
  50011=>"001000001",
  50012=>"101111101",
  50013=>"100110111",
  50014=>"101000011",
  50015=>"000010010",
  50016=>"011011001",
  50017=>"100110000",
  50018=>"000000010",
  50019=>"111000110",
  50020=>"110101101",
  50021=>"001001110",
  50022=>"001001000",
  50023=>"100001110",
  50024=>"011111001",
  50025=>"101100100",
  50026=>"001000010",
  50027=>"001010100",
  50028=>"001001110",
  50029=>"110101100",
  50030=>"101000101",
  50031=>"010011001",
  50032=>"101111011",
  50033=>"001100111",
  50034=>"111011000",
  50035=>"011101101",
  50036=>"000110101",
  50037=>"110110011",
  50038=>"000000001",
  50039=>"111001010",
  50040=>"101101100",
  50041=>"000111001",
  50042=>"100001010",
  50043=>"101100111",
  50044=>"011010111",
  50045=>"011101000",
  50046=>"001011111",
  50047=>"001010111",
  50048=>"000001101",
  50049=>"100101010",
  50050=>"011111011",
  50051=>"010000000",
  50052=>"001000001",
  50053=>"110011101",
  50054=>"011001101",
  50055=>"110010001",
  50056=>"001000101",
  50057=>"100010010",
  50058=>"001100000",
  50059=>"100011000",
  50060=>"011101001",
  50061=>"000000000",
  50062=>"011000101",
  50063=>"011111111",
  50064=>"011100111",
  50065=>"011100001",
  50066=>"000011011",
  50067=>"010100000",
  50068=>"000100100",
  50069=>"001011011",
  50070=>"001000010",
  50071=>"100011011",
  50072=>"101110111",
  50073=>"101000110",
  50074=>"100101000",
  50075=>"011000000",
  50076=>"010011111",
  50077=>"011000100",
  50078=>"101110110",
  50079=>"010000101",
  50080=>"000001110",
  50081=>"000010100",
  50082=>"001001101",
  50083=>"000100001",
  50084=>"000001110",
  50085=>"011110000",
  50086=>"001001001",
  50087=>"100010001",
  50088=>"000101111",
  50089=>"111101101",
  50090=>"100100011",
  50091=>"100010101",
  50092=>"110000000",
  50093=>"100100100",
  50094=>"000011000",
  50095=>"011110001",
  50096=>"001111010",
  50097=>"010111011",
  50098=>"100000001",
  50099=>"101111011",
  50100=>"011000100",
  50101=>"100010011",
  50102=>"110001010",
  50103=>"001100111",
  50104=>"111001011",
  50105=>"001010011",
  50106=>"100101100",
  50107=>"111011011",
  50108=>"101001000",
  50109=>"010000001",
  50110=>"001111011",
  50111=>"100100110",
  50112=>"011000100",
  50113=>"000010010",
  50114=>"101000010",
  50115=>"100110001",
  50116=>"001001111",
  50117=>"011111101",
  50118=>"001111000",
  50119=>"001101110",
  50120=>"001111010",
  50121=>"100000101",
  50122=>"100010111",
  50123=>"100001100",
  50124=>"111111111",
  50125=>"110101010",
  50126=>"111001100",
  50127=>"000110111",
  50128=>"101100100",
  50129=>"001101010",
  50130=>"111111001",
  50131=>"010100101",
  50132=>"011001010",
  50133=>"101110000",
  50134=>"111010011",
  50135=>"111000101",
  50136=>"101101101",
  50137=>"100101111",
  50138=>"111110101",
  50139=>"001110010",
  50140=>"000110010",
  50141=>"111001101",
  50142=>"111111100",
  50143=>"110110010",
  50144=>"010111100",
  50145=>"100101110",
  50146=>"001100110",
  50147=>"100010001",
  50148=>"100110100",
  50149=>"000100000",
  50150=>"111110111",
  50151=>"110100100",
  50152=>"000111010",
  50153=>"000101100",
  50154=>"010011000",
  50155=>"001001100",
  50156=>"011001010",
  50157=>"000110100",
  50158=>"111011110",
  50159=>"010110100",
  50160=>"010010010",
  50161=>"000100001",
  50162=>"101000000",
  50163=>"011101011",
  50164=>"000011101",
  50165=>"110100100",
  50166=>"101101111",
  50167=>"001111001",
  50168=>"101111000",
  50169=>"001001100",
  50170=>"011000010",
  50171=>"011111100",
  50172=>"001010000",
  50173=>"100000000",
  50174=>"110010111",
  50175=>"100001011",
  50176=>"010011111",
  50177=>"001110111",
  50178=>"010000101",
  50179=>"101010010",
  50180=>"010110011",
  50181=>"000011111",
  50182=>"000110001",
  50183=>"100110100",
  50184=>"111100001",
  50185=>"001000000",
  50186=>"000000101",
  50187=>"100101011",
  50188=>"000100111",
  50189=>"110101100",
  50190=>"011011000",
  50191=>"110100111",
  50192=>"000111000",
  50193=>"100000110",
  50194=>"100111100",
  50195=>"001101101",
  50196=>"100100101",
  50197=>"011001101",
  50198=>"100100111",
  50199=>"110010010",
  50200=>"100100010",
  50201=>"000010001",
  50202=>"101111100",
  50203=>"000000111",
  50204=>"100100000",
  50205=>"111010011",
  50206=>"100011011",
  50207=>"111111110",
  50208=>"101010110",
  50209=>"100101100",
  50210=>"010001110",
  50211=>"100100001",
  50212=>"101000000",
  50213=>"111010001",
  50214=>"001110101",
  50215=>"000010001",
  50216=>"011010111",
  50217=>"110000001",
  50218=>"100001101",
  50219=>"011111110",
  50220=>"010100110",
  50221=>"101111000",
  50222=>"101001010",
  50223=>"100001010",
  50224=>"000001101",
  50225=>"101000111",
  50226=>"010101001",
  50227=>"011001100",
  50228=>"000010011",
  50229=>"010000101",
  50230=>"000000110",
  50231=>"101111101",
  50232=>"000100001",
  50233=>"001000011",
  50234=>"000111111",
  50235=>"000101001",
  50236=>"000110111",
  50237=>"100111101",
  50238=>"010000010",
  50239=>"011100011",
  50240=>"101001110",
  50241=>"000000101",
  50242=>"110010110",
  50243=>"100010001",
  50244=>"001011001",
  50245=>"000101001",
  50246=>"010000010",
  50247=>"111101111",
  50248=>"111000010",
  50249=>"100111110",
  50250=>"000000100",
  50251=>"001110111",
  50252=>"011111100",
  50253=>"111010000",
  50254=>"011001110",
  50255=>"001111000",
  50256=>"101001101",
  50257=>"001110011",
  50258=>"110001100",
  50259=>"111001110",
  50260=>"000001100",
  50261=>"000100101",
  50262=>"001101000",
  50263=>"000010111",
  50264=>"110111000",
  50265=>"101110100",
  50266=>"111111100",
  50267=>"100100011",
  50268=>"100101100",
  50269=>"000111011",
  50270=>"001000001",
  50271=>"000011011",
  50272=>"100100010",
  50273=>"001100101",
  50274=>"101001101",
  50275=>"000001100",
  50276=>"100110111",
  50277=>"001101100",
  50278=>"000011100",
  50279=>"000101100",
  50280=>"001100100",
  50281=>"111101001",
  50282=>"101110001",
  50283=>"100100101",
  50284=>"111101100",
  50285=>"100000010",
  50286=>"100110011",
  50287=>"101001000",
  50288=>"110100000",
  50289=>"101101010",
  50290=>"110011111",
  50291=>"011011110",
  50292=>"100001001",
  50293=>"101001000",
  50294=>"111011011",
  50295=>"000111001",
  50296=>"101110100",
  50297=>"001011001",
  50298=>"100010110",
  50299=>"010111110",
  50300=>"100101010",
  50301=>"011100101",
  50302=>"000100001",
  50303=>"100001111",
  50304=>"011000011",
  50305=>"111101010",
  50306=>"000011001",
  50307=>"101100101",
  50308=>"010001110",
  50309=>"000000001",
  50310=>"010111011",
  50311=>"001110111",
  50312=>"101111001",
  50313=>"010000000",
  50314=>"110011010",
  50315=>"111001100",
  50316=>"100111110",
  50317=>"111110110",
  50318=>"011010110",
  50319=>"110001010",
  50320=>"010110110",
  50321=>"001111010",
  50322=>"110101000",
  50323=>"111001000",
  50324=>"101100011",
  50325=>"001110101",
  50326=>"010111100",
  50327=>"000000011",
  50328=>"111010001",
  50329=>"000011010",
  50330=>"001110110",
  50331=>"000011101",
  50332=>"101100100",
  50333=>"111010011",
  50334=>"010011111",
  50335=>"010111100",
  50336=>"001100011",
  50337=>"011110000",
  50338=>"010000101",
  50339=>"000001101",
  50340=>"000010101",
  50341=>"110111010",
  50342=>"000010110",
  50343=>"011010011",
  50344=>"110111101",
  50345=>"010010100",
  50346=>"011100010",
  50347=>"000010001",
  50348=>"000111001",
  50349=>"001101010",
  50350=>"101011101",
  50351=>"100100101",
  50352=>"000010000",
  50353=>"010110001",
  50354=>"010010000",
  50355=>"101110101",
  50356=>"110001000",
  50357=>"010110011",
  50358=>"000101000",
  50359=>"101011001",
  50360=>"000110010",
  50361=>"111000100",
  50362=>"111001011",
  50363=>"101110000",
  50364=>"010000010",
  50365=>"111000101",
  50366=>"001101110",
  50367=>"000111010",
  50368=>"001110010",
  50369=>"111001101",
  50370=>"111111000",
  50371=>"010000100",
  50372=>"011100010",
  50373=>"000000100",
  50374=>"101000101",
  50375=>"001100111",
  50376=>"010000100",
  50377=>"101101010",
  50378=>"011001101",
  50379=>"111010101",
  50380=>"111001011",
  50381=>"000010110",
  50382=>"001010001",
  50383=>"010001111",
  50384=>"111110101",
  50385=>"100111101",
  50386=>"101111000",
  50387=>"010010000",
  50388=>"000010010",
  50389=>"100101011",
  50390=>"011001000",
  50391=>"011001101",
  50392=>"010011101",
  50393=>"010100110",
  50394=>"011000010",
  50395=>"100001001",
  50396=>"100001100",
  50397=>"110000110",
  50398=>"001000100",
  50399=>"101011101",
  50400=>"100000000",
  50401=>"010000011",
  50402=>"111111011",
  50403=>"110100010",
  50404=>"010100011",
  50405=>"000110101",
  50406=>"011111000",
  50407=>"011000101",
  50408=>"100000101",
  50409=>"010011110",
  50410=>"010000010",
  50411=>"100000011",
  50412=>"110101101",
  50413=>"101110001",
  50414=>"000000001",
  50415=>"111000000",
  50416=>"001011100",
  50417=>"000010000",
  50418=>"100111000",
  50419=>"111001100",
  50420=>"001010110",
  50421=>"100101011",
  50422=>"110110111",
  50423=>"000001000",
  50424=>"000011111",
  50425=>"111111000",
  50426=>"110001011",
  50427=>"110000110",
  50428=>"111111010",
  50429=>"111001101",
  50430=>"110110111",
  50431=>"111001011",
  50432=>"100001110",
  50433=>"010101010",
  50434=>"001100001",
  50435=>"111101000",
  50436=>"011001110",
  50437=>"001001000",
  50438=>"010001111",
  50439=>"101111111",
  50440=>"011101000",
  50441=>"101010101",
  50442=>"011111110",
  50443=>"111011001",
  50444=>"000101001",
  50445=>"011001100",
  50446=>"101010101",
  50447=>"101010110",
  50448=>"110111110",
  50449=>"011101101",
  50450=>"101111100",
  50451=>"101000001",
  50452=>"011100011",
  50453=>"000101110",
  50454=>"001000000",
  50455=>"010000110",
  50456=>"011011010",
  50457=>"001001011",
  50458=>"010110110",
  50459=>"101111111",
  50460=>"101101111",
  50461=>"011100011",
  50462=>"011110110",
  50463=>"001101110",
  50464=>"000101001",
  50465=>"100100010",
  50466=>"101100101",
  50467=>"110110011",
  50468=>"010101001",
  50469=>"110101100",
  50470=>"010000000",
  50471=>"000101001",
  50472=>"111101001",
  50473=>"110010101",
  50474=>"011000111",
  50475=>"100111010",
  50476=>"110110010",
  50477=>"000100000",
  50478=>"100000100",
  50479=>"110101001",
  50480=>"001110100",
  50481=>"011101000",
  50482=>"101110111",
  50483=>"111100011",
  50484=>"110100101",
  50485=>"001011111",
  50486=>"000100100",
  50487=>"011101001",
  50488=>"011100001",
  50489=>"110011000",
  50490=>"000101000",
  50491=>"100110111",
  50492=>"100101111",
  50493=>"111000001",
  50494=>"011010000",
  50495=>"101001010",
  50496=>"011111111",
  50497=>"100001111",
  50498=>"101010100",
  50499=>"000111000",
  50500=>"110110101",
  50501=>"110011011",
  50502=>"001110101",
  50503=>"110011000",
  50504=>"001110011",
  50505=>"100000001",
  50506=>"000111011",
  50507=>"111000101",
  50508=>"011000111",
  50509=>"011111010",
  50510=>"010111101",
  50511=>"100100101",
  50512=>"100100000",
  50513=>"010011111",
  50514=>"011111100",
  50515=>"101101110",
  50516=>"101000000",
  50517=>"000111100",
  50518=>"111111000",
  50519=>"101001101",
  50520=>"100001000",
  50521=>"000100010",
  50522=>"011001110",
  50523=>"101101011",
  50524=>"111000100",
  50525=>"000111001",
  50526=>"001010001",
  50527=>"100001100",
  50528=>"111000001",
  50529=>"010110111",
  50530=>"110011111",
  50531=>"001100010",
  50532=>"100111101",
  50533=>"100001110",
  50534=>"010101100",
  50535=>"010001100",
  50536=>"010001110",
  50537=>"001011101",
  50538=>"100111000",
  50539=>"100110001",
  50540=>"111000011",
  50541=>"110101100",
  50542=>"100001101",
  50543=>"101101001",
  50544=>"000010000",
  50545=>"001000000",
  50546=>"100001011",
  50547=>"110100000",
  50548=>"111110101",
  50549=>"100001101",
  50550=>"010000000",
  50551=>"111000100",
  50552=>"011110110",
  50553=>"001010111",
  50554=>"101100001",
  50555=>"001111000",
  50556=>"111010101",
  50557=>"111100000",
  50558=>"100111110",
  50559=>"001010011",
  50560=>"110011101",
  50561=>"011111100",
  50562=>"011100011",
  50563=>"111000000",
  50564=>"000100110",
  50565=>"011101111",
  50566=>"101110100",
  50567=>"001011010",
  50568=>"101110111",
  50569=>"100001111",
  50570=>"011010011",
  50571=>"100011110",
  50572=>"001010100",
  50573=>"110011101",
  50574=>"100111001",
  50575=>"110001001",
  50576=>"100110010",
  50577=>"000000001",
  50578=>"000100000",
  50579=>"011000100",
  50580=>"100101000",
  50581=>"101111011",
  50582=>"000000011",
  50583=>"101100011",
  50584=>"101000111",
  50585=>"101001000",
  50586=>"010111101",
  50587=>"101000010",
  50588=>"011011001",
  50589=>"100011010",
  50590=>"000101110",
  50591=>"110100111",
  50592=>"100001000",
  50593=>"111010110",
  50594=>"001010111",
  50595=>"101001101",
  50596=>"000001001",
  50597=>"001011000",
  50598=>"110111111",
  50599=>"101010100",
  50600=>"111100101",
  50601=>"111011011",
  50602=>"000001000",
  50603=>"001000110",
  50604=>"011101100",
  50605=>"110010101",
  50606=>"000101000",
  50607=>"101000100",
  50608=>"111000000",
  50609=>"101001001",
  50610=>"100000001",
  50611=>"001010101",
  50612=>"000100001",
  50613=>"011101010",
  50614=>"010001100",
  50615=>"001001000",
  50616=>"000101000",
  50617=>"001010101",
  50618=>"001001000",
  50619=>"010011011",
  50620=>"100111111",
  50621=>"001110101",
  50622=>"100011011",
  50623=>"101111010",
  50624=>"101100101",
  50625=>"101000001",
  50626=>"001101010",
  50627=>"101000111",
  50628=>"110001111",
  50629=>"001000010",
  50630=>"000100000",
  50631=>"100000001",
  50632=>"111111011",
  50633=>"001001000",
  50634=>"110000101",
  50635=>"010011111",
  50636=>"010101000",
  50637=>"010011000",
  50638=>"100110001",
  50639=>"111011111",
  50640=>"010110001",
  50641=>"011011100",
  50642=>"101110101",
  50643=>"100010110",
  50644=>"110011000",
  50645=>"110010010",
  50646=>"001011101",
  50647=>"100000000",
  50648=>"000001100",
  50649=>"111000101",
  50650=>"111110110",
  50651=>"001000000",
  50652=>"001000000",
  50653=>"101001010",
  50654=>"110010111",
  50655=>"000100010",
  50656=>"001111000",
  50657=>"101011010",
  50658=>"110010000",
  50659=>"110000100",
  50660=>"100100100",
  50661=>"010001011",
  50662=>"101010101",
  50663=>"111101000",
  50664=>"111100011",
  50665=>"001101011",
  50666=>"101010110",
  50667=>"111110000",
  50668=>"101100000",
  50669=>"001101101",
  50670=>"001010111",
  50671=>"100010000",
  50672=>"001110000",
  50673=>"001000110",
  50674=>"011000011",
  50675=>"100011010",
  50676=>"011101100",
  50677=>"110100100",
  50678=>"111100111",
  50679=>"010100110",
  50680=>"000100100",
  50681=>"001100011",
  50682=>"000000010",
  50683=>"000111010",
  50684=>"001110000",
  50685=>"101010100",
  50686=>"110000010",
  50687=>"010000000",
  50688=>"011010111",
  50689=>"000001001",
  50690=>"111011000",
  50691=>"101010110",
  50692=>"110101100",
  50693=>"010011010",
  50694=>"101100001",
  50695=>"011011001",
  50696=>"000011100",
  50697=>"110000100",
  50698=>"011110100",
  50699=>"000000000",
  50700=>"001110111",
  50701=>"111011111",
  50702=>"000000000",
  50703=>"110010101",
  50704=>"101010100",
  50705=>"011110111",
  50706=>"100010001",
  50707=>"111100110",
  50708=>"000010011",
  50709=>"000011010",
  50710=>"001000111",
  50711=>"011000110",
  50712=>"101110011",
  50713=>"101111000",
  50714=>"110011100",
  50715=>"101010111",
  50716=>"111110001",
  50717=>"111010000",
  50718=>"101001101",
  50719=>"010010110",
  50720=>"010011111",
  50721=>"110010110",
  50722=>"011100000",
  50723=>"001001100",
  50724=>"101111100",
  50725=>"010100000",
  50726=>"100011011",
  50727=>"110111100",
  50728=>"100000100",
  50729=>"111001110",
  50730=>"110000101",
  50731=>"111000100",
  50732=>"001000100",
  50733=>"100111000",
  50734=>"000010101",
  50735=>"110010001",
  50736=>"000111110",
  50737=>"101100100",
  50738=>"000100010",
  50739=>"000011011",
  50740=>"100010111",
  50741=>"011011110",
  50742=>"111010100",
  50743=>"001000110",
  50744=>"001000011",
  50745=>"000001101",
  50746=>"010000010",
  50747=>"111100001",
  50748=>"000010100",
  50749=>"111100111",
  50750=>"000100100",
  50751=>"000110001",
  50752=>"000111000",
  50753=>"100010011",
  50754=>"001110011",
  50755=>"010010001",
  50756=>"000000100",
  50757=>"111100101",
  50758=>"100000101",
  50759=>"100111001",
  50760=>"010110000",
  50761=>"111100111",
  50762=>"011000001",
  50763=>"100111100",
  50764=>"110100110",
  50765=>"010101100",
  50766=>"110111100",
  50767=>"011011111",
  50768=>"110010010",
  50769=>"001000001",
  50770=>"000111111",
  50771=>"000000100",
  50772=>"111010111",
  50773=>"001001010",
  50774=>"000111011",
  50775=>"101110101",
  50776=>"011100101",
  50777=>"011011000",
  50778=>"010100100",
  50779=>"100000010",
  50780=>"001011101",
  50781=>"000100100",
  50782=>"001001101",
  50783=>"011010010",
  50784=>"010011110",
  50785=>"110011000",
  50786=>"010001111",
  50787=>"001000100",
  50788=>"011000010",
  50789=>"101101001",
  50790=>"010010101",
  50791=>"001011000",
  50792=>"110000101",
  50793=>"001011011",
  50794=>"111010000",
  50795=>"111000000",
  50796=>"001100111",
  50797=>"111010000",
  50798=>"100001100",
  50799=>"111101110",
  50800=>"111111001",
  50801=>"101100000",
  50802=>"011010111",
  50803=>"011110110",
  50804=>"010011101",
  50805=>"010111000",
  50806=>"100110001",
  50807=>"100110001",
  50808=>"110111111",
  50809=>"101001011",
  50810=>"100101111",
  50811=>"011111101",
  50812=>"100010101",
  50813=>"110111001",
  50814=>"001100100",
  50815=>"101011111",
  50816=>"010011101",
  50817=>"111011101",
  50818=>"000110011",
  50819=>"011011000",
  50820=>"001100111",
  50821=>"010010000",
  50822=>"010011100",
  50823=>"010111001",
  50824=>"101100011",
  50825=>"111001000",
  50826=>"101010011",
  50827=>"100100111",
  50828=>"100000000",
  50829=>"101000000",
  50830=>"011000010",
  50831=>"101000110",
  50832=>"110011011",
  50833=>"011100100",
  50834=>"111100111",
  50835=>"100001101",
  50836=>"000110010",
  50837=>"100011111",
  50838=>"111001000",
  50839=>"010111001",
  50840=>"010100110",
  50841=>"111100011",
  50842=>"000010100",
  50843=>"111010111",
  50844=>"000001010",
  50845=>"111101001",
  50846=>"011001001",
  50847=>"100001111",
  50848=>"001011001",
  50849=>"001111100",
  50850=>"001011010",
  50851=>"111111101",
  50852=>"010101111",
  50853=>"010001000",
  50854=>"001000000",
  50855=>"010100010",
  50856=>"011100000",
  50857=>"111010011",
  50858=>"000001100",
  50859=>"001101001",
  50860=>"110011111",
  50861=>"010101011",
  50862=>"101000110",
  50863=>"001011010",
  50864=>"010110110",
  50865=>"111111110",
  50866=>"111100001",
  50867=>"111110100",
  50868=>"111010100",
  50869=>"001111111",
  50870=>"100011000",
  50871=>"000100000",
  50872=>"011001010",
  50873=>"101110101",
  50874=>"001100010",
  50875=>"000000110",
  50876=>"100110111",
  50877=>"110011000",
  50878=>"000010100",
  50879=>"101011011",
  50880=>"000000111",
  50881=>"100011101",
  50882=>"000001010",
  50883=>"110101011",
  50884=>"001010100",
  50885=>"011011000",
  50886=>"011010001",
  50887=>"100111111",
  50888=>"111100000",
  50889=>"011110101",
  50890=>"110101000",
  50891=>"111001001",
  50892=>"010100001",
  50893=>"110011000",
  50894=>"100001111",
  50895=>"111101110",
  50896=>"110101100",
  50897=>"010011101",
  50898=>"110001011",
  50899=>"000000111",
  50900=>"010100010",
  50901=>"100001110",
  50902=>"001000110",
  50903=>"000111001",
  50904=>"000000111",
  50905=>"101111110",
  50906=>"001001000",
  50907=>"101110000",
  50908=>"110000000",
  50909=>"001000111",
  50910=>"101000111",
  50911=>"000110101",
  50912=>"011001110",
  50913=>"001100000",
  50914=>"100110100",
  50915=>"010111010",
  50916=>"111011011",
  50917=>"001011000",
  50918=>"100110000",
  50919=>"110101111",
  50920=>"010010100",
  50921=>"111000111",
  50922=>"110111110",
  50923=>"101110100",
  50924=>"010001001",
  50925=>"000110111",
  50926=>"110111011",
  50927=>"101101010",
  50928=>"111101101",
  50929=>"011100001",
  50930=>"011111110",
  50931=>"100110101",
  50932=>"100100101",
  50933=>"011000001",
  50934=>"000111011",
  50935=>"001010110",
  50936=>"010001101",
  50937=>"000010111",
  50938=>"010101110",
  50939=>"111010010",
  50940=>"011101111",
  50941=>"000000000",
  50942=>"000111010",
  50943=>"000111000",
  50944=>"001001110",
  50945=>"001000000",
  50946=>"000011110",
  50947=>"011100001",
  50948=>"100000101",
  50949=>"000100100",
  50950=>"011101011",
  50951=>"100000000",
  50952=>"011001010",
  50953=>"111001111",
  50954=>"001011111",
  50955=>"010101110",
  50956=>"001000100",
  50957=>"010010101",
  50958=>"010010001",
  50959=>"011111011",
  50960=>"001111110",
  50961=>"010100010",
  50962=>"111001101",
  50963=>"111001000",
  50964=>"000100110",
  50965=>"001010110",
  50966=>"011010101",
  50967=>"001101011",
  50968=>"000011100",
  50969=>"010100011",
  50970=>"000010101",
  50971=>"111010101",
  50972=>"110001100",
  50973=>"111100101",
  50974=>"010100001",
  50975=>"101001001",
  50976=>"010111001",
  50977=>"101001100",
  50978=>"111101011",
  50979=>"010100010",
  50980=>"101110100",
  50981=>"001000001",
  50982=>"000010011",
  50983=>"011111110",
  50984=>"101010011",
  50985=>"111000101",
  50986=>"100000000",
  50987=>"101001111",
  50988=>"010010100",
  50989=>"000000100",
  50990=>"000011000",
  50991=>"001111111",
  50992=>"000010011",
  50993=>"111010010",
  50994=>"001111000",
  50995=>"011111100",
  50996=>"100100000",
  50997=>"100100010",
  50998=>"100010010",
  50999=>"101100111",
  51000=>"111101010",
  51001=>"000010000",
  51002=>"101010100",
  51003=>"100100001",
  51004=>"011011001",
  51005=>"101001000",
  51006=>"010001000",
  51007=>"011010100",
  51008=>"100001000",
  51009=>"010111011",
  51010=>"100000111",
  51011=>"001000011",
  51012=>"000000000",
  51013=>"001101110",
  51014=>"101111100",
  51015=>"011011010",
  51016=>"001100000",
  51017=>"111111010",
  51018=>"011011010",
  51019=>"000110000",
  51020=>"001100100",
  51021=>"010111100",
  51022=>"000011100",
  51023=>"010101111",
  51024=>"010101111",
  51025=>"011110000",
  51026=>"000000100",
  51027=>"010011001",
  51028=>"111100000",
  51029=>"101101110",
  51030=>"000010000",
  51031=>"010010101",
  51032=>"100111011",
  51033=>"001000110",
  51034=>"011000001",
  51035=>"101000000",
  51036=>"010010100",
  51037=>"000000000",
  51038=>"111001010",
  51039=>"010001101",
  51040=>"101100110",
  51041=>"001010101",
  51042=>"000000010",
  51043=>"000111100",
  51044=>"000100010",
  51045=>"100000101",
  51046=>"000110011",
  51047=>"110010000",
  51048=>"101011000",
  51049=>"110011101",
  51050=>"100100100",
  51051=>"111001011",
  51052=>"010000111",
  51053=>"110010101",
  51054=>"100100001",
  51055=>"010010000",
  51056=>"010001110",
  51057=>"111011111",
  51058=>"101010010",
  51059=>"110110010",
  51060=>"000011010",
  51061=>"000010100",
  51062=>"110100000",
  51063=>"001000110",
  51064=>"101010010",
  51065=>"100101000",
  51066=>"100100111",
  51067=>"101101101",
  51068=>"010111101",
  51069=>"101001100",
  51070=>"111000101",
  51071=>"110011100",
  51072=>"010111100",
  51073=>"000111011",
  51074=>"111011011",
  51075=>"000011111",
  51076=>"101111100",
  51077=>"100001011",
  51078=>"101101111",
  51079=>"001100111",
  51080=>"110100001",
  51081=>"000010101",
  51082=>"110001111",
  51083=>"001010010",
  51084=>"111110101",
  51085=>"000100010",
  51086=>"011001110",
  51087=>"100011111",
  51088=>"100110110",
  51089=>"101001010",
  51090=>"101011001",
  51091=>"111000101",
  51092=>"101001100",
  51093=>"100101100",
  51094=>"111101011",
  51095=>"100010110",
  51096=>"111000001",
  51097=>"111010101",
  51098=>"000010100",
  51099=>"000101000",
  51100=>"101101000",
  51101=>"101100010",
  51102=>"000111101",
  51103=>"111000011",
  51104=>"100000111",
  51105=>"111000101",
  51106=>"000101100",
  51107=>"001100100",
  51108=>"010011010",
  51109=>"010111111",
  51110=>"101110101",
  51111=>"101011001",
  51112=>"100000101",
  51113=>"000111110",
  51114=>"011100110",
  51115=>"010111010",
  51116=>"010011111",
  51117=>"000101110",
  51118=>"011111110",
  51119=>"001010100",
  51120=>"110001101",
  51121=>"111000100",
  51122=>"010010000",
  51123=>"110001010",
  51124=>"010000010",
  51125=>"100110000",
  51126=>"110110111",
  51127=>"101110111",
  51128=>"011010100",
  51129=>"100010100",
  51130=>"100111110",
  51131=>"100110010",
  51132=>"101001100",
  51133=>"011000011",
  51134=>"010011000",
  51135=>"000101100",
  51136=>"111101111",
  51137=>"101001110",
  51138=>"111100000",
  51139=>"001011100",
  51140=>"011000010",
  51141=>"100010100",
  51142=>"101001001",
  51143=>"101001011",
  51144=>"000101100",
  51145=>"101001110",
  51146=>"111111011",
  51147=>"110011100",
  51148=>"101110001",
  51149=>"011000101",
  51150=>"001010100",
  51151=>"001111111",
  51152=>"011101000",
  51153=>"110000001",
  51154=>"011001101",
  51155=>"110010110",
  51156=>"000110000",
  51157=>"101111111",
  51158=>"011000110",
  51159=>"010000101",
  51160=>"000110111",
  51161=>"001111101",
  51162=>"001001011",
  51163=>"111111111",
  51164=>"100111000",
  51165=>"110110000",
  51166=>"110001111",
  51167=>"101101010",
  51168=>"101011110",
  51169=>"101110001",
  51170=>"101101001",
  51171=>"001001101",
  51172=>"000001001",
  51173=>"000110000",
  51174=>"010011100",
  51175=>"100101111",
  51176=>"011000010",
  51177=>"101010010",
  51178=>"100100001",
  51179=>"010000010",
  51180=>"000011110",
  51181=>"011010111",
  51182=>"101000101",
  51183=>"001100110",
  51184=>"000111001",
  51185=>"010110001",
  51186=>"111100111",
  51187=>"000111100",
  51188=>"110110111",
  51189=>"011111101",
  51190=>"011101101",
  51191=>"000111001",
  51192=>"000001111",
  51193=>"110111000",
  51194=>"001111001",
  51195=>"010101000",
  51196=>"001110101",
  51197=>"100000100",
  51198=>"011010010",
  51199=>"011111011",
  51200=>"001010001",
  51201=>"110100000",
  51202=>"110100011",
  51203=>"101011001",
  51204=>"011010111",
  51205=>"101100110",
  51206=>"110111100",
  51207=>"000000011",
  51208=>"100001011",
  51209=>"010111101",
  51210=>"011101000",
  51211=>"100111001",
  51212=>"101011001",
  51213=>"000110100",
  51214=>"011101001",
  51215=>"100100001",
  51216=>"111100111",
  51217=>"000011110",
  51218=>"110110110",
  51219=>"001100100",
  51220=>"100001010",
  51221=>"010101101",
  51222=>"100100000",
  51223=>"100001110",
  51224=>"101000000",
  51225=>"001111000",
  51226=>"100101111",
  51227=>"000111001",
  51228=>"000000101",
  51229=>"101000010",
  51230=>"011111101",
  51231=>"011010010",
  51232=>"110000010",
  51233=>"010000011",
  51234=>"110101111",
  51235=>"101010000",
  51236=>"101011000",
  51237=>"001001100",
  51238=>"001010101",
  51239=>"000100000",
  51240=>"000001001",
  51241=>"100010110",
  51242=>"100111100",
  51243=>"100100011",
  51244=>"100100101",
  51245=>"001001010",
  51246=>"110001010",
  51247=>"101001100",
  51248=>"000001101",
  51249=>"101101001",
  51250=>"011000110",
  51251=>"111101111",
  51252=>"101010010",
  51253=>"110011001",
  51254=>"011000000",
  51255=>"101011111",
  51256=>"110000010",
  51257=>"000001100",
  51258=>"101000110",
  51259=>"110011111",
  51260=>"110110111",
  51261=>"101001000",
  51262=>"000110001",
  51263=>"110010101",
  51264=>"101100111",
  51265=>"010100101",
  51266=>"000001101",
  51267=>"101101011",
  51268=>"100011011",
  51269=>"000010000",
  51270=>"001101101",
  51271=>"010101110",
  51272=>"100111100",
  51273=>"100010110",
  51274=>"011010110",
  51275=>"001000011",
  51276=>"101000100",
  51277=>"110001101",
  51278=>"011110010",
  51279=>"000000011",
  51280=>"101101001",
  51281=>"000010101",
  51282=>"001011011",
  51283=>"110111000",
  51284=>"010010110",
  51285=>"110011000",
  51286=>"011110001",
  51287=>"010000111",
  51288=>"001011011",
  51289=>"001100010",
  51290=>"101011111",
  51291=>"100100000",
  51292=>"011111111",
  51293=>"111000111",
  51294=>"010111111",
  51295=>"010000110",
  51296=>"101000011",
  51297=>"000000001",
  51298=>"001001110",
  51299=>"100001110",
  51300=>"001011110",
  51301=>"100011010",
  51302=>"000000000",
  51303=>"000000100",
  51304=>"110010010",
  51305=>"010001001",
  51306=>"010000101",
  51307=>"010010011",
  51308=>"000010101",
  51309=>"001001011",
  51310=>"110000111",
  51311=>"100111100",
  51312=>"010000001",
  51313=>"010111101",
  51314=>"101010100",
  51315=>"000101101",
  51316=>"010111110",
  51317=>"110101110",
  51318=>"011010011",
  51319=>"001001001",
  51320=>"101100001",
  51321=>"110011011",
  51322=>"000101100",
  51323=>"010000101",
  51324=>"011110000",
  51325=>"000010110",
  51326=>"001011111",
  51327=>"000010111",
  51328=>"001000001",
  51329=>"100001010",
  51330=>"010011111",
  51331=>"110110100",
  51332=>"101111000",
  51333=>"000111100",
  51334=>"000001110",
  51335=>"110010100",
  51336=>"111011111",
  51337=>"001000000",
  51338=>"010101100",
  51339=>"110001111",
  51340=>"000101110",
  51341=>"010011000",
  51342=>"001001100",
  51343=>"110110010",
  51344=>"111111111",
  51345=>"010110010",
  51346=>"000001011",
  51347=>"100011111",
  51348=>"000010001",
  51349=>"000101111",
  51350=>"001100001",
  51351=>"010101010",
  51352=>"001010001",
  51353=>"010001001",
  51354=>"001101000",
  51355=>"101000010",
  51356=>"000110000",
  51357=>"111111110",
  51358=>"110011000",
  51359=>"001111110",
  51360=>"101000100",
  51361=>"101110000",
  51362=>"100010100",
  51363=>"100000011",
  51364=>"100100000",
  51365=>"000101101",
  51366=>"001010100",
  51367=>"101110100",
  51368=>"010000001",
  51369=>"100100010",
  51370=>"001001000",
  51371=>"101100111",
  51372=>"011011000",
  51373=>"111000110",
  51374=>"000111001",
  51375=>"101000000",
  51376=>"100101101",
  51377=>"011001111",
  51378=>"101111000",
  51379=>"000011110",
  51380=>"110100001",
  51381=>"010110100",
  51382=>"100110000",
  51383=>"010001000",
  51384=>"100000100",
  51385=>"001011010",
  51386=>"101100100",
  51387=>"100111000",
  51388=>"101100011",
  51389=>"011001001",
  51390=>"100100000",
  51391=>"101001010",
  51392=>"011011010",
  51393=>"111111110",
  51394=>"010111001",
  51395=>"010110000",
  51396=>"100000111",
  51397=>"111111010",
  51398=>"011000110",
  51399=>"010111111",
  51400=>"111110010",
  51401=>"111011111",
  51402=>"011111110",
  51403=>"100100001",
  51404=>"100101101",
  51405=>"101111010",
  51406=>"111110001",
  51407=>"010101101",
  51408=>"101110111",
  51409=>"001100100",
  51410=>"001010001",
  51411=>"100000001",
  51412=>"011101010",
  51413=>"101011110",
  51414=>"011110101",
  51415=>"001111111",
  51416=>"101110001",
  51417=>"010110000",
  51418=>"000110110",
  51419=>"001001101",
  51420=>"001000100",
  51421=>"011100011",
  51422=>"100111110",
  51423=>"110001001",
  51424=>"011001011",
  51425=>"001110011",
  51426=>"101100101",
  51427=>"000010000",
  51428=>"011011101",
  51429=>"100011111",
  51430=>"001100000",
  51431=>"101011010",
  51432=>"100000010",
  51433=>"111110101",
  51434=>"111010110",
  51435=>"011110111",
  51436=>"000100110",
  51437=>"000001000",
  51438=>"110101111",
  51439=>"010000100",
  51440=>"110010011",
  51441=>"100010111",
  51442=>"011011010",
  51443=>"100011001",
  51444=>"000100100",
  51445=>"011101100",
  51446=>"011000100",
  51447=>"010000101",
  51448=>"100110101",
  51449=>"101101110",
  51450=>"101010000",
  51451=>"111000101",
  51452=>"100010010",
  51453=>"101000100",
  51454=>"110010100",
  51455=>"011001011",
  51456=>"010011010",
  51457=>"001101010",
  51458=>"011110111",
  51459=>"000010010",
  51460=>"011000011",
  51461=>"110011101",
  51462=>"011100001",
  51463=>"010010000",
  51464=>"101011101",
  51465=>"110111110",
  51466=>"010100011",
  51467=>"000000100",
  51468=>"100010001",
  51469=>"001000111",
  51470=>"101100100",
  51471=>"100010010",
  51472=>"101101111",
  51473=>"001001111",
  51474=>"100101010",
  51475=>"110000111",
  51476=>"010101101",
  51477=>"001000010",
  51478=>"100000110",
  51479=>"000101010",
  51480=>"110100000",
  51481=>"011101110",
  51482=>"101000011",
  51483=>"000010101",
  51484=>"001110100",
  51485=>"100110100",
  51486=>"010110000",
  51487=>"001000110",
  51488=>"111000001",
  51489=>"000101000",
  51490=>"001011010",
  51491=>"111101110",
  51492=>"101111110",
  51493=>"010101111",
  51494=>"011100001",
  51495=>"010111101",
  51496=>"110010001",
  51497=>"000111100",
  51498=>"110011100",
  51499=>"000011101",
  51500=>"100000000",
  51501=>"110101111",
  51502=>"000100011",
  51503=>"001100010",
  51504=>"101100110",
  51505=>"111001000",
  51506=>"101100001",
  51507=>"000111111",
  51508=>"011000111",
  51509=>"100010101",
  51510=>"010110000",
  51511=>"100101010",
  51512=>"111101101",
  51513=>"100100101",
  51514=>"000111101",
  51515=>"110101110",
  51516=>"100101001",
  51517=>"000010100",
  51518=>"001100111",
  51519=>"100001011",
  51520=>"111101100",
  51521=>"001111001",
  51522=>"001010000",
  51523=>"101000010",
  51524=>"110011100",
  51525=>"100110010",
  51526=>"000001011",
  51527=>"111010110",
  51528=>"011001100",
  51529=>"010001001",
  51530=>"011010001",
  51531=>"001000110",
  51532=>"001100011",
  51533=>"010011101",
  51534=>"100100000",
  51535=>"010101000",
  51536=>"111010000",
  51537=>"011111110",
  51538=>"100010101",
  51539=>"011101000",
  51540=>"100010101",
  51541=>"101001110",
  51542=>"101010000",
  51543=>"101100011",
  51544=>"000000100",
  51545=>"011100011",
  51546=>"011100001",
  51547=>"100011111",
  51548=>"111000011",
  51549=>"111000010",
  51550=>"010101010",
  51551=>"000010010",
  51552=>"001011101",
  51553=>"100011000",
  51554=>"001100101",
  51555=>"000011111",
  51556=>"111101000",
  51557=>"111110100",
  51558=>"001001111",
  51559=>"101001010",
  51560=>"010001001",
  51561=>"010110011",
  51562=>"010101000",
  51563=>"001001111",
  51564=>"100011100",
  51565=>"011000011",
  51566=>"001001110",
  51567=>"110111111",
  51568=>"011111011",
  51569=>"101000110",
  51570=>"110010000",
  51571=>"010000101",
  51572=>"001011010",
  51573=>"011100000",
  51574=>"011111001",
  51575=>"011010101",
  51576=>"111010100",
  51577=>"011110010",
  51578=>"011000000",
  51579=>"001001101",
  51580=>"000111001",
  51581=>"110110001",
  51582=>"100110010",
  51583=>"011011000",
  51584=>"111100000",
  51585=>"010001000",
  51586=>"100111111",
  51587=>"010110011",
  51588=>"011100001",
  51589=>"100111011",
  51590=>"111110110",
  51591=>"001111111",
  51592=>"100001101",
  51593=>"100001111",
  51594=>"010101010",
  51595=>"000000011",
  51596=>"000000000",
  51597=>"000110100",
  51598=>"001010011",
  51599=>"001110000",
  51600=>"001100001",
  51601=>"011000000",
  51602=>"100110000",
  51603=>"010100001",
  51604=>"100000000",
  51605=>"000100111",
  51606=>"000000000",
  51607=>"010111011",
  51608=>"000110000",
  51609=>"000010000",
  51610=>"010011110",
  51611=>"010000001",
  51612=>"010110000",
  51613=>"110101101",
  51614=>"110010010",
  51615=>"101111111",
  51616=>"101101010",
  51617=>"010111001",
  51618=>"010101110",
  51619=>"101000100",
  51620=>"100100000",
  51621=>"111010111",
  51622=>"001101110",
  51623=>"101000011",
  51624=>"011110000",
  51625=>"101011110",
  51626=>"000101011",
  51627=>"111101101",
  51628=>"100101101",
  51629=>"111101000",
  51630=>"110101100",
  51631=>"011110010",
  51632=>"000001110",
  51633=>"110111000",
  51634=>"010000111",
  51635=>"111111001",
  51636=>"111010010",
  51637=>"111110101",
  51638=>"111111110",
  51639=>"111110010",
  51640=>"101110000",
  51641=>"100110101",
  51642=>"101001000",
  51643=>"100101101",
  51644=>"110110000",
  51645=>"000001111",
  51646=>"001100001",
  51647=>"010010001",
  51648=>"110111011",
  51649=>"110111111",
  51650=>"000111010",
  51651=>"001010000",
  51652=>"001100010",
  51653=>"100111100",
  51654=>"000010001",
  51655=>"110001111",
  51656=>"010110100",
  51657=>"001111101",
  51658=>"111111111",
  51659=>"011011110",
  51660=>"111010001",
  51661=>"101011010",
  51662=>"100111111",
  51663=>"000101101",
  51664=>"100000001",
  51665=>"100000000",
  51666=>"111100000",
  51667=>"111010100",
  51668=>"100101100",
  51669=>"010010000",
  51670=>"000100010",
  51671=>"000001110",
  51672=>"111000111",
  51673=>"110110000",
  51674=>"000110100",
  51675=>"111000100",
  51676=>"011011010",
  51677=>"000110101",
  51678=>"000101001",
  51679=>"000100111",
  51680=>"001101000",
  51681=>"011001011",
  51682=>"000111011",
  51683=>"000001101",
  51684=>"011111000",
  51685=>"010010010",
  51686=>"110100111",
  51687=>"110101111",
  51688=>"110111111",
  51689=>"100000011",
  51690=>"000001111",
  51691=>"111100101",
  51692=>"101000101",
  51693=>"011001111",
  51694=>"001100100",
  51695=>"100100111",
  51696=>"001010111",
  51697=>"000010001",
  51698=>"110110010",
  51699=>"010011011",
  51700=>"111001100",
  51701=>"101011111",
  51702=>"110001101",
  51703=>"111100000",
  51704=>"001010111",
  51705=>"011110101",
  51706=>"100110100",
  51707=>"001100000",
  51708=>"100010100",
  51709=>"000100010",
  51710=>"000110101",
  51711=>"111100011",
  51712=>"001110100",
  51713=>"010011110",
  51714=>"100111101",
  51715=>"000010000",
  51716=>"001100110",
  51717=>"001111101",
  51718=>"101000110",
  51719=>"011001110",
  51720=>"000011100",
  51721=>"100011101",
  51722=>"010100011",
  51723=>"100010010",
  51724=>"011101001",
  51725=>"101101011",
  51726=>"010011000",
  51727=>"111000010",
  51728=>"110010101",
  51729=>"011001100",
  51730=>"110010100",
  51731=>"101111000",
  51732=>"110000011",
  51733=>"001111000",
  51734=>"011001001",
  51735=>"111101011",
  51736=>"010001111",
  51737=>"101011110",
  51738=>"001110011",
  51739=>"100111010",
  51740=>"010000001",
  51741=>"111000010",
  51742=>"101011111",
  51743=>"000111111",
  51744=>"110111010",
  51745=>"001101101",
  51746=>"010001010",
  51747=>"100101110",
  51748=>"111100100",
  51749=>"001011101",
  51750=>"101001010",
  51751=>"111001001",
  51752=>"010000011",
  51753=>"100101001",
  51754=>"001011011",
  51755=>"111001111",
  51756=>"100101110",
  51757=>"010001000",
  51758=>"101101110",
  51759=>"000000110",
  51760=>"111101101",
  51761=>"110101111",
  51762=>"000001111",
  51763=>"100010000",
  51764=>"000101011",
  51765=>"101010100",
  51766=>"000001101",
  51767=>"110110010",
  51768=>"010001111",
  51769=>"110000111",
  51770=>"000111011",
  51771=>"100100010",
  51772=>"000100010",
  51773=>"001011011",
  51774=>"011100101",
  51775=>"101000100",
  51776=>"111000100",
  51777=>"111110001",
  51778=>"101000011",
  51779=>"000001111",
  51780=>"110101101",
  51781=>"001110100",
  51782=>"101010101",
  51783=>"010000001",
  51784=>"011011001",
  51785=>"011101110",
  51786=>"000001010",
  51787=>"000011010",
  51788=>"001100100",
  51789=>"110011010",
  51790=>"001111101",
  51791=>"101001111",
  51792=>"110101101",
  51793=>"011001011",
  51794=>"001111000",
  51795=>"000111110",
  51796=>"100010110",
  51797=>"101100110",
  51798=>"101101100",
  51799=>"001000101",
  51800=>"001101001",
  51801=>"111100011",
  51802=>"101010100",
  51803=>"111101110",
  51804=>"000011010",
  51805=>"001110111",
  51806=>"111101001",
  51807=>"010010100",
  51808=>"101111101",
  51809=>"101110011",
  51810=>"111000111",
  51811=>"001101000",
  51812=>"111001010",
  51813=>"011101101",
  51814=>"000101010",
  51815=>"110010000",
  51816=>"100110011",
  51817=>"000110001",
  51818=>"001001110",
  51819=>"111000110",
  51820=>"100100011",
  51821=>"101000010",
  51822=>"100001110",
  51823=>"010000100",
  51824=>"110100011",
  51825=>"111000001",
  51826=>"100001010",
  51827=>"111100010",
  51828=>"101010111",
  51829=>"000100001",
  51830=>"100011110",
  51831=>"111100111",
  51832=>"001111111",
  51833=>"010111011",
  51834=>"000010010",
  51835=>"011010010",
  51836=>"110110011",
  51837=>"100001111",
  51838=>"110000101",
  51839=>"000000000",
  51840=>"001010100",
  51841=>"001111010",
  51842=>"011001110",
  51843=>"000011001",
  51844=>"011111111",
  51845=>"111000010",
  51846=>"001011110",
  51847=>"001100100",
  51848=>"011101010",
  51849=>"111010001",
  51850=>"111011000",
  51851=>"010101110",
  51852=>"110101111",
  51853=>"000001111",
  51854=>"010111001",
  51855=>"101010011",
  51856=>"011010010",
  51857=>"111101100",
  51858=>"101000001",
  51859=>"111110000",
  51860=>"001000011",
  51861=>"011100110",
  51862=>"010101011",
  51863=>"111110100",
  51864=>"000111101",
  51865=>"111111000",
  51866=>"000110101",
  51867=>"101100001",
  51868=>"100100110",
  51869=>"101001101",
  51870=>"100111111",
  51871=>"010110000",
  51872=>"000100000",
  51873=>"000000000",
  51874=>"110110111",
  51875=>"000101101",
  51876=>"111111100",
  51877=>"111100100",
  51878=>"100100111",
  51879=>"111000001",
  51880=>"100001000",
  51881=>"101001111",
  51882=>"111001011",
  51883=>"110100011",
  51884=>"001000100",
  51885=>"011011101",
  51886=>"010001000",
  51887=>"111010010",
  51888=>"001010010",
  51889=>"100000110",
  51890=>"000111111",
  51891=>"010011000",
  51892=>"110101011",
  51893=>"000111001",
  51894=>"010100011",
  51895=>"110011000",
  51896=>"111000111",
  51897=>"000000100",
  51898=>"100110001",
  51899=>"111010111",
  51900=>"001011010",
  51901=>"010110100",
  51902=>"100000110",
  51903=>"000111110",
  51904=>"100111110",
  51905=>"011111100",
  51906=>"000100101",
  51907=>"101111011",
  51908=>"010101110",
  51909=>"010010101",
  51910=>"100010010",
  51911=>"000100010",
  51912=>"001100001",
  51913=>"000000000",
  51914=>"110110111",
  51915=>"000010001",
  51916=>"111111100",
  51917=>"111101011",
  51918=>"111111001",
  51919=>"111100010",
  51920=>"110001010",
  51921=>"100111011",
  51922=>"010111010",
  51923=>"001001101",
  51924=>"001001011",
  51925=>"010000011",
  51926=>"011011001",
  51927=>"101111010",
  51928=>"001111011",
  51929=>"010101001",
  51930=>"101100011",
  51931=>"001101000",
  51932=>"100101101",
  51933=>"010111101",
  51934=>"111100011",
  51935=>"101100100",
  51936=>"001011010",
  51937=>"100000110",
  51938=>"110000000",
  51939=>"111000101",
  51940=>"000010110",
  51941=>"101110001",
  51942=>"110100110",
  51943=>"000111101",
  51944=>"001000010",
  51945=>"001111010",
  51946=>"111110010",
  51947=>"111011011",
  51948=>"010011111",
  51949=>"001111001",
  51950=>"000001111",
  51951=>"010111011",
  51952=>"011011010",
  51953=>"101010110",
  51954=>"010011011",
  51955=>"001111101",
  51956=>"101001111",
  51957=>"001110100",
  51958=>"101000110",
  51959=>"100111011",
  51960=>"011100011",
  51961=>"101010000",
  51962=>"001011111",
  51963=>"010010010",
  51964=>"000001000",
  51965=>"001101011",
  51966=>"010000001",
  51967=>"011111101",
  51968=>"000100011",
  51969=>"000110000",
  51970=>"001001111",
  51971=>"101101100",
  51972=>"101000100",
  51973=>"001000011",
  51974=>"101101011",
  51975=>"100101110",
  51976=>"010011000",
  51977=>"010111001",
  51978=>"000101001",
  51979=>"011000110",
  51980=>"001110101",
  51981=>"111000100",
  51982=>"000000111",
  51983=>"001110011",
  51984=>"011000011",
  51985=>"010101010",
  51986=>"101110000",
  51987=>"100110010",
  51988=>"111001101",
  51989=>"100000010",
  51990=>"100101000",
  51991=>"001101001",
  51992=>"011010110",
  51993=>"110001000",
  51994=>"100111101",
  51995=>"010011011",
  51996=>"100001100",
  51997=>"110101100",
  51998=>"001010010",
  51999=>"110000011",
  52000=>"001011111",
  52001=>"111000101",
  52002=>"001011101",
  52003=>"000111101",
  52004=>"010100100",
  52005=>"100100000",
  52006=>"000001101",
  52007=>"001001000",
  52008=>"100101000",
  52009=>"111010101",
  52010=>"110000001",
  52011=>"110011101",
  52012=>"001001010",
  52013=>"001100010",
  52014=>"001011101",
  52015=>"010001111",
  52016=>"000111010",
  52017=>"111001111",
  52018=>"001010010",
  52019=>"011100010",
  52020=>"000000101",
  52021=>"110001001",
  52022=>"010100000",
  52023=>"010001101",
  52024=>"101011001",
  52025=>"000111011",
  52026=>"010010100",
  52027=>"011111111",
  52028=>"001001110",
  52029=>"110001011",
  52030=>"001001000",
  52031=>"100010100",
  52032=>"010100010",
  52033=>"010100111",
  52034=>"110000010",
  52035=>"000010111",
  52036=>"110001010",
  52037=>"010000111",
  52038=>"110111000",
  52039=>"011111101",
  52040=>"111001000",
  52041=>"011110011",
  52042=>"010100110",
  52043=>"000001001",
  52044=>"000000101",
  52045=>"001011111",
  52046=>"101111111",
  52047=>"100010111",
  52048=>"100101010",
  52049=>"111000111",
  52050=>"111011010",
  52051=>"100111110",
  52052=>"011011100",
  52053=>"000010100",
  52054=>"000010010",
  52055=>"000011001",
  52056=>"010000000",
  52057=>"101011001",
  52058=>"100001011",
  52059=>"000011010",
  52060=>"101011111",
  52061=>"101101000",
  52062=>"010010011",
  52063=>"000011111",
  52064=>"010111011",
  52065=>"000101101",
  52066=>"110011100",
  52067=>"000100000",
  52068=>"011101110",
  52069=>"111000011",
  52070=>"011100011",
  52071=>"000001000",
  52072=>"101110011",
  52073=>"111011011",
  52074=>"101011010",
  52075=>"000111010",
  52076=>"100111011",
  52077=>"110000111",
  52078=>"111101001",
  52079=>"110111000",
  52080=>"001001010",
  52081=>"111000001",
  52082=>"110111100",
  52083=>"000101100",
  52084=>"111100011",
  52085=>"111001000",
  52086=>"011111001",
  52087=>"110000101",
  52088=>"000001110",
  52089=>"100000010",
  52090=>"101101100",
  52091=>"000110110",
  52092=>"001000000",
  52093=>"010000100",
  52094=>"011101011",
  52095=>"000111101",
  52096=>"110100001",
  52097=>"101011111",
  52098=>"100001101",
  52099=>"111100101",
  52100=>"110000000",
  52101=>"101101010",
  52102=>"111100010",
  52103=>"101000011",
  52104=>"111110100",
  52105=>"101001101",
  52106=>"111010110",
  52107=>"100011010",
  52108=>"011100110",
  52109=>"001011010",
  52110=>"110010010",
  52111=>"000111000",
  52112=>"000111111",
  52113=>"001110111",
  52114=>"001101010",
  52115=>"001010111",
  52116=>"110110101",
  52117=>"101011000",
  52118=>"010111101",
  52119=>"110001010",
  52120=>"011001110",
  52121=>"111010001",
  52122=>"001101111",
  52123=>"011100000",
  52124=>"001101101",
  52125=>"011111100",
  52126=>"101010001",
  52127=>"001111100",
  52128=>"111010110",
  52129=>"111100111",
  52130=>"110101010",
  52131=>"010101100",
  52132=>"000111101",
  52133=>"111010000",
  52134=>"110111000",
  52135=>"100000101",
  52136=>"010000111",
  52137=>"001010110",
  52138=>"111111000",
  52139=>"010001000",
  52140=>"101000010",
  52141=>"011111111",
  52142=>"010001100",
  52143=>"110101111",
  52144=>"011001011",
  52145=>"010110100",
  52146=>"111100011",
  52147=>"100110110",
  52148=>"011010010",
  52149=>"001101000",
  52150=>"110101000",
  52151=>"011101110",
  52152=>"011100111",
  52153=>"001110110",
  52154=>"011001010",
  52155=>"000010000",
  52156=>"100000010",
  52157=>"111001010",
  52158=>"100100000",
  52159=>"000011000",
  52160=>"011100110",
  52161=>"110100101",
  52162=>"010010110",
  52163=>"010000010",
  52164=>"101000101",
  52165=>"100000000",
  52166=>"100111001",
  52167=>"001101110",
  52168=>"000010001",
  52169=>"011011000",
  52170=>"110111100",
  52171=>"011111011",
  52172=>"101001100",
  52173=>"001100001",
  52174=>"000111001",
  52175=>"100110001",
  52176=>"000110010",
  52177=>"011001110",
  52178=>"000101010",
  52179=>"101001100",
  52180=>"111001000",
  52181=>"110100111",
  52182=>"101011100",
  52183=>"000011000",
  52184=>"101000110",
  52185=>"110110010",
  52186=>"011101101",
  52187=>"101000101",
  52188=>"011011100",
  52189=>"111011001",
  52190=>"110000011",
  52191=>"011010110",
  52192=>"001001000",
  52193=>"111110111",
  52194=>"010001000",
  52195=>"100011111",
  52196=>"000001110",
  52197=>"010110000",
  52198=>"100001000",
  52199=>"010110111",
  52200=>"111000011",
  52201=>"001110001",
  52202=>"110010011",
  52203=>"100000000",
  52204=>"010000110",
  52205=>"110011001",
  52206=>"001000101",
  52207=>"100011010",
  52208=>"011011000",
  52209=>"000111110",
  52210=>"010100000",
  52211=>"001010100",
  52212=>"010111010",
  52213=>"000101100",
  52214=>"000001100",
  52215=>"101000001",
  52216=>"100001011",
  52217=>"001010110",
  52218=>"011111000",
  52219=>"000000111",
  52220=>"000111110",
  52221=>"110111111",
  52222=>"001000011",
  52223=>"111000111",
  52224=>"111101100",
  52225=>"111111100",
  52226=>"010010101",
  52227=>"111100000",
  52228=>"000111111",
  52229=>"100011111",
  52230=>"101001010",
  52231=>"000010000",
  52232=>"001010011",
  52233=>"001111101",
  52234=>"100100010",
  52235=>"000111110",
  52236=>"110100000",
  52237=>"011111100",
  52238=>"000011010",
  52239=>"001011000",
  52240=>"110000110",
  52241=>"101001001",
  52242=>"100100000",
  52243=>"000001101",
  52244=>"100001100",
  52245=>"111101100",
  52246=>"001110100",
  52247=>"111000010",
  52248=>"011110001",
  52249=>"110110111",
  52250=>"101001010",
  52251=>"100100110",
  52252=>"111110111",
  52253=>"110011011",
  52254=>"111001100",
  52255=>"000001111",
  52256=>"000100001",
  52257=>"011000011",
  52258=>"010010010",
  52259=>"010011111",
  52260=>"000001110",
  52261=>"010111000",
  52262=>"110110001",
  52263=>"111011011",
  52264=>"110010011",
  52265=>"010101001",
  52266=>"001011111",
  52267=>"100011110",
  52268=>"110111100",
  52269=>"001010000",
  52270=>"111010001",
  52271=>"101011000",
  52272=>"001011000",
  52273=>"100000000",
  52274=>"111101100",
  52275=>"000110100",
  52276=>"001110000",
  52277=>"111010111",
  52278=>"100011010",
  52279=>"100011111",
  52280=>"000011010",
  52281=>"110101110",
  52282=>"101010100",
  52283=>"100000011",
  52284=>"001111111",
  52285=>"001111101",
  52286=>"001011000",
  52287=>"101111001",
  52288=>"111100110",
  52289=>"000001111",
  52290=>"101100111",
  52291=>"111010000",
  52292=>"001111100",
  52293=>"100001011",
  52294=>"110000001",
  52295=>"110010101",
  52296=>"101010000",
  52297=>"110101110",
  52298=>"101000110",
  52299=>"011100100",
  52300=>"111011001",
  52301=>"001010000",
  52302=>"011110111",
  52303=>"100010101",
  52304=>"000010010",
  52305=>"000000100",
  52306=>"001111101",
  52307=>"111100011",
  52308=>"000010110",
  52309=>"110110000",
  52310=>"011010101",
  52311=>"011110001",
  52312=>"101100000",
  52313=>"011100100",
  52314=>"101100010",
  52315=>"010111101",
  52316=>"101011111",
  52317=>"001101010",
  52318=>"001001001",
  52319=>"101100000",
  52320=>"001110100",
  52321=>"110110100",
  52322=>"111100111",
  52323=>"000111110",
  52324=>"011100000",
  52325=>"001100000",
  52326=>"110011001",
  52327=>"101110111",
  52328=>"011001000",
  52329=>"001101100",
  52330=>"001000101",
  52331=>"110000000",
  52332=>"110000010",
  52333=>"000111000",
  52334=>"010000101",
  52335=>"111101111",
  52336=>"000101011",
  52337=>"011100111",
  52338=>"000111010",
  52339=>"100110111",
  52340=>"111001011",
  52341=>"100111110",
  52342=>"110110010",
  52343=>"100011100",
  52344=>"111100111",
  52345=>"100010000",
  52346=>"111011010",
  52347=>"101111101",
  52348=>"101111111",
  52349=>"000011111",
  52350=>"111110110",
  52351=>"100110000",
  52352=>"100010011",
  52353=>"111110000",
  52354=>"000011100",
  52355=>"011000011",
  52356=>"111011000",
  52357=>"111111100",
  52358=>"011101011",
  52359=>"101110111",
  52360=>"010100001",
  52361=>"100100110",
  52362=>"001111000",
  52363=>"000010100",
  52364=>"111101100",
  52365=>"110000100",
  52366=>"101001010",
  52367=>"111101111",
  52368=>"111001110",
  52369=>"000000001",
  52370=>"111010010",
  52371=>"000011000",
  52372=>"111101111",
  52373=>"111000010",
  52374=>"011100110",
  52375=>"111100100",
  52376=>"010111100",
  52377=>"101101111",
  52378=>"010000010",
  52379=>"111001010",
  52380=>"001000001",
  52381=>"111010100",
  52382=>"010010000",
  52383=>"101010011",
  52384=>"111101111",
  52385=>"111010101",
  52386=>"111100011",
  52387=>"111001010",
  52388=>"101101000",
  52389=>"011000100",
  52390=>"000001110",
  52391=>"001110100",
  52392=>"001111010",
  52393=>"010111000",
  52394=>"011010000",
  52395=>"010101010",
  52396=>"000011011",
  52397=>"001001000",
  52398=>"011010111",
  52399=>"000101000",
  52400=>"010110100",
  52401=>"101000100",
  52402=>"001101001",
  52403=>"110010101",
  52404=>"110000111",
  52405=>"111001111",
  52406=>"001010100",
  52407=>"111111011",
  52408=>"111010010",
  52409=>"000000000",
  52410=>"101010000",
  52411=>"101100100",
  52412=>"111011001",
  52413=>"000100010",
  52414=>"101111111",
  52415=>"100101101",
  52416=>"111001110",
  52417=>"000100000",
  52418=>"111010111",
  52419=>"001110101",
  52420=>"000010111",
  52421=>"110100111",
  52422=>"101010011",
  52423=>"101001110",
  52424=>"100000111",
  52425=>"010010101",
  52426=>"101001000",
  52427=>"100101011",
  52428=>"101000001",
  52429=>"101110110",
  52430=>"111001100",
  52431=>"111100010",
  52432=>"111000001",
  52433=>"100110000",
  52434=>"000101010",
  52435=>"111001111",
  52436=>"000110010",
  52437=>"010100110",
  52438=>"110100001",
  52439=>"100001001",
  52440=>"100010100",
  52441=>"100011111",
  52442=>"111001110",
  52443=>"000111110",
  52444=>"101110000",
  52445=>"111101110",
  52446=>"000010010",
  52447=>"001011011",
  52448=>"010111000",
  52449=>"110101011",
  52450=>"000111111",
  52451=>"100000010",
  52452=>"011111111",
  52453=>"101000111",
  52454=>"100011111",
  52455=>"010010100",
  52456=>"001010100",
  52457=>"110001100",
  52458=>"101000010",
  52459=>"010111011",
  52460=>"011111100",
  52461=>"101010001",
  52462=>"100011000",
  52463=>"100010001",
  52464=>"010100000",
  52465=>"110100110",
  52466=>"111111001",
  52467=>"111010100",
  52468=>"111000011",
  52469=>"110100001",
  52470=>"100101001",
  52471=>"001001101",
  52472=>"101111011",
  52473=>"110111111",
  52474=>"000100110",
  52475=>"010001100",
  52476=>"010000010",
  52477=>"111111111",
  52478=>"010000000",
  52479=>"010101100",
  52480=>"011010100",
  52481=>"101001011",
  52482=>"101101000",
  52483=>"001100110",
  52484=>"101111110",
  52485=>"111000001",
  52486=>"101010110",
  52487=>"011000101",
  52488=>"101010111",
  52489=>"010111111",
  52490=>"100011110",
  52491=>"010100101",
  52492=>"111011110",
  52493=>"110101100",
  52494=>"000101101",
  52495=>"010010110",
  52496=>"011100010",
  52497=>"011001100",
  52498=>"100001010",
  52499=>"110101100",
  52500=>"100011111",
  52501=>"100101000",
  52502=>"000101110",
  52503=>"111011011",
  52504=>"010000000",
  52505=>"011111011",
  52506=>"011000111",
  52507=>"101000111",
  52508=>"110100110",
  52509=>"111100001",
  52510=>"101011001",
  52511=>"111000100",
  52512=>"010000110",
  52513=>"000010000",
  52514=>"011000101",
  52515=>"100000001",
  52516=>"101011000",
  52517=>"001110010",
  52518=>"011000000",
  52519=>"001010101",
  52520=>"010110110",
  52521=>"010101101",
  52522=>"100010010",
  52523=>"010111011",
  52524=>"110111010",
  52525=>"010001010",
  52526=>"101101111",
  52527=>"100011111",
  52528=>"111110101",
  52529=>"101001110",
  52530=>"010010011",
  52531=>"100000111",
  52532=>"011000100",
  52533=>"100110110",
  52534=>"100001111",
  52535=>"111111100",
  52536=>"101011010",
  52537=>"010100001",
  52538=>"000010100",
  52539=>"101111000",
  52540=>"010101101",
  52541=>"011111111",
  52542=>"000101010",
  52543=>"111100111",
  52544=>"001000001",
  52545=>"001101011",
  52546=>"010100000",
  52547=>"101100011",
  52548=>"111001100",
  52549=>"111010101",
  52550=>"011111110",
  52551=>"111111001",
  52552=>"011100000",
  52553=>"101011001",
  52554=>"111011011",
  52555=>"011100111",
  52556=>"010010010",
  52557=>"110010010",
  52558=>"001100001",
  52559=>"110001010",
  52560=>"110100010",
  52561=>"111000100",
  52562=>"010010100",
  52563=>"001101100",
  52564=>"001001000",
  52565=>"001010100",
  52566=>"110001101",
  52567=>"000101111",
  52568=>"111001110",
  52569=>"000010111",
  52570=>"010000001",
  52571=>"010000110",
  52572=>"001011101",
  52573=>"011100110",
  52574=>"010010111",
  52575=>"001011000",
  52576=>"011101110",
  52577=>"010001101",
  52578=>"011100101",
  52579=>"111001111",
  52580=>"101110101",
  52581=>"111011111",
  52582=>"100111101",
  52583=>"011000001",
  52584=>"101011001",
  52585=>"111110001",
  52586=>"111001010",
  52587=>"000000111",
  52588=>"011111010",
  52589=>"000000011",
  52590=>"011000110",
  52591=>"110000111",
  52592=>"000001110",
  52593=>"110111000",
  52594=>"001001011",
  52595=>"011011110",
  52596=>"001101111",
  52597=>"101011000",
  52598=>"000101010",
  52599=>"000111111",
  52600=>"011010011",
  52601=>"111111010",
  52602=>"110010010",
  52603=>"001001110",
  52604=>"010110110",
  52605=>"111100110",
  52606=>"011001000",
  52607=>"101001010",
  52608=>"111011011",
  52609=>"110110000",
  52610=>"011101101",
  52611=>"001000110",
  52612=>"110101100",
  52613=>"011110010",
  52614=>"100001000",
  52615=>"101011000",
  52616=>"100111001",
  52617=>"000111001",
  52618=>"010001000",
  52619=>"110100000",
  52620=>"000000110",
  52621=>"000000111",
  52622=>"000100101",
  52623=>"111010010",
  52624=>"110110001",
  52625=>"110101010",
  52626=>"010001010",
  52627=>"100110011",
  52628=>"001011111",
  52629=>"001011101",
  52630=>"000111001",
  52631=>"011001000",
  52632=>"111110110",
  52633=>"101001101",
  52634=>"101011111",
  52635=>"011110011",
  52636=>"011101111",
  52637=>"100111111",
  52638=>"001110100",
  52639=>"011011110",
  52640=>"001111111",
  52641=>"110011011",
  52642=>"111110110",
  52643=>"001010000",
  52644=>"001101011",
  52645=>"010100111",
  52646=>"010001000",
  52647=>"011000010",
  52648=>"001101000",
  52649=>"010100001",
  52650=>"010100111",
  52651=>"101001011",
  52652=>"000001010",
  52653=>"101001111",
  52654=>"011111000",
  52655=>"100100100",
  52656=>"000100010",
  52657=>"000011110",
  52658=>"100111100",
  52659=>"101010010",
  52660=>"000111111",
  52661=>"100000110",
  52662=>"111001111",
  52663=>"111011000",
  52664=>"101010100",
  52665=>"010011010",
  52666=>"001100010",
  52667=>"011010100",
  52668=>"110100111",
  52669=>"010011010",
  52670=>"001101111",
  52671=>"011001001",
  52672=>"110000111",
  52673=>"100111111",
  52674=>"111010010",
  52675=>"000010110",
  52676=>"111011111",
  52677=>"010000011",
  52678=>"001101110",
  52679=>"111000111",
  52680=>"111000101",
  52681=>"011000111",
  52682=>"111011110",
  52683=>"010101100",
  52684=>"101100110",
  52685=>"010000101",
  52686=>"111110101",
  52687=>"100100010",
  52688=>"011110110",
  52689=>"111111100",
  52690=>"011111001",
  52691=>"101111000",
  52692=>"100101111",
  52693=>"011011110",
  52694=>"110000011",
  52695=>"100100101",
  52696=>"110010101",
  52697=>"011000011",
  52698=>"111100110",
  52699=>"000100010",
  52700=>"000001110",
  52701=>"001111000",
  52702=>"100101000",
  52703=>"000100111",
  52704=>"101001000",
  52705=>"000001010",
  52706=>"000011101",
  52707=>"000001110",
  52708=>"000101001",
  52709=>"111111000",
  52710=>"111000100",
  52711=>"101110100",
  52712=>"010011111",
  52713=>"001011101",
  52714=>"000010101",
  52715=>"010001000",
  52716=>"011100100",
  52717=>"100001110",
  52718=>"111110110",
  52719=>"000000101",
  52720=>"000011101",
  52721=>"011000110",
  52722=>"101010100",
  52723=>"011110001",
  52724=>"111100011",
  52725=>"100111111",
  52726=>"111111111",
  52727=>"101100011",
  52728=>"001110111",
  52729=>"001110111",
  52730=>"010101001",
  52731=>"011010110",
  52732=>"001001100",
  52733=>"010111111",
  52734=>"010001101",
  52735=>"100010111",
  52736=>"110011001",
  52737=>"100100100",
  52738=>"101001101",
  52739=>"000110110",
  52740=>"101111110",
  52741=>"111011110",
  52742=>"010111010",
  52743=>"110110000",
  52744=>"000011000",
  52745=>"111001101",
  52746=>"000111010",
  52747=>"110011001",
  52748=>"101100100",
  52749=>"010101000",
  52750=>"100011111",
  52751=>"010011001",
  52752=>"100110010",
  52753=>"110111001",
  52754=>"010010001",
  52755=>"101111111",
  52756=>"110011100",
  52757=>"011100001",
  52758=>"111111000",
  52759=>"101001101",
  52760=>"000111010",
  52761=>"111100011",
  52762=>"111011100",
  52763=>"100111100",
  52764=>"111110001",
  52765=>"011111110",
  52766=>"111111011",
  52767=>"001001001",
  52768=>"100110010",
  52769=>"011011000",
  52770=>"011001000",
  52771=>"010110000",
  52772=>"011011000",
  52773=>"111011101",
  52774=>"110100011",
  52775=>"100111101",
  52776=>"001100100",
  52777=>"101110110",
  52778=>"001111100",
  52779=>"110011011",
  52780=>"100110000",
  52781=>"100000110",
  52782=>"010100110",
  52783=>"111101101",
  52784=>"010010110",
  52785=>"010001110",
  52786=>"111100011",
  52787=>"011011000",
  52788=>"010110100",
  52789=>"110001011",
  52790=>"110100100",
  52791=>"010010101",
  52792=>"100001000",
  52793=>"011101011",
  52794=>"000011100",
  52795=>"111110101",
  52796=>"100010111",
  52797=>"111101110",
  52798=>"101100100",
  52799=>"010011111",
  52800=>"100000110",
  52801=>"101000100",
  52802=>"001100011",
  52803=>"100111110",
  52804=>"001000001",
  52805=>"001101000",
  52806=>"101001110",
  52807=>"110011001",
  52808=>"100010100",
  52809=>"111101011",
  52810=>"101000000",
  52811=>"100100101",
  52812=>"000111001",
  52813=>"000001110",
  52814=>"011110110",
  52815=>"010110101",
  52816=>"110001010",
  52817=>"101001111",
  52818=>"100101000",
  52819=>"001001011",
  52820=>"010010010",
  52821=>"110001000",
  52822=>"100110101",
  52823=>"111000001",
  52824=>"101010001",
  52825=>"001010110",
  52826=>"111110101",
  52827=>"001000000",
  52828=>"110010100",
  52829=>"010011011",
  52830=>"111000110",
  52831=>"010000000",
  52832=>"001000100",
  52833=>"101011011",
  52834=>"110010111",
  52835=>"011110111",
  52836=>"011001010",
  52837=>"000011110",
  52838=>"010101110",
  52839=>"000001010",
  52840=>"011011100",
  52841=>"010101111",
  52842=>"101110101",
  52843=>"100110000",
  52844=>"010100010",
  52845=>"011001100",
  52846=>"000111010",
  52847=>"101100101",
  52848=>"100000100",
  52849=>"101101001",
  52850=>"010101000",
  52851=>"100000001",
  52852=>"110000111",
  52853=>"101000111",
  52854=>"000010110",
  52855=>"011000011",
  52856=>"110100111",
  52857=>"111101100",
  52858=>"000001110",
  52859=>"011110001",
  52860=>"000000100",
  52861=>"001000110",
  52862=>"110100111",
  52863=>"011101111",
  52864=>"100001111",
  52865=>"101010111",
  52866=>"100010111",
  52867=>"001011110",
  52868=>"011010100",
  52869=>"011100111",
  52870=>"100010010",
  52871=>"100110011",
  52872=>"111111001",
  52873=>"000101010",
  52874=>"110000011",
  52875=>"001010011",
  52876=>"101001100",
  52877=>"010000001",
  52878=>"111101000",
  52879=>"001011101",
  52880=>"110000000",
  52881=>"011111111",
  52882=>"010100000",
  52883=>"101101001",
  52884=>"000101101",
  52885=>"010101110",
  52886=>"001110011",
  52887=>"010110111",
  52888=>"001100110",
  52889=>"110001011",
  52890=>"000000111",
  52891=>"101011011",
  52892=>"011111011",
  52893=>"100101111",
  52894=>"101100010",
  52895=>"110101000",
  52896=>"010110001",
  52897=>"001111101",
  52898=>"000000010",
  52899=>"001001100",
  52900=>"111011101",
  52901=>"101111010",
  52902=>"111011100",
  52903=>"000100100",
  52904=>"101111101",
  52905=>"000100001",
  52906=>"101110100",
  52907=>"001011101",
  52908=>"110111111",
  52909=>"101110101",
  52910=>"100000011",
  52911=>"000010000",
  52912=>"100101110",
  52913=>"111001010",
  52914=>"001010000",
  52915=>"100001111",
  52916=>"001000011",
  52917=>"110101100",
  52918=>"101100010",
  52919=>"100001000",
  52920=>"000000000",
  52921=>"111011110",
  52922=>"101011001",
  52923=>"001011110",
  52924=>"000110000",
  52925=>"011010011",
  52926=>"000001101",
  52927=>"001101100",
  52928=>"000000011",
  52929=>"001001101",
  52930=>"011101011",
  52931=>"101100011",
  52932=>"011001100",
  52933=>"111010111",
  52934=>"010001000",
  52935=>"111111001",
  52936=>"011110100",
  52937=>"000110000",
  52938=>"111100010",
  52939=>"100010001",
  52940=>"110001101",
  52941=>"001000011",
  52942=>"000001000",
  52943=>"000000101",
  52944=>"100110110",
  52945=>"000100110",
  52946=>"101110001",
  52947=>"110001011",
  52948=>"011010011",
  52949=>"100000110",
  52950=>"001100110",
  52951=>"000000011",
  52952=>"000100100",
  52953=>"000100101",
  52954=>"101000111",
  52955=>"110111000",
  52956=>"111111110",
  52957=>"100100001",
  52958=>"000111011",
  52959=>"010001111",
  52960=>"100101000",
  52961=>"100011010",
  52962=>"011101010",
  52963=>"011000101",
  52964=>"101110011",
  52965=>"100100100",
  52966=>"010110011",
  52967=>"111001011",
  52968=>"000011111",
  52969=>"101010000",
  52970=>"010100011",
  52971=>"001001000",
  52972=>"000111101",
  52973=>"010100101",
  52974=>"011111110",
  52975=>"111011101",
  52976=>"001010011",
  52977=>"000000100",
  52978=>"010000000",
  52979=>"011001100",
  52980=>"010101000",
  52981=>"000110101",
  52982=>"010110111",
  52983=>"111001100",
  52984=>"001111010",
  52985=>"100110010",
  52986=>"010111100",
  52987=>"010101000",
  52988=>"110010101",
  52989=>"111111111",
  52990=>"101111000",
  52991=>"110110010",
  52992=>"001000000",
  52993=>"110110011",
  52994=>"000001100",
  52995=>"101100010",
  52996=>"110110011",
  52997=>"010000000",
  52998=>"011111010",
  52999=>"100110001",
  53000=>"000010010",
  53001=>"101011100",
  53002=>"111001001",
  53003=>"001000111",
  53004=>"011001000",
  53005=>"101010111",
  53006=>"101011101",
  53007=>"010111100",
  53008=>"110011110",
  53009=>"101001001",
  53010=>"000000000",
  53011=>"101011011",
  53012=>"110001001",
  53013=>"110010111",
  53014=>"000100001",
  53015=>"011001000",
  53016=>"001101101",
  53017=>"001111010",
  53018=>"000101101",
  53019=>"110111111",
  53020=>"110111111",
  53021=>"111110111",
  53022=>"111101100",
  53023=>"010010000",
  53024=>"001111111",
  53025=>"101010001",
  53026=>"010101000",
  53027=>"111011011",
  53028=>"010110100",
  53029=>"111011011",
  53030=>"100111111",
  53031=>"100000101",
  53032=>"111011100",
  53033=>"110001110",
  53034=>"011011110",
  53035=>"000100111",
  53036=>"001100100",
  53037=>"010100011",
  53038=>"001000000",
  53039=>"010000010",
  53040=>"011111000",
  53041=>"111010001",
  53042=>"011101100",
  53043=>"011100111",
  53044=>"101110001",
  53045=>"100001001",
  53046=>"000010100",
  53047=>"001010011",
  53048=>"011010011",
  53049=>"001000101",
  53050=>"100100100",
  53051=>"111111000",
  53052=>"110010110",
  53053=>"101111110",
  53054=>"100110001",
  53055=>"010001000",
  53056=>"101100111",
  53057=>"100100010",
  53058=>"011010000",
  53059=>"001110110",
  53060=>"101100110",
  53061=>"100111010",
  53062=>"000001111",
  53063=>"101010110",
  53064=>"010010111",
  53065=>"011101000",
  53066=>"000100100",
  53067=>"101001010",
  53068=>"101011110",
  53069=>"111101001",
  53070=>"010010010",
  53071=>"101110101",
  53072=>"111101110",
  53073=>"000110111",
  53074=>"111001111",
  53075=>"110100000",
  53076=>"000110000",
  53077=>"010010011",
  53078=>"100110101",
  53079=>"010110110",
  53080=>"011000110",
  53081=>"011100001",
  53082=>"100101011",
  53083=>"000110001",
  53084=>"100101100",
  53085=>"011010001",
  53086=>"010001001",
  53087=>"111011010",
  53088=>"101110110",
  53089=>"111110111",
  53090=>"111100110",
  53091=>"011100001",
  53092=>"011001111",
  53093=>"011101000",
  53094=>"010011110",
  53095=>"000111000",
  53096=>"011111001",
  53097=>"000111110",
  53098=>"111110000",
  53099=>"111101110",
  53100=>"010001000",
  53101=>"100000111",
  53102=>"011010100",
  53103=>"100100001",
  53104=>"101010110",
  53105=>"111101000",
  53106=>"101011001",
  53107=>"011110111",
  53108=>"011111001",
  53109=>"010100001",
  53110=>"101111000",
  53111=>"110110101",
  53112=>"000111101",
  53113=>"000010000",
  53114=>"011010101",
  53115=>"101010000",
  53116=>"100000100",
  53117=>"011011100",
  53118=>"110001000",
  53119=>"111100011",
  53120=>"100001111",
  53121=>"110000000",
  53122=>"011100001",
  53123=>"000010011",
  53124=>"010101010",
  53125=>"010100011",
  53126=>"101001011",
  53127=>"110010010",
  53128=>"011011100",
  53129=>"111001100",
  53130=>"111101000",
  53131=>"111111100",
  53132=>"101100101",
  53133=>"001101001",
  53134=>"010001011",
  53135=>"110100100",
  53136=>"111011000",
  53137=>"001101110",
  53138=>"110001000",
  53139=>"110001111",
  53140=>"001001010",
  53141=>"011011001",
  53142=>"010111111",
  53143=>"111111001",
  53144=>"011101100",
  53145=>"001011000",
  53146=>"100101101",
  53147=>"010001111",
  53148=>"110011010",
  53149=>"101010010",
  53150=>"011000000",
  53151=>"100101001",
  53152=>"111011101",
  53153=>"010000100",
  53154=>"100001001",
  53155=>"100100001",
  53156=>"101001001",
  53157=>"101101001",
  53158=>"011110000",
  53159=>"001011100",
  53160=>"001010010",
  53161=>"000000001",
  53162=>"101111111",
  53163=>"011101001",
  53164=>"011011101",
  53165=>"101011000",
  53166=>"100001111",
  53167=>"110101001",
  53168=>"101111001",
  53169=>"000100011",
  53170=>"100100110",
  53171=>"101011101",
  53172=>"110000111",
  53173=>"100010111",
  53174=>"101001101",
  53175=>"100100110",
  53176=>"000100100",
  53177=>"000010100",
  53178=>"001011001",
  53179=>"000001111",
  53180=>"010000100",
  53181=>"111001101",
  53182=>"101111111",
  53183=>"101101001",
  53184=>"011110010",
  53185=>"011101011",
  53186=>"001000110",
  53187=>"000000100",
  53188=>"000101010",
  53189=>"101000001",
  53190=>"011111100",
  53191=>"011000111",
  53192=>"110100001",
  53193=>"100011101",
  53194=>"010000110",
  53195=>"010010111",
  53196=>"001000011",
  53197=>"011111001",
  53198=>"101011010",
  53199=>"000010010",
  53200=>"000011101",
  53201=>"000010000",
  53202=>"001110100",
  53203=>"101100101",
  53204=>"001010100",
  53205=>"100011111",
  53206=>"001001011",
  53207=>"000111100",
  53208=>"011010110",
  53209=>"111111001",
  53210=>"000011011",
  53211=>"100001110",
  53212=>"001110000",
  53213=>"001001000",
  53214=>"111010001",
  53215=>"000001000",
  53216=>"110010111",
  53217=>"101110110",
  53218=>"000100001",
  53219=>"111010111",
  53220=>"100011110",
  53221=>"110010100",
  53222=>"011110111",
  53223=>"000001101",
  53224=>"100110100",
  53225=>"001000101",
  53226=>"011000111",
  53227=>"001010111",
  53228=>"010010101",
  53229=>"001000000",
  53230=>"100000010",
  53231=>"010001101",
  53232=>"001111010",
  53233=>"101011010",
  53234=>"100001011",
  53235=>"110010000",
  53236=>"011010001",
  53237=>"111001001",
  53238=>"100100100",
  53239=>"110111001",
  53240=>"101110000",
  53241=>"000101011",
  53242=>"010101111",
  53243=>"100001011",
  53244=>"111101100",
  53245=>"000010111",
  53246=>"111101010",
  53247=>"011101001",
  53248=>"001010001",
  53249=>"010101101",
  53250=>"011011011",
  53251=>"000001011",
  53252=>"100011110",
  53253=>"000011101",
  53254=>"101111101",
  53255=>"000001000",
  53256=>"001011100",
  53257=>"100011000",
  53258=>"101011111",
  53259=>"000001111",
  53260=>"001011100",
  53261=>"001101100",
  53262=>"010100001",
  53263=>"011101011",
  53264=>"001001001",
  53265=>"010110110",
  53266=>"000000100",
  53267=>"011101110",
  53268=>"110010000",
  53269=>"101010111",
  53270=>"001010011",
  53271=>"101000110",
  53272=>"001000001",
  53273=>"000101110",
  53274=>"010110111",
  53275=>"000000010",
  53276=>"011110010",
  53277=>"111111100",
  53278=>"101000111",
  53279=>"100011001",
  53280=>"011101001",
  53281=>"111001100",
  53282=>"101111100",
  53283=>"101000100",
  53284=>"101000000",
  53285=>"001101010",
  53286=>"110101010",
  53287=>"010101001",
  53288=>"111101011",
  53289=>"011000101",
  53290=>"111101110",
  53291=>"101111111",
  53292=>"000000011",
  53293=>"110011111",
  53294=>"001000001",
  53295=>"100101011",
  53296=>"000010010",
  53297=>"000011001",
  53298=>"110111001",
  53299=>"100011010",
  53300=>"100011100",
  53301=>"001110100",
  53302=>"101010001",
  53303=>"111000111",
  53304=>"001000100",
  53305=>"000111111",
  53306=>"101100101",
  53307=>"111100101",
  53308=>"001000101",
  53309=>"011011111",
  53310=>"000001010",
  53311=>"011111111",
  53312=>"000111000",
  53313=>"010001111",
  53314=>"111111010",
  53315=>"110111110",
  53316=>"100011101",
  53317=>"010100100",
  53318=>"100111001",
  53319=>"111010111",
  53320=>"001001000",
  53321=>"110111110",
  53322=>"111101101",
  53323=>"101111110",
  53324=>"001111111",
  53325=>"010110000",
  53326=>"101111000",
  53327=>"010000110",
  53328=>"011001111",
  53329=>"101011111",
  53330=>"111011101",
  53331=>"111100111",
  53332=>"110000100",
  53333=>"100101011",
  53334=>"101011010",
  53335=>"011100011",
  53336=>"100001001",
  53337=>"010001110",
  53338=>"010000000",
  53339=>"010000000",
  53340=>"000111111",
  53341=>"111011101",
  53342=>"111000011",
  53343=>"110000111",
  53344=>"010101100",
  53345=>"011100111",
  53346=>"100111000",
  53347=>"111110111",
  53348=>"000100001",
  53349=>"110010010",
  53350=>"000010011",
  53351=>"011111011",
  53352=>"001001110",
  53353=>"000000110",
  53354=>"001000110",
  53355=>"110001111",
  53356=>"000111010",
  53357=>"010110110",
  53358=>"011000100",
  53359=>"010101110",
  53360=>"101001011",
  53361=>"110010100",
  53362=>"100000001",
  53363=>"101100100",
  53364=>"000011111",
  53365=>"110100111",
  53366=>"001111111",
  53367=>"001110110",
  53368=>"000011111",
  53369=>"101011100",
  53370=>"000100010",
  53371=>"001110100",
  53372=>"011010001",
  53373=>"100011001",
  53374=>"110010001",
  53375=>"000111000",
  53376=>"000000000",
  53377=>"011010011",
  53378=>"010100111",
  53379=>"101010110",
  53380=>"000010000",
  53381=>"000001000",
  53382=>"101001000",
  53383=>"010001111",
  53384=>"010101110",
  53385=>"101001011",
  53386=>"110000100",
  53387=>"101111110",
  53388=>"011000110",
  53389=>"111110101",
  53390=>"110010000",
  53391=>"101110100",
  53392=>"001111011",
  53393=>"101001000",
  53394=>"111100101",
  53395=>"000100110",
  53396=>"001000010",
  53397=>"110001101",
  53398=>"100100111",
  53399=>"000101010",
  53400=>"011011010",
  53401=>"111110001",
  53402=>"000101001",
  53403=>"111000100",
  53404=>"101001001",
  53405=>"000100000",
  53406=>"100000111",
  53407=>"011100111",
  53408=>"000011100",
  53409=>"110100010",
  53410=>"010001011",
  53411=>"101000111",
  53412=>"010001100",
  53413=>"110001100",
  53414=>"011000100",
  53415=>"100001101",
  53416=>"100000011",
  53417=>"000001000",
  53418=>"010111100",
  53419=>"111010111",
  53420=>"000100101",
  53421=>"001111001",
  53422=>"111101110",
  53423=>"100000110",
  53424=>"001110101",
  53425=>"001001101",
  53426=>"011001111",
  53427=>"000110110",
  53428=>"000010110",
  53429=>"000011100",
  53430=>"010001001",
  53431=>"010100000",
  53432=>"010101111",
  53433=>"111001111",
  53434=>"011001011",
  53435=>"101011000",
  53436=>"000110000",
  53437=>"000101100",
  53438=>"110100001",
  53439=>"010110110",
  53440=>"110010010",
  53441=>"010011001",
  53442=>"111010110",
  53443=>"011001111",
  53444=>"101100010",
  53445=>"100011011",
  53446=>"101100111",
  53447=>"000101110",
  53448=>"101010111",
  53449=>"111101001",
  53450=>"000101101",
  53451=>"011011010",
  53452=>"100110101",
  53453=>"000000000",
  53454=>"110000011",
  53455=>"000111100",
  53456=>"100011010",
  53457=>"100100001",
  53458=>"000001101",
  53459=>"010010000",
  53460=>"011001000",
  53461=>"011000100",
  53462=>"010010000",
  53463=>"000100011",
  53464=>"010000100",
  53465=>"011100111",
  53466=>"010001111",
  53467=>"010000010",
  53468=>"101101010",
  53469=>"010010110",
  53470=>"101011110",
  53471=>"001110111",
  53472=>"011001100",
  53473=>"000011001",
  53474=>"100000101",
  53475=>"011101111",
  53476=>"010111111",
  53477=>"111001110",
  53478=>"010010110",
  53479=>"101101111",
  53480=>"011101110",
  53481=>"111110001",
  53482=>"000000111",
  53483=>"101010011",
  53484=>"100011011",
  53485=>"011000010",
  53486=>"111010010",
  53487=>"111010101",
  53488=>"000010000",
  53489=>"110101100",
  53490=>"011001001",
  53491=>"011000000",
  53492=>"110001000",
  53493=>"100101110",
  53494=>"100010010",
  53495=>"000100111",
  53496=>"101001010",
  53497=>"010000100",
  53498=>"000011011",
  53499=>"000000100",
  53500=>"110001010",
  53501=>"000101011",
  53502=>"110101100",
  53503=>"001111111",
  53504=>"100111010",
  53505=>"011111000",
  53506=>"100011111",
  53507=>"111011111",
  53508=>"010010111",
  53509=>"010011111",
  53510=>"111001100",
  53511=>"001100010",
  53512=>"011011000",
  53513=>"101100011",
  53514=>"010110111",
  53515=>"011101101",
  53516=>"011011001",
  53517=>"110001100",
  53518=>"010001011",
  53519=>"010111011",
  53520=>"001111010",
  53521=>"100101110",
  53522=>"101001110",
  53523=>"101010111",
  53524=>"110111101",
  53525=>"111101111",
  53526=>"001010001",
  53527=>"010000101",
  53528=>"011011101",
  53529=>"010001001",
  53530=>"011001000",
  53531=>"001010010",
  53532=>"110100011",
  53533=>"010101101",
  53534=>"110000110",
  53535=>"001101011",
  53536=>"000000001",
  53537=>"111111110",
  53538=>"001000000",
  53539=>"011100100",
  53540=>"000010011",
  53541=>"111100110",
  53542=>"101100110",
  53543=>"111011011",
  53544=>"110011011",
  53545=>"000110011",
  53546=>"000100000",
  53547=>"011110100",
  53548=>"000001010",
  53549=>"010001110",
  53550=>"111111111",
  53551=>"101111111",
  53552=>"011111111",
  53553=>"100110111",
  53554=>"110101001",
  53555=>"010110111",
  53556=>"010000100",
  53557=>"010101001",
  53558=>"110010110",
  53559=>"101000010",
  53560=>"101011011",
  53561=>"111100111",
  53562=>"110101111",
  53563=>"100000100",
  53564=>"001010101",
  53565=>"101000111",
  53566=>"100001001",
  53567=>"101110100",
  53568=>"011001111",
  53569=>"111111110",
  53570=>"100111110",
  53571=>"100100011",
  53572=>"100110001",
  53573=>"000000110",
  53574=>"101001110",
  53575=>"101101111",
  53576=>"101000110",
  53577=>"010000101",
  53578=>"101001000",
  53579=>"001011100",
  53580=>"110011001",
  53581=>"010010111",
  53582=>"101101111",
  53583=>"110111111",
  53584=>"001011101",
  53585=>"000010011",
  53586=>"000010011",
  53587=>"011001100",
  53588=>"101100011",
  53589=>"110001101",
  53590=>"110011111",
  53591=>"110010100",
  53592=>"101110000",
  53593=>"001111100",
  53594=>"000011010",
  53595=>"011111011",
  53596=>"100000000",
  53597=>"100001011",
  53598=>"111000010",
  53599=>"101110101",
  53600=>"001001100",
  53601=>"100000111",
  53602=>"010010010",
  53603=>"010010100",
  53604=>"010001010",
  53605=>"000111011",
  53606=>"100111111",
  53607=>"011101000",
  53608=>"011000000",
  53609=>"010100001",
  53610=>"011100000",
  53611=>"010010001",
  53612=>"110111010",
  53613=>"001000110",
  53614=>"000001111",
  53615=>"101111111",
  53616=>"000100011",
  53617=>"110011000",
  53618=>"100010000",
  53619=>"101011101",
  53620=>"111000100",
  53621=>"100010100",
  53622=>"101001100",
  53623=>"011001010",
  53624=>"110100100",
  53625=>"011010000",
  53626=>"100010111",
  53627=>"100110100",
  53628=>"011000101",
  53629=>"100000001",
  53630=>"101011100",
  53631=>"100011111",
  53632=>"101000111",
  53633=>"101010101",
  53634=>"110111010",
  53635=>"101001010",
  53636=>"001101111",
  53637=>"111001100",
  53638=>"011001010",
  53639=>"111110111",
  53640=>"000010100",
  53641=>"010101110",
  53642=>"001100010",
  53643=>"101001111",
  53644=>"111001000",
  53645=>"011110000",
  53646=>"011110011",
  53647=>"010111110",
  53648=>"101110001",
  53649=>"001011000",
  53650=>"011111000",
  53651=>"000111100",
  53652=>"010110100",
  53653=>"001100001",
  53654=>"000110110",
  53655=>"011110111",
  53656=>"111100010",
  53657=>"001100011",
  53658=>"111110010",
  53659=>"000010000",
  53660=>"001101100",
  53661=>"101100010",
  53662=>"101011011",
  53663=>"101101100",
  53664=>"111110000",
  53665=>"110000001",
  53666=>"011100010",
  53667=>"001000010",
  53668=>"101100010",
  53669=>"011011001",
  53670=>"011110010",
  53671=>"000011110",
  53672=>"011000000",
  53673=>"101100000",
  53674=>"000011101",
  53675=>"100100000",
  53676=>"011010101",
  53677=>"111001110",
  53678=>"010010011",
  53679=>"100001111",
  53680=>"100001000",
  53681=>"000111011",
  53682=>"100011010",
  53683=>"011010001",
  53684=>"110010001",
  53685=>"000111000",
  53686=>"000111010",
  53687=>"010011001",
  53688=>"001100010",
  53689=>"000000110",
  53690=>"111101011",
  53691=>"111110011",
  53692=>"101101100",
  53693=>"001111000",
  53694=>"011111100",
  53695=>"110100010",
  53696=>"010010000",
  53697=>"111010011",
  53698=>"100111110",
  53699=>"011010110",
  53700=>"001000000",
  53701=>"001010000",
  53702=>"001000000",
  53703=>"010100000",
  53704=>"111111001",
  53705=>"110111010",
  53706=>"111010001",
  53707=>"011100000",
  53708=>"011100011",
  53709=>"001101000",
  53710=>"100110100",
  53711=>"000110010",
  53712=>"110101111",
  53713=>"011010110",
  53714=>"101000101",
  53715=>"110100110",
  53716=>"001011010",
  53717=>"111101100",
  53718=>"111000110",
  53719=>"110101100",
  53720=>"110011101",
  53721=>"010101000",
  53722=>"111001000",
  53723=>"001110101",
  53724=>"011001100",
  53725=>"000010010",
  53726=>"001001111",
  53727=>"010101110",
  53728=>"101001011",
  53729=>"110110111",
  53730=>"010010010",
  53731=>"111101111",
  53732=>"010101000",
  53733=>"010001100",
  53734=>"100001100",
  53735=>"100010110",
  53736=>"101110110",
  53737=>"011101100",
  53738=>"000001001",
  53739=>"001111010",
  53740=>"110101011",
  53741=>"010011111",
  53742=>"000001101",
  53743=>"001110001",
  53744=>"010110001",
  53745=>"011001000",
  53746=>"110011000",
  53747=>"111010111",
  53748=>"001000101",
  53749=>"011110111",
  53750=>"100101111",
  53751=>"000100110",
  53752=>"100000110",
  53753=>"100100010",
  53754=>"101000001",
  53755=>"110111101",
  53756=>"000001011",
  53757=>"111010001",
  53758=>"010100111",
  53759=>"111011011",
  53760=>"001001101",
  53761=>"001110001",
  53762=>"000110111",
  53763=>"101111011",
  53764=>"010110011",
  53765=>"100010111",
  53766=>"111001111",
  53767=>"101100111",
  53768=>"000100110",
  53769=>"001100001",
  53770=>"110100111",
  53771=>"100001101",
  53772=>"100101101",
  53773=>"000000101",
  53774=>"000001110",
  53775=>"000101001",
  53776=>"100100101",
  53777=>"011000101",
  53778=>"000101110",
  53779=>"101011100",
  53780=>"100110110",
  53781=>"001111001",
  53782=>"011001011",
  53783=>"000011110",
  53784=>"100011110",
  53785=>"000000110",
  53786=>"111011101",
  53787=>"011110111",
  53788=>"001111110",
  53789=>"001010000",
  53790=>"010100111",
  53791=>"110101110",
  53792=>"001000010",
  53793=>"101001101",
  53794=>"111100001",
  53795=>"110101100",
  53796=>"010000000",
  53797=>"100111011",
  53798=>"111100100",
  53799=>"010101110",
  53800=>"111001011",
  53801=>"000111110",
  53802=>"100010100",
  53803=>"101101101",
  53804=>"101011110",
  53805=>"011010100",
  53806=>"111001001",
  53807=>"111100011",
  53808=>"111010010",
  53809=>"001000100",
  53810=>"101110001",
  53811=>"111111111",
  53812=>"110110001",
  53813=>"001110111",
  53814=>"100001110",
  53815=>"101111111",
  53816=>"001101101",
  53817=>"110101111",
  53818=>"101111101",
  53819=>"101011010",
  53820=>"000100010",
  53821=>"111000100",
  53822=>"111110001",
  53823=>"010011111",
  53824=>"110100110",
  53825=>"010010101",
  53826=>"010111011",
  53827=>"110100001",
  53828=>"010010101",
  53829=>"000100001",
  53830=>"001100000",
  53831=>"001111001",
  53832=>"001001100",
  53833=>"100101011",
  53834=>"001001111",
  53835=>"111001010",
  53836=>"000000000",
  53837=>"110111011",
  53838=>"010110100",
  53839=>"000000010",
  53840=>"010011100",
  53841=>"011111111",
  53842=>"011100111",
  53843=>"010100110",
  53844=>"010110111",
  53845=>"010110101",
  53846=>"110001111",
  53847=>"101011110",
  53848=>"101110110",
  53849=>"101101011",
  53850=>"110101101",
  53851=>"111011001",
  53852=>"010100001",
  53853=>"000000101",
  53854=>"010100011",
  53855=>"011101011",
  53856=>"100011001",
  53857=>"000110101",
  53858=>"110111010",
  53859=>"010010010",
  53860=>"110011100",
  53861=>"011111110",
  53862=>"110110111",
  53863=>"000010001",
  53864=>"001001011",
  53865=>"110000000",
  53866=>"100000100",
  53867=>"010100110",
  53868=>"101000011",
  53869=>"001000010",
  53870=>"001101101",
  53871=>"101001110",
  53872=>"011001011",
  53873=>"101110111",
  53874=>"000000011",
  53875=>"000010110",
  53876=>"100100010",
  53877=>"001100110",
  53878=>"110010101",
  53879=>"011111101",
  53880=>"001100001",
  53881=>"101000010",
  53882=>"000010100",
  53883=>"010001110",
  53884=>"111100000",
  53885=>"111111010",
  53886=>"110110000",
  53887=>"010111111",
  53888=>"110001000",
  53889=>"111110111",
  53890=>"111001111",
  53891=>"111100111",
  53892=>"011000111",
  53893=>"110100110",
  53894=>"100000011",
  53895=>"011100110",
  53896=>"111000111",
  53897=>"101001011",
  53898=>"111101000",
  53899=>"011100100",
  53900=>"000100100",
  53901=>"000101011",
  53902=>"110100100",
  53903=>"101010010",
  53904=>"101000010",
  53905=>"011000000",
  53906=>"101111100",
  53907=>"101001111",
  53908=>"001100011",
  53909=>"001100101",
  53910=>"110101101",
  53911=>"000000111",
  53912=>"111101111",
  53913=>"000001100",
  53914=>"011001000",
  53915=>"011111001",
  53916=>"100110100",
  53917=>"111101101",
  53918=>"010010000",
  53919=>"000010110",
  53920=>"010111110",
  53921=>"000001001",
  53922=>"010010110",
  53923=>"010010101",
  53924=>"110110110",
  53925=>"110101011",
  53926=>"001000000",
  53927=>"111101111",
  53928=>"010000101",
  53929=>"000110011",
  53930=>"100010001",
  53931=>"110000011",
  53932=>"111101111",
  53933=>"000010000",
  53934=>"100110010",
  53935=>"010001100",
  53936=>"001110001",
  53937=>"000000111",
  53938=>"000110111",
  53939=>"101111111",
  53940=>"111100110",
  53941=>"010101100",
  53942=>"011110010",
  53943=>"011111001",
  53944=>"111111010",
  53945=>"100100101",
  53946=>"001011010",
  53947=>"101100110",
  53948=>"101111110",
  53949=>"100111111",
  53950=>"011000000",
  53951=>"101011111",
  53952=>"100000001",
  53953=>"010000101",
  53954=>"111111110",
  53955=>"111011110",
  53956=>"100111011",
  53957=>"000000110",
  53958=>"010001000",
  53959=>"000011010",
  53960=>"111000100",
  53961=>"001000001",
  53962=>"011011111",
  53963=>"010111001",
  53964=>"111111011",
  53965=>"110111000",
  53966=>"110000001",
  53967=>"000001010",
  53968=>"110011110",
  53969=>"010100111",
  53970=>"011100000",
  53971=>"101001011",
  53972=>"000001010",
  53973=>"111011011",
  53974=>"111110001",
  53975=>"000100110",
  53976=>"100111111",
  53977=>"101100100",
  53978=>"110011010",
  53979=>"001101101",
  53980=>"111101000",
  53981=>"000101000",
  53982=>"110101110",
  53983=>"110000111",
  53984=>"011100101",
  53985=>"101111111",
  53986=>"101010001",
  53987=>"010000011",
  53988=>"111111011",
  53989=>"111111001",
  53990=>"011101000",
  53991=>"011101100",
  53992=>"110001101",
  53993=>"101010000",
  53994=>"101110111",
  53995=>"100111100",
  53996=>"100010001",
  53997=>"000101010",
  53998=>"111100110",
  53999=>"001001011",
  54000=>"111000010",
  54001=>"101001111",
  54002=>"001000000",
  54003=>"111100111",
  54004=>"101111101",
  54005=>"010000101",
  54006=>"000001000",
  54007=>"111001101",
  54008=>"011001101",
  54009=>"000101010",
  54010=>"111100000",
  54011=>"011100100",
  54012=>"010010011",
  54013=>"010110011",
  54014=>"101101100",
  54015=>"111000101",
  54016=>"011010100",
  54017=>"000011010",
  54018=>"001001100",
  54019=>"110101001",
  54020=>"110111111",
  54021=>"101001110",
  54022=>"101111011",
  54023=>"011101100",
  54024=>"001010110",
  54025=>"011110110",
  54026=>"011110111",
  54027=>"010000001",
  54028=>"011100101",
  54029=>"111010111",
  54030=>"101110011",
  54031=>"101001011",
  54032=>"110011110",
  54033=>"101100000",
  54034=>"101000010",
  54035=>"111101110",
  54036=>"110001011",
  54037=>"000101001",
  54038=>"010010011",
  54039=>"001100101",
  54040=>"000011011",
  54041=>"100010001",
  54042=>"110011001",
  54043=>"010000001",
  54044=>"000001101",
  54045=>"000111000",
  54046=>"100110111",
  54047=>"001010001",
  54048=>"000101101",
  54049=>"101000111",
  54050=>"111000000",
  54051=>"000001010",
  54052=>"111110010",
  54053=>"001000111",
  54054=>"100110000",
  54055=>"101011100",
  54056=>"101001111",
  54057=>"110101001",
  54058=>"100001101",
  54059=>"000000000",
  54060=>"101110011",
  54061=>"001000011",
  54062=>"100111110",
  54063=>"111011011",
  54064=>"010000001",
  54065=>"101011000",
  54066=>"010110001",
  54067=>"000110101",
  54068=>"000100100",
  54069=>"111000000",
  54070=>"010001110",
  54071=>"010101010",
  54072=>"111111011",
  54073=>"100010111",
  54074=>"010110010",
  54075=>"010000001",
  54076=>"111101111",
  54077=>"000110001",
  54078=>"001111011",
  54079=>"011110001",
  54080=>"000100001",
  54081=>"000011110",
  54082=>"110010001",
  54083=>"010001010",
  54084=>"100101111",
  54085=>"100111101",
  54086=>"110000010",
  54087=>"100110010",
  54088=>"001010000",
  54089=>"001100110",
  54090=>"110110111",
  54091=>"110000000",
  54092=>"011010100",
  54093=>"000101010",
  54094=>"111010101",
  54095=>"000011001",
  54096=>"000101111",
  54097=>"000110100",
  54098=>"010101110",
  54099=>"000010001",
  54100=>"000110010",
  54101=>"101000100",
  54102=>"001000110",
  54103=>"001111000",
  54104=>"111000010",
  54105=>"101011011",
  54106=>"010010010",
  54107=>"101010011",
  54108=>"000101000",
  54109=>"110001111",
  54110=>"010011100",
  54111=>"000111110",
  54112=>"001010110",
  54113=>"000101011",
  54114=>"111010111",
  54115=>"000000111",
  54116=>"001110111",
  54117=>"100010000",
  54118=>"000010011",
  54119=>"101011001",
  54120=>"010010100",
  54121=>"100011010",
  54122=>"000000100",
  54123=>"000010011",
  54124=>"000100100",
  54125=>"110001000",
  54126=>"000011010",
  54127=>"111101110",
  54128=>"110111011",
  54129=>"100100001",
  54130=>"110111000",
  54131=>"011101101",
  54132=>"100111111",
  54133=>"001111010",
  54134=>"000001111",
  54135=>"111010000",
  54136=>"100000000",
  54137=>"001101110",
  54138=>"010000111",
  54139=>"010001000",
  54140=>"010111111",
  54141=>"010101101",
  54142=>"001100000",
  54143=>"111111010",
  54144=>"111101111",
  54145=>"110110011",
  54146=>"010001111",
  54147=>"000110000",
  54148=>"100101111",
  54149=>"001001000",
  54150=>"010000111",
  54151=>"100001011",
  54152=>"011011110",
  54153=>"001111110",
  54154=>"100111111",
  54155=>"101000000",
  54156=>"100101001",
  54157=>"110011011",
  54158=>"111111101",
  54159=>"110001011",
  54160=>"100111011",
  54161=>"100001100",
  54162=>"000010111",
  54163=>"000010000",
  54164=>"110010101",
  54165=>"100111110",
  54166=>"101010111",
  54167=>"110011001",
  54168=>"111001100",
  54169=>"000101111",
  54170=>"110011101",
  54171=>"001101110",
  54172=>"011111101",
  54173=>"000110101",
  54174=>"110100101",
  54175=>"010101011",
  54176=>"100100110",
  54177=>"110010100",
  54178=>"011101000",
  54179=>"100001111",
  54180=>"111100010",
  54181=>"011110101",
  54182=>"101100010",
  54183=>"100111010",
  54184=>"011000110",
  54185=>"011100101",
  54186=>"100011111",
  54187=>"000010000",
  54188=>"110001010",
  54189=>"000011111",
  54190=>"010111000",
  54191=>"011001011",
  54192=>"011100100",
  54193=>"011000010",
  54194=>"110001110",
  54195=>"100010000",
  54196=>"111101101",
  54197=>"001001001",
  54198=>"000110000",
  54199=>"010100001",
  54200=>"011100000",
  54201=>"111100001",
  54202=>"100011000",
  54203=>"110000000",
  54204=>"110010000",
  54205=>"001100001",
  54206=>"111110111",
  54207=>"000001101",
  54208=>"101010111",
  54209=>"010001000",
  54210=>"101101111",
  54211=>"000001010",
  54212=>"011001110",
  54213=>"010100001",
  54214=>"001111011",
  54215=>"111001000",
  54216=>"110100000",
  54217=>"101011100",
  54218=>"111100010",
  54219=>"111001101",
  54220=>"101010101",
  54221=>"110000001",
  54222=>"101000101",
  54223=>"001010101",
  54224=>"010001011",
  54225=>"101101000",
  54226=>"111001001",
  54227=>"001010011",
  54228=>"011111001",
  54229=>"010000111",
  54230=>"001010101",
  54231=>"001101100",
  54232=>"110111100",
  54233=>"110000111",
  54234=>"110010111",
  54235=>"001010100",
  54236=>"110110010",
  54237=>"010011111",
  54238=>"110100111",
  54239=>"100010011",
  54240=>"010101001",
  54241=>"101011111",
  54242=>"111111111",
  54243=>"010100011",
  54244=>"010110111",
  54245=>"100010101",
  54246=>"101100000",
  54247=>"000100101",
  54248=>"011110111",
  54249=>"110111011",
  54250=>"101011000",
  54251=>"011000000",
  54252=>"000011001",
  54253=>"110101000",
  54254=>"010100011",
  54255=>"110000000",
  54256=>"011010011",
  54257=>"101101000",
  54258=>"001001001",
  54259=>"110111010",
  54260=>"001010011",
  54261=>"110101100",
  54262=>"110100110",
  54263=>"001000011",
  54264=>"111100000",
  54265=>"001010101",
  54266=>"101101111",
  54267=>"110101000",
  54268=>"000111011",
  54269=>"100010011",
  54270=>"100010000",
  54271=>"011011011",
  54272=>"100100101",
  54273=>"011100110",
  54274=>"011110000",
  54275=>"001100100",
  54276=>"011110101",
  54277=>"001100001",
  54278=>"100101010",
  54279=>"110101011",
  54280=>"100010101",
  54281=>"001010001",
  54282=>"010000010",
  54283=>"001101101",
  54284=>"000000000",
  54285=>"010111101",
  54286=>"101000100",
  54287=>"111000101",
  54288=>"000110111",
  54289=>"111110011",
  54290=>"010100010",
  54291=>"001110001",
  54292=>"011000111",
  54293=>"001110011",
  54294=>"100111101",
  54295=>"100100100",
  54296=>"000010101",
  54297=>"101011110",
  54298=>"110001011",
  54299=>"110010001",
  54300=>"111010001",
  54301=>"111101010",
  54302=>"101110100",
  54303=>"111101110",
  54304=>"111011010",
  54305=>"110101100",
  54306=>"010110110",
  54307=>"011011000",
  54308=>"001000000",
  54309=>"000100001",
  54310=>"010110101",
  54311=>"000010001",
  54312=>"011011000",
  54313=>"110110100",
  54314=>"110111101",
  54315=>"000110101",
  54316=>"111111001",
  54317=>"010111111",
  54318=>"101110111",
  54319=>"101111010",
  54320=>"010101011",
  54321=>"110101010",
  54322=>"011010010",
  54323=>"111111010",
  54324=>"011100001",
  54325=>"111100101",
  54326=>"000001101",
  54327=>"100100001",
  54328=>"000010111",
  54329=>"001010110",
  54330=>"110011101",
  54331=>"111101110",
  54332=>"110011000",
  54333=>"100010101",
  54334=>"010011010",
  54335=>"111000010",
  54336=>"101011111",
  54337=>"001100110",
  54338=>"001101100",
  54339=>"001101111",
  54340=>"100001101",
  54341=>"011011001",
  54342=>"001011110",
  54343=>"111001101",
  54344=>"100000111",
  54345=>"000000011",
  54346=>"000011001",
  54347=>"010000011",
  54348=>"000110110",
  54349=>"111000100",
  54350=>"000010010",
  54351=>"010000110",
  54352=>"110010000",
  54353=>"010111010",
  54354=>"000100110",
  54355=>"010001101",
  54356=>"101100110",
  54357=>"000110011",
  54358=>"011100111",
  54359=>"101110000",
  54360=>"110011111",
  54361=>"000100010",
  54362=>"011101111",
  54363=>"100001011",
  54364=>"101001000",
  54365=>"000010111",
  54366=>"100100001",
  54367=>"011100000",
  54368=>"000100111",
  54369=>"000001110",
  54370=>"111100011",
  54371=>"011100010",
  54372=>"111010100",
  54373=>"010110000",
  54374=>"000011011",
  54375=>"001110110",
  54376=>"110001010",
  54377=>"011100100",
  54378=>"010000010",
  54379=>"011000011",
  54380=>"000010001",
  54381=>"010110110",
  54382=>"010001000",
  54383=>"111010101",
  54384=>"001001000",
  54385=>"010110110",
  54386=>"101111110",
  54387=>"111111011",
  54388=>"001011100",
  54389=>"110111000",
  54390=>"100101000",
  54391=>"011111100",
  54392=>"010110011",
  54393=>"100000100",
  54394=>"001010010",
  54395=>"101110001",
  54396=>"110110101",
  54397=>"001100111",
  54398=>"000001011",
  54399=>"011011000",
  54400=>"110101000",
  54401=>"010110001",
  54402=>"110000011",
  54403=>"101001000",
  54404=>"110111011",
  54405=>"010011100",
  54406=>"101101001",
  54407=>"000010001",
  54408=>"001111000",
  54409=>"011010000",
  54410=>"110101011",
  54411=>"101000110",
  54412=>"001100110",
  54413=>"100100100",
  54414=>"011101110",
  54415=>"000110000",
  54416=>"111100111",
  54417=>"011111111",
  54418=>"111110111",
  54419=>"111111100",
  54420=>"111001110",
  54421=>"110101111",
  54422=>"110000001",
  54423=>"011000011",
  54424=>"111001011",
  54425=>"101100011",
  54426=>"011101100",
  54427=>"000001001",
  54428=>"101100011",
  54429=>"010100110",
  54430=>"101001011",
  54431=>"110100010",
  54432=>"110000100",
  54433=>"011110011",
  54434=>"010100111",
  54435=>"001111101",
  54436=>"111111100",
  54437=>"111100001",
  54438=>"111110001",
  54439=>"110010010",
  54440=>"100101000",
  54441=>"011100101",
  54442=>"100101101",
  54443=>"100101010",
  54444=>"010111011",
  54445=>"101111011",
  54446=>"000000000",
  54447=>"011000111",
  54448=>"110000010",
  54449=>"001100011",
  54450=>"111000100",
  54451=>"000010011",
  54452=>"101111111",
  54453=>"110111010",
  54454=>"110011010",
  54455=>"100101010",
  54456=>"001000011",
  54457=>"010010000",
  54458=>"110011101",
  54459=>"001110111",
  54460=>"111110000",
  54461=>"100001000",
  54462=>"010101010",
  54463=>"100011111",
  54464=>"010000111",
  54465=>"010010010",
  54466=>"101010011",
  54467=>"011100101",
  54468=>"010000011",
  54469=>"000000100",
  54470=>"110101101",
  54471=>"010100010",
  54472=>"001000110",
  54473=>"111101111",
  54474=>"111111010",
  54475=>"011011010",
  54476=>"110101011",
  54477=>"111101001",
  54478=>"000001011",
  54479=>"101010000",
  54480=>"000101111",
  54481=>"000100111",
  54482=>"110010010",
  54483=>"101001101",
  54484=>"011001010",
  54485=>"001101010",
  54486=>"100101101",
  54487=>"110111010",
  54488=>"011100101",
  54489=>"000101001",
  54490=>"110101101",
  54491=>"100110101",
  54492=>"111100001",
  54493=>"111111101",
  54494=>"001100000",
  54495=>"110000001",
  54496=>"000011101",
  54497=>"010101100",
  54498=>"001011111",
  54499=>"001100100",
  54500=>"000000111",
  54501=>"011010100",
  54502=>"111010111",
  54503=>"011000010",
  54504=>"110011011",
  54505=>"001001000",
  54506=>"000100111",
  54507=>"100110001",
  54508=>"100011000",
  54509=>"111000110",
  54510=>"010110011",
  54511=>"010010100",
  54512=>"100101111",
  54513=>"101001000",
  54514=>"100101110",
  54515=>"000011000",
  54516=>"000011110",
  54517=>"101101110",
  54518=>"110010010",
  54519=>"001101111",
  54520=>"000010110",
  54521=>"110001001",
  54522=>"101100001",
  54523=>"010111101",
  54524=>"000110001",
  54525=>"010110101",
  54526=>"111010010",
  54527=>"111111111",
  54528=>"111110111",
  54529=>"100001011",
  54530=>"010011101",
  54531=>"000101001",
  54532=>"101110100",
  54533=>"100110011",
  54534=>"010010110",
  54535=>"100010110",
  54536=>"011111101",
  54537=>"111110000",
  54538=>"111111011",
  54539=>"010110001",
  54540=>"101001100",
  54541=>"100100101",
  54542=>"010000111",
  54543=>"000000011",
  54544=>"111010111",
  54545=>"001110010",
  54546=>"010101111",
  54547=>"110011010",
  54548=>"001000001",
  54549=>"101010011",
  54550=>"001011110",
  54551=>"010001010",
  54552=>"101010011",
  54553=>"010111101",
  54554=>"100010010",
  54555=>"100000011",
  54556=>"111100000",
  54557=>"010110010",
  54558=>"010110101",
  54559=>"100011110",
  54560=>"000001100",
  54561=>"100110100",
  54562=>"010101011",
  54563=>"110011001",
  54564=>"010000110",
  54565=>"010010111",
  54566=>"010010011",
  54567=>"010011000",
  54568=>"101101011",
  54569=>"000010011",
  54570=>"101101100",
  54571=>"111101101",
  54572=>"100010110",
  54573=>"000001100",
  54574=>"000000000",
  54575=>"001111111",
  54576=>"100111000",
  54577=>"110101010",
  54578=>"111010101",
  54579=>"001001001",
  54580=>"011000101",
  54581=>"010110001",
  54582=>"000100001",
  54583=>"000110010",
  54584=>"101001111",
  54585=>"111111110",
  54586=>"101101100",
  54587=>"111000000",
  54588=>"000100010",
  54589=>"110100011",
  54590=>"011010001",
  54591=>"010101000",
  54592=>"001000010",
  54593=>"111110000",
  54594=>"111010101",
  54595=>"111100110",
  54596=>"100000111",
  54597=>"000011110",
  54598=>"001100101",
  54599=>"110010010",
  54600=>"010110110",
  54601=>"111010010",
  54602=>"100000011",
  54603=>"100001001",
  54604=>"100111110",
  54605=>"111001010",
  54606=>"100001100",
  54607=>"111011000",
  54608=>"100010111",
  54609=>"110101011",
  54610=>"010101001",
  54611=>"111010011",
  54612=>"001000101",
  54613=>"010001011",
  54614=>"000100101",
  54615=>"110111101",
  54616=>"011011011",
  54617=>"001011111",
  54618=>"100001100",
  54619=>"001001000",
  54620=>"100100010",
  54621=>"000001010",
  54622=>"100010101",
  54623=>"000100101",
  54624=>"110111001",
  54625=>"000011101",
  54626=>"111000111",
  54627=>"000101001",
  54628=>"111111101",
  54629=>"111000111",
  54630=>"010011011",
  54631=>"110011001",
  54632=>"101111111",
  54633=>"011100000",
  54634=>"001001010",
  54635=>"101110111",
  54636=>"001001001",
  54637=>"010000000",
  54638=>"011111011",
  54639=>"011001000",
  54640=>"100010101",
  54641=>"010001011",
  54642=>"001010111",
  54643=>"111010100",
  54644=>"001001001",
  54645=>"011101000",
  54646=>"101011010",
  54647=>"011101110",
  54648=>"010001111",
  54649=>"100100000",
  54650=>"110011100",
  54651=>"111111011",
  54652=>"111101111",
  54653=>"000110101",
  54654=>"110110100",
  54655=>"000001110",
  54656=>"000010010",
  54657=>"100000101",
  54658=>"111000100",
  54659=>"110110111",
  54660=>"001000111",
  54661=>"111111100",
  54662=>"111000001",
  54663=>"001110011",
  54664=>"100000011",
  54665=>"010011100",
  54666=>"100111010",
  54667=>"110100001",
  54668=>"000101111",
  54669=>"101000110",
  54670=>"100011001",
  54671=>"001100001",
  54672=>"000110000",
  54673=>"011000011",
  54674=>"110110101",
  54675=>"001111101",
  54676=>"011101011",
  54677=>"110000111",
  54678=>"011010001",
  54679=>"100100100",
  54680=>"011101011",
  54681=>"000010001",
  54682=>"000000011",
  54683=>"000111010",
  54684=>"001011111",
  54685=>"101111111",
  54686=>"011100000",
  54687=>"010000101",
  54688=>"101000011",
  54689=>"011000100",
  54690=>"010011001",
  54691=>"101111101",
  54692=>"111010111",
  54693=>"110010001",
  54694=>"010110110",
  54695=>"000001000",
  54696=>"000000100",
  54697=>"111100110",
  54698=>"101110111",
  54699=>"000111000",
  54700=>"110110000",
  54701=>"110011110",
  54702=>"001000100",
  54703=>"001110000",
  54704=>"111110111",
  54705=>"101001010",
  54706=>"000110001",
  54707=>"110110011",
  54708=>"001000101",
  54709=>"100111001",
  54710=>"010001101",
  54711=>"100000001",
  54712=>"001001100",
  54713=>"001100111",
  54714=>"101000000",
  54715=>"111001000",
  54716=>"011101001",
  54717=>"100011011",
  54718=>"001100110",
  54719=>"011101010",
  54720=>"000110001",
  54721=>"111101011",
  54722=>"111110100",
  54723=>"001010001",
  54724=>"101110011",
  54725=>"110101010",
  54726=>"010111100",
  54727=>"110100010",
  54728=>"001011010",
  54729=>"110001111",
  54730=>"101101011",
  54731=>"010000100",
  54732=>"111111111",
  54733=>"000011010",
  54734=>"111001110",
  54735=>"001000001",
  54736=>"111000111",
  54737=>"110111110",
  54738=>"100101011",
  54739=>"110101010",
  54740=>"011101011",
  54741=>"011000101",
  54742=>"101110101",
  54743=>"111010010",
  54744=>"101000010",
  54745=>"110001101",
  54746=>"001000101",
  54747=>"101011100",
  54748=>"111000110",
  54749=>"111111011",
  54750=>"010011110",
  54751=>"111101100",
  54752=>"001010100",
  54753=>"100111110",
  54754=>"010011011",
  54755=>"010011100",
  54756=>"000111100",
  54757=>"100101110",
  54758=>"000000100",
  54759=>"000010100",
  54760=>"111011110",
  54761=>"010110001",
  54762=>"100111001",
  54763=>"101110100",
  54764=>"001110110",
  54765=>"011111101",
  54766=>"111101101",
  54767=>"001001001",
  54768=>"010000111",
  54769=>"111000101",
  54770=>"000110011",
  54771=>"111101011",
  54772=>"101110010",
  54773=>"011111001",
  54774=>"001101011",
  54775=>"000110110",
  54776=>"001110111",
  54777=>"101110101",
  54778=>"011111010",
  54779=>"011001010",
  54780=>"001101110",
  54781=>"100010110",
  54782=>"011011100",
  54783=>"100010000",
  54784=>"110101010",
  54785=>"100101111",
  54786=>"100101100",
  54787=>"010000101",
  54788=>"111011000",
  54789=>"000001110",
  54790=>"110010001",
  54791=>"101110011",
  54792=>"110101000",
  54793=>"010111011",
  54794=>"000010101",
  54795=>"000101001",
  54796=>"010001011",
  54797=>"100110101",
  54798=>"100000101",
  54799=>"110110110",
  54800=>"010111110",
  54801=>"011011000",
  54802=>"110101110",
  54803=>"100010111",
  54804=>"011010110",
  54805=>"101110110",
  54806=>"110011010",
  54807=>"000001110",
  54808=>"010000110",
  54809=>"111001010",
  54810=>"110110001",
  54811=>"011000101",
  54812=>"000010001",
  54813=>"100001011",
  54814=>"101000011",
  54815=>"110010100",
  54816=>"110011010",
  54817=>"011100010",
  54818=>"110111111",
  54819=>"101100001",
  54820=>"110001011",
  54821=>"001010111",
  54822=>"001110110",
  54823=>"111001100",
  54824=>"101111000",
  54825=>"110101011",
  54826=>"000111000",
  54827=>"101100010",
  54828=>"010111111",
  54829=>"001111011",
  54830=>"011101111",
  54831=>"110110000",
  54832=>"000100101",
  54833=>"110010000",
  54834=>"111111010",
  54835=>"101101100",
  54836=>"111000001",
  54837=>"001010110",
  54838=>"011111010",
  54839=>"100000111",
  54840=>"111111001",
  54841=>"110000110",
  54842=>"000111110",
  54843=>"010100010",
  54844=>"000110010",
  54845=>"000000010",
  54846=>"010011110",
  54847=>"110100100",
  54848=>"100001011",
  54849=>"010100101",
  54850=>"100111101",
  54851=>"001000000",
  54852=>"010100110",
  54853=>"111111101",
  54854=>"011001000",
  54855=>"110011010",
  54856=>"000011110",
  54857=>"110000110",
  54858=>"101100000",
  54859=>"001010001",
  54860=>"000010111",
  54861=>"111110010",
  54862=>"101100111",
  54863=>"101100101",
  54864=>"011101001",
  54865=>"111101000",
  54866=>"110100011",
  54867=>"001011001",
  54868=>"110100011",
  54869=>"001000011",
  54870=>"100111110",
  54871=>"101010110",
  54872=>"010110101",
  54873=>"001100011",
  54874=>"101010111",
  54875=>"100010011",
  54876=>"110110010",
  54877=>"000010001",
  54878=>"011011110",
  54879=>"111100100",
  54880=>"010110100",
  54881=>"000011000",
  54882=>"010111110",
  54883=>"011100110",
  54884=>"110011001",
  54885=>"001100100",
  54886=>"111101001",
  54887=>"101100000",
  54888=>"100110101",
  54889=>"100000000",
  54890=>"111001011",
  54891=>"010010101",
  54892=>"010011011",
  54893=>"011011001",
  54894=>"000110100",
  54895=>"011000100",
  54896=>"111011001",
  54897=>"100001000",
  54898=>"101011111",
  54899=>"011000001",
  54900=>"001000011",
  54901=>"101011001",
  54902=>"010000110",
  54903=>"010111100",
  54904=>"101000001",
  54905=>"011111011",
  54906=>"111111001",
  54907=>"001010001",
  54908=>"000001111",
  54909=>"100001001",
  54910=>"001101011",
  54911=>"111000100",
  54912=>"100010101",
  54913=>"000010011",
  54914=>"101101101",
  54915=>"111011000",
  54916=>"111011011",
  54917=>"111111101",
  54918=>"010100001",
  54919=>"011101000",
  54920=>"111011111",
  54921=>"100001100",
  54922=>"100010000",
  54923=>"111101101",
  54924=>"000100000",
  54925=>"111001100",
  54926=>"111100111",
  54927=>"111010111",
  54928=>"001110000",
  54929=>"101110110",
  54930=>"000101100",
  54931=>"101111010",
  54932=>"101011011",
  54933=>"001000101",
  54934=>"010110101",
  54935=>"011101010",
  54936=>"011010101",
  54937=>"000110111",
  54938=>"011100011",
  54939=>"110001001",
  54940=>"010110111",
  54941=>"101001001",
  54942=>"110110010",
  54943=>"000110000",
  54944=>"001110101",
  54945=>"011011110",
  54946=>"010110100",
  54947=>"111011100",
  54948=>"001101000",
  54949=>"011100110",
  54950=>"110001111",
  54951=>"010110000",
  54952=>"000101111",
  54953=>"001000101",
  54954=>"101000110",
  54955=>"101011001",
  54956=>"010001100",
  54957=>"011111111",
  54958=>"101111010",
  54959=>"011111111",
  54960=>"000110101",
  54961=>"000010110",
  54962=>"101000101",
  54963=>"101011010",
  54964=>"111001111",
  54965=>"100101111",
  54966=>"011010101",
  54967=>"011101011",
  54968=>"000100001",
  54969=>"000100100",
  54970=>"001111100",
  54971=>"011101100",
  54972=>"010100101",
  54973=>"001101100",
  54974=>"111000010",
  54975=>"101011010",
  54976=>"011101100",
  54977=>"111001110",
  54978=>"000101001",
  54979=>"010100111",
  54980=>"010010110",
  54981=>"101010111",
  54982=>"010101001",
  54983=>"001110000",
  54984=>"011110010",
  54985=>"101011010",
  54986=>"100111000",
  54987=>"111000110",
  54988=>"001110100",
  54989=>"110100111",
  54990=>"100001101",
  54991=>"001010100",
  54992=>"110100111",
  54993=>"111010000",
  54994=>"011011110",
  54995=>"111001011",
  54996=>"100100110",
  54997=>"101110010",
  54998=>"011111010",
  54999=>"111011011",
  55000=>"101111111",
  55001=>"000010001",
  55002=>"011001000",
  55003=>"101000010",
  55004=>"000110000",
  55005=>"010111011",
  55006=>"101110101",
  55007=>"100001011",
  55008=>"011111110",
  55009=>"110010011",
  55010=>"101000100",
  55011=>"100111111",
  55012=>"001000110",
  55013=>"111111101",
  55014=>"100010000",
  55015=>"011110100",
  55016=>"011011011",
  55017=>"111001001",
  55018=>"101001000",
  55019=>"001101111",
  55020=>"000110001",
  55021=>"110111000",
  55022=>"000110001",
  55023=>"011001111",
  55024=>"011011010",
  55025=>"100101000",
  55026=>"111111011",
  55027=>"111011010",
  55028=>"101001010",
  55029=>"100001100",
  55030=>"010101011",
  55031=>"110011011",
  55032=>"101010000",
  55033=>"011000101",
  55034=>"111101000",
  55035=>"000000110",
  55036=>"110101111",
  55037=>"010000101",
  55038=>"111110111",
  55039=>"110000000",
  55040=>"101101101",
  55041=>"111010000",
  55042=>"111110011",
  55043=>"010110011",
  55044=>"110001000",
  55045=>"100111110",
  55046=>"011110000",
  55047=>"001000000",
  55048=>"110101101",
  55049=>"110101000",
  55050=>"101110010",
  55051=>"111101101",
  55052=>"000110100",
  55053=>"110001010",
  55054=>"100010111",
  55055=>"101110110",
  55056=>"100000100",
  55057=>"110000101",
  55058=>"101011000",
  55059=>"100101001",
  55060=>"000011101",
  55061=>"110100010",
  55062=>"011101011",
  55063=>"100100110",
  55064=>"101100001",
  55065=>"000101100",
  55066=>"000000101",
  55067=>"001110111",
  55068=>"111000101",
  55069=>"110101100",
  55070=>"000100010",
  55071=>"011110001",
  55072=>"101111111",
  55073=>"110110010",
  55074=>"110110011",
  55075=>"111011111",
  55076=>"011010000",
  55077=>"010000101",
  55078=>"000100101",
  55079=>"101101010",
  55080=>"110100010",
  55081=>"010111010",
  55082=>"111111000",
  55083=>"011011101",
  55084=>"001100000",
  55085=>"000000101",
  55086=>"010110001",
  55087=>"111110111",
  55088=>"111010110",
  55089=>"101110000",
  55090=>"100100110",
  55091=>"100000111",
  55092=>"000001000",
  55093=>"111101011",
  55094=>"011010110",
  55095=>"100000101",
  55096=>"110001101",
  55097=>"001000011",
  55098=>"000001010",
  55099=>"010101100",
  55100=>"000000111",
  55101=>"110100101",
  55102=>"000101101",
  55103=>"110000011",
  55104=>"101100111",
  55105=>"010000000",
  55106=>"110010111",
  55107=>"101100000",
  55108=>"110100111",
  55109=>"111001111",
  55110=>"000101100",
  55111=>"000100001",
  55112=>"010011100",
  55113=>"001100000",
  55114=>"011100001",
  55115=>"000001101",
  55116=>"011001100",
  55117=>"010100111",
  55118=>"100111111",
  55119=>"101101011",
  55120=>"100101111",
  55121=>"101001010",
  55122=>"010110011",
  55123=>"010011111",
  55124=>"010100110",
  55125=>"111111010",
  55126=>"001011100",
  55127=>"010110111",
  55128=>"110100110",
  55129=>"111100100",
  55130=>"100001001",
  55131=>"011000000",
  55132=>"000001000",
  55133=>"011011110",
  55134=>"110101001",
  55135=>"010101001",
  55136=>"010101000",
  55137=>"101111101",
  55138=>"100010000",
  55139=>"110100100",
  55140=>"111001011",
  55141=>"111000001",
  55142=>"110111100",
  55143=>"010101010",
  55144=>"011111010",
  55145=>"101111010",
  55146=>"001000111",
  55147=>"100111000",
  55148=>"110110000",
  55149=>"110000101",
  55150=>"001111110",
  55151=>"010100101",
  55152=>"011011011",
  55153=>"111000010",
  55154=>"110101110",
  55155=>"111110100",
  55156=>"010000110",
  55157=>"110101100",
  55158=>"100101001",
  55159=>"110001010",
  55160=>"110110011",
  55161=>"011010010",
  55162=>"010110010",
  55163=>"100011010",
  55164=>"000101111",
  55165=>"100010010",
  55166=>"110111111",
  55167=>"111001001",
  55168=>"010011110",
  55169=>"101011000",
  55170=>"111110110",
  55171=>"101011010",
  55172=>"110010000",
  55173=>"111111001",
  55174=>"100000111",
  55175=>"110000011",
  55176=>"110101000",
  55177=>"111000001",
  55178=>"111110011",
  55179=>"100010100",
  55180=>"000001010",
  55181=>"000010000",
  55182=>"110110111",
  55183=>"110101010",
  55184=>"110111100",
  55185=>"100000010",
  55186=>"000110111",
  55187=>"100101100",
  55188=>"101001100",
  55189=>"101100000",
  55190=>"001100100",
  55191=>"110010110",
  55192=>"000000001",
  55193=>"100110001",
  55194=>"101111100",
  55195=>"010001110",
  55196=>"010110111",
  55197=>"100010111",
  55198=>"110111011",
  55199=>"111100011",
  55200=>"000011000",
  55201=>"001010001",
  55202=>"101101010",
  55203=>"001010110",
  55204=>"101101110",
  55205=>"010010111",
  55206=>"110101100",
  55207=>"000010111",
  55208=>"010111011",
  55209=>"010100100",
  55210=>"101010011",
  55211=>"110001011",
  55212=>"010000011",
  55213=>"010111011",
  55214=>"101011101",
  55215=>"010000100",
  55216=>"010000001",
  55217=>"110101100",
  55218=>"011101001",
  55219=>"100100100",
  55220=>"010111010",
  55221=>"110110011",
  55222=>"000111111",
  55223=>"000000101",
  55224=>"111110000",
  55225=>"011010111",
  55226=>"010001010",
  55227=>"111101001",
  55228=>"100111101",
  55229=>"010110000",
  55230=>"000001000",
  55231=>"000101001",
  55232=>"111110010",
  55233=>"000100010",
  55234=>"001000100",
  55235=>"000000100",
  55236=>"111101000",
  55237=>"011111000",
  55238=>"010101111",
  55239=>"001001010",
  55240=>"001010111",
  55241=>"100111000",
  55242=>"101000010",
  55243=>"010011100",
  55244=>"000010011",
  55245=>"000111001",
  55246=>"110010000",
  55247=>"010010100",
  55248=>"100100011",
  55249=>"110110010",
  55250=>"000000100",
  55251=>"100000011",
  55252=>"000010100",
  55253=>"101011111",
  55254=>"001001111",
  55255=>"101011110",
  55256=>"001001100",
  55257=>"100101010",
  55258=>"110110111",
  55259=>"010110011",
  55260=>"010000110",
  55261=>"001001011",
  55262=>"100011011",
  55263=>"111110101",
  55264=>"010011100",
  55265=>"110001100",
  55266=>"111000100",
  55267=>"001101001",
  55268=>"101111100",
  55269=>"000010101",
  55270=>"001101111",
  55271=>"000100110",
  55272=>"101101000",
  55273=>"010100101",
  55274=>"101000100",
  55275=>"011000000",
  55276=>"100010111",
  55277=>"110100010",
  55278=>"000010000",
  55279=>"000001010",
  55280=>"110001010",
  55281=>"110001100",
  55282=>"010011000",
  55283=>"000111000",
  55284=>"011001001",
  55285=>"110011101",
  55286=>"101110100",
  55287=>"110111011",
  55288=>"000001001",
  55289=>"101011010",
  55290=>"010010101",
  55291=>"011000000",
  55292=>"011000000",
  55293=>"000010001",
  55294=>"011101101",
  55295=>"111011111",
  55296=>"010001011",
  55297=>"001001001",
  55298=>"110001110",
  55299=>"111010111",
  55300=>"011111111",
  55301=>"110011000",
  55302=>"010011110",
  55303=>"001011010",
  55304=>"011001110",
  55305=>"010101101",
  55306=>"101010001",
  55307=>"100010000",
  55308=>"010100000",
  55309=>"000010100",
  55310=>"001111001",
  55311=>"000110110",
  55312=>"110001101",
  55313=>"111000000",
  55314=>"000100011",
  55315=>"010110010",
  55316=>"000100000",
  55317=>"101101100",
  55318=>"001111100",
  55319=>"100001100",
  55320=>"100011111",
  55321=>"011010010",
  55322=>"000101110",
  55323=>"111101001",
  55324=>"011100111",
  55325=>"101001111",
  55326=>"011000000",
  55327=>"010110110",
  55328=>"100110010",
  55329=>"001110001",
  55330=>"101100100",
  55331=>"111011000",
  55332=>"111011111",
  55333=>"001111000",
  55334=>"101111100",
  55335=>"001110000",
  55336=>"000101001",
  55337=>"011000000",
  55338=>"010101110",
  55339=>"000101001",
  55340=>"101000101",
  55341=>"100011011",
  55342=>"111001000",
  55343=>"000101110",
  55344=>"001001001",
  55345=>"011000101",
  55346=>"111010110",
  55347=>"111110010",
  55348=>"001000101",
  55349=>"000111100",
  55350=>"010111111",
  55351=>"111011101",
  55352=>"001100101",
  55353=>"101001110",
  55354=>"111111011",
  55355=>"001111110",
  55356=>"110110110",
  55357=>"011101110",
  55358=>"000101000",
  55359=>"000001001",
  55360=>"000010011",
  55361=>"100001000",
  55362=>"011111110",
  55363=>"101011100",
  55364=>"101001000",
  55365=>"000001110",
  55366=>"110001111",
  55367=>"011001001",
  55368=>"000000111",
  55369=>"111111010",
  55370=>"100011101",
  55371=>"110111101",
  55372=>"011111010",
  55373=>"110001011",
  55374=>"100100011",
  55375=>"101101001",
  55376=>"100001010",
  55377=>"111000110",
  55378=>"111100101",
  55379=>"000001111",
  55380=>"011001010",
  55381=>"101101111",
  55382=>"010001000",
  55383=>"011011011",
  55384=>"111000000",
  55385=>"000101110",
  55386=>"010000011",
  55387=>"100100111",
  55388=>"100000000",
  55389=>"000000011",
  55390=>"000000110",
  55391=>"010000011",
  55392=>"101000101",
  55393=>"001111101",
  55394=>"111101001",
  55395=>"100010100",
  55396=>"010100011",
  55397=>"001011110",
  55398=>"001010100",
  55399=>"000000011",
  55400=>"001000010",
  55401=>"000110111",
  55402=>"100010100",
  55403=>"100001001",
  55404=>"010000110",
  55405=>"000101111",
  55406=>"001100000",
  55407=>"101011001",
  55408=>"011110111",
  55409=>"101111100",
  55410=>"100001011",
  55411=>"111101000",
  55412=>"101100011",
  55413=>"001010101",
  55414=>"100110011",
  55415=>"110010111",
  55416=>"100110110",
  55417=>"110000111",
  55418=>"110000010",
  55419=>"111011000",
  55420=>"010101110",
  55421=>"101100011",
  55422=>"000010001",
  55423=>"100001000",
  55424=>"010110011",
  55425=>"110100000",
  55426=>"000000010",
  55427=>"001110100",
  55428=>"010111100",
  55429=>"001010101",
  55430=>"110011110",
  55431=>"001000001",
  55432=>"101000011",
  55433=>"001101011",
  55434=>"100000111",
  55435=>"100010100",
  55436=>"001111111",
  55437=>"001100000",
  55438=>"110110100",
  55439=>"110010011",
  55440=>"010110111",
  55441=>"100010111",
  55442=>"001001001",
  55443=>"111100110",
  55444=>"010110110",
  55445=>"011110100",
  55446=>"001000110",
  55447=>"000001100",
  55448=>"000000100",
  55449=>"000111010",
  55450=>"110001100",
  55451=>"111011110",
  55452=>"111011000",
  55453=>"010010100",
  55454=>"011111010",
  55455=>"010110011",
  55456=>"000101001",
  55457=>"010100100",
  55458=>"110110011",
  55459=>"001101000",
  55460=>"000110011",
  55461=>"100001111",
  55462=>"110010110",
  55463=>"001100010",
  55464=>"100001001",
  55465=>"001111101",
  55466=>"100011001",
  55467=>"111110110",
  55468=>"101111101",
  55469=>"011111100",
  55470=>"111001010",
  55471=>"010010100",
  55472=>"110001100",
  55473=>"111101111",
  55474=>"000111100",
  55475=>"001011000",
  55476=>"110011100",
  55477=>"011100111",
  55478=>"101010001",
  55479=>"011001000",
  55480=>"001010000",
  55481=>"000001011",
  55482=>"011000101",
  55483=>"111000101",
  55484=>"011111111",
  55485=>"101000000",
  55486=>"101110011",
  55487=>"011100110",
  55488=>"110000100",
  55489=>"111001011",
  55490=>"001000111",
  55491=>"100110100",
  55492=>"111010001",
  55493=>"000010011",
  55494=>"111111101",
  55495=>"111011100",
  55496=>"000001010",
  55497=>"001100010",
  55498=>"010110110",
  55499=>"010100000",
  55500=>"100011010",
  55501=>"100100101",
  55502=>"011001110",
  55503=>"111110111",
  55504=>"001101000",
  55505=>"001000010",
  55506=>"100001010",
  55507=>"110100011",
  55508=>"110100000",
  55509=>"110010010",
  55510=>"101011110",
  55511=>"110000000",
  55512=>"111000001",
  55513=>"110010010",
  55514=>"100000010",
  55515=>"001110001",
  55516=>"010100000",
  55517=>"001000000",
  55518=>"011101001",
  55519=>"111110111",
  55520=>"010001011",
  55521=>"010010110",
  55522=>"101000000",
  55523=>"000011011",
  55524=>"110101101",
  55525=>"000001101",
  55526=>"010011000",
  55527=>"000010000",
  55528=>"010011101",
  55529=>"100001111",
  55530=>"101011010",
  55531=>"010000110",
  55532=>"001010001",
  55533=>"100011011",
  55534=>"100000010",
  55535=>"111010111",
  55536=>"100000110",
  55537=>"011001110",
  55538=>"001000001",
  55539=>"101011100",
  55540=>"101101110",
  55541=>"110000100",
  55542=>"111100000",
  55543=>"001001000",
  55544=>"001010010",
  55545=>"110011101",
  55546=>"010111001",
  55547=>"010010001",
  55548=>"001100001",
  55549=>"110111101",
  55550=>"110000100",
  55551=>"100000010",
  55552=>"011110101",
  55553=>"100110100",
  55554=>"011001111",
  55555=>"101111100",
  55556=>"100001110",
  55557=>"010011110",
  55558=>"100110000",
  55559=>"011000110",
  55560=>"010111111",
  55561=>"100100111",
  55562=>"000011110",
  55563=>"110000010",
  55564=>"010111100",
  55565=>"000000010",
  55566=>"001000111",
  55567=>"110010110",
  55568=>"101101110",
  55569=>"111110001",
  55570=>"110110100",
  55571=>"111000101",
  55572=>"100011101",
  55573=>"111101111",
  55574=>"111110011",
  55575=>"110010111",
  55576=>"000101101",
  55577=>"011011110",
  55578=>"100000001",
  55579=>"111100111",
  55580=>"011001000",
  55581=>"100111011",
  55582=>"000011110",
  55583=>"000000011",
  55584=>"010001100",
  55585=>"001100010",
  55586=>"100100101",
  55587=>"011010111",
  55588=>"000111110",
  55589=>"101100101",
  55590=>"100110010",
  55591=>"111011000",
  55592=>"101100111",
  55593=>"010000101",
  55594=>"001010000",
  55595=>"011111001",
  55596=>"101101100",
  55597=>"000100011",
  55598=>"100101010",
  55599=>"001011000",
  55600=>"111010011",
  55601=>"010101111",
  55602=>"001011011",
  55603=>"010010011",
  55604=>"000010101",
  55605=>"011011000",
  55606=>"100010010",
  55607=>"101111010",
  55608=>"011100100",
  55609=>"110100011",
  55610=>"001001010",
  55611=>"010100000",
  55612=>"110000101",
  55613=>"001111100",
  55614=>"101011001",
  55615=>"111100101",
  55616=>"100100000",
  55617=>"010000101",
  55618=>"010001010",
  55619=>"111101101",
  55620=>"101111101",
  55621=>"000011110",
  55622=>"011000011",
  55623=>"101101000",
  55624=>"000110011",
  55625=>"001010001",
  55626=>"000001010",
  55627=>"000110111",
  55628=>"011010110",
  55629=>"111111010",
  55630=>"011000110",
  55631=>"111101100",
  55632=>"110110000",
  55633=>"011001011",
  55634=>"101101001",
  55635=>"100010011",
  55636=>"110111100",
  55637=>"000101010",
  55638=>"001001111",
  55639=>"011000011",
  55640=>"001000010",
  55641=>"000110011",
  55642=>"000101011",
  55643=>"101001011",
  55644=>"011100110",
  55645=>"001101100",
  55646=>"111101011",
  55647=>"110100101",
  55648=>"010000101",
  55649=>"101110111",
  55650=>"010010011",
  55651=>"001001011",
  55652=>"111001001",
  55653=>"111110011",
  55654=>"000111010",
  55655=>"000001011",
  55656=>"000111000",
  55657=>"000010110",
  55658=>"110100101",
  55659=>"111111000",
  55660=>"011100111",
  55661=>"001011111",
  55662=>"010100001",
  55663=>"000010110",
  55664=>"011100111",
  55665=>"101000110",
  55666=>"101100011",
  55667=>"011110111",
  55668=>"101110000",
  55669=>"010111110",
  55670=>"111100111",
  55671=>"001111101",
  55672=>"101011010",
  55673=>"001001101",
  55674=>"000010000",
  55675=>"000111001",
  55676=>"100011110",
  55677=>"111011010",
  55678=>"100100010",
  55679=>"000001100",
  55680=>"100111010",
  55681=>"000100101",
  55682=>"001010010",
  55683=>"100000011",
  55684=>"011100011",
  55685=>"111110100",
  55686=>"101100110",
  55687=>"000000100",
  55688=>"000101111",
  55689=>"111100011",
  55690=>"010110111",
  55691=>"111010010",
  55692=>"010101110",
  55693=>"001000110",
  55694=>"110010010",
  55695=>"001101011",
  55696=>"101001010",
  55697=>"100001111",
  55698=>"110100010",
  55699=>"010111010",
  55700=>"011001011",
  55701=>"000110000",
  55702=>"010111011",
  55703=>"001001111",
  55704=>"101101000",
  55705=>"001110111",
  55706=>"110000100",
  55707=>"000011110",
  55708=>"111001110",
  55709=>"111001111",
  55710=>"000110010",
  55711=>"111111011",
  55712=>"100001110",
  55713=>"111110011",
  55714=>"001101100",
  55715=>"001100001",
  55716=>"101100110",
  55717=>"010000000",
  55718=>"010110111",
  55719=>"111110010",
  55720=>"001111010",
  55721=>"000001111",
  55722=>"010100011",
  55723=>"110101111",
  55724=>"000001111",
  55725=>"111010111",
  55726=>"100010111",
  55727=>"000110001",
  55728=>"000010011",
  55729=>"100010001",
  55730=>"101001001",
  55731=>"110100111",
  55732=>"010111111",
  55733=>"000110011",
  55734=>"001100100",
  55735=>"101111010",
  55736=>"010011101",
  55737=>"110010010",
  55738=>"000101001",
  55739=>"011110101",
  55740=>"111011110",
  55741=>"001101100",
  55742=>"100111001",
  55743=>"001010111",
  55744=>"010001010",
  55745=>"000001000",
  55746=>"001101111",
  55747=>"001111101",
  55748=>"010010101",
  55749=>"011000100",
  55750=>"110011110",
  55751=>"111000011",
  55752=>"011010000",
  55753=>"010100110",
  55754=>"111101001",
  55755=>"100011001",
  55756=>"011000100",
  55757=>"011001100",
  55758=>"011001011",
  55759=>"010100010",
  55760=>"110110101",
  55761=>"011101000",
  55762=>"110110001",
  55763=>"010000111",
  55764=>"100001010",
  55765=>"010110111",
  55766=>"110010101",
  55767=>"010010000",
  55768=>"010010010",
  55769=>"101111001",
  55770=>"001111111",
  55771=>"011011010",
  55772=>"001010001",
  55773=>"110011001",
  55774=>"100000001",
  55775=>"110001000",
  55776=>"010000010",
  55777=>"110111011",
  55778=>"010111010",
  55779=>"001100100",
  55780=>"010011100",
  55781=>"111010111",
  55782=>"001001110",
  55783=>"101010000",
  55784=>"001110010",
  55785=>"000010000",
  55786=>"111110101",
  55787=>"100000110",
  55788=>"001010010",
  55789=>"000010101",
  55790=>"000001101",
  55791=>"001001010",
  55792=>"110101110",
  55793=>"100111100",
  55794=>"111100000",
  55795=>"011011101",
  55796=>"101100011",
  55797=>"111011111",
  55798=>"100000001",
  55799=>"010000000",
  55800=>"100101000",
  55801=>"000100001",
  55802=>"111001100",
  55803=>"110000010",
  55804=>"001001101",
  55805=>"010101111",
  55806=>"101110001",
  55807=>"111011100",
  55808=>"111100101",
  55809=>"110001001",
  55810=>"101000001",
  55811=>"100010010",
  55812=>"110110111",
  55813=>"111000110",
  55814=>"111111001",
  55815=>"000111100",
  55816=>"000100101",
  55817=>"100100000",
  55818=>"000100010",
  55819=>"110101100",
  55820=>"101001100",
  55821=>"000010101",
  55822=>"111000111",
  55823=>"011001000",
  55824=>"110011000",
  55825=>"010011110",
  55826=>"001100001",
  55827=>"000111100",
  55828=>"011000101",
  55829=>"101111111",
  55830=>"001111111",
  55831=>"111100111",
  55832=>"111010111",
  55833=>"110010010",
  55834=>"000011010",
  55835=>"101011000",
  55836=>"000001110",
  55837=>"111110011",
  55838=>"001011011",
  55839=>"010100110",
  55840=>"001011000",
  55841=>"010000110",
  55842=>"110100111",
  55843=>"000000010",
  55844=>"101100101",
  55845=>"100010000",
  55846=>"001100111",
  55847=>"011111110",
  55848=>"000101000",
  55849=>"001111010",
  55850=>"110000011",
  55851=>"110110010",
  55852=>"010100010",
  55853=>"001100010",
  55854=>"010000011",
  55855=>"001101010",
  55856=>"000010011",
  55857=>"110001100",
  55858=>"110110110",
  55859=>"000011001",
  55860=>"010000110",
  55861=>"001101001",
  55862=>"001001110",
  55863=>"111100001",
  55864=>"111001010",
  55865=>"101101010",
  55866=>"000111010",
  55867=>"000101110",
  55868=>"010110100",
  55869=>"010011111",
  55870=>"100000000",
  55871=>"011011011",
  55872=>"000100001",
  55873=>"111001000",
  55874=>"110111101",
  55875=>"011000101",
  55876=>"001000100",
  55877=>"111111110",
  55878=>"000000000",
  55879=>"010000000",
  55880=>"101100001",
  55881=>"000101011",
  55882=>"010010111",
  55883=>"010101101",
  55884=>"100011101",
  55885=>"001011010",
  55886=>"111111110",
  55887=>"000001110",
  55888=>"011010111",
  55889=>"101110001",
  55890=>"001000100",
  55891=>"001100101",
  55892=>"001111000",
  55893=>"111110101",
  55894=>"110110100",
  55895=>"001101101",
  55896=>"011110101",
  55897=>"110000001",
  55898=>"111000110",
  55899=>"000110111",
  55900=>"101101111",
  55901=>"001011011",
  55902=>"111111010",
  55903=>"001101100",
  55904=>"011011011",
  55905=>"100111001",
  55906=>"111010111",
  55907=>"011111001",
  55908=>"000111010",
  55909=>"001100100",
  55910=>"000111101",
  55911=>"101110000",
  55912=>"101010111",
  55913=>"001101100",
  55914=>"101100111",
  55915=>"100111000",
  55916=>"111000110",
  55917=>"111010110",
  55918=>"111000101",
  55919=>"101001010",
  55920=>"001101101",
  55921=>"110100111",
  55922=>"111100101",
  55923=>"100100100",
  55924=>"000010011",
  55925=>"111111101",
  55926=>"100010010",
  55927=>"101011101",
  55928=>"101110000",
  55929=>"100001111",
  55930=>"000001111",
  55931=>"101100011",
  55932=>"101100011",
  55933=>"101001100",
  55934=>"101001111",
  55935=>"001111011",
  55936=>"110110001",
  55937=>"000111111",
  55938=>"100001000",
  55939=>"010001111",
  55940=>"011001001",
  55941=>"100000111",
  55942=>"001101111",
  55943=>"111101001",
  55944=>"000111101",
  55945=>"110110111",
  55946=>"101111010",
  55947=>"001100111",
  55948=>"000101001",
  55949=>"111101000",
  55950=>"110010011",
  55951=>"010001001",
  55952=>"000001110",
  55953=>"000101011",
  55954=>"110000101",
  55955=>"011000001",
  55956=>"011001100",
  55957=>"001101011",
  55958=>"100011011",
  55959=>"100000110",
  55960=>"110100000",
  55961=>"101101100",
  55962=>"110000111",
  55963=>"100110000",
  55964=>"000100001",
  55965=>"110101010",
  55966=>"101111001",
  55967=>"011000001",
  55968=>"011101001",
  55969=>"011011110",
  55970=>"111010001",
  55971=>"010011010",
  55972=>"001100010",
  55973=>"110101001",
  55974=>"010001011",
  55975=>"101100111",
  55976=>"111011110",
  55977=>"001010000",
  55978=>"010100000",
  55979=>"110111001",
  55980=>"100110010",
  55981=>"000001001",
  55982=>"000101011",
  55983=>"111010111",
  55984=>"001010110",
  55985=>"010011001",
  55986=>"011111000",
  55987=>"000010000",
  55988=>"001001100",
  55989=>"111110011",
  55990=>"010100111",
  55991=>"001010001",
  55992=>"101011101",
  55993=>"010111000",
  55994=>"100001111",
  55995=>"011111110",
  55996=>"111011011",
  55997=>"011010000",
  55998=>"001111110",
  55999=>"001010111",
  56000=>"101000001",
  56001=>"010100101",
  56002=>"011010110",
  56003=>"000100001",
  56004=>"111001010",
  56005=>"010111110",
  56006=>"011010010",
  56007=>"111011001",
  56008=>"001000000",
  56009=>"111100100",
  56010=>"111011111",
  56011=>"100001010",
  56012=>"010010010",
  56013=>"101000011",
  56014=>"101001001",
  56015=>"110000101",
  56016=>"010100010",
  56017=>"111110001",
  56018=>"100101011",
  56019=>"000111000",
  56020=>"110111101",
  56021=>"011110110",
  56022=>"101010011",
  56023=>"100011001",
  56024=>"000001101",
  56025=>"110001100",
  56026=>"111111110",
  56027=>"001101010",
  56028=>"110110110",
  56029=>"101110101",
  56030=>"110011110",
  56031=>"111010100",
  56032=>"001101100",
  56033=>"110000101",
  56034=>"000100000",
  56035=>"000000001",
  56036=>"111001110",
  56037=>"110111111",
  56038=>"101110000",
  56039=>"111000011",
  56040=>"001001000",
  56041=>"010101000",
  56042=>"101010100",
  56043=>"000110111",
  56044=>"010011101",
  56045=>"011100101",
  56046=>"100101100",
  56047=>"010010000",
  56048=>"100011011",
  56049=>"000000011",
  56050=>"101000010",
  56051=>"111101010",
  56052=>"000010010",
  56053=>"100000101",
  56054=>"010110000",
  56055=>"000001110",
  56056=>"100010001",
  56057=>"101111100",
  56058=>"101000010",
  56059=>"001101111",
  56060=>"110111011",
  56061=>"111010101",
  56062=>"010001001",
  56063=>"010011010",
  56064=>"100110101",
  56065=>"110111101",
  56066=>"100100111",
  56067=>"111011001",
  56068=>"111111111",
  56069=>"011000111",
  56070=>"110100001",
  56071=>"010001010",
  56072=>"011101001",
  56073=>"101000111",
  56074=>"000011000",
  56075=>"100101111",
  56076=>"100100010",
  56077=>"100000110",
  56078=>"010001001",
  56079=>"101010000",
  56080=>"111101010",
  56081=>"001000011",
  56082=>"100101010",
  56083=>"011110001",
  56084=>"011101011",
  56085=>"100010001",
  56086=>"110101010",
  56087=>"001000110",
  56088=>"111011101",
  56089=>"001100111",
  56090=>"100000100",
  56091=>"110100001",
  56092=>"111110010",
  56093=>"110000001",
  56094=>"111001011",
  56095=>"100101011",
  56096=>"111100000",
  56097=>"110100010",
  56098=>"100111101",
  56099=>"111100000",
  56100=>"001010101",
  56101=>"111101001",
  56102=>"100101010",
  56103=>"100010100",
  56104=>"000001000",
  56105=>"000101001",
  56106=>"111001000",
  56107=>"101011000",
  56108=>"001001100",
  56109=>"000101110",
  56110=>"010101010",
  56111=>"000101110",
  56112=>"000000101",
  56113=>"000111010",
  56114=>"101000110",
  56115=>"011000100",
  56116=>"000111111",
  56117=>"100100001",
  56118=>"000110111",
  56119=>"001001111",
  56120=>"001111001",
  56121=>"010100000",
  56122=>"011000001",
  56123=>"010111100",
  56124=>"001111011",
  56125=>"110011101",
  56126=>"010010010",
  56127=>"110011111",
  56128=>"111101100",
  56129=>"111010011",
  56130=>"000100100",
  56131=>"100011101",
  56132=>"101000110",
  56133=>"001000100",
  56134=>"101011011",
  56135=>"011001001",
  56136=>"100101110",
  56137=>"110111010",
  56138=>"000001110",
  56139=>"101111110",
  56140=>"001010110",
  56141=>"010110110",
  56142=>"110010100",
  56143=>"111001111",
  56144=>"010010111",
  56145=>"001001100",
  56146=>"010001100",
  56147=>"101010100",
  56148=>"011011101",
  56149=>"001000001",
  56150=>"000100111",
  56151=>"001001000",
  56152=>"101001000",
  56153=>"101010000",
  56154=>"011010000",
  56155=>"101001000",
  56156=>"111011110",
  56157=>"000000011",
  56158=>"011110010",
  56159=>"111101100",
  56160=>"001001111",
  56161=>"101111010",
  56162=>"110001101",
  56163=>"011101110",
  56164=>"111001100",
  56165=>"010101111",
  56166=>"000010010",
  56167=>"001001110",
  56168=>"100111100",
  56169=>"000011100",
  56170=>"000101111",
  56171=>"010001010",
  56172=>"000000100",
  56173=>"000101010",
  56174=>"101000010",
  56175=>"110111000",
  56176=>"111001111",
  56177=>"010100111",
  56178=>"100011001",
  56179=>"100101000",
  56180=>"110110101",
  56181=>"010110010",
  56182=>"110101101",
  56183=>"110001000",
  56184=>"010110010",
  56185=>"111111100",
  56186=>"101101101",
  56187=>"110110011",
  56188=>"111110100",
  56189=>"011110101",
  56190=>"010111101",
  56191=>"010000101",
  56192=>"110101111",
  56193=>"101110101",
  56194=>"011010111",
  56195=>"000010001",
  56196=>"000001000",
  56197=>"011101001",
  56198=>"101000001",
  56199=>"101000110",
  56200=>"000101100",
  56201=>"011011101",
  56202=>"110111101",
  56203=>"101110010",
  56204=>"001011111",
  56205=>"111101111",
  56206=>"000000001",
  56207=>"000101001",
  56208=>"001111010",
  56209=>"000000000",
  56210=>"111111001",
  56211=>"110011110",
  56212=>"100010010",
  56213=>"101011100",
  56214=>"001100010",
  56215=>"111111110",
  56216=>"100010110",
  56217=>"101101000",
  56218=>"011000000",
  56219=>"011100001",
  56220=>"000111010",
  56221=>"011000011",
  56222=>"111100111",
  56223=>"110100010",
  56224=>"001010110",
  56225=>"110001001",
  56226=>"111110101",
  56227=>"000011010",
  56228=>"000100110",
  56229=>"100101000",
  56230=>"010101010",
  56231=>"111000001",
  56232=>"001110011",
  56233=>"111111010",
  56234=>"110100110",
  56235=>"011001111",
  56236=>"000110110",
  56237=>"101001100",
  56238=>"010100100",
  56239=>"010010101",
  56240=>"000001010",
  56241=>"110000000",
  56242=>"000000110",
  56243=>"010110011",
  56244=>"011011011",
  56245=>"111100011",
  56246=>"110010010",
  56247=>"001101010",
  56248=>"101111010",
  56249=>"101011010",
  56250=>"101101100",
  56251=>"011110000",
  56252=>"011100001",
  56253=>"111001000",
  56254=>"011000010",
  56255=>"101110110",
  56256=>"101100111",
  56257=>"010110000",
  56258=>"111000101",
  56259=>"111011000",
  56260=>"011101011",
  56261=>"101001101",
  56262=>"110011010",
  56263=>"110000000",
  56264=>"110111110",
  56265=>"000000010",
  56266=>"010010100",
  56267=>"011001100",
  56268=>"011010100",
  56269=>"010010000",
  56270=>"100001101",
  56271=>"011001111",
  56272=>"001101100",
  56273=>"101111010",
  56274=>"111111001",
  56275=>"010110111",
  56276=>"100100101",
  56277=>"000011000",
  56278=>"100000000",
  56279=>"101001100",
  56280=>"010010000",
  56281=>"001111100",
  56282=>"010110101",
  56283=>"001110100",
  56284=>"111010111",
  56285=>"000110101",
  56286=>"011100110",
  56287=>"000001001",
  56288=>"000011111",
  56289=>"111011010",
  56290=>"010011100",
  56291=>"110111101",
  56292=>"100001001",
  56293=>"000010000",
  56294=>"010010111",
  56295=>"101000000",
  56296=>"001110001",
  56297=>"111111001",
  56298=>"010000011",
  56299=>"100001001",
  56300=>"011111111",
  56301=>"110100101",
  56302=>"110110111",
  56303=>"110100001",
  56304=>"010011001",
  56305=>"100100011",
  56306=>"111010101",
  56307=>"111001000",
  56308=>"010010001",
  56309=>"111101010",
  56310=>"111110001",
  56311=>"010010011",
  56312=>"100010000",
  56313=>"000000100",
  56314=>"010100100",
  56315=>"000010010",
  56316=>"110001001",
  56317=>"000001001",
  56318=>"100100100",
  56319=>"111000001",
  56320=>"010010011",
  56321=>"011101010",
  56322=>"000100101",
  56323=>"010101101",
  56324=>"000100100",
  56325=>"110111110",
  56326=>"001101000",
  56327=>"100001101",
  56328=>"110000110",
  56329=>"110100111",
  56330=>"111010000",
  56331=>"001100101",
  56332=>"001111011",
  56333=>"011011010",
  56334=>"011001000",
  56335=>"111001110",
  56336=>"010001010",
  56337=>"011011000",
  56338=>"010001100",
  56339=>"001101100",
  56340=>"010001111",
  56341=>"010011001",
  56342=>"010010000",
  56343=>"001111100",
  56344=>"000010100",
  56345=>"111100110",
  56346=>"100101000",
  56347=>"000011001",
  56348=>"100011100",
  56349=>"101101111",
  56350=>"001010111",
  56351=>"110000010",
  56352=>"001000010",
  56353=>"010110010",
  56354=>"011001100",
  56355=>"010000100",
  56356=>"010111100",
  56357=>"000001001",
  56358=>"000001000",
  56359=>"100101010",
  56360=>"100101111",
  56361=>"010010000",
  56362=>"111011110",
  56363=>"110110001",
  56364=>"101111110",
  56365=>"000110010",
  56366=>"010001010",
  56367=>"101101010",
  56368=>"110110011",
  56369=>"111010000",
  56370=>"010100000",
  56371=>"000001000",
  56372=>"100101111",
  56373=>"011110001",
  56374=>"001100111",
  56375=>"110111100",
  56376=>"111001011",
  56377=>"110000001",
  56378=>"010010001",
  56379=>"010111111",
  56380=>"010000011",
  56381=>"101001001",
  56382=>"011011000",
  56383=>"011001100",
  56384=>"110100011",
  56385=>"011100000",
  56386=>"010010111",
  56387=>"011101110",
  56388=>"010100010",
  56389=>"111100000",
  56390=>"100011000",
  56391=>"101001011",
  56392=>"001010010",
  56393=>"111110011",
  56394=>"100000101",
  56395=>"100011001",
  56396=>"010000101",
  56397=>"000101101",
  56398=>"000111010",
  56399=>"101110111",
  56400=>"011111000",
  56401=>"100101110",
  56402=>"110110111",
  56403=>"100100001",
  56404=>"010011101",
  56405=>"001110110",
  56406=>"000111100",
  56407=>"011110001",
  56408=>"110000111",
  56409=>"011011111",
  56410=>"110001111",
  56411=>"111101111",
  56412=>"100110010",
  56413=>"010101101",
  56414=>"001001110",
  56415=>"100001100",
  56416=>"110010101",
  56417=>"001111111",
  56418=>"110000000",
  56419=>"010011010",
  56420=>"101101100",
  56421=>"100111011",
  56422=>"010110010",
  56423=>"010010101",
  56424=>"101011011",
  56425=>"110100100",
  56426=>"111101100",
  56427=>"001011111",
  56428=>"110110000",
  56429=>"000010010",
  56430=>"010101100",
  56431=>"100000111",
  56432=>"110000110",
  56433=>"100000000",
  56434=>"001101101",
  56435=>"101000101",
  56436=>"110011010",
  56437=>"011111001",
  56438=>"010111101",
  56439=>"011111100",
  56440=>"100111000",
  56441=>"011010011",
  56442=>"001101011",
  56443=>"011000011",
  56444=>"010001100",
  56445=>"011111101",
  56446=>"111111101",
  56447=>"110111100",
  56448=>"101100101",
  56449=>"101111001",
  56450=>"111100010",
  56451=>"110000101",
  56452=>"111011001",
  56453=>"000001010",
  56454=>"100111011",
  56455=>"000111100",
  56456=>"000001000",
  56457=>"000000001",
  56458=>"001011011",
  56459=>"001010111",
  56460=>"101100000",
  56461=>"010111010",
  56462=>"101100111",
  56463=>"011101110",
  56464=>"101000110",
  56465=>"000010000",
  56466=>"001100000",
  56467=>"000110101",
  56468=>"110001000",
  56469=>"011110011",
  56470=>"011111111",
  56471=>"100110100",
  56472=>"101011010",
  56473=>"001101111",
  56474=>"110110100",
  56475=>"100000010",
  56476=>"010100000",
  56477=>"001010100",
  56478=>"000101110",
  56479=>"011001010",
  56480=>"100001101",
  56481=>"111100000",
  56482=>"011101001",
  56483=>"011101000",
  56484=>"110010010",
  56485=>"001101101",
  56486=>"010101010",
  56487=>"000110101",
  56488=>"001111110",
  56489=>"100100100",
  56490=>"100110000",
  56491=>"010101101",
  56492=>"011100010",
  56493=>"010001000",
  56494=>"110010011",
  56495=>"001010001",
  56496=>"001101000",
  56497=>"011000100",
  56498=>"011111000",
  56499=>"111110110",
  56500=>"010111101",
  56501=>"011011000",
  56502=>"011100001",
  56503=>"110111011",
  56504=>"001101001",
  56505=>"011101000",
  56506=>"110111001",
  56507=>"110001111",
  56508=>"000011000",
  56509=>"110100001",
  56510=>"111000101",
  56511=>"010000000",
  56512=>"010100101",
  56513=>"001010110",
  56514=>"100000011",
  56515=>"110111000",
  56516=>"000111011",
  56517=>"001111010",
  56518=>"000010111",
  56519=>"110100111",
  56520=>"001010100",
  56521=>"111100010",
  56522=>"001111000",
  56523=>"010100000",
  56524=>"000011001",
  56525=>"100101100",
  56526=>"100100001",
  56527=>"011001100",
  56528=>"110101101",
  56529=>"011111010",
  56530=>"010000010",
  56531=>"000101010",
  56532=>"110000011",
  56533=>"000011111",
  56534=>"000001111",
  56535=>"101111001",
  56536=>"011111011",
  56537=>"100111011",
  56538=>"111110000",
  56539=>"001110110",
  56540=>"111010101",
  56541=>"010000001",
  56542=>"010011010",
  56543=>"010010001",
  56544=>"010100010",
  56545=>"111100010",
  56546=>"111100100",
  56547=>"000110010",
  56548=>"011111001",
  56549=>"101100111",
  56550=>"110100000",
  56551=>"101101100",
  56552=>"111110000",
  56553=>"100001000",
  56554=>"100111111",
  56555=>"010001010",
  56556=>"010111111",
  56557=>"111110001",
  56558=>"110100001",
  56559=>"100101000",
  56560=>"001001000",
  56561=>"011101001",
  56562=>"010101001",
  56563=>"110000001",
  56564=>"101000001",
  56565=>"000011011",
  56566=>"010111011",
  56567=>"010010011",
  56568=>"101000100",
  56569=>"111101110",
  56570=>"001011010",
  56571=>"000110100",
  56572=>"011110010",
  56573=>"001010011",
  56574=>"111001101",
  56575=>"110001111",
  56576=>"001001100",
  56577=>"111111111",
  56578=>"001101111",
  56579=>"101100001",
  56580=>"000111110",
  56581=>"010011111",
  56582=>"010111011",
  56583=>"110000000",
  56584=>"001000110",
  56585=>"001011111",
  56586=>"000100100",
  56587=>"111111111",
  56588=>"011100010",
  56589=>"000100110",
  56590=>"111000101",
  56591=>"100110100",
  56592=>"101001101",
  56593=>"111011111",
  56594=>"010001100",
  56595=>"000111100",
  56596=>"010111000",
  56597=>"100101001",
  56598=>"110000100",
  56599=>"111100111",
  56600=>"110000000",
  56601=>"101101100",
  56602=>"011000111",
  56603=>"100100101",
  56604=>"000000010",
  56605=>"111001011",
  56606=>"101000100",
  56607=>"110111110",
  56608=>"010110010",
  56609=>"000001100",
  56610=>"100000111",
  56611=>"110100011",
  56612=>"000011111",
  56613=>"100100100",
  56614=>"111110011",
  56615=>"010111000",
  56616=>"101101101",
  56617=>"000100011",
  56618=>"110100010",
  56619=>"100101110",
  56620=>"111011111",
  56621=>"111010100",
  56622=>"011001101",
  56623=>"011000110",
  56624=>"101111000",
  56625=>"111000101",
  56626=>"100100010",
  56627=>"000000011",
  56628=>"101011101",
  56629=>"110011001",
  56630=>"110111111",
  56631=>"001110110",
  56632=>"110001111",
  56633=>"110001011",
  56634=>"010011010",
  56635=>"000000000",
  56636=>"001011001",
  56637=>"111000100",
  56638=>"010111011",
  56639=>"010100100",
  56640=>"110110000",
  56641=>"110000011",
  56642=>"111000001",
  56643=>"110111000",
  56644=>"100000110",
  56645=>"101101111",
  56646=>"001111010",
  56647=>"100011100",
  56648=>"111110110",
  56649=>"001001000",
  56650=>"111111111",
  56651=>"001011011",
  56652=>"010101100",
  56653=>"101000110",
  56654=>"001100011",
  56655=>"011100110",
  56656=>"110101001",
  56657=>"001100100",
  56658=>"111111101",
  56659=>"000100001",
  56660=>"010100101",
  56661=>"111110111",
  56662=>"000010011",
  56663=>"000001000",
  56664=>"110110000",
  56665=>"001010000",
  56666=>"111010111",
  56667=>"000000101",
  56668=>"010001010",
  56669=>"001010001",
  56670=>"111100110",
  56671=>"011110001",
  56672=>"101001111",
  56673=>"011000101",
  56674=>"101000100",
  56675=>"000100110",
  56676=>"000101010",
  56677=>"101001101",
  56678=>"001000000",
  56679=>"001110000",
  56680=>"010101001",
  56681=>"000000100",
  56682=>"001100001",
  56683=>"000001011",
  56684=>"010100000",
  56685=>"000111010",
  56686=>"110100001",
  56687=>"010010110",
  56688=>"110100011",
  56689=>"000000001",
  56690=>"100111001",
  56691=>"010110100",
  56692=>"110011101",
  56693=>"001110111",
  56694=>"110100111",
  56695=>"010100111",
  56696=>"001000000",
  56697=>"001001111",
  56698=>"110111111",
  56699=>"100100110",
  56700=>"001010111",
  56701=>"000111101",
  56702=>"100000101",
  56703=>"011010011",
  56704=>"001011101",
  56705=>"100101100",
  56706=>"010011101",
  56707=>"100100001",
  56708=>"011010100",
  56709=>"010000001",
  56710=>"100000111",
  56711=>"111101000",
  56712=>"000111111",
  56713=>"111101001",
  56714=>"111111011",
  56715=>"000000101",
  56716=>"011010110",
  56717=>"110100010",
  56718=>"000100011",
  56719=>"011000100",
  56720=>"001111011",
  56721=>"111111110",
  56722=>"000101110",
  56723=>"010011011",
  56724=>"110100010",
  56725=>"011000010",
  56726=>"010110000",
  56727=>"110000000",
  56728=>"000110100",
  56729=>"110000111",
  56730=>"100110000",
  56731=>"111101011",
  56732=>"000000010",
  56733=>"111100110",
  56734=>"100011110",
  56735=>"111010101",
  56736=>"010011101",
  56737=>"011011010",
  56738=>"010001001",
  56739=>"100101010",
  56740=>"110110011",
  56741=>"001100011",
  56742=>"110111100",
  56743=>"101100001",
  56744=>"111111010",
  56745=>"110010100",
  56746=>"001110110",
  56747=>"010110111",
  56748=>"101111010",
  56749=>"011101110",
  56750=>"101001100",
  56751=>"111100000",
  56752=>"101000100",
  56753=>"011111011",
  56754=>"111101101",
  56755=>"011000100",
  56756=>"011100011",
  56757=>"110110110",
  56758=>"000101110",
  56759=>"110010111",
  56760=>"110110011",
  56761=>"100111001",
  56762=>"000100011",
  56763=>"100001010",
  56764=>"011010010",
  56765=>"110100001",
  56766=>"110000100",
  56767=>"111101111",
  56768=>"110010111",
  56769=>"001111100",
  56770=>"001110011",
  56771=>"000001001",
  56772=>"100001011",
  56773=>"111101010",
  56774=>"000001111",
  56775=>"110100000",
  56776=>"100101011",
  56777=>"101010001",
  56778=>"110100101",
  56779=>"101111111",
  56780=>"100101001",
  56781=>"100010100",
  56782=>"010001001",
  56783=>"100011111",
  56784=>"101110011",
  56785=>"001010111",
  56786=>"101010011",
  56787=>"010111010",
  56788=>"110010100",
  56789=>"000110101",
  56790=>"111110000",
  56791=>"111101100",
  56792=>"010110110",
  56793=>"000000111",
  56794=>"000111111",
  56795=>"111010100",
  56796=>"000010101",
  56797=>"000100100",
  56798=>"111010111",
  56799=>"000101110",
  56800=>"000111110",
  56801=>"110101000",
  56802=>"011010110",
  56803=>"000111001",
  56804=>"100001011",
  56805=>"011111001",
  56806=>"010000111",
  56807=>"011101000",
  56808=>"110100010",
  56809=>"010101110",
  56810=>"001100100",
  56811=>"110011000",
  56812=>"011000111",
  56813=>"000110011",
  56814=>"010100111",
  56815=>"010100010",
  56816=>"101010001",
  56817=>"010011110",
  56818=>"100100111",
  56819=>"101111101",
  56820=>"110111001",
  56821=>"010111101",
  56822=>"000011010",
  56823=>"001100010",
  56824=>"100111010",
  56825=>"111101001",
  56826=>"110111011",
  56827=>"011110001",
  56828=>"001001001",
  56829=>"110111001",
  56830=>"111100001",
  56831=>"001000100",
  56832=>"001001110",
  56833=>"011010101",
  56834=>"111111000",
  56835=>"111101100",
  56836=>"011111110",
  56837=>"011000111",
  56838=>"100001001",
  56839=>"110101101",
  56840=>"110011100",
  56841=>"110111101",
  56842=>"100101100",
  56843=>"100111001",
  56844=>"011111101",
  56845=>"010001011",
  56846=>"010010110",
  56847=>"001000001",
  56848=>"011001111",
  56849=>"001011101",
  56850=>"111001110",
  56851=>"010100111",
  56852=>"110011100",
  56853=>"101000000",
  56854=>"000101100",
  56855=>"101111101",
  56856=>"111011100",
  56857=>"001111111",
  56858=>"111111111",
  56859=>"010110011",
  56860=>"001011111",
  56861=>"100011011",
  56862=>"111100111",
  56863=>"001100100",
  56864=>"001001010",
  56865=>"111111111",
  56866=>"000011001",
  56867=>"010011110",
  56868=>"111111110",
  56869=>"001000111",
  56870=>"001001110",
  56871=>"001101000",
  56872=>"110001100",
  56873=>"101011010",
  56874=>"010101010",
  56875=>"000100101",
  56876=>"100100011",
  56877=>"111000010",
  56878=>"000011111",
  56879=>"000101010",
  56880=>"011011010",
  56881=>"001100011",
  56882=>"100100100",
  56883=>"000110100",
  56884=>"101100100",
  56885=>"011001010",
  56886=>"010101011",
  56887=>"010001000",
  56888=>"001101000",
  56889=>"111111001",
  56890=>"001101110",
  56891=>"010101000",
  56892=>"011101000",
  56893=>"011111100",
  56894=>"001011100",
  56895=>"011000111",
  56896=>"101000101",
  56897=>"010010000",
  56898=>"011101011",
  56899=>"011101101",
  56900=>"111000110",
  56901=>"010001010",
  56902=>"111100101",
  56903=>"110100010",
  56904=>"111111001",
  56905=>"001000001",
  56906=>"111101111",
  56907=>"001100101",
  56908=>"001100011",
  56909=>"011100111",
  56910=>"100111010",
  56911=>"100110101",
  56912=>"111111011",
  56913=>"001100000",
  56914=>"011010000",
  56915=>"110001110",
  56916=>"010100111",
  56917=>"100001100",
  56918=>"000000101",
  56919=>"101011111",
  56920=>"000000000",
  56921=>"101010100",
  56922=>"000111000",
  56923=>"000110001",
  56924=>"100100010",
  56925=>"100100000",
  56926=>"110001011",
  56927=>"111000110",
  56928=>"001011110",
  56929=>"100110000",
  56930=>"000110101",
  56931=>"110110111",
  56932=>"111101011",
  56933=>"011111111",
  56934=>"001010011",
  56935=>"111100011",
  56936=>"001111101",
  56937=>"000011110",
  56938=>"000001010",
  56939=>"101110111",
  56940=>"100010010",
  56941=>"110010000",
  56942=>"000010001",
  56943=>"001001110",
  56944=>"110010011",
  56945=>"000100111",
  56946=>"010000100",
  56947=>"010111011",
  56948=>"000010000",
  56949=>"001001111",
  56950=>"011111110",
  56951=>"110010010",
  56952=>"111111100",
  56953=>"110011010",
  56954=>"101010011",
  56955=>"110010111",
  56956=>"101011100",
  56957=>"101001100",
  56958=>"010110011",
  56959=>"011000010",
  56960=>"110011101",
  56961=>"110101001",
  56962=>"011110100",
  56963=>"111111010",
  56964=>"111001001",
  56965=>"001000110",
  56966=>"010101010",
  56967=>"010111000",
  56968=>"100101111",
  56969=>"111010101",
  56970=>"110110010",
  56971=>"100101010",
  56972=>"010001110",
  56973=>"000000010",
  56974=>"101000000",
  56975=>"001011100",
  56976=>"100101011",
  56977=>"000101101",
  56978=>"101110111",
  56979=>"110000001",
  56980=>"100010010",
  56981=>"101011011",
  56982=>"000000001",
  56983=>"101100110",
  56984=>"011001010",
  56985=>"100011011",
  56986=>"010101100",
  56987=>"110000110",
  56988=>"101011011",
  56989=>"010011010",
  56990=>"010110111",
  56991=>"100010101",
  56992=>"100001100",
  56993=>"110101010",
  56994=>"111101111",
  56995=>"101000001",
  56996=>"110000100",
  56997=>"010010011",
  56998=>"110101001",
  56999=>"000101010",
  57000=>"001101100",
  57001=>"000001010",
  57002=>"100101100",
  57003=>"111011110",
  57004=>"100111111",
  57005=>"100100011",
  57006=>"111000100",
  57007=>"101010111",
  57008=>"101101001",
  57009=>"000101101",
  57010=>"100110111",
  57011=>"100101110",
  57012=>"010011101",
  57013=>"110110111",
  57014=>"101101001",
  57015=>"011000100",
  57016=>"010000001",
  57017=>"110110001",
  57018=>"001000111",
  57019=>"001011100",
  57020=>"110010101",
  57021=>"011100101",
  57022=>"111111101",
  57023=>"011111000",
  57024=>"111011111",
  57025=>"100010000",
  57026=>"101111110",
  57027=>"010101001",
  57028=>"011100101",
  57029=>"110000100",
  57030=>"011011000",
  57031=>"011010111",
  57032=>"010111011",
  57033=>"101101011",
  57034=>"111101100",
  57035=>"000110111",
  57036=>"110100101",
  57037=>"000100101",
  57038=>"000101110",
  57039=>"011001010",
  57040=>"100111011",
  57041=>"110010010",
  57042=>"110000001",
  57043=>"110101101",
  57044=>"000000110",
  57045=>"011110010",
  57046=>"001111011",
  57047=>"100110011",
  57048=>"111111100",
  57049=>"001111100",
  57050=>"001000010",
  57051=>"111101011",
  57052=>"101111100",
  57053=>"101110010",
  57054=>"100111100",
  57055=>"110111101",
  57056=>"010000111",
  57057=>"001011010",
  57058=>"001011000",
  57059=>"100110011",
  57060=>"110111001",
  57061=>"101010000",
  57062=>"110010111",
  57063=>"011011100",
  57064=>"101100111",
  57065=>"111110101",
  57066=>"110100101",
  57067=>"001110110",
  57068=>"011011100",
  57069=>"111110100",
  57070=>"000110001",
  57071=>"111110111",
  57072=>"111101000",
  57073=>"001101110",
  57074=>"001011110",
  57075=>"101000001",
  57076=>"101100000",
  57077=>"100000101",
  57078=>"000110101",
  57079=>"001110110",
  57080=>"110010011",
  57081=>"010010000",
  57082=>"100011011",
  57083=>"010010011",
  57084=>"111100101",
  57085=>"010101000",
  57086=>"111110101",
  57087=>"100010000",
  57088=>"101111000",
  57089=>"101101111",
  57090=>"101100011",
  57091=>"000110001",
  57092=>"000001111",
  57093=>"001101111",
  57094=>"011101111",
  57095=>"011010011",
  57096=>"000111101",
  57097=>"011101111",
  57098=>"100110110",
  57099=>"110010000",
  57100=>"011110010",
  57101=>"101010010",
  57102=>"101001000",
  57103=>"111010110",
  57104=>"110011010",
  57105=>"110101111",
  57106=>"000000100",
  57107=>"010011011",
  57108=>"100001100",
  57109=>"111110101",
  57110=>"001101010",
  57111=>"000100001",
  57112=>"010010000",
  57113=>"100100011",
  57114=>"001111111",
  57115=>"100001010",
  57116=>"011000011",
  57117=>"111011111",
  57118=>"000100010",
  57119=>"111111100",
  57120=>"100011110",
  57121=>"101101101",
  57122=>"101000110",
  57123=>"000100001",
  57124=>"100100110",
  57125=>"111101001",
  57126=>"101010111",
  57127=>"100100100",
  57128=>"010001111",
  57129=>"101111001",
  57130=>"101001011",
  57131=>"001001111",
  57132=>"001000111",
  57133=>"010100010",
  57134=>"000100011",
  57135=>"001000110",
  57136=>"110110011",
  57137=>"101001010",
  57138=>"010111010",
  57139=>"110101101",
  57140=>"001010111",
  57141=>"101010000",
  57142=>"011110011",
  57143=>"100111011",
  57144=>"111111011",
  57145=>"000100010",
  57146=>"001010011",
  57147=>"011110001",
  57148=>"010111011",
  57149=>"000000000",
  57150=>"110010111",
  57151=>"000111001",
  57152=>"100010111",
  57153=>"100000110",
  57154=>"111110101",
  57155=>"000001100",
  57156=>"000101101",
  57157=>"011010111",
  57158=>"100100101",
  57159=>"100000110",
  57160=>"111011110",
  57161=>"111011000",
  57162=>"000101110",
  57163=>"000110010",
  57164=>"111011001",
  57165=>"100100101",
  57166=>"110101110",
  57167=>"000000001",
  57168=>"100100100",
  57169=>"011101001",
  57170=>"001001101",
  57171=>"000001111",
  57172=>"100000000",
  57173=>"111111001",
  57174=>"001100000",
  57175=>"101110101",
  57176=>"111001111",
  57177=>"001000010",
  57178=>"111110101",
  57179=>"101010000",
  57180=>"110000110",
  57181=>"110000001",
  57182=>"010010010",
  57183=>"010110011",
  57184=>"010010111",
  57185=>"111011000",
  57186=>"100111010",
  57187=>"010111100",
  57188=>"010101010",
  57189=>"001001011",
  57190=>"000110010",
  57191=>"110000011",
  57192=>"101100110",
  57193=>"110010101",
  57194=>"111001111",
  57195=>"100101101",
  57196=>"010001110",
  57197=>"111010110",
  57198=>"100001101",
  57199=>"010010001",
  57200=>"001110011",
  57201=>"110001001",
  57202=>"100001101",
  57203=>"100100011",
  57204=>"011010111",
  57205=>"011110110",
  57206=>"000000000",
  57207=>"111001001",
  57208=>"100011000",
  57209=>"000111110",
  57210=>"000011001",
  57211=>"000111101",
  57212=>"100000001",
  57213=>"001001110",
  57214=>"100101100",
  57215=>"111010011",
  57216=>"001110001",
  57217=>"100010111",
  57218=>"011001100",
  57219=>"110111010",
  57220=>"101000001",
  57221=>"100000010",
  57222=>"000101110",
  57223=>"000110100",
  57224=>"111101010",
  57225=>"000011001",
  57226=>"000010000",
  57227=>"010001110",
  57228=>"101011010",
  57229=>"101101110",
  57230=>"000110001",
  57231=>"101011110",
  57232=>"010000001",
  57233=>"100001110",
  57234=>"111111100",
  57235=>"000110111",
  57236=>"011000000",
  57237=>"000100010",
  57238=>"000101111",
  57239=>"010111010",
  57240=>"101100010",
  57241=>"000000111",
  57242=>"110010101",
  57243=>"011100010",
  57244=>"100100111",
  57245=>"010100011",
  57246=>"001011011",
  57247=>"000011110",
  57248=>"101111011",
  57249=>"011101111",
  57250=>"000110111",
  57251=>"100101010",
  57252=>"110001010",
  57253=>"011010010",
  57254=>"010010100",
  57255=>"010010011",
  57256=>"010001001",
  57257=>"001110000",
  57258=>"111110110",
  57259=>"011110111",
  57260=>"101010000",
  57261=>"010110011",
  57262=>"010010101",
  57263=>"011111111",
  57264=>"010001110",
  57265=>"010111000",
  57266=>"001111010",
  57267=>"000011000",
  57268=>"101000010",
  57269=>"001001001",
  57270=>"110011011",
  57271=>"001011001",
  57272=>"001111010",
  57273=>"000100000",
  57274=>"111011101",
  57275=>"101100101",
  57276=>"111111110",
  57277=>"011101111",
  57278=>"001100000",
  57279=>"001000110",
  57280=>"100111000",
  57281=>"010010011",
  57282=>"001111111",
  57283=>"010010011",
  57284=>"010000100",
  57285=>"001011000",
  57286=>"100000101",
  57287=>"111110001",
  57288=>"111110001",
  57289=>"100010000",
  57290=>"111110111",
  57291=>"011101111",
  57292=>"111010111",
  57293=>"000011100",
  57294=>"000100100",
  57295=>"110010111",
  57296=>"111100111",
  57297=>"110010011",
  57298=>"001111111",
  57299=>"111111111",
  57300=>"011001001",
  57301=>"110101101",
  57302=>"010011101",
  57303=>"010011100",
  57304=>"111011000",
  57305=>"000111011",
  57306=>"101010010",
  57307=>"011001000",
  57308=>"111100111",
  57309=>"100001011",
  57310=>"100001101",
  57311=>"000101100",
  57312=>"000111111",
  57313=>"011101111",
  57314=>"111111110",
  57315=>"110110100",
  57316=>"011000011",
  57317=>"111001111",
  57318=>"101110011",
  57319=>"000100100",
  57320=>"000001010",
  57321=>"010001110",
  57322=>"010100101",
  57323=>"110000001",
  57324=>"010010110",
  57325=>"111011010",
  57326=>"000100000",
  57327=>"010011100",
  57328=>"101111111",
  57329=>"111001100",
  57330=>"101011110",
  57331=>"001101111",
  57332=>"000010101",
  57333=>"011010011",
  57334=>"011101110",
  57335=>"011011110",
  57336=>"111000010",
  57337=>"001001111",
  57338=>"000111110",
  57339=>"000100010",
  57340=>"011101000",
  57341=>"011100001",
  57342=>"011111101",
  57343=>"100011001",
  57344=>"111001110",
  57345=>"001100011",
  57346=>"100000100",
  57347=>"111001001",
  57348=>"000000101",
  57349=>"100001011",
  57350=>"100001101",
  57351=>"010111111",
  57352=>"010000011",
  57353=>"000001001",
  57354=>"001001111",
  57355=>"110100000",
  57356=>"111011110",
  57357=>"100010111",
  57358=>"011010000",
  57359=>"111101000",
  57360=>"010001001",
  57361=>"110000111",
  57362=>"010110100",
  57363=>"011100110",
  57364=>"111111111",
  57365=>"100010101",
  57366=>"011001110",
  57367=>"011111000",
  57368=>"100011000",
  57369=>"101000001",
  57370=>"000011101",
  57371=>"110110101",
  57372=>"110100000",
  57373=>"101010111",
  57374=>"001000001",
  57375=>"011000000",
  57376=>"101000001",
  57377=>"000010000",
  57378=>"100110001",
  57379=>"111010011",
  57380=>"010101010",
  57381=>"011001001",
  57382=>"001000111",
  57383=>"111001011",
  57384=>"111000100",
  57385=>"111000101",
  57386=>"100100001",
  57387=>"110110010",
  57388=>"000100000",
  57389=>"101010110",
  57390=>"101010111",
  57391=>"000111001",
  57392=>"110110011",
  57393=>"001001111",
  57394=>"010100011",
  57395=>"100110101",
  57396=>"001110000",
  57397=>"001111010",
  57398=>"001000100",
  57399=>"000001101",
  57400=>"011011111",
  57401=>"001010001",
  57402=>"000100101",
  57403=>"101100011",
  57404=>"010111010",
  57405=>"001101010",
  57406=>"110000001",
  57407=>"011010100",
  57408=>"111010111",
  57409=>"100111010",
  57410=>"101001010",
  57411=>"100100100",
  57412=>"101011110",
  57413=>"110100111",
  57414=>"001110111",
  57415=>"100010000",
  57416=>"111001001",
  57417=>"110001110",
  57418=>"001011011",
  57419=>"000001010",
  57420=>"001110000",
  57421=>"000100000",
  57422=>"000001000",
  57423=>"101001101",
  57424=>"010111001",
  57425=>"010000000",
  57426=>"011000010",
  57427=>"010110000",
  57428=>"101110011",
  57429=>"110111110",
  57430=>"101100011",
  57431=>"010010010",
  57432=>"110001010",
  57433=>"011001000",
  57434=>"101001111",
  57435=>"101010001",
  57436=>"011010001",
  57437=>"011010101",
  57438=>"001111101",
  57439=>"010011011",
  57440=>"010010010",
  57441=>"111011111",
  57442=>"111010001",
  57443=>"001110010",
  57444=>"000111001",
  57445=>"110110001",
  57446=>"101110011",
  57447=>"101011000",
  57448=>"000100110",
  57449=>"000111100",
  57450=>"111100101",
  57451=>"111101010",
  57452=>"111101111",
  57453=>"011000010",
  57454=>"011101001",
  57455=>"011010010",
  57456=>"001010000",
  57457=>"000101100",
  57458=>"000010100",
  57459=>"001000110",
  57460=>"100111110",
  57461=>"110001100",
  57462=>"000001000",
  57463=>"000111110",
  57464=>"011110110",
  57465=>"111111000",
  57466=>"000111101",
  57467=>"001010001",
  57468=>"001010110",
  57469=>"101110011",
  57470=>"010110000",
  57471=>"101100100",
  57472=>"101110010",
  57473=>"011010111",
  57474=>"000010011",
  57475=>"000000010",
  57476=>"101101111",
  57477=>"110010010",
  57478=>"000100111",
  57479=>"100100101",
  57480=>"011100111",
  57481=>"111111101",
  57482=>"010110011",
  57483=>"111111000",
  57484=>"001011000",
  57485=>"001011100",
  57486=>"110100111",
  57487=>"010001001",
  57488=>"011100101",
  57489=>"010111011",
  57490=>"011010101",
  57491=>"011111101",
  57492=>"000111001",
  57493=>"010001101",
  57494=>"010001001",
  57495=>"011100111",
  57496=>"111111101",
  57497=>"111011111",
  57498=>"011101101",
  57499=>"101101011",
  57500=>"110000010",
  57501=>"111111001",
  57502=>"110100100",
  57503=>"110001110",
  57504=>"000000000",
  57505=>"011000001",
  57506=>"000111100",
  57507=>"110110101",
  57508=>"011010111",
  57509=>"111010100",
  57510=>"100111011",
  57511=>"001111100",
  57512=>"101101010",
  57513=>"101111101",
  57514=>"111110111",
  57515=>"000000011",
  57516=>"110000100",
  57517=>"101100011",
  57518=>"011110110",
  57519=>"011111110",
  57520=>"000001111",
  57521=>"010001110",
  57522=>"110010110",
  57523=>"110111001",
  57524=>"001101001",
  57525=>"000010010",
  57526=>"010011010",
  57527=>"110111111",
  57528=>"010100001",
  57529=>"111001111",
  57530=>"101011011",
  57531=>"000110100",
  57532=>"111110001",
  57533=>"111111111",
  57534=>"101001101",
  57535=>"010110000",
  57536=>"100100101",
  57537=>"010011111",
  57538=>"111011000",
  57539=>"111111010",
  57540=>"001110011",
  57541=>"101110110",
  57542=>"001010110",
  57543=>"011111110",
  57544=>"111110011",
  57545=>"001101111",
  57546=>"000011101",
  57547=>"111001010",
  57548=>"001101011",
  57549=>"010011001",
  57550=>"000111000",
  57551=>"001101100",
  57552=>"010010100",
  57553=>"100101001",
  57554=>"100111110",
  57555=>"100000110",
  57556=>"100110011",
  57557=>"110111000",
  57558=>"000100111",
  57559=>"100111111",
  57560=>"010001000",
  57561=>"101010001",
  57562=>"100101001",
  57563=>"100100010",
  57564=>"010001001",
  57565=>"100010100",
  57566=>"110000001",
  57567=>"000110111",
  57568=>"110111010",
  57569=>"111000001",
  57570=>"010000111",
  57571=>"110011010",
  57572=>"100101100",
  57573=>"010100100",
  57574=>"010101010",
  57575=>"000111111",
  57576=>"110111100",
  57577=>"100011100",
  57578=>"001111100",
  57579=>"010001010",
  57580=>"000001010",
  57581=>"111111001",
  57582=>"001111000",
  57583=>"111010101",
  57584=>"010101111",
  57585=>"100001001",
  57586=>"011000000",
  57587=>"000111000",
  57588=>"001110111",
  57589=>"010000001",
  57590=>"111110111",
  57591=>"101001001",
  57592=>"100110110",
  57593=>"111000011",
  57594=>"000010001",
  57595=>"001000101",
  57596=>"111101011",
  57597=>"010001111",
  57598=>"000001001",
  57599=>"001111000",
  57600=>"101111001",
  57601=>"111001100",
  57602=>"011011111",
  57603=>"101100010",
  57604=>"110110100",
  57605=>"011110110",
  57606=>"111001000",
  57607=>"110111011",
  57608=>"011000010",
  57609=>"001101010",
  57610=>"001010010",
  57611=>"010000110",
  57612=>"010000001",
  57613=>"010000100",
  57614=>"111101010",
  57615=>"000110000",
  57616=>"111111111",
  57617=>"110000001",
  57618=>"111000100",
  57619=>"000000011",
  57620=>"111001111",
  57621=>"110111111",
  57622=>"000001111",
  57623=>"010111100",
  57624=>"111101100",
  57625=>"101000010",
  57626=>"110010011",
  57627=>"001001011",
  57628=>"100010101",
  57629=>"100001111",
  57630=>"110100000",
  57631=>"111110110",
  57632=>"000001010",
  57633=>"100000110",
  57634=>"111110100",
  57635=>"001111101",
  57636=>"111000000",
  57637=>"000101011",
  57638=>"011000100",
  57639=>"010000011",
  57640=>"100011011",
  57641=>"001101011",
  57642=>"110111101",
  57643=>"100100000",
  57644=>"111110111",
  57645=>"010101000",
  57646=>"011000101",
  57647=>"101000000",
  57648=>"011011100",
  57649=>"001000101",
  57650=>"110111111",
  57651=>"011000000",
  57652=>"011101011",
  57653=>"001010111",
  57654=>"100001011",
  57655=>"110110001",
  57656=>"011111000",
  57657=>"110010001",
  57658=>"000010110",
  57659=>"110001110",
  57660=>"101010110",
  57661=>"111001101",
  57662=>"100100010",
  57663=>"111001010",
  57664=>"100110010",
  57665=>"001111111",
  57666=>"111010100",
  57667=>"101011111",
  57668=>"100001101",
  57669=>"000000101",
  57670=>"000001011",
  57671=>"000111010",
  57672=>"010100011",
  57673=>"000011101",
  57674=>"000101000",
  57675=>"110001000",
  57676=>"111000010",
  57677=>"100010101",
  57678=>"001101100",
  57679=>"111010101",
  57680=>"000011000",
  57681=>"100011101",
  57682=>"011010110",
  57683=>"010100000",
  57684=>"011110000",
  57685=>"110000111",
  57686=>"001000101",
  57687=>"001010110",
  57688=>"010000011",
  57689=>"011000111",
  57690=>"011111111",
  57691=>"111010101",
  57692=>"100011001",
  57693=>"011000101",
  57694=>"111111111",
  57695=>"101111010",
  57696=>"110100001",
  57697=>"100001011",
  57698=>"100000010",
  57699=>"011111000",
  57700=>"111001001",
  57701=>"011011110",
  57702=>"101111100",
  57703=>"001111000",
  57704=>"111100101",
  57705=>"010101000",
  57706=>"010111000",
  57707=>"000100001",
  57708=>"011101010",
  57709=>"000000111",
  57710=>"101000100",
  57711=>"000110110",
  57712=>"001001111",
  57713=>"001101101",
  57714=>"010100111",
  57715=>"110100111",
  57716=>"100101101",
  57717=>"111001111",
  57718=>"111111111",
  57719=>"000100010",
  57720=>"010011011",
  57721=>"100100101",
  57722=>"000100101",
  57723=>"001100000",
  57724=>"111111110",
  57725=>"000000101",
  57726=>"010101011",
  57727=>"100110110",
  57728=>"001011100",
  57729=>"110011010",
  57730=>"011111101",
  57731=>"100101010",
  57732=>"001000110",
  57733=>"000001000",
  57734=>"111101100",
  57735=>"111011100",
  57736=>"011110000",
  57737=>"100000110",
  57738=>"110101011",
  57739=>"100001001",
  57740=>"001010100",
  57741=>"111000010",
  57742=>"000100001",
  57743=>"001101111",
  57744=>"111110110",
  57745=>"001000000",
  57746=>"001011110",
  57747=>"001100101",
  57748=>"101101100",
  57749=>"011111110",
  57750=>"010011011",
  57751=>"101000000",
  57752=>"001010100",
  57753=>"010101011",
  57754=>"111001010",
  57755=>"000101000",
  57756=>"101101101",
  57757=>"111100011",
  57758=>"101111000",
  57759=>"000101010",
  57760=>"011100000",
  57761=>"110000011",
  57762=>"111000011",
  57763=>"101100001",
  57764=>"000101101",
  57765=>"101100001",
  57766=>"110101010",
  57767=>"000110000",
  57768=>"101100010",
  57769=>"101001110",
  57770=>"010000111",
  57771=>"010011101",
  57772=>"011100010",
  57773=>"110001110",
  57774=>"010000101",
  57775=>"001000001",
  57776=>"111011000",
  57777=>"010001011",
  57778=>"110001111",
  57779=>"010110110",
  57780=>"010000001",
  57781=>"011000011",
  57782=>"100000001",
  57783=>"101110000",
  57784=>"011001010",
  57785=>"000011000",
  57786=>"001000111",
  57787=>"100010001",
  57788=>"101011011",
  57789=>"100111110",
  57790=>"100100010",
  57791=>"010110110",
  57792=>"010010111",
  57793=>"101100011",
  57794=>"111100011",
  57795=>"100010000",
  57796=>"110100011",
  57797=>"110000000",
  57798=>"111000101",
  57799=>"111011111",
  57800=>"101000011",
  57801=>"101111011",
  57802=>"010011000",
  57803=>"111110101",
  57804=>"000100111",
  57805=>"001000110",
  57806=>"000011011",
  57807=>"001000000",
  57808=>"010010000",
  57809=>"011000111",
  57810=>"111001100",
  57811=>"000000010",
  57812=>"100100100",
  57813=>"111101000",
  57814=>"000001110",
  57815=>"101101001",
  57816=>"010111110",
  57817=>"010000100",
  57818=>"100110111",
  57819=>"011011011",
  57820=>"000010100",
  57821=>"001111111",
  57822=>"101110110",
  57823=>"001000111",
  57824=>"011011011",
  57825=>"001100111",
  57826=>"111000011",
  57827=>"000100110",
  57828=>"101101000",
  57829=>"111000001",
  57830=>"011010110",
  57831=>"100000001",
  57832=>"111101110",
  57833=>"001010110",
  57834=>"000010000",
  57835=>"100110000",
  57836=>"100100111",
  57837=>"110010000",
  57838=>"101011101",
  57839=>"110100001",
  57840=>"010011100",
  57841=>"000001001",
  57842=>"001010011",
  57843=>"011101111",
  57844=>"101011100",
  57845=>"001111011",
  57846=>"111000001",
  57847=>"111011110",
  57848=>"101110101",
  57849=>"111001111",
  57850=>"011111001",
  57851=>"010111010",
  57852=>"000011100",
  57853=>"111100000",
  57854=>"000000101",
  57855=>"011111111",
  57856=>"001011101",
  57857=>"101100111",
  57858=>"110101000",
  57859=>"001001111",
  57860=>"111100110",
  57861=>"100100100",
  57862=>"110000101",
  57863=>"101110110",
  57864=>"111110111",
  57865=>"101001000",
  57866=>"111001100",
  57867=>"111001100",
  57868=>"011111110",
  57869=>"110100100",
  57870=>"010001000",
  57871=>"111110001",
  57872=>"001010100",
  57873=>"101111100",
  57874=>"111101010",
  57875=>"101101011",
  57876=>"000000011",
  57877=>"100111100",
  57878=>"011010110",
  57879=>"111001011",
  57880=>"101111111",
  57881=>"111001011",
  57882=>"110110000",
  57883=>"000010100",
  57884=>"110001110",
  57885=>"101010010",
  57886=>"100101110",
  57887=>"010010010",
  57888=>"010001010",
  57889=>"001111010",
  57890=>"111110001",
  57891=>"010111100",
  57892=>"001110111",
  57893=>"011110111",
  57894=>"110101100",
  57895=>"101001101",
  57896=>"010010101",
  57897=>"100100100",
  57898=>"010110011",
  57899=>"110011111",
  57900=>"100101000",
  57901=>"010100001",
  57902=>"111100110",
  57903=>"110001110",
  57904=>"010000111",
  57905=>"111111000",
  57906=>"111101100",
  57907=>"101111000",
  57908=>"011101011",
  57909=>"000010001",
  57910=>"000011010",
  57911=>"010010001",
  57912=>"011101010",
  57913=>"111011001",
  57914=>"101000110",
  57915=>"011011100",
  57916=>"111011110",
  57917=>"001001000",
  57918=>"111001101",
  57919=>"111100110",
  57920=>"000111001",
  57921=>"011110111",
  57922=>"011111111",
  57923=>"101110001",
  57924=>"110001001",
  57925=>"010000101",
  57926=>"000000000",
  57927=>"111000111",
  57928=>"011101010",
  57929=>"111001111",
  57930=>"111011111",
  57931=>"111000001",
  57932=>"000010100",
  57933=>"111011011",
  57934=>"100100110",
  57935=>"110111111",
  57936=>"001100010",
  57937=>"010110111",
  57938=>"000000110",
  57939=>"100101001",
  57940=>"100111101",
  57941=>"000100001",
  57942=>"000011100",
  57943=>"011101011",
  57944=>"111100101",
  57945=>"001011111",
  57946=>"100101001",
  57947=>"001000011",
  57948=>"111100101",
  57949=>"000001001",
  57950=>"110100000",
  57951=>"110111001",
  57952=>"100110111",
  57953=>"000000011",
  57954=>"001101110",
  57955=>"101000011",
  57956=>"001000000",
  57957=>"010001001",
  57958=>"011110010",
  57959=>"111111111",
  57960=>"010101010",
  57961=>"100000011",
  57962=>"000011000",
  57963=>"011111010",
  57964=>"101000000",
  57965=>"010101101",
  57966=>"001001000",
  57967=>"010001100",
  57968=>"011010110",
  57969=>"000100011",
  57970=>"000101100",
  57971=>"101001111",
  57972=>"100011000",
  57973=>"110110000",
  57974=>"111001010",
  57975=>"111011111",
  57976=>"010010001",
  57977=>"101001110",
  57978=>"111000000",
  57979=>"010111000",
  57980=>"011101000",
  57981=>"011001010",
  57982=>"000010011",
  57983=>"000011111",
  57984=>"100001010",
  57985=>"110100011",
  57986=>"110011000",
  57987=>"010110101",
  57988=>"101001000",
  57989=>"100110100",
  57990=>"010010001",
  57991=>"101101000",
  57992=>"110011000",
  57993=>"101000001",
  57994=>"000111101",
  57995=>"100100100",
  57996=>"111111010",
  57997=>"001001000",
  57998=>"111110110",
  57999=>"111001011",
  58000=>"001001011",
  58001=>"111011101",
  58002=>"100011101",
  58003=>"000001100",
  58004=>"001101100",
  58005=>"101001101",
  58006=>"011000101",
  58007=>"011110110",
  58008=>"010100111",
  58009=>"000111111",
  58010=>"001011100",
  58011=>"000011010",
  58012=>"000101011",
  58013=>"100001000",
  58014=>"000011110",
  58015=>"101101101",
  58016=>"001110011",
  58017=>"111110101",
  58018=>"010000101",
  58019=>"101001001",
  58020=>"000101000",
  58021=>"110000100",
  58022=>"111101100",
  58023=>"000011000",
  58024=>"110110010",
  58025=>"011000100",
  58026=>"011000001",
  58027=>"001000111",
  58028=>"011011000",
  58029=>"010101110",
  58030=>"100100111",
  58031=>"010111111",
  58032=>"101111111",
  58033=>"101101111",
  58034=>"111110101",
  58035=>"111001010",
  58036=>"111100010",
  58037=>"001000011",
  58038=>"010110101",
  58039=>"110111110",
  58040=>"100111101",
  58041=>"011011010",
  58042=>"111010010",
  58043=>"110110100",
  58044=>"111111000",
  58045=>"110111101",
  58046=>"111101010",
  58047=>"111000100",
  58048=>"010000110",
  58049=>"000010110",
  58050=>"000000101",
  58051=>"011001011",
  58052=>"111000110",
  58053=>"000110100",
  58054=>"100100110",
  58055=>"010001100",
  58056=>"011010000",
  58057=>"010100001",
  58058=>"010001100",
  58059=>"101101010",
  58060=>"000110111",
  58061=>"011011010",
  58062=>"001110000",
  58063=>"111100111",
  58064=>"110111101",
  58065=>"000010100",
  58066=>"111010000",
  58067=>"100011001",
  58068=>"011110000",
  58069=>"111110000",
  58070=>"101001001",
  58071=>"110111111",
  58072=>"011001001",
  58073=>"001011010",
  58074=>"000001000",
  58075=>"000101110",
  58076=>"010011111",
  58077=>"011011100",
  58078=>"100001100",
  58079=>"100110011",
  58080=>"100010010",
  58081=>"010000110",
  58082=>"101111100",
  58083=>"101100110",
  58084=>"011010001",
  58085=>"000000000",
  58086=>"101001110",
  58087=>"111111101",
  58088=>"111110101",
  58089=>"111110110",
  58090=>"100101001",
  58091=>"010010000",
  58092=>"000100010",
  58093=>"011110111",
  58094=>"101010000",
  58095=>"000000001",
  58096=>"001001111",
  58097=>"110001110",
  58098=>"001011001",
  58099=>"111110100",
  58100=>"100011001",
  58101=>"101001100",
  58102=>"110010010",
  58103=>"000010000",
  58104=>"111001101",
  58105=>"110111011",
  58106=>"100000110",
  58107=>"100011000",
  58108=>"110111100",
  58109=>"010100001",
  58110=>"111110000",
  58111=>"000100111",
  58112=>"000001100",
  58113=>"011001101",
  58114=>"001100100",
  58115=>"000000001",
  58116=>"010100000",
  58117=>"000111101",
  58118=>"101010011",
  58119=>"001001110",
  58120=>"100000000",
  58121=>"110000011",
  58122=>"100010011",
  58123=>"111101000",
  58124=>"110110001",
  58125=>"001011100",
  58126=>"000000101",
  58127=>"110001101",
  58128=>"101110010",
  58129=>"010111011",
  58130=>"010001001",
  58131=>"011111101",
  58132=>"111010110",
  58133=>"010001000",
  58134=>"110000000",
  58135=>"111111010",
  58136=>"010011101",
  58137=>"100110001",
  58138=>"101101110",
  58139=>"110001011",
  58140=>"001000010",
  58141=>"100111011",
  58142=>"101110000",
  58143=>"000111100",
  58144=>"110110011",
  58145=>"100110110",
  58146=>"111110110",
  58147=>"110000000",
  58148=>"111111001",
  58149=>"001011001",
  58150=>"101000001",
  58151=>"111000101",
  58152=>"101011111",
  58153=>"111011001",
  58154=>"000111100",
  58155=>"110111010",
  58156=>"000101110",
  58157=>"000100100",
  58158=>"100100011",
  58159=>"110001010",
  58160=>"011110011",
  58161=>"101110110",
  58162=>"101001101",
  58163=>"011111110",
  58164=>"011000010",
  58165=>"000000011",
  58166=>"101111110",
  58167=>"000001011",
  58168=>"111110000",
  58169=>"010000000",
  58170=>"111111000",
  58171=>"110101001",
  58172=>"100110101",
  58173=>"000001001",
  58174=>"010111100",
  58175=>"111000100",
  58176=>"110100010",
  58177=>"001111000",
  58178=>"101010101",
  58179=>"101100001",
  58180=>"000000001",
  58181=>"110110010",
  58182=>"000011010",
  58183=>"010001000",
  58184=>"111100111",
  58185=>"111111011",
  58186=>"010100100",
  58187=>"001010000",
  58188=>"100100101",
  58189=>"001000101",
  58190=>"010100010",
  58191=>"101000000",
  58192=>"010000001",
  58193=>"111101001",
  58194=>"010101100",
  58195=>"000110010",
  58196=>"110010000",
  58197=>"101110011",
  58198=>"101110010",
  58199=>"000100010",
  58200=>"000111010",
  58201=>"000001000",
  58202=>"100110101",
  58203=>"011011111",
  58204=>"000010110",
  58205=>"001100000",
  58206=>"011000010",
  58207=>"111111000",
  58208=>"011101110",
  58209=>"110000101",
  58210=>"010000000",
  58211=>"100000100",
  58212=>"011011111",
  58213=>"110011100",
  58214=>"000001100",
  58215=>"100000010",
  58216=>"101010100",
  58217=>"000101111",
  58218=>"000001111",
  58219=>"111101110",
  58220=>"000111000",
  58221=>"111000111",
  58222=>"001011011",
  58223=>"111100000",
  58224=>"001001111",
  58225=>"001011010",
  58226=>"100111110",
  58227=>"100001111",
  58228=>"000001001",
  58229=>"110010001",
  58230=>"010010011",
  58231=>"110111001",
  58232=>"111000000",
  58233=>"010010001",
  58234=>"111000100",
  58235=>"100001001",
  58236=>"001010011",
  58237=>"001010101",
  58238=>"011010100",
  58239=>"101111111",
  58240=>"000100110",
  58241=>"000100001",
  58242=>"100110111",
  58243=>"111011110",
  58244=>"011001101",
  58245=>"010000010",
  58246=>"011010110",
  58247=>"011011101",
  58248=>"110011010",
  58249=>"110101100",
  58250=>"000001000",
  58251=>"111101111",
  58252=>"010100101",
  58253=>"111011100",
  58254=>"001000111",
  58255=>"001110011",
  58256=>"001110110",
  58257=>"100101101",
  58258=>"000100011",
  58259=>"111111001",
  58260=>"000010100",
  58261=>"000000101",
  58262=>"010101100",
  58263=>"110000110",
  58264=>"011110110",
  58265=>"111110111",
  58266=>"000100101",
  58267=>"000000011",
  58268=>"010110001",
  58269=>"001000000",
  58270=>"101000100",
  58271=>"000011110",
  58272=>"101111010",
  58273=>"101101110",
  58274=>"110001000",
  58275=>"010110001",
  58276=>"001001110",
  58277=>"010111011",
  58278=>"110001110",
  58279=>"101110010",
  58280=>"010001000",
  58281=>"111001101",
  58282=>"011110001",
  58283=>"101101110",
  58284=>"101111010",
  58285=>"000011000",
  58286=>"010001001",
  58287=>"111001110",
  58288=>"000110110",
  58289=>"010010001",
  58290=>"001000101",
  58291=>"100001010",
  58292=>"101100000",
  58293=>"101001101",
  58294=>"000100101",
  58295=>"010010011",
  58296=>"010100111",
  58297=>"100111111",
  58298=>"101100111",
  58299=>"010101010",
  58300=>"111011000",
  58301=>"101001110",
  58302=>"100010010",
  58303=>"000100000",
  58304=>"000100101",
  58305=>"110101010",
  58306=>"010110111",
  58307=>"011000111",
  58308=>"011101100",
  58309=>"100101011",
  58310=>"010010000",
  58311=>"010011110",
  58312=>"100110100",
  58313=>"011110100",
  58314=>"001010010",
  58315=>"111111101",
  58316=>"010101001",
  58317=>"001000001",
  58318=>"111101010",
  58319=>"111010100",
  58320=>"011011011",
  58321=>"010111111",
  58322=>"110101011",
  58323=>"000011110",
  58324=>"000000000",
  58325=>"111001110",
  58326=>"100010010",
  58327=>"111000000",
  58328=>"010011000",
  58329=>"100010011",
  58330=>"101101110",
  58331=>"000100110",
  58332=>"000100111",
  58333=>"101111000",
  58334=>"111101011",
  58335=>"000001110",
  58336=>"010010101",
  58337=>"100100000",
  58338=>"000011000",
  58339=>"000001000",
  58340=>"100111010",
  58341=>"101101101",
  58342=>"111110010",
  58343=>"100000100",
  58344=>"001101110",
  58345=>"111000011",
  58346=>"011010101",
  58347=>"110111100",
  58348=>"101100000",
  58349=>"000100000",
  58350=>"100110101",
  58351=>"000011011",
  58352=>"011100001",
  58353=>"111101011",
  58354=>"010010011",
  58355=>"110000001",
  58356=>"111011011",
  58357=>"001110101",
  58358=>"101000111",
  58359=>"001111101",
  58360=>"101000001",
  58361=>"001010111",
  58362=>"000111100",
  58363=>"000010101",
  58364=>"000000010",
  58365=>"111010111",
  58366=>"110111101",
  58367=>"011110101",
  58368=>"010100110",
  58369=>"110100010",
  58370=>"110010001",
  58371=>"111000001",
  58372=>"011111101",
  58373=>"001100010",
  58374=>"001100011",
  58375=>"101101000",
  58376=>"011001100",
  58377=>"001001000",
  58378=>"001000110",
  58379=>"001100001",
  58380=>"111100110",
  58381=>"010001001",
  58382=>"101111001",
  58383=>"100001000",
  58384=>"001011101",
  58385=>"110101101",
  58386=>"011100110",
  58387=>"111100110",
  58388=>"000000101",
  58389=>"011111001",
  58390=>"101000000",
  58391=>"000000000",
  58392=>"011100010",
  58393=>"000000000",
  58394=>"111000101",
  58395=>"001011001",
  58396=>"101100100",
  58397=>"110011000",
  58398=>"011101110",
  58399=>"011000100",
  58400=>"110101011",
  58401=>"001111001",
  58402=>"010100101",
  58403=>"101010011",
  58404=>"001101110",
  58405=>"100000011",
  58406=>"101011111",
  58407=>"001001100",
  58408=>"100110000",
  58409=>"010100001",
  58410=>"101001100",
  58411=>"100000010",
  58412=>"011100111",
  58413=>"000010101",
  58414=>"101111000",
  58415=>"101011001",
  58416=>"000010111",
  58417=>"011000000",
  58418=>"000000001",
  58419=>"011101001",
  58420=>"000000001",
  58421=>"011000010",
  58422=>"101100010",
  58423=>"011111100",
  58424=>"010100111",
  58425=>"100010010",
  58426=>"000011101",
  58427=>"110111111",
  58428=>"100000010",
  58429=>"011100001",
  58430=>"000101100",
  58431=>"101001100",
  58432=>"000010111",
  58433=>"010010010",
  58434=>"010011001",
  58435=>"010000100",
  58436=>"101110110",
  58437=>"000100101",
  58438=>"111100111",
  58439=>"001000111",
  58440=>"000111111",
  58441=>"010111010",
  58442=>"111000000",
  58443=>"001000001",
  58444=>"001101110",
  58445=>"000100110",
  58446=>"011101000",
  58447=>"111110000",
  58448=>"100111101",
  58449=>"000011101",
  58450=>"110111110",
  58451=>"101011000",
  58452=>"100111110",
  58453=>"001011010",
  58454=>"110000110",
  58455=>"000101110",
  58456=>"101010010",
  58457=>"100111100",
  58458=>"110000010",
  58459=>"001000001",
  58460=>"001101111",
  58461=>"111111110",
  58462=>"101001001",
  58463=>"000011101",
  58464=>"110000001",
  58465=>"001001000",
  58466=>"100111101",
  58467=>"101111000",
  58468=>"010100111",
  58469=>"111110000",
  58470=>"100010010",
  58471=>"011011111",
  58472=>"000111000",
  58473=>"011111010",
  58474=>"101000110",
  58475=>"000001010",
  58476=>"111000101",
  58477=>"101011010",
  58478=>"001011101",
  58479=>"000000011",
  58480=>"011101011",
  58481=>"100101111",
  58482=>"001010111",
  58483=>"110111110",
  58484=>"000100011",
  58485=>"001110110",
  58486=>"011100111",
  58487=>"101100100",
  58488=>"000011100",
  58489=>"100000010",
  58490=>"010000000",
  58491=>"000101010",
  58492=>"101001000",
  58493=>"010001010",
  58494=>"100000001",
  58495=>"010110001",
  58496=>"001011000",
  58497=>"011000001",
  58498=>"010100010",
  58499=>"100000000",
  58500=>"000010011",
  58501=>"000001100",
  58502=>"110100110",
  58503=>"000101010",
  58504=>"010100101",
  58505=>"100010010",
  58506=>"010100011",
  58507=>"100110110",
  58508=>"011111011",
  58509=>"001010000",
  58510=>"110010000",
  58511=>"000101101",
  58512=>"100111010",
  58513=>"101111011",
  58514=>"101110000",
  58515=>"101111001",
  58516=>"001111010",
  58517=>"010101100",
  58518=>"101001110",
  58519=>"111110010",
  58520=>"111000100",
  58521=>"001011100",
  58522=>"011011100",
  58523=>"111111111",
  58524=>"110010111",
  58525=>"100110111",
  58526=>"110111101",
  58527=>"010010011",
  58528=>"000000000",
  58529=>"000111010",
  58530=>"001100000",
  58531=>"001011000",
  58532=>"111011011",
  58533=>"010011111",
  58534=>"010100001",
  58535=>"010011111",
  58536=>"100101000",
  58537=>"100011101",
  58538=>"010011000",
  58539=>"000010010",
  58540=>"111000010",
  58541=>"000000001",
  58542=>"010100100",
  58543=>"001100100",
  58544=>"100010111",
  58545=>"011001011",
  58546=>"110100111",
  58547=>"100000111",
  58548=>"010100110",
  58549=>"000001011",
  58550=>"101000011",
  58551=>"000110000",
  58552=>"010001001",
  58553=>"010000100",
  58554=>"101010011",
  58555=>"011101010",
  58556=>"101110010",
  58557=>"001100111",
  58558=>"000110111",
  58559=>"111110001",
  58560=>"111000101",
  58561=>"000100000",
  58562=>"100000011",
  58563=>"000000101",
  58564=>"001101000",
  58565=>"101101001",
  58566=>"001010010",
  58567=>"010110110",
  58568=>"111010100",
  58569=>"100001000",
  58570=>"011001001",
  58571=>"010000011",
  58572=>"001011100",
  58573=>"111100111",
  58574=>"101100111",
  58575=>"011111101",
  58576=>"100101001",
  58577=>"000110101",
  58578=>"110110010",
  58579=>"000111010",
  58580=>"100100100",
  58581=>"010110010",
  58582=>"101100000",
  58583=>"000001010",
  58584=>"010100110",
  58585=>"001011000",
  58586=>"000100111",
  58587=>"010100000",
  58588=>"010100100",
  58589=>"011010111",
  58590=>"011000111",
  58591=>"101011111",
  58592=>"000011000",
  58593=>"010000100",
  58594=>"010110110",
  58595=>"000011110",
  58596=>"101110100",
  58597=>"101010000",
  58598=>"101000010",
  58599=>"101101111",
  58600=>"001100001",
  58601=>"101001000",
  58602=>"010010101",
  58603=>"111010010",
  58604=>"000110100",
  58605=>"101010000",
  58606=>"110000001",
  58607=>"010110010",
  58608=>"110010010",
  58609=>"100000110",
  58610=>"100111111",
  58611=>"011100111",
  58612=>"011110010",
  58613=>"011100101",
  58614=>"100111000",
  58615=>"001011111",
  58616=>"100011010",
  58617=>"011101010",
  58618=>"010001000",
  58619=>"001100000",
  58620=>"010010111",
  58621=>"011111001",
  58622=>"010111001",
  58623=>"100001011",
  58624=>"010010100",
  58625=>"110000111",
  58626=>"100101100",
  58627=>"000110011",
  58628=>"011001100",
  58629=>"100110101",
  58630=>"111010010",
  58631=>"001101001",
  58632=>"010010000",
  58633=>"100001101",
  58634=>"011011000",
  58635=>"100100110",
  58636=>"000010000",
  58637=>"001000101",
  58638=>"100000011",
  58639=>"100011100",
  58640=>"110001101",
  58641=>"000111011",
  58642=>"001100000",
  58643=>"100001111",
  58644=>"000100001",
  58645=>"111110110",
  58646=>"111111111",
  58647=>"110101100",
  58648=>"100101110",
  58649=>"011111000",
  58650=>"000001110",
  58651=>"111111111",
  58652=>"010000000",
  58653=>"001111000",
  58654=>"100011001",
  58655=>"010000110",
  58656=>"001001110",
  58657=>"001101100",
  58658=>"000010001",
  58659=>"010110101",
  58660=>"111001101",
  58661=>"011101011",
  58662=>"110110010",
  58663=>"100000101",
  58664=>"111100001",
  58665=>"110011111",
  58666=>"100111101",
  58667=>"101101010",
  58668=>"100001001",
  58669=>"111011111",
  58670=>"111001011",
  58671=>"110101001",
  58672=>"111101000",
  58673=>"101110011",
  58674=>"111111001",
  58675=>"000101110",
  58676=>"001011000",
  58677=>"000010111",
  58678=>"011000111",
  58679=>"010000000",
  58680=>"000011110",
  58681=>"001111111",
  58682=>"101010101",
  58683=>"011011101",
  58684=>"100000011",
  58685=>"011111101",
  58686=>"011000011",
  58687=>"000110100",
  58688=>"000001000",
  58689=>"110100000",
  58690=>"111100101",
  58691=>"111000110",
  58692=>"111111001",
  58693=>"111001001",
  58694=>"010011001",
  58695=>"011100000",
  58696=>"100001000",
  58697=>"110110111",
  58698=>"111101010",
  58699=>"110101011",
  58700=>"000001110",
  58701=>"110100101",
  58702=>"000000111",
  58703=>"011011101",
  58704=>"101001110",
  58705=>"000111101",
  58706=>"011101100",
  58707=>"000011111",
  58708=>"010011111",
  58709=>"011111011",
  58710=>"000110000",
  58711=>"011001111",
  58712=>"100001001",
  58713=>"111110111",
  58714=>"001011010",
  58715=>"111110100",
  58716=>"101001011",
  58717=>"010011010",
  58718=>"011010001",
  58719=>"001110001",
  58720=>"001010010",
  58721=>"010110001",
  58722=>"110110101",
  58723=>"000010010",
  58724=>"111110110",
  58725=>"101111110",
  58726=>"101100110",
  58727=>"000010100",
  58728=>"110010100",
  58729=>"000000110",
  58730=>"011011000",
  58731=>"100010010",
  58732=>"010001010",
  58733=>"000101011",
  58734=>"111001101",
  58735=>"010110100",
  58736=>"100110001",
  58737=>"111111110",
  58738=>"001010100",
  58739=>"100011010",
  58740=>"111110001",
  58741=>"110101000",
  58742=>"101111001",
  58743=>"100001000",
  58744=>"111000001",
  58745=>"010110110",
  58746=>"010110000",
  58747=>"101100001",
  58748=>"110001010",
  58749=>"000110111",
  58750=>"010110111",
  58751=>"100110000",
  58752=>"000001011",
  58753=>"000000010",
  58754=>"111001011",
  58755=>"111110000",
  58756=>"100011111",
  58757=>"001000011",
  58758=>"001110110",
  58759=>"110001111",
  58760=>"101001100",
  58761=>"011010111",
  58762=>"000001010",
  58763=>"010001001",
  58764=>"000011011",
  58765=>"010110111",
  58766=>"010011101",
  58767=>"000010111",
  58768=>"101000101",
  58769=>"001011000",
  58770=>"000101010",
  58771=>"111001000",
  58772=>"000000110",
  58773=>"010110010",
  58774=>"101111111",
  58775=>"110001100",
  58776=>"001011011",
  58777=>"101101100",
  58778=>"001001001",
  58779=>"000000000",
  58780=>"011111001",
  58781=>"000010011",
  58782=>"000100001",
  58783=>"100011001",
  58784=>"111100111",
  58785=>"011111111",
  58786=>"000111100",
  58787=>"100010010",
  58788=>"001011100",
  58789=>"001011110",
  58790=>"100000100",
  58791=>"100110101",
  58792=>"010111010",
  58793=>"111110100",
  58794=>"010101100",
  58795=>"001101000",
  58796=>"100011100",
  58797=>"011000110",
  58798=>"011011110",
  58799=>"010111100",
  58800=>"000000000",
  58801=>"100011011",
  58802=>"100110000",
  58803=>"100110111",
  58804=>"111011010",
  58805=>"010010100",
  58806=>"111101110",
  58807=>"010111010",
  58808=>"100001010",
  58809=>"001001010",
  58810=>"000111000",
  58811=>"110011010",
  58812=>"011100111",
  58813=>"010110111",
  58814=>"010100011",
  58815=>"110100110",
  58816=>"000101000",
  58817=>"001010001",
  58818=>"110110100",
  58819=>"100000000",
  58820=>"000101100",
  58821=>"111101100",
  58822=>"010111100",
  58823=>"101000000",
  58824=>"111001000",
  58825=>"000000110",
  58826=>"100000100",
  58827=>"010110101",
  58828=>"001010101",
  58829=>"110111110",
  58830=>"111101111",
  58831=>"111011000",
  58832=>"010100000",
  58833=>"001111101",
  58834=>"001110100",
  58835=>"010000000",
  58836=>"110110100",
  58837=>"010000010",
  58838=>"001101010",
  58839=>"001110010",
  58840=>"111101101",
  58841=>"011010000",
  58842=>"100010100",
  58843=>"001111001",
  58844=>"001010100",
  58845=>"100001010",
  58846=>"001111101",
  58847=>"000110110",
  58848=>"011001101",
  58849=>"010001110",
  58850=>"011010010",
  58851=>"101000101",
  58852=>"010011110",
  58853=>"011101100",
  58854=>"011010010",
  58855=>"101001000",
  58856=>"011000010",
  58857=>"101000011",
  58858=>"000011111",
  58859=>"000010000",
  58860=>"011111000",
  58861=>"000000111",
  58862=>"000010101",
  58863=>"010101011",
  58864=>"101001001",
  58865=>"110111001",
  58866=>"011010000",
  58867=>"011010101",
  58868=>"001001110",
  58869=>"110010110",
  58870=>"001010010",
  58871=>"010101111",
  58872=>"010000101",
  58873=>"101100001",
  58874=>"010111110",
  58875=>"111000111",
  58876=>"100100011",
  58877=>"100011101",
  58878=>"011100110",
  58879=>"111100100",
  58880=>"000010011",
  58881=>"100011010",
  58882=>"000011010",
  58883=>"010000000",
  58884=>"100000100",
  58885=>"110110000",
  58886=>"111001000",
  58887=>"100001011",
  58888=>"000001101",
  58889=>"101100101",
  58890=>"000100010",
  58891=>"111010100",
  58892=>"100000010",
  58893=>"111010110",
  58894=>"011101101",
  58895=>"010010100",
  58896=>"010100101",
  58897=>"110000101",
  58898=>"101001010",
  58899=>"111010011",
  58900=>"000001101",
  58901=>"011100000",
  58902=>"011100010",
  58903=>"110111111",
  58904=>"110001011",
  58905=>"000001011",
  58906=>"101101111",
  58907=>"000010010",
  58908=>"110110101",
  58909=>"101010000",
  58910=>"110111110",
  58911=>"010110101",
  58912=>"000010010",
  58913=>"011110001",
  58914=>"100101010",
  58915=>"010001010",
  58916=>"101111111",
  58917=>"011101100",
  58918=>"100101000",
  58919=>"010000001",
  58920=>"000101000",
  58921=>"010011010",
  58922=>"011010000",
  58923=>"000000001",
  58924=>"001010001",
  58925=>"000010100",
  58926=>"110001010",
  58927=>"010110100",
  58928=>"110111010",
  58929=>"001000101",
  58930=>"010010000",
  58931=>"110111010",
  58932=>"100011111",
  58933=>"001000111",
  58934=>"110000000",
  58935=>"011110000",
  58936=>"111000101",
  58937=>"010000011",
  58938=>"111100001",
  58939=>"101111100",
  58940=>"001101010",
  58941=>"001011110",
  58942=>"100110110",
  58943=>"100100101",
  58944=>"000100100",
  58945=>"100100011",
  58946=>"110101011",
  58947=>"100001101",
  58948=>"010100111",
  58949=>"000011111",
  58950=>"001110000",
  58951=>"111000011",
  58952=>"110010110",
  58953=>"000000001",
  58954=>"111101111",
  58955=>"001101100",
  58956=>"011100000",
  58957=>"010001000",
  58958=>"011111001",
  58959=>"110011100",
  58960=>"110010101",
  58961=>"011011011",
  58962=>"000001001",
  58963=>"000001111",
  58964=>"100011000",
  58965=>"000010110",
  58966=>"010110100",
  58967=>"111010101",
  58968=>"110011000",
  58969=>"100111111",
  58970=>"101111101",
  58971=>"111111110",
  58972=>"111111100",
  58973=>"000001001",
  58974=>"010110101",
  58975=>"011100011",
  58976=>"010001011",
  58977=>"001101100",
  58978=>"011000111",
  58979=>"001000001",
  58980=>"100000000",
  58981=>"000010101",
  58982=>"000001101",
  58983=>"000101110",
  58984=>"000001001",
  58985=>"101101010",
  58986=>"110111111",
  58987=>"011011111",
  58988=>"000011010",
  58989=>"011010100",
  58990=>"011101011",
  58991=>"101100100",
  58992=>"111101110",
  58993=>"101011001",
  58994=>"100001001",
  58995=>"010000110",
  58996=>"001100110",
  58997=>"010001110",
  58998=>"010110011",
  58999=>"011000001",
  59000=>"010000111",
  59001=>"100011011",
  59002=>"110010100",
  59003=>"101011101",
  59004=>"101000001",
  59005=>"011101011",
  59006=>"001000010",
  59007=>"000011101",
  59008=>"011010111",
  59009=>"010110111",
  59010=>"100101011",
  59011=>"101010111",
  59012=>"000000000",
  59013=>"011101000",
  59014=>"101000000",
  59015=>"101100111",
  59016=>"011000000",
  59017=>"100010001",
  59018=>"001011010",
  59019=>"010101110",
  59020=>"111111111",
  59021=>"011100101",
  59022=>"101011001",
  59023=>"100001010",
  59024=>"000110111",
  59025=>"001101100",
  59026=>"011101000",
  59027=>"010101100",
  59028=>"001101001",
  59029=>"010001000",
  59030=>"101001001",
  59031=>"101000110",
  59032=>"000000111",
  59033=>"110111010",
  59034=>"000010100",
  59035=>"110010110",
  59036=>"100000110",
  59037=>"110110010",
  59038=>"111110011",
  59039=>"001100010",
  59040=>"010101111",
  59041=>"011010100",
  59042=>"010111100",
  59043=>"111100000",
  59044=>"100101100",
  59045=>"111010001",
  59046=>"010000100",
  59047=>"100001011",
  59048=>"010100001",
  59049=>"011110011",
  59050=>"010110011",
  59051=>"010100110",
  59052=>"000010010",
  59053=>"101111100",
  59054=>"011111011",
  59055=>"111111001",
  59056=>"000001101",
  59057=>"011000000",
  59058=>"100110001",
  59059=>"011000101",
  59060=>"011011011",
  59061=>"111011011",
  59062=>"000110101",
  59063=>"011100011",
  59064=>"110000110",
  59065=>"111110110",
  59066=>"110110001",
  59067=>"010001110",
  59068=>"011000011",
  59069=>"000001110",
  59070=>"000101110",
  59071=>"001100110",
  59072=>"000111101",
  59073=>"101001110",
  59074=>"001000011",
  59075=>"000011000",
  59076=>"000000000",
  59077=>"010101011",
  59078=>"011000101",
  59079=>"111001110",
  59080=>"101010001",
  59081=>"101011100",
  59082=>"011110111",
  59083=>"000101010",
  59084=>"110011001",
  59085=>"111001110",
  59086=>"000111010",
  59087=>"010011111",
  59088=>"110010010",
  59089=>"011010101",
  59090=>"010110100",
  59091=>"110001111",
  59092=>"010010100",
  59093=>"110100000",
  59094=>"100110101",
  59095=>"100110011",
  59096=>"110111001",
  59097=>"110101101",
  59098=>"010110101",
  59099=>"111101100",
  59100=>"111000001",
  59101=>"101111111",
  59102=>"111110111",
  59103=>"000001000",
  59104=>"111001001",
  59105=>"001001000",
  59106=>"111110100",
  59107=>"110101010",
  59108=>"100101110",
  59109=>"101000010",
  59110=>"111110111",
  59111=>"110110001",
  59112=>"100001011",
  59113=>"101111011",
  59114=>"000100111",
  59115=>"010111000",
  59116=>"000100101",
  59117=>"100010010",
  59118=>"110110111",
  59119=>"001100001",
  59120=>"000011101",
  59121=>"111101001",
  59122=>"001000001",
  59123=>"000010010",
  59124=>"110101001",
  59125=>"010010110",
  59126=>"010000001",
  59127=>"101000001",
  59128=>"000101000",
  59129=>"100110011",
  59130=>"001010101",
  59131=>"000010000",
  59132=>"111000001",
  59133=>"100011010",
  59134=>"100011110",
  59135=>"001000001",
  59136=>"011000001",
  59137=>"011110000",
  59138=>"110010000",
  59139=>"101001001",
  59140=>"010010111",
  59141=>"110010000",
  59142=>"001100010",
  59143=>"110100100",
  59144=>"101100001",
  59145=>"001000000",
  59146=>"011011010",
  59147=>"110110101",
  59148=>"100001000",
  59149=>"111111111",
  59150=>"100101010",
  59151=>"000010100",
  59152=>"111000001",
  59153=>"111110000",
  59154=>"000111010",
  59155=>"111101001",
  59156=>"101001110",
  59157=>"000001111",
  59158=>"011101001",
  59159=>"111100101",
  59160=>"101000110",
  59161=>"000000000",
  59162=>"000000000",
  59163=>"101011110",
  59164=>"011100011",
  59165=>"011100011",
  59166=>"010110010",
  59167=>"001010001",
  59168=>"010001010",
  59169=>"000010001",
  59170=>"110010011",
  59171=>"100111111",
  59172=>"111101110",
  59173=>"001000001",
  59174=>"001011100",
  59175=>"010001100",
  59176=>"010110110",
  59177=>"101101100",
  59178=>"101000011",
  59179=>"000011111",
  59180=>"010001001",
  59181=>"101111000",
  59182=>"000100110",
  59183=>"111011011",
  59184=>"010111001",
  59185=>"101101010",
  59186=>"010001000",
  59187=>"111111101",
  59188=>"101001110",
  59189=>"111000010",
  59190=>"100111100",
  59191=>"100011111",
  59192=>"101101000",
  59193=>"001001111",
  59194=>"000011111",
  59195=>"011001011",
  59196=>"100101010",
  59197=>"101001000",
  59198=>"100100110",
  59199=>"110110110",
  59200=>"011100001",
  59201=>"101011111",
  59202=>"110000001",
  59203=>"010001110",
  59204=>"000011000",
  59205=>"011110110",
  59206=>"000000001",
  59207=>"001001111",
  59208=>"101001111",
  59209=>"010010110",
  59210=>"001100010",
  59211=>"010110110",
  59212=>"100011001",
  59213=>"101001000",
  59214=>"011001010",
  59215=>"110111110",
  59216=>"101000001",
  59217=>"111011001",
  59218=>"110100000",
  59219=>"101010000",
  59220=>"010101111",
  59221=>"110101011",
  59222=>"111111101",
  59223=>"100010011",
  59224=>"100101111",
  59225=>"111011100",
  59226=>"111101011",
  59227=>"010111101",
  59228=>"111111001",
  59229=>"110001101",
  59230=>"100000101",
  59231=>"000010100",
  59232=>"010110001",
  59233=>"011110001",
  59234=>"111010001",
  59235=>"000110100",
  59236=>"010100111",
  59237=>"111100011",
  59238=>"001001010",
  59239=>"001010111",
  59240=>"001101100",
  59241=>"011001010",
  59242=>"010111001",
  59243=>"110111100",
  59244=>"110111001",
  59245=>"000100110",
  59246=>"001010000",
  59247=>"100011010",
  59248=>"000010101",
  59249=>"101000101",
  59250=>"000001001",
  59251=>"110011010",
  59252=>"111100010",
  59253=>"000001000",
  59254=>"000101001",
  59255=>"111111111",
  59256=>"000110111",
  59257=>"001000000",
  59258=>"001000111",
  59259=>"010001000",
  59260=>"111100110",
  59261=>"110001101",
  59262=>"011010110",
  59263=>"110101100",
  59264=>"110000100",
  59265=>"001000110",
  59266=>"111100111",
  59267=>"001000101",
  59268=>"110000001",
  59269=>"011000010",
  59270=>"110111101",
  59271=>"000001011",
  59272=>"100010101",
  59273=>"011100110",
  59274=>"001011011",
  59275=>"011001010",
  59276=>"010111001",
  59277=>"101111110",
  59278=>"110011111",
  59279=>"000000101",
  59280=>"010000011",
  59281=>"110010000",
  59282=>"011010101",
  59283=>"000111001",
  59284=>"100000001",
  59285=>"001001010",
  59286=>"010011010",
  59287=>"000111101",
  59288=>"100110111",
  59289=>"000110111",
  59290=>"000011100",
  59291=>"011110111",
  59292=>"101110101",
  59293=>"010110101",
  59294=>"000001001",
  59295=>"100001010",
  59296=>"010110010",
  59297=>"000111101",
  59298=>"110110101",
  59299=>"101100010",
  59300=>"000101100",
  59301=>"001011011",
  59302=>"111110010",
  59303=>"010110100",
  59304=>"000010010",
  59305=>"001111100",
  59306=>"111100010",
  59307=>"010111011",
  59308=>"100000000",
  59309=>"011100100",
  59310=>"100011011",
  59311=>"011111111",
  59312=>"010000001",
  59313=>"010111011",
  59314=>"111010000",
  59315=>"100000100",
  59316=>"001110010",
  59317=>"010101001",
  59318=>"101100101",
  59319=>"001000001",
  59320=>"010101100",
  59321=>"111001001",
  59322=>"000000011",
  59323=>"110011100",
  59324=>"100000000",
  59325=>"001110001",
  59326=>"010000011",
  59327=>"010001001",
  59328=>"110110010",
  59329=>"101110001",
  59330=>"010011000",
  59331=>"011010000",
  59332=>"110000000",
  59333=>"000000100",
  59334=>"110101000",
  59335=>"010000111",
  59336=>"111100001",
  59337=>"011111101",
  59338=>"010001110",
  59339=>"000101010",
  59340=>"101001010",
  59341=>"111110111",
  59342=>"101000010",
  59343=>"000100001",
  59344=>"000101011",
  59345=>"011010000",
  59346=>"110101110",
  59347=>"011000100",
  59348=>"100000011",
  59349=>"100101100",
  59350=>"111101000",
  59351=>"111000010",
  59352=>"100100101",
  59353=>"111110111",
  59354=>"000010111",
  59355=>"100010111",
  59356=>"101111011",
  59357=>"001100111",
  59358=>"101000111",
  59359=>"001011111",
  59360=>"011111010",
  59361=>"010001101",
  59362=>"100110010",
  59363=>"000100010",
  59364=>"010101110",
  59365=>"001010001",
  59366=>"111101111",
  59367=>"110100001",
  59368=>"111110111",
  59369=>"010100100",
  59370=>"001001110",
  59371=>"100110011",
  59372=>"000001001",
  59373=>"010101110",
  59374=>"001000111",
  59375=>"101001001",
  59376=>"010010000",
  59377=>"011000010",
  59378=>"000010111",
  59379=>"001011010",
  59380=>"000100100",
  59381=>"111111001",
  59382=>"011100111",
  59383=>"001011100",
  59384=>"101010110",
  59385=>"111000011",
  59386=>"110100011",
  59387=>"000000000",
  59388=>"001011111",
  59389=>"011100010",
  59390=>"001000000",
  59391=>"100110110",
  59392=>"111011001",
  59393=>"011010001",
  59394=>"111100101",
  59395=>"011000010",
  59396=>"111000010",
  59397=>"110011000",
  59398=>"010100111",
  59399=>"001110000",
  59400=>"111001100",
  59401=>"100100001",
  59402=>"110000110",
  59403=>"010011011",
  59404=>"110100100",
  59405=>"011001101",
  59406=>"100000000",
  59407=>"000101101",
  59408=>"001100110",
  59409=>"011010010",
  59410=>"110011011",
  59411=>"110110111",
  59412=>"111000111",
  59413=>"111010011",
  59414=>"000110100",
  59415=>"011001011",
  59416=>"001011001",
  59417=>"001001100",
  59418=>"110101100",
  59419=>"101011011",
  59420=>"000110101",
  59421=>"010010010",
  59422=>"111000111",
  59423=>"100101100",
  59424=>"011000000",
  59425=>"101100111",
  59426=>"000000110",
  59427=>"100011000",
  59428=>"000101100",
  59429=>"101010101",
  59430=>"111010001",
  59431=>"101111001",
  59432=>"111100010",
  59433=>"110010001",
  59434=>"010000011",
  59435=>"110011010",
  59436=>"010001101",
  59437=>"011100000",
  59438=>"000010001",
  59439=>"000000101",
  59440=>"110010010",
  59441=>"110000000",
  59442=>"011001101",
  59443=>"101111001",
  59444=>"011101001",
  59445=>"100110000",
  59446=>"000011001",
  59447=>"010011111",
  59448=>"011010000",
  59449=>"101101010",
  59450=>"000101011",
  59451=>"111010001",
  59452=>"001111000",
  59453=>"111000001",
  59454=>"000111000",
  59455=>"000010100",
  59456=>"111001011",
  59457=>"000001101",
  59458=>"101010010",
  59459=>"111111110",
  59460=>"011100100",
  59461=>"001110111",
  59462=>"001110111",
  59463=>"011010000",
  59464=>"001100001",
  59465=>"001000101",
  59466=>"010011100",
  59467=>"001100010",
  59468=>"101111011",
  59469=>"111001111",
  59470=>"101011000",
  59471=>"010101000",
  59472=>"110100110",
  59473=>"011010011",
  59474=>"101001000",
  59475=>"101010011",
  59476=>"101101010",
  59477=>"110110101",
  59478=>"001000111",
  59479=>"011101111",
  59480=>"001110110",
  59481=>"100011010",
  59482=>"011011110",
  59483=>"101100001",
  59484=>"000111000",
  59485=>"010011001",
  59486=>"000011110",
  59487=>"011000101",
  59488=>"001000011",
  59489=>"101010101",
  59490=>"110111000",
  59491=>"010011001",
  59492=>"001000010",
  59493=>"010101011",
  59494=>"111111001",
  59495=>"110111111",
  59496=>"111110011",
  59497=>"110010011",
  59498=>"000011001",
  59499=>"110110110",
  59500=>"011111001",
  59501=>"011101100",
  59502=>"001001110",
  59503=>"111110101",
  59504=>"110101011",
  59505=>"010101101",
  59506=>"011010111",
  59507=>"010111100",
  59508=>"100111101",
  59509=>"010001010",
  59510=>"011110111",
  59511=>"111010001",
  59512=>"100110100",
  59513=>"000000100",
  59514=>"100011101",
  59515=>"101101111",
  59516=>"100001110",
  59517=>"000100110",
  59518=>"110101001",
  59519=>"011101010",
  59520=>"010001100",
  59521=>"101110111",
  59522=>"100101001",
  59523=>"000000001",
  59524=>"101100011",
  59525=>"111111101",
  59526=>"100001000",
  59527=>"100001000",
  59528=>"011011110",
  59529=>"000001111",
  59530=>"101010001",
  59531=>"001011000",
  59532=>"010101110",
  59533=>"011010001",
  59534=>"111000010",
  59535=>"100000000",
  59536=>"011111011",
  59537=>"011010010",
  59538=>"000110100",
  59539=>"110011100",
  59540=>"101001010",
  59541=>"110000010",
  59542=>"011100010",
  59543=>"010001100",
  59544=>"011101010",
  59545=>"110101000",
  59546=>"000111100",
  59547=>"011110110",
  59548=>"010110100",
  59549=>"110010001",
  59550=>"000111001",
  59551=>"010100101",
  59552=>"011000011",
  59553=>"110100111",
  59554=>"101000000",
  59555=>"000101011",
  59556=>"100000110",
  59557=>"111010011",
  59558=>"000011000",
  59559=>"010101111",
  59560=>"100110001",
  59561=>"001000111",
  59562=>"000110110",
  59563=>"011010110",
  59564=>"000111110",
  59565=>"110101110",
  59566=>"110001000",
  59567=>"000000101",
  59568=>"011001101",
  59569=>"001111001",
  59570=>"100011000",
  59571=>"100110110",
  59572=>"001111011",
  59573=>"011110111",
  59574=>"001001110",
  59575=>"001000100",
  59576=>"011011010",
  59577=>"000001010",
  59578=>"001100111",
  59579=>"010000010",
  59580=>"010110001",
  59581=>"000010111",
  59582=>"101100110",
  59583=>"011010010",
  59584=>"010010110",
  59585=>"111110000",
  59586=>"000110110",
  59587=>"111000000",
  59588=>"111110001",
  59589=>"100011000",
  59590=>"101100001",
  59591=>"000101011",
  59592=>"000011100",
  59593=>"101110000",
  59594=>"110001101",
  59595=>"111011101",
  59596=>"011010000",
  59597=>"111110101",
  59598=>"001000110",
  59599=>"101000111",
  59600=>"100111001",
  59601=>"111011001",
  59602=>"010001100",
  59603=>"110111111",
  59604=>"100110101",
  59605=>"001010101",
  59606=>"011010000",
  59607=>"010110100",
  59608=>"010110000",
  59609=>"100010100",
  59610=>"111011010",
  59611=>"000000100",
  59612=>"000011100",
  59613=>"101010110",
  59614=>"011101010",
  59615=>"100100010",
  59616=>"101001100",
  59617=>"000010101",
  59618=>"110101000",
  59619=>"000101111",
  59620=>"001101010",
  59621=>"101000001",
  59622=>"000010111",
  59623=>"000101001",
  59624=>"000000010",
  59625=>"100100111",
  59626=>"001101111",
  59627=>"010101110",
  59628=>"100110010",
  59629=>"001011101",
  59630=>"101001001",
  59631=>"010000000",
  59632=>"110101111",
  59633=>"111111101",
  59634=>"100010011",
  59635=>"100011011",
  59636=>"100101111",
  59637=>"010010010",
  59638=>"010000010",
  59639=>"110111000",
  59640=>"000101101",
  59641=>"010100101",
  59642=>"100001011",
  59643=>"111001100",
  59644=>"001100001",
  59645=>"011111101",
  59646=>"101001011",
  59647=>"011001000",
  59648=>"000010010",
  59649=>"010001111",
  59650=>"101001000",
  59651=>"100011101",
  59652=>"100101011",
  59653=>"001111100",
  59654=>"100111001",
  59655=>"011110101",
  59656=>"000111001",
  59657=>"111110101",
  59658=>"101111000",
  59659=>"000010110",
  59660=>"111010001",
  59661=>"000001010",
  59662=>"000010101",
  59663=>"011010001",
  59664=>"010000110",
  59665=>"100000001",
  59666=>"101111111",
  59667=>"111101000",
  59668=>"001111111",
  59669=>"000010001",
  59670=>"000110010",
  59671=>"001000001",
  59672=>"101100111",
  59673=>"110010100",
  59674=>"111000110",
  59675=>"111111010",
  59676=>"100011100",
  59677=>"101111110",
  59678=>"111000000",
  59679=>"111100011",
  59680=>"000100101",
  59681=>"001010001",
  59682=>"101011111",
  59683=>"110101110",
  59684=>"100110100",
  59685=>"011111111",
  59686=>"000100010",
  59687=>"110111101",
  59688=>"111111010",
  59689=>"111001100",
  59690=>"101000101",
  59691=>"011101110",
  59692=>"010000101",
  59693=>"111110110",
  59694=>"000000000",
  59695=>"000100001",
  59696=>"001001010",
  59697=>"010110111",
  59698=>"010001111",
  59699=>"100111101",
  59700=>"001110110",
  59701=>"000110010",
  59702=>"100100011",
  59703=>"111110110",
  59704=>"001000000",
  59705=>"001010001",
  59706=>"101100100",
  59707=>"111101101",
  59708=>"011001011",
  59709=>"000000101",
  59710=>"000010010",
  59711=>"011100001",
  59712=>"000100111",
  59713=>"000010010",
  59714=>"000100000",
  59715=>"111010100",
  59716=>"101110111",
  59717=>"001001101",
  59718=>"101000101",
  59719=>"110110001",
  59720=>"101001010",
  59721=>"000101000",
  59722=>"110110101",
  59723=>"010100011",
  59724=>"001101100",
  59725=>"100110000",
  59726=>"001000001",
  59727=>"100111001",
  59728=>"101000100",
  59729=>"101011101",
  59730=>"001001110",
  59731=>"011110111",
  59732=>"101000100",
  59733=>"000001101",
  59734=>"011101010",
  59735=>"110001101",
  59736=>"001000010",
  59737=>"100110111",
  59738=>"011111110",
  59739=>"101011010",
  59740=>"011010000",
  59741=>"101001000",
  59742=>"101110011",
  59743=>"110011101",
  59744=>"100110010",
  59745=>"001011101",
  59746=>"100001011",
  59747=>"001111001",
  59748=>"010011000",
  59749=>"010110101",
  59750=>"101000000",
  59751=>"101110000",
  59752=>"100100101",
  59753=>"011100101",
  59754=>"010111000",
  59755=>"100100111",
  59756=>"111111111",
  59757=>"010111000",
  59758=>"101110110",
  59759=>"010010000",
  59760=>"001000100",
  59761=>"110001111",
  59762=>"011101000",
  59763=>"110111100",
  59764=>"001111111",
  59765=>"001010011",
  59766=>"100011001",
  59767=>"100000011",
  59768=>"001010010",
  59769=>"101000001",
  59770=>"010011011",
  59771=>"101110010",
  59772=>"000011010",
  59773=>"111110110",
  59774=>"001000111",
  59775=>"011101000",
  59776=>"111011101",
  59777=>"111000100",
  59778=>"111101111",
  59779=>"111111111",
  59780=>"000000000",
  59781=>"000001011",
  59782=>"100001000",
  59783=>"110111011",
  59784=>"011101001",
  59785=>"111001011",
  59786=>"011111110",
  59787=>"111001101",
  59788=>"100101011",
  59789=>"111111111",
  59790=>"000010011",
  59791=>"111101111",
  59792=>"110011001",
  59793=>"111010110",
  59794=>"001101010",
  59795=>"011001011",
  59796=>"011100010",
  59797=>"010000011",
  59798=>"000000001",
  59799=>"111011010",
  59800=>"110001011",
  59801=>"001000101",
  59802=>"110001011",
  59803=>"100100100",
  59804=>"100110010",
  59805=>"001110001",
  59806=>"011110110",
  59807=>"101001011",
  59808=>"100100100",
  59809=>"000000101",
  59810=>"100110000",
  59811=>"100100010",
  59812=>"011110011",
  59813=>"110000001",
  59814=>"010101101",
  59815=>"001110110",
  59816=>"100101110",
  59817=>"101100100",
  59818=>"001100001",
  59819=>"110111110",
  59820=>"001101100",
  59821=>"000101100",
  59822=>"110100100",
  59823=>"011011011",
  59824=>"100000101",
  59825=>"111111011",
  59826=>"001101110",
  59827=>"001000001",
  59828=>"001111110",
  59829=>"011001010",
  59830=>"010010110",
  59831=>"010101010",
  59832=>"000001101",
  59833=>"101000010",
  59834=>"111101000",
  59835=>"111100111",
  59836=>"110100111",
  59837=>"100110110",
  59838=>"010110100",
  59839=>"111000111",
  59840=>"101000010",
  59841=>"001111010",
  59842=>"001011000",
  59843=>"111010011",
  59844=>"110101111",
  59845=>"010010000",
  59846=>"101101000",
  59847=>"100011010",
  59848=>"101010100",
  59849=>"001110100",
  59850=>"111110110",
  59851=>"100001100",
  59852=>"100101101",
  59853=>"101111011",
  59854=>"000111101",
  59855=>"010100001",
  59856=>"101010111",
  59857=>"110001110",
  59858=>"010110001",
  59859=>"000100000",
  59860=>"001001010",
  59861=>"010011110",
  59862=>"010110011",
  59863=>"011101101",
  59864=>"010011101",
  59865=>"000101101",
  59866=>"000110100",
  59867=>"110000110",
  59868=>"000100101",
  59869=>"101101101",
  59870=>"001011011",
  59871=>"100110011",
  59872=>"111010111",
  59873=>"111011001",
  59874=>"111110111",
  59875=>"001110110",
  59876=>"110000001",
  59877=>"000100011",
  59878=>"101111010",
  59879=>"000001101",
  59880=>"100110000",
  59881=>"010001100",
  59882=>"000000000",
  59883=>"111110111",
  59884=>"010110101",
  59885=>"011001000",
  59886=>"100010101",
  59887=>"010100000",
  59888=>"000110000",
  59889=>"010110011",
  59890=>"101011101",
  59891=>"001101100",
  59892=>"111011110",
  59893=>"111010011",
  59894=>"100111000",
  59895=>"110011011",
  59896=>"110000001",
  59897=>"001100110",
  59898=>"111111101",
  59899=>"101010011",
  59900=>"001000110",
  59901=>"010000010",
  59902=>"110100010",
  59903=>"100110011",
  59904=>"001010011",
  59905=>"001001010",
  59906=>"100000011",
  59907=>"010001011",
  59908=>"111101011",
  59909=>"001000000",
  59910=>"000011001",
  59911=>"001011101",
  59912=>"111011001",
  59913=>"011100001",
  59914=>"100110110",
  59915=>"001010001",
  59916=>"010111011",
  59917=>"011010011",
  59918=>"101010011",
  59919=>"100101100",
  59920=>"010100110",
  59921=>"101100001",
  59922=>"100011100",
  59923=>"011100011",
  59924=>"011111010",
  59925=>"001111000",
  59926=>"011000010",
  59927=>"111100011",
  59928=>"010110000",
  59929=>"110010111",
  59930=>"010010010",
  59931=>"101000000",
  59932=>"000100000",
  59933=>"001111010",
  59934=>"000111110",
  59935=>"000010111",
  59936=>"011000100",
  59937=>"001110011",
  59938=>"001000110",
  59939=>"001110110",
  59940=>"011011111",
  59941=>"111101010",
  59942=>"100111000",
  59943=>"101000100",
  59944=>"101010111",
  59945=>"101111111",
  59946=>"000110010",
  59947=>"101101001",
  59948=>"101001111",
  59949=>"110000110",
  59950=>"101110010",
  59951=>"110110001",
  59952=>"111111101",
  59953=>"011010001",
  59954=>"100100010",
  59955=>"110010101",
  59956=>"000000011",
  59957=>"011100000",
  59958=>"100111101",
  59959=>"101101010",
  59960=>"110011010",
  59961=>"000111011",
  59962=>"101000011",
  59963=>"000110100",
  59964=>"110100100",
  59965=>"100000010",
  59966=>"000100000",
  59967=>"111110101",
  59968=>"001110001",
  59969=>"000000001",
  59970=>"000100011",
  59971=>"011010111",
  59972=>"011110100",
  59973=>"111001010",
  59974=>"000010011",
  59975=>"010011110",
  59976=>"011010100",
  59977=>"110101101",
  59978=>"001100010",
  59979=>"101100100",
  59980=>"110011101",
  59981=>"100100001",
  59982=>"110101100",
  59983=>"010110100",
  59984=>"010001110",
  59985=>"000111000",
  59986=>"100000011",
  59987=>"001001110",
  59988=>"001010111",
  59989=>"110100000",
  59990=>"011101111",
  59991=>"011011010",
  59992=>"111001101",
  59993=>"000011000",
  59994=>"110101111",
  59995=>"110111001",
  59996=>"000000111",
  59997=>"111111010",
  59998=>"111110111",
  59999=>"100100111",
  60000=>"100110110",
  60001=>"001100000",
  60002=>"110110000",
  60003=>"111010111",
  60004=>"100010100",
  60005=>"001100100",
  60006=>"100000010",
  60007=>"001000100",
  60008=>"100111110",
  60009=>"011000110",
  60010=>"001010001",
  60011=>"010010000",
  60012=>"010101011",
  60013=>"010011010",
  60014=>"100010111",
  60015=>"011011010",
  60016=>"011110000",
  60017=>"010000110",
  60018=>"111101101",
  60019=>"011010010",
  60020=>"100100001",
  60021=>"100111001",
  60022=>"110000000",
  60023=>"101110110",
  60024=>"111011101",
  60025=>"000000110",
  60026=>"000110000",
  60027=>"001001000",
  60028=>"110111100",
  60029=>"111000011",
  60030=>"000011001",
  60031=>"000100011",
  60032=>"100100000",
  60033=>"001011000",
  60034=>"100011000",
  60035=>"111100101",
  60036=>"000111110",
  60037=>"111101000",
  60038=>"011010001",
  60039=>"101100100",
  60040=>"001010110",
  60041=>"011101100",
  60042=>"000100110",
  60043=>"101011111",
  60044=>"010000010",
  60045=>"001000101",
  60046=>"110011011",
  60047=>"111000111",
  60048=>"011100000",
  60049=>"101001111",
  60050=>"001111101",
  60051=>"110100000",
  60052=>"001110101",
  60053=>"011111111",
  60054=>"010011000",
  60055=>"100111101",
  60056=>"011010110",
  60057=>"100011110",
  60058=>"000110011",
  60059=>"111111000",
  60060=>"010111000",
  60061=>"110110111",
  60062=>"010101101",
  60063=>"001111010",
  60064=>"111000000",
  60065=>"111100111",
  60066=>"111000000",
  60067=>"100000111",
  60068=>"111111011",
  60069=>"111111011",
  60070=>"111001010",
  60071=>"000100001",
  60072=>"001110000",
  60073=>"111011010",
  60074=>"111010001",
  60075=>"111100010",
  60076=>"001101110",
  60077=>"111111110",
  60078=>"100110110",
  60079=>"110001101",
  60080=>"010001010",
  60081=>"011011011",
  60082=>"100100101",
  60083=>"001110100",
  60084=>"111111101",
  60085=>"010001001",
  60086=>"110001110",
  60087=>"011101000",
  60088=>"010000101",
  60089=>"111111111",
  60090=>"010100011",
  60091=>"100011101",
  60092=>"000010101",
  60093=>"101110001",
  60094=>"110111101",
  60095=>"101101101",
  60096=>"101000011",
  60097=>"000011011",
  60098=>"101010010",
  60099=>"001100110",
  60100=>"110000000",
  60101=>"001000010",
  60102=>"011111010",
  60103=>"001010110",
  60104=>"000001010",
  60105=>"001101010",
  60106=>"010000101",
  60107=>"111010101",
  60108=>"101111100",
  60109=>"111011010",
  60110=>"000000111",
  60111=>"000001101",
  60112=>"111111110",
  60113=>"111111100",
  60114=>"100101001",
  60115=>"100011010",
  60116=>"101111011",
  60117=>"001011100",
  60118=>"101101100",
  60119=>"110101101",
  60120=>"010101101",
  60121=>"101110100",
  60122=>"101011100",
  60123=>"101011000",
  60124=>"011111101",
  60125=>"101111000",
  60126=>"111100011",
  60127=>"100111110",
  60128=>"001111111",
  60129=>"101011001",
  60130=>"001011010",
  60131=>"101011111",
  60132=>"010100011",
  60133=>"001100001",
  60134=>"111010010",
  60135=>"101000000",
  60136=>"110010111",
  60137=>"100100000",
  60138=>"001100001",
  60139=>"111001010",
  60140=>"100100010",
  60141=>"000111111",
  60142=>"000001010",
  60143=>"101011011",
  60144=>"011001110",
  60145=>"010100001",
  60146=>"100000100",
  60147=>"101111000",
  60148=>"011011000",
  60149=>"111011001",
  60150=>"110111111",
  60151=>"111110100",
  60152=>"001110001",
  60153=>"111101100",
  60154=>"110010010",
  60155=>"000010000",
  60156=>"010111100",
  60157=>"000110001",
  60158=>"000011000",
  60159=>"101111010",
  60160=>"000010010",
  60161=>"010001000",
  60162=>"000010010",
  60163=>"101100000",
  60164=>"100101010",
  60165=>"100100110",
  60166=>"010001000",
  60167=>"001001010",
  60168=>"011010000",
  60169=>"000100101",
  60170=>"001110000",
  60171=>"100110101",
  60172=>"100000110",
  60173=>"111000111",
  60174=>"111000000",
  60175=>"101001000",
  60176=>"101110011",
  60177=>"001011100",
  60178=>"011100000",
  60179=>"001001011",
  60180=>"011101101",
  60181=>"101100001",
  60182=>"110110100",
  60183=>"101011101",
  60184=>"001001011",
  60185=>"001010010",
  60186=>"001000001",
  60187=>"100011010",
  60188=>"010000100",
  60189=>"110111100",
  60190=>"001001000",
  60191=>"010001001",
  60192=>"100001110",
  60193=>"000010001",
  60194=>"100011011",
  60195=>"100100000",
  60196=>"111100010",
  60197=>"000001000",
  60198=>"001000100",
  60199=>"101010110",
  60200=>"111101000",
  60201=>"110101100",
  60202=>"010000100",
  60203=>"011111111",
  60204=>"010000100",
  60205=>"111111111",
  60206=>"101111100",
  60207=>"111011110",
  60208=>"000001000",
  60209=>"000101011",
  60210=>"000001010",
  60211=>"010011100",
  60212=>"110001000",
  60213=>"010011000",
  60214=>"110010010",
  60215=>"111111100",
  60216=>"010100001",
  60217=>"000101010",
  60218=>"001011000",
  60219=>"010000110",
  60220=>"101111100",
  60221=>"111010100",
  60222=>"010000100",
  60223=>"011101110",
  60224=>"010000011",
  60225=>"000001110",
  60226=>"000011100",
  60227=>"001101000",
  60228=>"011011000",
  60229=>"000000011",
  60230=>"111001011",
  60231=>"100111111",
  60232=>"000110110",
  60233=>"110111100",
  60234=>"001110011",
  60235=>"011000101",
  60236=>"010010110",
  60237=>"100101100",
  60238=>"101101001",
  60239=>"111011101",
  60240=>"101011000",
  60241=>"000000111",
  60242=>"001011001",
  60243=>"001010010",
  60244=>"101110010",
  60245=>"001000100",
  60246=>"001001011",
  60247=>"010011010",
  60248=>"011000000",
  60249=>"100110011",
  60250=>"001000110",
  60251=>"110111110",
  60252=>"010100000",
  60253=>"110000101",
  60254=>"001110110",
  60255=>"101100001",
  60256=>"100010000",
  60257=>"101111001",
  60258=>"100011111",
  60259=>"000010000",
  60260=>"010010101",
  60261=>"110010000",
  60262=>"000011111",
  60263=>"111000111",
  60264=>"100100001",
  60265=>"011000001",
  60266=>"110010110",
  60267=>"010011001",
  60268=>"000001001",
  60269=>"111001100",
  60270=>"101101000",
  60271=>"010001011",
  60272=>"000001001",
  60273=>"100001101",
  60274=>"110000101",
  60275=>"001001001",
  60276=>"101101100",
  60277=>"000010000",
  60278=>"001011110",
  60279=>"101101001",
  60280=>"111001111",
  60281=>"110000101",
  60282=>"111110010",
  60283=>"010110101",
  60284=>"110100010",
  60285=>"001001100",
  60286=>"100000000",
  60287=>"110001100",
  60288=>"101000011",
  60289=>"101000001",
  60290=>"010111101",
  60291=>"010010001",
  60292=>"100000100",
  60293=>"111111101",
  60294=>"011011000",
  60295=>"011000100",
  60296=>"001100110",
  60297=>"110111010",
  60298=>"100110111",
  60299=>"000101010",
  60300=>"100111000",
  60301=>"000001001",
  60302=>"111000101",
  60303=>"111110110",
  60304=>"110101001",
  60305=>"110010000",
  60306=>"000000000",
  60307=>"101111011",
  60308=>"100001101",
  60309=>"110110101",
  60310=>"000000001",
  60311=>"100000001",
  60312=>"101100111",
  60313=>"001000011",
  60314=>"100111101",
  60315=>"010100011",
  60316=>"001010111",
  60317=>"011111000",
  60318=>"001000111",
  60319=>"001111110",
  60320=>"111011100",
  60321=>"010101111",
  60322=>"001001110",
  60323=>"011110010",
  60324=>"010001101",
  60325=>"010100101",
  60326=>"010000011",
  60327=>"101101111",
  60328=>"000000111",
  60329=>"111110100",
  60330=>"100110011",
  60331=>"110110000",
  60332=>"000000000",
  60333=>"111111011",
  60334=>"001010011",
  60335=>"101111010",
  60336=>"101110111",
  60337=>"110000000",
  60338=>"101101111",
  60339=>"000010110",
  60340=>"001111101",
  60341=>"100110100",
  60342=>"100001110",
  60343=>"101011000",
  60344=>"111111011",
  60345=>"100010100",
  60346=>"000000111",
  60347=>"110000110",
  60348=>"101000101",
  60349=>"111011111",
  60350=>"110011100",
  60351=>"011010100",
  60352=>"110111110",
  60353=>"000000001",
  60354=>"001100000",
  60355=>"100001000",
  60356=>"001001110",
  60357=>"100011001",
  60358=>"111011011",
  60359=>"111101010",
  60360=>"100010000",
  60361=>"111100000",
  60362=>"010010010",
  60363=>"011011111",
  60364=>"001000110",
  60365=>"100000010",
  60366=>"101101100",
  60367=>"101001001",
  60368=>"101100011",
  60369=>"000110111",
  60370=>"010000011",
  60371=>"100100101",
  60372=>"100010100",
  60373=>"100000011",
  60374=>"000010001",
  60375=>"100101110",
  60376=>"001111110",
  60377=>"001110111",
  60378=>"000100011",
  60379=>"101110000",
  60380=>"100000111",
  60381=>"101010100",
  60382=>"110000001",
  60383=>"001001100",
  60384=>"011010000",
  60385=>"011110101",
  60386=>"001000110",
  60387=>"111001100",
  60388=>"001001000",
  60389=>"101000000",
  60390=>"111100100",
  60391=>"001111111",
  60392=>"000100011",
  60393=>"100011110",
  60394=>"001110010",
  60395=>"000100000",
  60396=>"000110110",
  60397=>"101010110",
  60398=>"101100001",
  60399=>"000110111",
  60400=>"001000000",
  60401=>"110010110",
  60402=>"001100000",
  60403=>"001001011",
  60404=>"011111110",
  60405=>"110010111",
  60406=>"011010100",
  60407=>"000011001",
  60408=>"110000011",
  60409=>"011111101",
  60410=>"110000000",
  60411=>"000101000",
  60412=>"000011111",
  60413=>"001111001",
  60414=>"100001001",
  60415=>"101000011",
  60416=>"011010011",
  60417=>"100110101",
  60418=>"010011110",
  60419=>"011100000",
  60420=>"001011001",
  60421=>"001111000",
  60422=>"100100100",
  60423=>"110001111",
  60424=>"100101100",
  60425=>"011100111",
  60426=>"111111011",
  60427=>"110001010",
  60428=>"000011101",
  60429=>"011101101",
  60430=>"001010100",
  60431=>"010111101",
  60432=>"001000001",
  60433=>"101101011",
  60434=>"010100110",
  60435=>"110110001",
  60436=>"111001110",
  60437=>"110000011",
  60438=>"111101111",
  60439=>"000110101",
  60440=>"010000110",
  60441=>"001010100",
  60442=>"100011000",
  60443=>"110100100",
  60444=>"000011000",
  60445=>"111000011",
  60446=>"001101011",
  60447=>"110111010",
  60448=>"110110111",
  60449=>"100001011",
  60450=>"010101000",
  60451=>"001101000",
  60452=>"010000110",
  60453=>"011111010",
  60454=>"110001001",
  60455=>"111000001",
  60456=>"010110110",
  60457=>"110110110",
  60458=>"111010001",
  60459=>"101111111",
  60460=>"000101011",
  60461=>"010100011",
  60462=>"111111110",
  60463=>"011110100",
  60464=>"110111100",
  60465=>"011011001",
  60466=>"011110100",
  60467=>"001100111",
  60468=>"010011000",
  60469=>"101110010",
  60470=>"000001010",
  60471=>"001011011",
  60472=>"000010000",
  60473=>"011001111",
  60474=>"110001000",
  60475=>"100000000",
  60476=>"001111011",
  60477=>"110110010",
  60478=>"010100111",
  60479=>"001100011",
  60480=>"111010100",
  60481=>"110111000",
  60482=>"000010011",
  60483=>"000100111",
  60484=>"100011011",
  60485=>"000111111",
  60486=>"110000100",
  60487=>"011011011",
  60488=>"001001010",
  60489=>"100100111",
  60490=>"100000000",
  60491=>"011110000",
  60492=>"001100010",
  60493=>"001100000",
  60494=>"111111111",
  60495=>"100001110",
  60496=>"011101000",
  60497=>"001100000",
  60498=>"111011111",
  60499=>"010001010",
  60500=>"010011101",
  60501=>"010010111",
  60502=>"011001111",
  60503=>"010001100",
  60504=>"000001010",
  60505=>"110010000",
  60506=>"110111100",
  60507=>"000011010",
  60508=>"001000110",
  60509=>"111010010",
  60510=>"000011110",
  60511=>"000001000",
  60512=>"010110001",
  60513=>"001000100",
  60514=>"000001010",
  60515=>"000110100",
  60516=>"110110001",
  60517=>"001111011",
  60518=>"000000010",
  60519=>"100011001",
  60520=>"110000000",
  60521=>"010110111",
  60522=>"000000000",
  60523=>"110101110",
  60524=>"000001000",
  60525=>"111011000",
  60526=>"110001010",
  60527=>"001100111",
  60528=>"010001111",
  60529=>"001110101",
  60530=>"110000001",
  60531=>"001001000",
  60532=>"001011011",
  60533=>"111011011",
  60534=>"110101011",
  60535=>"100101111",
  60536=>"000101100",
  60537=>"101001101",
  60538=>"100000111",
  60539=>"010111011",
  60540=>"110101111",
  60541=>"010000000",
  60542=>"110101001",
  60543=>"000100001",
  60544=>"110101101",
  60545=>"000001110",
  60546=>"000001101",
  60547=>"101011110",
  60548=>"001001110",
  60549=>"111100000",
  60550=>"100111111",
  60551=>"010101100",
  60552=>"100111111",
  60553=>"100100010",
  60554=>"000110001",
  60555=>"101110001",
  60556=>"101111111",
  60557=>"011001001",
  60558=>"100010010",
  60559=>"011011101",
  60560=>"001001101",
  60561=>"001011001",
  60562=>"101010110",
  60563=>"011101101",
  60564=>"101010110",
  60565=>"100101011",
  60566=>"100010000",
  60567=>"101111010",
  60568=>"011000101",
  60569=>"100000000",
  60570=>"011110000",
  60571=>"111111100",
  60572=>"010110001",
  60573=>"000111101",
  60574=>"101100101",
  60575=>"001001101",
  60576=>"001011000",
  60577=>"000111110",
  60578=>"110100010",
  60579=>"000111010",
  60580=>"000100000",
  60581=>"011010000",
  60582=>"010101000",
  60583=>"100110000",
  60584=>"011111000",
  60585=>"001111101",
  60586=>"000101100",
  60587=>"110011101",
  60588=>"001010001",
  60589=>"100101101",
  60590=>"011111010",
  60591=>"000111100",
  60592=>"001111010",
  60593=>"100110111",
  60594=>"010010111",
  60595=>"110010110",
  60596=>"010010101",
  60597=>"010010101",
  60598=>"101100100",
  60599=>"011101110",
  60600=>"000110101",
  60601=>"110110110",
  60602=>"111111111",
  60603=>"001001101",
  60604=>"111111101",
  60605=>"110110110",
  60606=>"001000111",
  60607=>"000000011",
  60608=>"110100001",
  60609=>"010011110",
  60610=>"001100100",
  60611=>"100101110",
  60612=>"110111000",
  60613=>"100101111",
  60614=>"110000011",
  60615=>"011000000",
  60616=>"001101110",
  60617=>"011010111",
  60618=>"001000011",
  60619=>"101000110",
  60620=>"100111000",
  60621=>"001111101",
  60622=>"001111111",
  60623=>"100110100",
  60624=>"101001101",
  60625=>"011011110",
  60626=>"100001010",
  60627=>"110010111",
  60628=>"101011011",
  60629=>"110001001",
  60630=>"111011010",
  60631=>"100101100",
  60632=>"000011010",
  60633=>"000000101",
  60634=>"010001000",
  60635=>"000000101",
  60636=>"010101000",
  60637=>"011000011",
  60638=>"100000101",
  60639=>"010000111",
  60640=>"001101011",
  60641=>"111110010",
  60642=>"101001100",
  60643=>"111001010",
  60644=>"100100010",
  60645=>"111111011",
  60646=>"000011010",
  60647=>"000111011",
  60648=>"010110001",
  60649=>"011111110",
  60650=>"110010000",
  60651=>"000110011",
  60652=>"111010111",
  60653=>"111010010",
  60654=>"111010000",
  60655=>"001011001",
  60656=>"111110011",
  60657=>"001100001",
  60658=>"110101100",
  60659=>"001110000",
  60660=>"100111011",
  60661=>"100001111",
  60662=>"001110011",
  60663=>"001110100",
  60664=>"011100110",
  60665=>"110111100",
  60666=>"100010000",
  60667=>"100101100",
  60668=>"010010000",
  60669=>"010101110",
  60670=>"001000100",
  60671=>"100100111",
  60672=>"000001100",
  60673=>"010001001",
  60674=>"011111110",
  60675=>"001011110",
  60676=>"001100110",
  60677=>"010101000",
  60678=>"111111100",
  60679=>"011100010",
  60680=>"000110110",
  60681=>"001110100",
  60682=>"011110010",
  60683=>"010100100",
  60684=>"010001110",
  60685=>"001111011",
  60686=>"000110100",
  60687=>"100110010",
  60688=>"111110001",
  60689=>"000011110",
  60690=>"111100011",
  60691=>"010000000",
  60692=>"011100001",
  60693=>"011101001",
  60694=>"010011010",
  60695=>"101100100",
  60696=>"111010001",
  60697=>"110001111",
  60698=>"001101001",
  60699=>"010101011",
  60700=>"010010110",
  60701=>"111010110",
  60702=>"110111100",
  60703=>"101111101",
  60704=>"100011101",
  60705=>"000011101",
  60706=>"101110001",
  60707=>"110010011",
  60708=>"011110001",
  60709=>"110000000",
  60710=>"011000010",
  60711=>"011011010",
  60712=>"010010001",
  60713=>"100011110",
  60714=>"000001001",
  60715=>"111111011",
  60716=>"111010110",
  60717=>"011110110",
  60718=>"111110111",
  60719=>"011111110",
  60720=>"110101110",
  60721=>"101011110",
  60722=>"011101010",
  60723=>"100111000",
  60724=>"100100100",
  60725=>"011111011",
  60726=>"111111101",
  60727=>"111001111",
  60728=>"101011000",
  60729=>"110110010",
  60730=>"011100000",
  60731=>"010100010",
  60732=>"101000111",
  60733=>"100001100",
  60734=>"010010110",
  60735=>"010000110",
  60736=>"100100001",
  60737=>"111011101",
  60738=>"001010000",
  60739=>"100010011",
  60740=>"011111111",
  60741=>"100010110",
  60742=>"001100101",
  60743=>"000100001",
  60744=>"100111110",
  60745=>"010011110",
  60746=>"111111010",
  60747=>"011111000",
  60748=>"110100000",
  60749=>"011010100",
  60750=>"001110010",
  60751=>"111001001",
  60752=>"011101011",
  60753=>"001110000",
  60754=>"100110000",
  60755=>"111111011",
  60756=>"011100011",
  60757=>"001110010",
  60758=>"000101011",
  60759=>"100001000",
  60760=>"010000001",
  60761=>"000000110",
  60762=>"010000011",
  60763=>"011100101",
  60764=>"001011101",
  60765=>"000000010",
  60766=>"100001010",
  60767=>"100011101",
  60768=>"011001110",
  60769=>"100000111",
  60770=>"010110100",
  60771=>"100010110",
  60772=>"111000010",
  60773=>"001111100",
  60774=>"000011110",
  60775=>"100100100",
  60776=>"101000000",
  60777=>"100101010",
  60778=>"001000010",
  60779=>"110111110",
  60780=>"000010110",
  60781=>"000000111",
  60782=>"010010111",
  60783=>"001111101",
  60784=>"110001101",
  60785=>"000101010",
  60786=>"101011000",
  60787=>"110010100",
  60788=>"110111110",
  60789=>"111100110",
  60790=>"010110101",
  60791=>"101011100",
  60792=>"011101100",
  60793=>"001010001",
  60794=>"011011111",
  60795=>"001111111",
  60796=>"110101010",
  60797=>"110101001",
  60798=>"000110000",
  60799=>"001110001",
  60800=>"110100110",
  60801=>"101001100",
  60802=>"011011011",
  60803=>"001110011",
  60804=>"001101010",
  60805=>"000110000",
  60806=>"001110101",
  60807=>"010001110",
  60808=>"001000101",
  60809=>"001010011",
  60810=>"001010010",
  60811=>"000000011",
  60812=>"111010011",
  60813=>"000100000",
  60814=>"111100101",
  60815=>"000110001",
  60816=>"001000001",
  60817=>"001001101",
  60818=>"000101000",
  60819=>"100111111",
  60820=>"100001010",
  60821=>"010000001",
  60822=>"111000010",
  60823=>"100111101",
  60824=>"001101010",
  60825=>"110010001",
  60826=>"101011001",
  60827=>"001110001",
  60828=>"010010101",
  60829=>"010000000",
  60830=>"101101110",
  60831=>"001010110",
  60832=>"100111100",
  60833=>"100000110",
  60834=>"000111010",
  60835=>"000010100",
  60836=>"100110000",
  60837=>"010001111",
  60838=>"001111101",
  60839=>"010000000",
  60840=>"110100010",
  60841=>"111101011",
  60842=>"001100001",
  60843=>"010111000",
  60844=>"001100000",
  60845=>"000100101",
  60846=>"101111011",
  60847=>"000001110",
  60848=>"000110101",
  60849=>"011110010",
  60850=>"110110100",
  60851=>"001100110",
  60852=>"000100101",
  60853=>"110010001",
  60854=>"000010000",
  60855=>"000111000",
  60856=>"011011110",
  60857=>"111110101",
  60858=>"101011010",
  60859=>"011101111",
  60860=>"000010011",
  60861=>"000000010",
  60862=>"001111010",
  60863=>"000001111",
  60864=>"111001000",
  60865=>"011110000",
  60866=>"011011101",
  60867=>"101111001",
  60868=>"010000011",
  60869=>"101110110",
  60870=>"011001101",
  60871=>"000101110",
  60872=>"111101000",
  60873=>"000110001",
  60874=>"011100000",
  60875=>"111101111",
  60876=>"101011000",
  60877=>"110010101",
  60878=>"101010101",
  60879=>"101111100",
  60880=>"010001100",
  60881=>"101011101",
  60882=>"000111101",
  60883=>"011110100",
  60884=>"111111111",
  60885=>"001111011",
  60886=>"101011101",
  60887=>"111111000",
  60888=>"111000101",
  60889=>"101001000",
  60890=>"001111100",
  60891=>"000010111",
  60892=>"110110001",
  60893=>"001100001",
  60894=>"011111011",
  60895=>"111100101",
  60896=>"011010011",
  60897=>"101110000",
  60898=>"001000111",
  60899=>"100101111",
  60900=>"101101111",
  60901=>"101100110",
  60902=>"000110011",
  60903=>"001111001",
  60904=>"011011110",
  60905=>"011111111",
  60906=>"110110110",
  60907=>"111011010",
  60908=>"111110111",
  60909=>"101111001",
  60910=>"000101010",
  60911=>"010100000",
  60912=>"001001111",
  60913=>"111100111",
  60914=>"100000011",
  60915=>"100101011",
  60916=>"001000000",
  60917=>"101000100",
  60918=>"110101001",
  60919=>"110111001",
  60920=>"000001111",
  60921=>"100011110",
  60922=>"010110001",
  60923=>"001110001",
  60924=>"000100000",
  60925=>"111011110",
  60926=>"110110010",
  60927=>"000101001",
  60928=>"100000011",
  60929=>"111111101",
  60930=>"010011110",
  60931=>"000011010",
  60932=>"000011100",
  60933=>"000110000",
  60934=>"110110010",
  60935=>"000110111",
  60936=>"000111001",
  60937=>"100000001",
  60938=>"101110111",
  60939=>"011101010",
  60940=>"111000110",
  60941=>"100111110",
  60942=>"110011111",
  60943=>"111111100",
  60944=>"111111011",
  60945=>"101000000",
  60946=>"001111011",
  60947=>"001011001",
  60948=>"010101110",
  60949=>"101001001",
  60950=>"010110101",
  60951=>"100000001",
  60952=>"100001010",
  60953=>"010111111",
  60954=>"011000110",
  60955=>"110011110",
  60956=>"111011111",
  60957=>"000011110",
  60958=>"100010001",
  60959=>"011111110",
  60960=>"001110110",
  60961=>"110110100",
  60962=>"100110101",
  60963=>"010110101",
  60964=>"001010111",
  60965=>"111111010",
  60966=>"011000011",
  60967=>"100110000",
  60968=>"100100001",
  60969=>"001110010",
  60970=>"001010111",
  60971=>"011110101",
  60972=>"110110000",
  60973=>"000010000",
  60974=>"011110000",
  60975=>"101110110",
  60976=>"011110101",
  60977=>"010001110",
  60978=>"110111111",
  60979=>"100001101",
  60980=>"010011001",
  60981=>"101111110",
  60982=>"001100101",
  60983=>"101100111",
  60984=>"111111011",
  60985=>"100001111",
  60986=>"010111000",
  60987=>"010101111",
  60988=>"001011110",
  60989=>"011011111",
  60990=>"101000011",
  60991=>"001111101",
  60992=>"100110110",
  60993=>"011101101",
  60994=>"011110000",
  60995=>"110000101",
  60996=>"101001101",
  60997=>"010001111",
  60998=>"011000010",
  60999=>"101110010",
  61000=>"101001111",
  61001=>"100000100",
  61002=>"001110101",
  61003=>"010010101",
  61004=>"011011100",
  61005=>"000000111",
  61006=>"010000000",
  61007=>"101100001",
  61008=>"100100101",
  61009=>"101110010",
  61010=>"001101000",
  61011=>"111101101",
  61012=>"011110010",
  61013=>"111001110",
  61014=>"100100010",
  61015=>"110110111",
  61016=>"101011111",
  61017=>"000101111",
  61018=>"101000010",
  61019=>"001011101",
  61020=>"110001111",
  61021=>"011111111",
  61022=>"011001001",
  61023=>"000110111",
  61024=>"100001001",
  61025=>"100100000",
  61026=>"001101001",
  61027=>"011000100",
  61028=>"100000010",
  61029=>"100100001",
  61030=>"001101010",
  61031=>"111101100",
  61032=>"011010100",
  61033=>"000111011",
  61034=>"111010010",
  61035=>"011011001",
  61036=>"100101010",
  61037=>"110110010",
  61038=>"000101011",
  61039=>"011001101",
  61040=>"101100000",
  61041=>"001110011",
  61042=>"110000001",
  61043=>"111110101",
  61044=>"100011001",
  61045=>"010100001",
  61046=>"101001001",
  61047=>"011110101",
  61048=>"100100100",
  61049=>"001100101",
  61050=>"010110100",
  61051=>"100100011",
  61052=>"011110110",
  61053=>"101100100",
  61054=>"011011110",
  61055=>"101010001",
  61056=>"111011001",
  61057=>"100101000",
  61058=>"111111000",
  61059=>"011111110",
  61060=>"101111100",
  61061=>"111101110",
  61062=>"011000011",
  61063=>"011101101",
  61064=>"100110111",
  61065=>"100100011",
  61066=>"111110001",
  61067=>"010100001",
  61068=>"000110101",
  61069=>"010100010",
  61070=>"010010010",
  61071=>"111011011",
  61072=>"101111101",
  61073=>"100011111",
  61074=>"001011110",
  61075=>"101010101",
  61076=>"001011010",
  61077=>"000010111",
  61078=>"000001000",
  61079=>"101011110",
  61080=>"100001010",
  61081=>"010111001",
  61082=>"110100110",
  61083=>"011110011",
  61084=>"111010011",
  61085=>"110101100",
  61086=>"111011110",
  61087=>"011010000",
  61088=>"101000010",
  61089=>"000000001",
  61090=>"001001001",
  61091=>"101110000",
  61092=>"111110001",
  61093=>"011010101",
  61094=>"000000111",
  61095=>"100000000",
  61096=>"001101100",
  61097=>"000110111",
  61098=>"011011010",
  61099=>"110010011",
  61100=>"110110101",
  61101=>"001100001",
  61102=>"011000111",
  61103=>"011011000",
  61104=>"001111000",
  61105=>"110110000",
  61106=>"010000001",
  61107=>"101110101",
  61108=>"111100000",
  61109=>"000100110",
  61110=>"011100000",
  61111=>"101111000",
  61112=>"110101111",
  61113=>"110110011",
  61114=>"100100110",
  61115=>"000111010",
  61116=>"101001111",
  61117=>"010001000",
  61118=>"000010000",
  61119=>"000000001",
  61120=>"000100010",
  61121=>"001001000",
  61122=>"110010110",
  61123=>"001100001",
  61124=>"110111000",
  61125=>"011011010",
  61126=>"101000101",
  61127=>"111110010",
  61128=>"100101000",
  61129=>"000010010",
  61130=>"111010010",
  61131=>"101110100",
  61132=>"010100111",
  61133=>"011001110",
  61134=>"111100110",
  61135=>"101001011",
  61136=>"010010001",
  61137=>"111010111",
  61138=>"010110011",
  61139=>"111000110",
  61140=>"010000111",
  61141=>"011110001",
  61142=>"100100111",
  61143=>"101101100",
  61144=>"100101001",
  61145=>"100011111",
  61146=>"100010001",
  61147=>"100010011",
  61148=>"011110011",
  61149=>"100110101",
  61150=>"000000000",
  61151=>"101111100",
  61152=>"111000100",
  61153=>"100100000",
  61154=>"101100111",
  61155=>"100101110",
  61156=>"001001011",
  61157=>"111001111",
  61158=>"100101101",
  61159=>"110011111",
  61160=>"000010111",
  61161=>"110011100",
  61162=>"100111001",
  61163=>"111101011",
  61164=>"001100000",
  61165=>"001011011",
  61166=>"111011001",
  61167=>"000111100",
  61168=>"011001011",
  61169=>"101010001",
  61170=>"001010111",
  61171=>"100110011",
  61172=>"000110000",
  61173=>"101100111",
  61174=>"100011100",
  61175=>"001011011",
  61176=>"100010001",
  61177=>"011000110",
  61178=>"001000000",
  61179=>"001111101",
  61180=>"011101101",
  61181=>"001000111",
  61182=>"011011011",
  61183=>"110111111",
  61184=>"010010100",
  61185=>"111000000",
  61186=>"101100100",
  61187=>"010011011",
  61188=>"010000010",
  61189=>"010011100",
  61190=>"000001001",
  61191=>"011010011",
  61192=>"010001101",
  61193=>"111111000",
  61194=>"011110101",
  61195=>"101011011",
  61196=>"010111111",
  61197=>"010111111",
  61198=>"101111001",
  61199=>"001100011",
  61200=>"100011001",
  61201=>"001000110",
  61202=>"100000100",
  61203=>"000011000",
  61204=>"011001101",
  61205=>"001000001",
  61206=>"101010110",
  61207=>"010000100",
  61208=>"101111011",
  61209=>"000110111",
  61210=>"111111011",
  61211=>"001010001",
  61212=>"111111010",
  61213=>"001000101",
  61214=>"001101111",
  61215=>"110111000",
  61216=>"100111100",
  61217=>"100110011",
  61218=>"100111110",
  61219=>"001000011",
  61220=>"000000000",
  61221=>"100000110",
  61222=>"111000101",
  61223=>"110111111",
  61224=>"001010100",
  61225=>"000011010",
  61226=>"111111101",
  61227=>"000100110",
  61228=>"101101101",
  61229=>"111000010",
  61230=>"100010001",
  61231=>"100010011",
  61232=>"111111000",
  61233=>"101100001",
  61234=>"110000010",
  61235=>"110010001",
  61236=>"110110101",
  61237=>"111110101",
  61238=>"000010101",
  61239=>"100111110",
  61240=>"001110000",
  61241=>"010000000",
  61242=>"000000010",
  61243=>"011000011",
  61244=>"000001100",
  61245=>"111001101",
  61246=>"101011011",
  61247=>"000000011",
  61248=>"000000000",
  61249=>"100111100",
  61250=>"100010100",
  61251=>"000010101",
  61252=>"100100000",
  61253=>"000011110",
  61254=>"000011011",
  61255=>"001100010",
  61256=>"001001100",
  61257=>"110111011",
  61258=>"101101101",
  61259=>"001111101",
  61260=>"000110101",
  61261=>"110010101",
  61262=>"001010011",
  61263=>"010110011",
  61264=>"010111010",
  61265=>"111000011",
  61266=>"001000100",
  61267=>"101110101",
  61268=>"100001100",
  61269=>"110100111",
  61270=>"101110111",
  61271=>"110001001",
  61272=>"000101111",
  61273=>"000111010",
  61274=>"101010101",
  61275=>"011000010",
  61276=>"111110010",
  61277=>"111001010",
  61278=>"001111111",
  61279=>"010011000",
  61280=>"011011010",
  61281=>"111000101",
  61282=>"000100100",
  61283=>"100010001",
  61284=>"100010100",
  61285=>"111101111",
  61286=>"011011101",
  61287=>"101001101",
  61288=>"101011110",
  61289=>"000110111",
  61290=>"011110001",
  61291=>"010010110",
  61292=>"111111001",
  61293=>"011101110",
  61294=>"010100100",
  61295=>"001010011",
  61296=>"110000110",
  61297=>"011001110",
  61298=>"110110110",
  61299=>"000010000",
  61300=>"100111101",
  61301=>"111110000",
  61302=>"101110000",
  61303=>"000011010",
  61304=>"010000101",
  61305=>"001011011",
  61306=>"111101101",
  61307=>"011110011",
  61308=>"010010000",
  61309=>"011101001",
  61310=>"010011111",
  61311=>"011100100",
  61312=>"000011010",
  61313=>"000001010",
  61314=>"110010010",
  61315=>"000110000",
  61316=>"111011000",
  61317=>"111101110",
  61318=>"100110001",
  61319=>"010111111",
  61320=>"011110100",
  61321=>"010111101",
  61322=>"110101110",
  61323=>"101011111",
  61324=>"000110001",
  61325=>"000110000",
  61326=>"000010010",
  61327=>"001110001",
  61328=>"110000000",
  61329=>"111100111",
  61330=>"000001010",
  61331=>"101111101",
  61332=>"001000000",
  61333=>"010100011",
  61334=>"001101010",
  61335=>"111001011",
  61336=>"000110111",
  61337=>"001110000",
  61338=>"010100000",
  61339=>"100011101",
  61340=>"101101000",
  61341=>"011111000",
  61342=>"111100111",
  61343=>"100100011",
  61344=>"110001101",
  61345=>"100010001",
  61346=>"011111110",
  61347=>"011111110",
  61348=>"110011110",
  61349=>"101110101",
  61350=>"001001101",
  61351=>"101110001",
  61352=>"110100100",
  61353=>"011000111",
  61354=>"111010110",
  61355=>"111100001",
  61356=>"000100100",
  61357=>"100001001",
  61358=>"100010101",
  61359=>"110110111",
  61360=>"100001011",
  61361=>"101111111",
  61362=>"010111101",
  61363=>"011110100",
  61364=>"010110100",
  61365=>"100101100",
  61366=>"100100001",
  61367=>"010100101",
  61368=>"110010101",
  61369=>"011110100",
  61370=>"111010110",
  61371=>"100000001",
  61372=>"111111010",
  61373=>"111101011",
  61374=>"001110100",
  61375=>"011111100",
  61376=>"110101100",
  61377=>"001010000",
  61378=>"111010001",
  61379=>"100011010",
  61380=>"010011000",
  61381=>"001100011",
  61382=>"010011010",
  61383=>"010011101",
  61384=>"011100110",
  61385=>"000011111",
  61386=>"000100010",
  61387=>"011111011",
  61388=>"011111010",
  61389=>"111110111",
  61390=>"000001101",
  61391=>"000010011",
  61392=>"111110100",
  61393=>"000110001",
  61394=>"011110111",
  61395=>"101111010",
  61396=>"011100111",
  61397=>"101100001",
  61398=>"011000100",
  61399=>"011011001",
  61400=>"011111100",
  61401=>"111111111",
  61402=>"110001010",
  61403=>"111100011",
  61404=>"111110000",
  61405=>"101101101",
  61406=>"101100011",
  61407=>"011010000",
  61408=>"111101110",
  61409=>"001011111",
  61410=>"011100000",
  61411=>"001111001",
  61412=>"011100100",
  61413=>"111010001",
  61414=>"110011001",
  61415=>"110101010",
  61416=>"110101001",
  61417=>"010011010",
  61418=>"001111100",
  61419=>"111001000",
  61420=>"000111110",
  61421=>"000101100",
  61422=>"001111011",
  61423=>"001001010",
  61424=>"011111010",
  61425=>"100010010",
  61426=>"000000001",
  61427=>"111110010",
  61428=>"011010000",
  61429=>"011111110",
  61430=>"000110000",
  61431=>"011011101",
  61432=>"010111011",
  61433=>"001001111",
  61434=>"111100000",
  61435=>"000100111",
  61436=>"111100000",
  61437=>"011110110",
  61438=>"000001001",
  61439=>"011011111",
  61440=>"100000001",
  61441=>"100000101",
  61442=>"011011101",
  61443=>"010000011",
  61444=>"100100001",
  61445=>"101011011",
  61446=>"111001110",
  61447=>"100001111",
  61448=>"110000011",
  61449=>"011110101",
  61450=>"000100110",
  61451=>"010111000",
  61452=>"001011100",
  61453=>"000111100",
  61454=>"000101100",
  61455=>"101010110",
  61456=>"011011010",
  61457=>"011011110",
  61458=>"011111011",
  61459=>"011110100",
  61460=>"010001101",
  61461=>"110000001",
  61462=>"111010110",
  61463=>"000100100",
  61464=>"001011110",
  61465=>"101111001",
  61466=>"000000100",
  61467=>"011101111",
  61468=>"101000111",
  61469=>"010000111",
  61470=>"111011010",
  61471=>"111101001",
  61472=>"011001001",
  61473=>"100011101",
  61474=>"000000011",
  61475=>"000001110",
  61476=>"001111011",
  61477=>"011100011",
  61478=>"110010011",
  61479=>"011001100",
  61480=>"100001001",
  61481=>"111110010",
  61482=>"100101111",
  61483=>"101010000",
  61484=>"111111011",
  61485=>"101101011",
  61486=>"000001001",
  61487=>"000101001",
  61488=>"011101101",
  61489=>"011010110",
  61490=>"110011011",
  61491=>"001110011",
  61492=>"111100111",
  61493=>"100111101",
  61494=>"011111001",
  61495=>"000100010",
  61496=>"111000110",
  61497=>"000010100",
  61498=>"001010110",
  61499=>"010101001",
  61500=>"010101000",
  61501=>"100001110",
  61502=>"100011000",
  61503=>"111001100",
  61504=>"100011100",
  61505=>"011100111",
  61506=>"110001100",
  61507=>"011111001",
  61508=>"111111110",
  61509=>"101101100",
  61510=>"110000010",
  61511=>"000111101",
  61512=>"000101011",
  61513=>"111101011",
  61514=>"001011001",
  61515=>"100011101",
  61516=>"001000001",
  61517=>"100111110",
  61518=>"001011000",
  61519=>"100011010",
  61520=>"100010001",
  61521=>"111010110",
  61522=>"100101010",
  61523=>"010000001",
  61524=>"111111000",
  61525=>"010000101",
  61526=>"010110101",
  61527=>"010101111",
  61528=>"001111110",
  61529=>"010000110",
  61530=>"110011011",
  61531=>"011111110",
  61532=>"000000000",
  61533=>"110011111",
  61534=>"001000100",
  61535=>"111110010",
  61536=>"011101111",
  61537=>"101011110",
  61538=>"010001000",
  61539=>"110011100",
  61540=>"000010100",
  61541=>"100111010",
  61542=>"000011001",
  61543=>"100001011",
  61544=>"100100100",
  61545=>"100000110",
  61546=>"111010101",
  61547=>"010000001",
  61548=>"101101110",
  61549=>"000010110",
  61550=>"010010110",
  61551=>"101110110",
  61552=>"001100001",
  61553=>"101110010",
  61554=>"010100100",
  61555=>"111011110",
  61556=>"011100001",
  61557=>"101010001",
  61558=>"101101100",
  61559=>"000000000",
  61560=>"010001011",
  61561=>"110100000",
  61562=>"000011011",
  61563=>"111101011",
  61564=>"000100111",
  61565=>"111010101",
  61566=>"001101010",
  61567=>"101100010",
  61568=>"001000100",
  61569=>"011010000",
  61570=>"111110110",
  61571=>"011100000",
  61572=>"100000110",
  61573=>"000000010",
  61574=>"011100011",
  61575=>"000110000",
  61576=>"100001101",
  61577=>"011110000",
  61578=>"111100111",
  61579=>"100111011",
  61580=>"111100110",
  61581=>"100010010",
  61582=>"001000010",
  61583=>"110010010",
  61584=>"100100000",
  61585=>"001000000",
  61586=>"011101001",
  61587=>"010101101",
  61588=>"001000100",
  61589=>"001010110",
  61590=>"001000100",
  61591=>"100001000",
  61592=>"000011111",
  61593=>"101001110",
  61594=>"110000011",
  61595=>"000011011",
  61596=>"010010110",
  61597=>"010101110",
  61598=>"001000000",
  61599=>"111101000",
  61600=>"101100110",
  61601=>"111101111",
  61602=>"100100110",
  61603=>"001011110",
  61604=>"010010101",
  61605=>"100000110",
  61606=>"110001011",
  61607=>"100000001",
  61608=>"101010000",
  61609=>"010110010",
  61610=>"110011100",
  61611=>"111110111",
  61612=>"100111001",
  61613=>"010100110",
  61614=>"110101111",
  61615=>"101101110",
  61616=>"011000010",
  61617=>"110101000",
  61618=>"100110000",
  61619=>"000010010",
  61620=>"000101000",
  61621=>"100100110",
  61622=>"001101111",
  61623=>"111101001",
  61624=>"001000100",
  61625=>"100010100",
  61626=>"001001110",
  61627=>"110010000",
  61628=>"111011010",
  61629=>"001101100",
  61630=>"011010010",
  61631=>"000010011",
  61632=>"011101011",
  61633=>"100110101",
  61634=>"101001010",
  61635=>"110010101",
  61636=>"001000111",
  61637=>"010110011",
  61638=>"110000100",
  61639=>"110111001",
  61640=>"011010011",
  61641=>"011110001",
  61642=>"011011110",
  61643=>"111110100",
  61644=>"101111010",
  61645=>"110000011",
  61646=>"010000100",
  61647=>"010000000",
  61648=>"111101011",
  61649=>"011010101",
  61650=>"101011010",
  61651=>"100110111",
  61652=>"000000111",
  61653=>"010110111",
  61654=>"001111010",
  61655=>"000000001",
  61656=>"001000010",
  61657=>"111101011",
  61658=>"110000000",
  61659=>"010001111",
  61660=>"101100011",
  61661=>"110000111",
  61662=>"010000000",
  61663=>"000111111",
  61664=>"000100000",
  61665=>"110001100",
  61666=>"011100000",
  61667=>"110010110",
  61668=>"001110110",
  61669=>"101111101",
  61670=>"101011001",
  61671=>"000001110",
  61672=>"010101000",
  61673=>"000111111",
  61674=>"011100011",
  61675=>"100010011",
  61676=>"100100000",
  61677=>"110010010",
  61678=>"111010110",
  61679=>"111101101",
  61680=>"000000000",
  61681=>"011110011",
  61682=>"000001011",
  61683=>"010010101",
  61684=>"010011100",
  61685=>"011101010",
  61686=>"110111101",
  61687=>"001100100",
  61688=>"101011101",
  61689=>"110000000",
  61690=>"100111110",
  61691=>"011000000",
  61692=>"100101111",
  61693=>"001001111",
  61694=>"100101011",
  61695=>"101001010",
  61696=>"011010010",
  61697=>"010100111",
  61698=>"001011101",
  61699=>"100111101",
  61700=>"101000000",
  61701=>"110111011",
  61702=>"111100001",
  61703=>"001110011",
  61704=>"000111000",
  61705=>"110111000",
  61706=>"001011001",
  61707=>"000100110",
  61708=>"001110101",
  61709=>"000111011",
  61710=>"010101101",
  61711=>"111111011",
  61712=>"001000011",
  61713=>"101101111",
  61714=>"111101110",
  61715=>"110010010",
  61716=>"000010001",
  61717=>"000111110",
  61718=>"001010010",
  61719=>"000000011",
  61720=>"101001001",
  61721=>"000001100",
  61722=>"000000011",
  61723=>"101001000",
  61724=>"010100001",
  61725=>"100111000",
  61726=>"110101001",
  61727=>"010011101",
  61728=>"100001101",
  61729=>"101000011",
  61730=>"100101110",
  61731=>"111110001",
  61732=>"001110101",
  61733=>"000100111",
  61734=>"111100111",
  61735=>"110001011",
  61736=>"101001001",
  61737=>"101110000",
  61738=>"010010110",
  61739=>"001110001",
  61740=>"000001010",
  61741=>"011101110",
  61742=>"010010010",
  61743=>"100011111",
  61744=>"110000110",
  61745=>"000010010",
  61746=>"111110111",
  61747=>"111110110",
  61748=>"000001010",
  61749=>"011101100",
  61750=>"110011111",
  61751=>"100011011",
  61752=>"110000001",
  61753=>"001101100",
  61754=>"100000110",
  61755=>"111111010",
  61756=>"111101111",
  61757=>"110011011",
  61758=>"100101101",
  61759=>"101111011",
  61760=>"110111101",
  61761=>"011100001",
  61762=>"111100011",
  61763=>"110010010",
  61764=>"110101100",
  61765=>"100000011",
  61766=>"010000000",
  61767=>"111101111",
  61768=>"001111001",
  61769=>"100010111",
  61770=>"100001011",
  61771=>"111101011",
  61772=>"001110110",
  61773=>"000001111",
  61774=>"010001011",
  61775=>"101000001",
  61776=>"111110100",
  61777=>"011100111",
  61778=>"111101111",
  61779=>"111001111",
  61780=>"111010011",
  61781=>"110000111",
  61782=>"100110110",
  61783=>"010111101",
  61784=>"000111001",
  61785=>"101011101",
  61786=>"111001111",
  61787=>"001000001",
  61788=>"111101011",
  61789=>"000000110",
  61790=>"000111110",
  61791=>"010011000",
  61792=>"011001000",
  61793=>"101110110",
  61794=>"101101101",
  61795=>"100001000",
  61796=>"010101110",
  61797=>"111111100",
  61798=>"100001000",
  61799=>"011101011",
  61800=>"101101110",
  61801=>"000010001",
  61802=>"010011101",
  61803=>"111110011",
  61804=>"101010010",
  61805=>"100101110",
  61806=>"000100000",
  61807=>"110101100",
  61808=>"111110001",
  61809=>"110100111",
  61810=>"001100001",
  61811=>"100000101",
  61812=>"000110100",
  61813=>"101111011",
  61814=>"111110110",
  61815=>"010110111",
  61816=>"111011101",
  61817=>"100000010",
  61818=>"011111111",
  61819=>"110111010",
  61820=>"100101011",
  61821=>"010000011",
  61822=>"100010101",
  61823=>"010111100",
  61824=>"001011101",
  61825=>"101101010",
  61826=>"011110101",
  61827=>"101100011",
  61828=>"101110011",
  61829=>"110010100",
  61830=>"001111110",
  61831=>"111110010",
  61832=>"101010100",
  61833=>"001001101",
  61834=>"100101111",
  61835=>"100110000",
  61836=>"100001110",
  61837=>"000010110",
  61838=>"110000100",
  61839=>"010010111",
  61840=>"010001100",
  61841=>"010111001",
  61842=>"010011101",
  61843=>"010100000",
  61844=>"100010000",
  61845=>"100110100",
  61846=>"010010000",
  61847=>"111100101",
  61848=>"110101000",
  61849=>"010011011",
  61850=>"100111111",
  61851=>"110010011",
  61852=>"111011010",
  61853=>"000101010",
  61854=>"101001101",
  61855=>"000111101",
  61856=>"110111011",
  61857=>"011110100",
  61858=>"010000010",
  61859=>"010100100",
  61860=>"111101100",
  61861=>"110000000",
  61862=>"111110100",
  61863=>"011101011",
  61864=>"101100011",
  61865=>"100011101",
  61866=>"000000011",
  61867=>"111110011",
  61868=>"101010001",
  61869=>"000000011",
  61870=>"111111101",
  61871=>"101011011",
  61872=>"101001001",
  61873=>"110001100",
  61874=>"010010111",
  61875=>"000101111",
  61876=>"000011100",
  61877=>"001000001",
  61878=>"011001110",
  61879=>"011011101",
  61880=>"011111001",
  61881=>"001011111",
  61882=>"100111011",
  61883=>"101011001",
  61884=>"001111101",
  61885=>"010101000",
  61886=>"000001010",
  61887=>"000101011",
  61888=>"011001001",
  61889=>"000010101",
  61890=>"111111001",
  61891=>"011001101",
  61892=>"011010100",
  61893=>"000111000",
  61894=>"011010110",
  61895=>"010100000",
  61896=>"101100011",
  61897=>"010111011",
  61898=>"110000100",
  61899=>"110110111",
  61900=>"111001111",
  61901=>"001010110",
  61902=>"000100111",
  61903=>"000010101",
  61904=>"110100000",
  61905=>"011000110",
  61906=>"111110011",
  61907=>"110011100",
  61908=>"010010010",
  61909=>"110111001",
  61910=>"111111111",
  61911=>"011010100",
  61912=>"000101010",
  61913=>"100110101",
  61914=>"101011101",
  61915=>"111001010",
  61916=>"100101001",
  61917=>"011001011",
  61918=>"101001101",
  61919=>"110001111",
  61920=>"100010100",
  61921=>"110010111",
  61922=>"011010101",
  61923=>"010001001",
  61924=>"000101010",
  61925=>"010001011",
  61926=>"001011110",
  61927=>"001111010",
  61928=>"111101001",
  61929=>"100010011",
  61930=>"101000100",
  61931=>"101100101",
  61932=>"001001011",
  61933=>"010010011",
  61934=>"100101011",
  61935=>"111100000",
  61936=>"001110100",
  61937=>"010001001",
  61938=>"101101101",
  61939=>"101110100",
  61940=>"001000011",
  61941=>"011111100",
  61942=>"010100101",
  61943=>"110110001",
  61944=>"000010001",
  61945=>"000011010",
  61946=>"100000110",
  61947=>"101000110",
  61948=>"001110111",
  61949=>"100010101",
  61950=>"101111111",
  61951=>"101000101",
  61952=>"100010100",
  61953=>"010111001",
  61954=>"001110000",
  61955=>"111011101",
  61956=>"111001100",
  61957=>"000010000",
  61958=>"010100011",
  61959=>"100010110",
  61960=>"011000100",
  61961=>"001110101",
  61962=>"101111111",
  61963=>"101010000",
  61964=>"101111010",
  61965=>"001111110",
  61966=>"100111111",
  61967=>"100011111",
  61968=>"110001101",
  61969=>"010111111",
  61970=>"110010010",
  61971=>"011001101",
  61972=>"010000011",
  61973=>"110100001",
  61974=>"011110011",
  61975=>"001001001",
  61976=>"001100001",
  61977=>"011011001",
  61978=>"010011111",
  61979=>"101100001",
  61980=>"100011000",
  61981=>"100000100",
  61982=>"010000110",
  61983=>"000001101",
  61984=>"001101011",
  61985=>"101110011",
  61986=>"000001101",
  61987=>"110101010",
  61988=>"101010110",
  61989=>"011111001",
  61990=>"000000010",
  61991=>"010010000",
  61992=>"001000000",
  61993=>"111011010",
  61994=>"001101111",
  61995=>"010000101",
  61996=>"001100000",
  61997=>"011000011",
  61998=>"011011001",
  61999=>"011000010",
  62000=>"001100101",
  62001=>"111101000",
  62002=>"010110101",
  62003=>"001011001",
  62004=>"110000000",
  62005=>"101000100",
  62006=>"010010101",
  62007=>"000001010",
  62008=>"111011110",
  62009=>"110001001",
  62010=>"100001110",
  62011=>"111101100",
  62012=>"100100100",
  62013=>"101100011",
  62014=>"011010010",
  62015=>"111011101",
  62016=>"001000000",
  62017=>"000101111",
  62018=>"111010101",
  62019=>"010011100",
  62020=>"100010111",
  62021=>"000111001",
  62022=>"110100000",
  62023=>"101000011",
  62024=>"000001001",
  62025=>"011110001",
  62026=>"111110011",
  62027=>"011100101",
  62028=>"000100001",
  62029=>"100111100",
  62030=>"011011111",
  62031=>"000001010",
  62032=>"111001000",
  62033=>"010111101",
  62034=>"000001001",
  62035=>"011000110",
  62036=>"010000110",
  62037=>"100010111",
  62038=>"000001000",
  62039=>"111111111",
  62040=>"000111111",
  62041=>"001000001",
  62042=>"010000110",
  62043=>"001101011",
  62044=>"010101001",
  62045=>"000000100",
  62046=>"000100001",
  62047=>"011001111",
  62048=>"001011110",
  62049=>"111110100",
  62050=>"010111011",
  62051=>"101010110",
  62052=>"101001100",
  62053=>"001000110",
  62054=>"100111100",
  62055=>"110111111",
  62056=>"111000011",
  62057=>"000101100",
  62058=>"011101110",
  62059=>"010101100",
  62060=>"101110011",
  62061=>"100010001",
  62062=>"010011111",
  62063=>"101100001",
  62064=>"100011110",
  62065=>"101001111",
  62066=>"111001010",
  62067=>"000000100",
  62068=>"010111100",
  62069=>"110011111",
  62070=>"100100100",
  62071=>"001011010",
  62072=>"101001010",
  62073=>"001000000",
  62074=>"001100001",
  62075=>"110011011",
  62076=>"110111011",
  62077=>"100010000",
  62078=>"011011100",
  62079=>"001011110",
  62080=>"000010001",
  62081=>"100111111",
  62082=>"000000010",
  62083=>"100010010",
  62084=>"100110111",
  62085=>"100001110",
  62086=>"011010111",
  62087=>"101110100",
  62088=>"011001101",
  62089=>"110000011",
  62090=>"001011101",
  62091=>"000011011",
  62092=>"010000110",
  62093=>"111110101",
  62094=>"010001000",
  62095=>"010000011",
  62096=>"100100100",
  62097=>"110100000",
  62098=>"110011110",
  62099=>"100111011",
  62100=>"111100101",
  62101=>"101111000",
  62102=>"000010110",
  62103=>"001010001",
  62104=>"111011001",
  62105=>"110010000",
  62106=>"101101010",
  62107=>"110000001",
  62108=>"000101001",
  62109=>"000000011",
  62110=>"000000110",
  62111=>"001100000",
  62112=>"100101111",
  62113=>"000100000",
  62114=>"100100100",
  62115=>"100001110",
  62116=>"011101111",
  62117=>"000111000",
  62118=>"000100000",
  62119=>"010100010",
  62120=>"110001100",
  62121=>"101100000",
  62122=>"101001111",
  62123=>"001110000",
  62124=>"100011110",
  62125=>"001000000",
  62126=>"101110001",
  62127=>"110011110",
  62128=>"010111001",
  62129=>"001000011",
  62130=>"000001100",
  62131=>"010001100",
  62132=>"000000001",
  62133=>"010001011",
  62134=>"010111100",
  62135=>"010001101",
  62136=>"000110011",
  62137=>"001110001",
  62138=>"100010100",
  62139=>"001000110",
  62140=>"000011100",
  62141=>"001100000",
  62142=>"010110111",
  62143=>"011001100",
  62144=>"010100101",
  62145=>"100100111",
  62146=>"110011011",
  62147=>"110010100",
  62148=>"000000011",
  62149=>"000100111",
  62150=>"101110110",
  62151=>"000011101",
  62152=>"001111001",
  62153=>"000101110",
  62154=>"110101001",
  62155=>"101100011",
  62156=>"000100000",
  62157=>"110011101",
  62158=>"010000000",
  62159=>"000110101",
  62160=>"011001000",
  62161=>"010000111",
  62162=>"011110011",
  62163=>"010001001",
  62164=>"110000111",
  62165=>"100010100",
  62166=>"010100100",
  62167=>"111011111",
  62168=>"001000100",
  62169=>"000000100",
  62170=>"111111001",
  62171=>"100111010",
  62172=>"111100111",
  62173=>"111100011",
  62174=>"001010101",
  62175=>"111111011",
  62176=>"000111100",
  62177=>"110110101",
  62178=>"110110010",
  62179=>"110111011",
  62180=>"000101001",
  62181=>"111101010",
  62182=>"101101000",
  62183=>"000000001",
  62184=>"010110100",
  62185=>"110101101",
  62186=>"001110010",
  62187=>"101000100",
  62188=>"000110100",
  62189=>"001101110",
  62190=>"100000110",
  62191=>"011111100",
  62192=>"001001110",
  62193=>"001100101",
  62194=>"011110001",
  62195=>"000100110",
  62196=>"110101110",
  62197=>"010100011",
  62198=>"000011101",
  62199=>"110000100",
  62200=>"010000110",
  62201=>"101100010",
  62202=>"111101010",
  62203=>"000000010",
  62204=>"110110101",
  62205=>"111010001",
  62206=>"100101111",
  62207=>"001110111",
  62208=>"000110101",
  62209=>"001110010",
  62210=>"110110010",
  62211=>"101010110",
  62212=>"000101100",
  62213=>"101000010",
  62214=>"111100001",
  62215=>"100101100",
  62216=>"010111111",
  62217=>"000010000",
  62218=>"001010001",
  62219=>"011011111",
  62220=>"000000001",
  62221=>"110110110",
  62222=>"100001001",
  62223=>"100011011",
  62224=>"100111110",
  62225=>"000011101",
  62226=>"100000111",
  62227=>"001111111",
  62228=>"010110000",
  62229=>"101000111",
  62230=>"100101000",
  62231=>"010101001",
  62232=>"010110011",
  62233=>"000001100",
  62234=>"000010011",
  62235=>"111000100",
  62236=>"000110011",
  62237=>"100111011",
  62238=>"000100111",
  62239=>"100000100",
  62240=>"101111111",
  62241=>"111000000",
  62242=>"111110011",
  62243=>"111010101",
  62244=>"111101111",
  62245=>"110101111",
  62246=>"011110111",
  62247=>"110111100",
  62248=>"011010001",
  62249=>"000100101",
  62250=>"001100110",
  62251=>"111001100",
  62252=>"110111011",
  62253=>"111011101",
  62254=>"001000001",
  62255=>"111010110",
  62256=>"010101100",
  62257=>"100111101",
  62258=>"001100100",
  62259=>"011111111",
  62260=>"000001110",
  62261=>"100010001",
  62262=>"101000000",
  62263=>"110100111",
  62264=>"011100111",
  62265=>"010011110",
  62266=>"010110101",
  62267=>"001100000",
  62268=>"100101000",
  62269=>"000010111",
  62270=>"000110111",
  62271=>"100000101",
  62272=>"100001111",
  62273=>"111110011",
  62274=>"101111110",
  62275=>"110000111",
  62276=>"101100000",
  62277=>"001010101",
  62278=>"110110001",
  62279=>"100101011",
  62280=>"100100110",
  62281=>"100101110",
  62282=>"000111011",
  62283=>"111101100",
  62284=>"001001010",
  62285=>"011101011",
  62286=>"100000011",
  62287=>"110111111",
  62288=>"000001011",
  62289=>"011111001",
  62290=>"011100000",
  62291=>"000000011",
  62292=>"011101111",
  62293=>"001000001",
  62294=>"111101001",
  62295=>"100010010",
  62296=>"000110011",
  62297=>"101110011",
  62298=>"111000111",
  62299=>"100111101",
  62300=>"111000011",
  62301=>"100110001",
  62302=>"100101110",
  62303=>"010011100",
  62304=>"110100000",
  62305=>"001101110",
  62306=>"100100100",
  62307=>"100001010",
  62308=>"100001111",
  62309=>"110100001",
  62310=>"100110010",
  62311=>"100010001",
  62312=>"111111111",
  62313=>"000110111",
  62314=>"011111011",
  62315=>"101101111",
  62316=>"010000001",
  62317=>"000000010",
  62318=>"100011001",
  62319=>"101001011",
  62320=>"001011100",
  62321=>"000100111",
  62322=>"011011010",
  62323=>"100101000",
  62324=>"001001010",
  62325=>"000010001",
  62326=>"001111110",
  62327=>"010101010",
  62328=>"011000010",
  62329=>"100100011",
  62330=>"111101100",
  62331=>"011011010",
  62332=>"000000111",
  62333=>"011111111",
  62334=>"011000110",
  62335=>"111100110",
  62336=>"011110001",
  62337=>"010100101",
  62338=>"101010111",
  62339=>"100000001",
  62340=>"010010100",
  62341=>"001101101",
  62342=>"010110001",
  62343=>"001010001",
  62344=>"010100010",
  62345=>"010010010",
  62346=>"101101010",
  62347=>"101111111",
  62348=>"010100100",
  62349=>"011110000",
  62350=>"010110111",
  62351=>"000100010",
  62352=>"011001001",
  62353=>"011111101",
  62354=>"000010101",
  62355=>"111110100",
  62356=>"100011000",
  62357=>"011010111",
  62358=>"000101011",
  62359=>"111100001",
  62360=>"011101111",
  62361=>"100111111",
  62362=>"101011000",
  62363=>"010010001",
  62364=>"111010101",
  62365=>"100101000",
  62366=>"011011100",
  62367=>"001011101",
  62368=>"101110010",
  62369=>"111000100",
  62370=>"101111000",
  62371=>"001101111",
  62372=>"010010010",
  62373=>"011101010",
  62374=>"101001100",
  62375=>"101001000",
  62376=>"000101001",
  62377=>"111110011",
  62378=>"010000010",
  62379=>"101010001",
  62380=>"011000010",
  62381=>"001010001",
  62382=>"011101001",
  62383=>"000000010",
  62384=>"110100000",
  62385=>"101110000",
  62386=>"000000001",
  62387=>"000000110",
  62388=>"101101001",
  62389=>"011100100",
  62390=>"011110111",
  62391=>"000001100",
  62392=>"110001101",
  62393=>"110001111",
  62394=>"010111000",
  62395=>"101110000",
  62396=>"110111000",
  62397=>"100101100",
  62398=>"000100000",
  62399=>"001101010",
  62400=>"101111111",
  62401=>"011100010",
  62402=>"100000101",
  62403=>"001101001",
  62404=>"010111100",
  62405=>"000000101",
  62406=>"100011001",
  62407=>"011111010",
  62408=>"001010000",
  62409=>"111110111",
  62410=>"001001000",
  62411=>"011110101",
  62412=>"111001010",
  62413=>"110001000",
  62414=>"110101101",
  62415=>"011001011",
  62416=>"111000110",
  62417=>"011101000",
  62418=>"000101100",
  62419=>"001101000",
  62420=>"101010001",
  62421=>"101101000",
  62422=>"110100100",
  62423=>"011000011",
  62424=>"000101100",
  62425=>"100110110",
  62426=>"100110111",
  62427=>"111001111",
  62428=>"010010001",
  62429=>"101101000",
  62430=>"010011100",
  62431=>"110111110",
  62432=>"101111010",
  62433=>"001110111",
  62434=>"110101111",
  62435=>"110111011",
  62436=>"001001110",
  62437=>"001000011",
  62438=>"010100001",
  62439=>"010011101",
  62440=>"101100110",
  62441=>"000001111",
  62442=>"000001101",
  62443=>"001010011",
  62444=>"110010001",
  62445=>"000000001",
  62446=>"101111001",
  62447=>"000101000",
  62448=>"000010001",
  62449=>"110011000",
  62450=>"101010110",
  62451=>"010101000",
  62452=>"111110010",
  62453=>"000101011",
  62454=>"100111110",
  62455=>"010010001",
  62456=>"111111101",
  62457=>"010110101",
  62458=>"110000001",
  62459=>"110011001",
  62460=>"100101001",
  62461=>"101101101",
  62462=>"010101011",
  62463=>"110110111",
  62464=>"010111101",
  62465=>"000101000",
  62466=>"001100110",
  62467=>"110011010",
  62468=>"101101100",
  62469=>"110110010",
  62470=>"100001011",
  62471=>"011111100",
  62472=>"110101011",
  62473=>"000111011",
  62474=>"001101011",
  62475=>"010100110",
  62476=>"011001101",
  62477=>"000001101",
  62478=>"011011111",
  62479=>"111101111",
  62480=>"100101100",
  62481=>"100110111",
  62482=>"011100000",
  62483=>"011110100",
  62484=>"101101110",
  62485=>"100111011",
  62486=>"100101101",
  62487=>"001101101",
  62488=>"011110110",
  62489=>"111011000",
  62490=>"010100110",
  62491=>"100101011",
  62492=>"100110001",
  62493=>"010100101",
  62494=>"010001101",
  62495=>"111000110",
  62496=>"001110001",
  62497=>"000110011",
  62498=>"100000000",
  62499=>"100100101",
  62500=>"000000001",
  62501=>"000000110",
  62502=>"101001001",
  62503=>"110010010",
  62504=>"111000100",
  62505=>"000001101",
  62506=>"111101010",
  62507=>"101011100",
  62508=>"100000001",
  62509=>"101110100",
  62510=>"110000100",
  62511=>"101011010",
  62512=>"101101111",
  62513=>"100111100",
  62514=>"011111011",
  62515=>"001001111",
  62516=>"111011001",
  62517=>"001110000",
  62518=>"000001101",
  62519=>"101010111",
  62520=>"000011100",
  62521=>"011101000",
  62522=>"100111000",
  62523=>"010001100",
  62524=>"100100000",
  62525=>"011001101",
  62526=>"111000001",
  62527=>"110110110",
  62528=>"101000111",
  62529=>"110111001",
  62530=>"100111100",
  62531=>"110110001",
  62532=>"100110100",
  62533=>"100010101",
  62534=>"001101111",
  62535=>"001100111",
  62536=>"010000010",
  62537=>"001001010",
  62538=>"001101100",
  62539=>"101101101",
  62540=>"000110101",
  62541=>"100101001",
  62542=>"000000010",
  62543=>"110101101",
  62544=>"011101110",
  62545=>"001111111",
  62546=>"101011000",
  62547=>"000101100",
  62548=>"000110000",
  62549=>"011010001",
  62550=>"110100101",
  62551=>"000100101",
  62552=>"010010011",
  62553=>"010111001",
  62554=>"101111110",
  62555=>"100001110",
  62556=>"111111110",
  62557=>"111110100",
  62558=>"011010101",
  62559=>"110110111",
  62560=>"001111101",
  62561=>"111110101",
  62562=>"100010111",
  62563=>"110111111",
  62564=>"000100001",
  62565=>"111100110",
  62566=>"001001110",
  62567=>"100010100",
  62568=>"100100110",
  62569=>"110111111",
  62570=>"000011100",
  62571=>"001111010",
  62572=>"101000110",
  62573=>"111101001",
  62574=>"011001001",
  62575=>"010001101",
  62576=>"011111001",
  62577=>"011111111",
  62578=>"111101101",
  62579=>"000111010",
  62580=>"111110111",
  62581=>"101011101",
  62582=>"011111110",
  62583=>"100100100",
  62584=>"111110011",
  62585=>"110111011",
  62586=>"000111111",
  62587=>"101101111",
  62588=>"101100100",
  62589=>"110001110",
  62590=>"110001011",
  62591=>"101111011",
  62592=>"011101011",
  62593=>"110001001",
  62594=>"100100010",
  62595=>"111101000",
  62596=>"101000010",
  62597=>"101111001",
  62598=>"001000101",
  62599=>"001010010",
  62600=>"001001011",
  62601=>"010000111",
  62602=>"100100000",
  62603=>"110100100",
  62604=>"100010010",
  62605=>"000101101",
  62606=>"010101101",
  62607=>"110010100",
  62608=>"000000111",
  62609=>"011001011",
  62610=>"000001011",
  62611=>"111100110",
  62612=>"011001001",
  62613=>"111111110",
  62614=>"101010111",
  62615=>"010000000",
  62616=>"000101000",
  62617=>"010010010",
  62618=>"011111001",
  62619=>"010111100",
  62620=>"110110000",
  62621=>"000000010",
  62622=>"101100101",
  62623=>"110101001",
  62624=>"001111110",
  62625=>"110010101",
  62626=>"001001101",
  62627=>"000010101",
  62628=>"101110100",
  62629=>"001101110",
  62630=>"110101100",
  62631=>"001001110",
  62632=>"011011100",
  62633=>"011111010",
  62634=>"100111110",
  62635=>"011010000",
  62636=>"111011011",
  62637=>"110101100",
  62638=>"011001000",
  62639=>"000100011",
  62640=>"010011011",
  62641=>"100011000",
  62642=>"111110100",
  62643=>"100100101",
  62644=>"000000000",
  62645=>"000000010",
  62646=>"010111111",
  62647=>"111000100",
  62648=>"011000111",
  62649=>"110100000",
  62650=>"111011001",
  62651=>"010100111",
  62652=>"000000100",
  62653=>"001010000",
  62654=>"000100000",
  62655=>"001100000",
  62656=>"010000000",
  62657=>"010000011",
  62658=>"000100101",
  62659=>"111111101",
  62660=>"010101101",
  62661=>"010101110",
  62662=>"111100100",
  62663=>"011001111",
  62664=>"001000100",
  62665=>"010111000",
  62666=>"010100100",
  62667=>"011110000",
  62668=>"001111000",
  62669=>"011000111",
  62670=>"111000010",
  62671=>"010101110",
  62672=>"111011101",
  62673=>"010110000",
  62674=>"101111010",
  62675=>"111010110",
  62676=>"100000100",
  62677=>"100101111",
  62678=>"100011101",
  62679=>"011010101",
  62680=>"111011011",
  62681=>"001101001",
  62682=>"011100000",
  62683=>"000000101",
  62684=>"010011111",
  62685=>"111001011",
  62686=>"100000000",
  62687=>"000111001",
  62688=>"110000010",
  62689=>"000010001",
  62690=>"101111011",
  62691=>"101101110",
  62692=>"011100010",
  62693=>"000110001",
  62694=>"010110100",
  62695=>"111111100",
  62696=>"111101011",
  62697=>"010000100",
  62698=>"010010111",
  62699=>"100100100",
  62700=>"100000010",
  62701=>"000000001",
  62702=>"101011011",
  62703=>"101111111",
  62704=>"011000110",
  62705=>"001111000",
  62706=>"110110011",
  62707=>"010111011",
  62708=>"111001100",
  62709=>"000110101",
  62710=>"011000000",
  62711=>"001000000",
  62712=>"101111111",
  62713=>"100110110",
  62714=>"011000010",
  62715=>"010101000",
  62716=>"111100111",
  62717=>"010011001",
  62718=>"100110001",
  62719=>"100101110",
  62720=>"110011001",
  62721=>"010110111",
  62722=>"111000000",
  62723=>"011001101",
  62724=>"101010001",
  62725=>"110011110",
  62726=>"010111101",
  62727=>"110000001",
  62728=>"011001000",
  62729=>"110101110",
  62730=>"110110100",
  62731=>"011010010",
  62732=>"101110100",
  62733=>"010110111",
  62734=>"100001100",
  62735=>"011101000",
  62736=>"001101100",
  62737=>"111111000",
  62738=>"010101001",
  62739=>"010010011",
  62740=>"101101101",
  62741=>"111011011",
  62742=>"110101101",
  62743=>"101111010",
  62744=>"100011000",
  62745=>"101011110",
  62746=>"100010000",
  62747=>"101010000",
  62748=>"000000010",
  62749=>"100101011",
  62750=>"010011010",
  62751=>"011111011",
  62752=>"010000001",
  62753=>"100010000",
  62754=>"010110000",
  62755=>"010100011",
  62756=>"110011100",
  62757=>"011000000",
  62758=>"100010000",
  62759=>"110001000",
  62760=>"001001011",
  62761=>"011010111",
  62762=>"010111111",
  62763=>"111011111",
  62764=>"010000011",
  62765=>"010010100",
  62766=>"010101000",
  62767=>"000110111",
  62768=>"110100101",
  62769=>"010111011",
  62770=>"100000001",
  62771=>"101001011",
  62772=>"110111101",
  62773=>"000001100",
  62774=>"110100100",
  62775=>"010011100",
  62776=>"010100010",
  62777=>"001010011",
  62778=>"100010011",
  62779=>"010110010",
  62780=>"110001011",
  62781=>"101100111",
  62782=>"010100000",
  62783=>"101100101",
  62784=>"110001000",
  62785=>"001001110",
  62786=>"000101000",
  62787=>"100110011",
  62788=>"111001101",
  62789=>"011001111",
  62790=>"101000111",
  62791=>"111011111",
  62792=>"110001010",
  62793=>"100100111",
  62794=>"101100000",
  62795=>"101111101",
  62796=>"110001000",
  62797=>"101000110",
  62798=>"101110110",
  62799=>"001111100",
  62800=>"001110110",
  62801=>"101100111",
  62802=>"111111011",
  62803=>"011101001",
  62804=>"000101001",
  62805=>"001111100",
  62806=>"110011100",
  62807=>"101110000",
  62808=>"111111101",
  62809=>"001111100",
  62810=>"110011101",
  62811=>"101000110",
  62812=>"111011100",
  62813=>"100010000",
  62814=>"110101001",
  62815=>"001100011",
  62816=>"000000100",
  62817=>"000011111",
  62818=>"000000001",
  62819=>"010000011",
  62820=>"000111100",
  62821=>"000000011",
  62822=>"100000110",
  62823=>"010000110",
  62824=>"000111101",
  62825=>"011010011",
  62826=>"110010111",
  62827=>"110001101",
  62828=>"001000110",
  62829=>"100001111",
  62830=>"111010111",
  62831=>"000110011",
  62832=>"010000011",
  62833=>"010101011",
  62834=>"000101000",
  62835=>"110000100",
  62836=>"010011000",
  62837=>"011111010",
  62838=>"111000001",
  62839=>"000110101",
  62840=>"100011101",
  62841=>"110111001",
  62842=>"000100000",
  62843=>"110011110",
  62844=>"111000000",
  62845=>"110111011",
  62846=>"011101011",
  62847=>"100000100",
  62848=>"000001111",
  62849=>"010000000",
  62850=>"000101001",
  62851=>"001110000",
  62852=>"100100011",
  62853=>"010111011",
  62854=>"110110100",
  62855=>"100000000",
  62856=>"100000101",
  62857=>"010100100",
  62858=>"011010101",
  62859=>"111010001",
  62860=>"010011100",
  62861=>"100000000",
  62862=>"101001111",
  62863=>"000111011",
  62864=>"100101011",
  62865=>"001011110",
  62866=>"011010011",
  62867=>"011110010",
  62868=>"110010010",
  62869=>"111001011",
  62870=>"000110010",
  62871=>"011101110",
  62872=>"000000001",
  62873=>"110000101",
  62874=>"110100010",
  62875=>"011001111",
  62876=>"011110000",
  62877=>"000000011",
  62878=>"100001100",
  62879=>"011011101",
  62880=>"100001001",
  62881=>"111000111",
  62882=>"001111111",
  62883=>"010010001",
  62884=>"101000000",
  62885=>"001000100",
  62886=>"111000000",
  62887=>"010101100",
  62888=>"001011110",
  62889=>"011000101",
  62890=>"000000010",
  62891=>"101000010",
  62892=>"100001101",
  62893=>"000011001",
  62894=>"111000011",
  62895=>"110110011",
  62896=>"100101000",
  62897=>"000000100",
  62898=>"001110111",
  62899=>"011010111",
  62900=>"011110010",
  62901=>"010111010",
  62902=>"100111011",
  62903=>"000100100",
  62904=>"100001111",
  62905=>"111101101",
  62906=>"101010110",
  62907=>"101101000",
  62908=>"100110000",
  62909=>"000111101",
  62910=>"110000001",
  62911=>"110010100",
  62912=>"010110111",
  62913=>"101011000",
  62914=>"111100110",
  62915=>"000100101",
  62916=>"000111001",
  62917=>"011010100",
  62918=>"000001110",
  62919=>"100101101",
  62920=>"111010111",
  62921=>"010000011",
  62922=>"000001110",
  62923=>"110010111",
  62924=>"111111001",
  62925=>"110110100",
  62926=>"000000011",
  62927=>"101000011",
  62928=>"110111001",
  62929=>"001110111",
  62930=>"001011101",
  62931=>"011001010",
  62932=>"000101010",
  62933=>"110100000",
  62934=>"100001010",
  62935=>"000000110",
  62936=>"000010000",
  62937=>"110111010",
  62938=>"101101100",
  62939=>"101001000",
  62940=>"110111001",
  62941=>"111101111",
  62942=>"110111101",
  62943=>"010010001",
  62944=>"111100011",
  62945=>"111110011",
  62946=>"011011111",
  62947=>"011010100",
  62948=>"111101001",
  62949=>"000010001",
  62950=>"110000101",
  62951=>"011000001",
  62952=>"101101110",
  62953=>"110100101",
  62954=>"100001011",
  62955=>"011011000",
  62956=>"101010101",
  62957=>"011100010",
  62958=>"000110101",
  62959=>"110100100",
  62960=>"000100100",
  62961=>"100000000",
  62962=>"110001111",
  62963=>"010010111",
  62964=>"101000011",
  62965=>"011000010",
  62966=>"010010001",
  62967=>"011000000",
  62968=>"000011100",
  62969=>"010101000",
  62970=>"000010110",
  62971=>"111000001",
  62972=>"000110110",
  62973=>"010111001",
  62974=>"110110000",
  62975=>"001010110",
  62976=>"101011100",
  62977=>"010100000",
  62978=>"010101101",
  62979=>"111111111",
  62980=>"101011110",
  62981=>"000110110",
  62982=>"100110011",
  62983=>"101000001",
  62984=>"010010000",
  62985=>"011111001",
  62986=>"111111110",
  62987=>"101000101",
  62988=>"100100010",
  62989=>"001110001",
  62990=>"000000101",
  62991=>"000111111",
  62992=>"101000111",
  62993=>"000100010",
  62994=>"110011000",
  62995=>"010010110",
  62996=>"010110001",
  62997=>"001000111",
  62998=>"110111001",
  62999=>"011010010",
  63000=>"101110000",
  63001=>"011011001",
  63002=>"011111101",
  63003=>"111001100",
  63004=>"000111111",
  63005=>"000001000",
  63006=>"000101000",
  63007=>"000100000",
  63008=>"011010110",
  63009=>"100101000",
  63010=>"001011110",
  63011=>"111000010",
  63012=>"001110010",
  63013=>"001000110",
  63014=>"111000101",
  63015=>"011000000",
  63016=>"101000111",
  63017=>"110110110",
  63018=>"011101110",
  63019=>"100111000",
  63020=>"010101000",
  63021=>"010010011",
  63022=>"000001011",
  63023=>"000011010",
  63024=>"011101001",
  63025=>"001101111",
  63026=>"101001110",
  63027=>"000100001",
  63028=>"001100001",
  63029=>"010000110",
  63030=>"100010101",
  63031=>"111011011",
  63032=>"010101100",
  63033=>"100001000",
  63034=>"001101010",
  63035=>"111101101",
  63036=>"111010010",
  63037=>"101001011",
  63038=>"110110011",
  63039=>"001100000",
  63040=>"111110001",
  63041=>"101001100",
  63042=>"010111011",
  63043=>"101110110",
  63044=>"110010000",
  63045=>"101111101",
  63046=>"010100011",
  63047=>"110011011",
  63048=>"111111000",
  63049=>"111010010",
  63050=>"100101100",
  63051=>"110001001",
  63052=>"000001011",
  63053=>"000011100",
  63054=>"100110101",
  63055=>"110010100",
  63056=>"001001111",
  63057=>"101101001",
  63058=>"011000110",
  63059=>"100110101",
  63060=>"100010111",
  63061=>"101111011",
  63062=>"101111001",
  63063=>"001001101",
  63064=>"101111100",
  63065=>"010011111",
  63066=>"111011001",
  63067=>"010010110",
  63068=>"000110011",
  63069=>"101010100",
  63070=>"101100110",
  63071=>"001010111",
  63072=>"010010010",
  63073=>"000101000",
  63074=>"000000010",
  63075=>"000000001",
  63076=>"100111010",
  63077=>"011110111",
  63078=>"110001111",
  63079=>"111000000",
  63080=>"011100010",
  63081=>"000001010",
  63082=>"101110111",
  63083=>"001100011",
  63084=>"001110111",
  63085=>"100011110",
  63086=>"000110101",
  63087=>"111001100",
  63088=>"010110010",
  63089=>"010000100",
  63090=>"111000101",
  63091=>"000000000",
  63092=>"000011011",
  63093=>"101101001",
  63094=>"110001100",
  63095=>"110000010",
  63096=>"011101100",
  63097=>"010010110",
  63098=>"101000001",
  63099=>"001000011",
  63100=>"010010101",
  63101=>"110000111",
  63102=>"001010101",
  63103=>"010010001",
  63104=>"110000000",
  63105=>"111010011",
  63106=>"000011010",
  63107=>"011010001",
  63108=>"110001111",
  63109=>"110101001",
  63110=>"101111001",
  63111=>"010011110",
  63112=>"100000110",
  63113=>"010010000",
  63114=>"100110101",
  63115=>"101111011",
  63116=>"000010011",
  63117=>"100111001",
  63118=>"001100001",
  63119=>"100011111",
  63120=>"100101001",
  63121=>"101010010",
  63122=>"111011100",
  63123=>"110011111",
  63124=>"011110110",
  63125=>"101011011",
  63126=>"111000000",
  63127=>"111111010",
  63128=>"011000011",
  63129=>"001110001",
  63130=>"001101011",
  63131=>"100111101",
  63132=>"010010100",
  63133=>"000111000",
  63134=>"000101000",
  63135=>"011000101",
  63136=>"000100110",
  63137=>"000001001",
  63138=>"110010110",
  63139=>"000100111",
  63140=>"111111111",
  63141=>"011000011",
  63142=>"011000100",
  63143=>"010111101",
  63144=>"110111010",
  63145=>"100111111",
  63146=>"111010000",
  63147=>"001100111",
  63148=>"111010001",
  63149=>"011011000",
  63150=>"111000001",
  63151=>"010110011",
  63152=>"100111101",
  63153=>"111100100",
  63154=>"100000010",
  63155=>"101000001",
  63156=>"011101000",
  63157=>"101101001",
  63158=>"011000010",
  63159=>"101101111",
  63160=>"000010011",
  63161=>"110100001",
  63162=>"110110000",
  63163=>"110100111",
  63164=>"110010001",
  63165=>"001111111",
  63166=>"010111100",
  63167=>"100100011",
  63168=>"111010001",
  63169=>"111110101",
  63170=>"111111011",
  63171=>"110111111",
  63172=>"001011101",
  63173=>"001111000",
  63174=>"111101110",
  63175=>"110100010",
  63176=>"001000000",
  63177=>"000010000",
  63178=>"011101110",
  63179=>"100101111",
  63180=>"001001110",
  63181=>"101000000",
  63182=>"000010001",
  63183=>"111011000",
  63184=>"000100011",
  63185=>"000000111",
  63186=>"100001001",
  63187=>"000000010",
  63188=>"100100111",
  63189=>"111111111",
  63190=>"111100101",
  63191=>"101001110",
  63192=>"100010000",
  63193=>"101001011",
  63194=>"000000110",
  63195=>"110110001",
  63196=>"010100101",
  63197=>"000000011",
  63198=>"111001100",
  63199=>"111010110",
  63200=>"001101111",
  63201=>"110100111",
  63202=>"000101111",
  63203=>"000100000",
  63204=>"000110011",
  63205=>"010001001",
  63206=>"111101110",
  63207=>"010100100",
  63208=>"100010000",
  63209=>"010100000",
  63210=>"101001111",
  63211=>"010110000",
  63212=>"011010111",
  63213=>"111011010",
  63214=>"111100110",
  63215=>"000101011",
  63216=>"110010010",
  63217=>"010011001",
  63218=>"100101000",
  63219=>"010110011",
  63220=>"001101110",
  63221=>"101011110",
  63222=>"110110011",
  63223=>"010101110",
  63224=>"011001001",
  63225=>"010110000",
  63226=>"001101001",
  63227=>"101010000",
  63228=>"110100011",
  63229=>"000011101",
  63230=>"001010110",
  63231=>"111011101",
  63232=>"111111110",
  63233=>"010000101",
  63234=>"010110111",
  63235=>"000100110",
  63236=>"011111111",
  63237=>"011101001",
  63238=>"011001000",
  63239=>"110011001",
  63240=>"101101000",
  63241=>"000100011",
  63242=>"111110110",
  63243=>"110111100",
  63244=>"010111010",
  63245=>"001011100",
  63246=>"100000101",
  63247=>"111101000",
  63248=>"100111110",
  63249=>"001111111",
  63250=>"111001000",
  63251=>"100010111",
  63252=>"011110110",
  63253=>"011101110",
  63254=>"000101101",
  63255=>"111101111",
  63256=>"000100101",
  63257=>"001101001",
  63258=>"110010100",
  63259=>"111000001",
  63260=>"101111001",
  63261=>"000110001",
  63262=>"010011010",
  63263=>"011010101",
  63264=>"000000000",
  63265=>"101000111",
  63266=>"010000100",
  63267=>"011011010",
  63268=>"101111000",
  63269=>"111100011",
  63270=>"111111100",
  63271=>"110110000",
  63272=>"011011111",
  63273=>"001100110",
  63274=>"011100101",
  63275=>"011010110",
  63276=>"011111111",
  63277=>"100110111",
  63278=>"001000101",
  63279=>"000001111",
  63280=>"001100010",
  63281=>"011111001",
  63282=>"010110001",
  63283=>"001101100",
  63284=>"101010000",
  63285=>"011110010",
  63286=>"111011110",
  63287=>"110100101",
  63288=>"100001101",
  63289=>"000111001",
  63290=>"100001100",
  63291=>"101001100",
  63292=>"000111101",
  63293=>"001100101",
  63294=>"000111101",
  63295=>"110010011",
  63296=>"001100101",
  63297=>"011001101",
  63298=>"010101011",
  63299=>"100101011",
  63300=>"100001001",
  63301=>"000101101",
  63302=>"101101100",
  63303=>"011110010",
  63304=>"101101100",
  63305=>"111111100",
  63306=>"001001000",
  63307=>"100100110",
  63308=>"011110000",
  63309=>"010000101",
  63310=>"001000110",
  63311=>"010100011",
  63312=>"000100000",
  63313=>"101010000",
  63314=>"010011111",
  63315=>"111111000",
  63316=>"101101101",
  63317=>"101110100",
  63318=>"011011110",
  63319=>"100111001",
  63320=>"110100110",
  63321=>"110000000",
  63322=>"101001011",
  63323=>"001011111",
  63324=>"101000011",
  63325=>"010111111",
  63326=>"011110100",
  63327=>"001000011",
  63328=>"111101111",
  63329=>"000011000",
  63330=>"001010011",
  63331=>"001010111",
  63332=>"011101101",
  63333=>"100011000",
  63334=>"110100000",
  63335=>"101000100",
  63336=>"100010100",
  63337=>"101110100",
  63338=>"000011100",
  63339=>"100010101",
  63340=>"101110001",
  63341=>"100111011",
  63342=>"111101111",
  63343=>"010101101",
  63344=>"010001010",
  63345=>"010110000",
  63346=>"001000111",
  63347=>"100011010",
  63348=>"001101110",
  63349=>"111010011",
  63350=>"000001110",
  63351=>"001000010",
  63352=>"110010001",
  63353=>"111111001",
  63354=>"110011001",
  63355=>"001001011",
  63356=>"101100111",
  63357=>"010010110",
  63358=>"010111111",
  63359=>"011101001",
  63360=>"011011110",
  63361=>"001011111",
  63362=>"000001010",
  63363=>"010010101",
  63364=>"100110101",
  63365=>"100010011",
  63366=>"000100000",
  63367=>"000001100",
  63368=>"111001100",
  63369=>"010101101",
  63370=>"011010111",
  63371=>"011001010",
  63372=>"000100011",
  63373=>"111000001",
  63374=>"011110100",
  63375=>"010010101",
  63376=>"001001101",
  63377=>"110000000",
  63378=>"000100101",
  63379=>"011110001",
  63380=>"000010010",
  63381=>"111110001",
  63382=>"000000010",
  63383=>"111111111",
  63384=>"110101111",
  63385=>"010100100",
  63386=>"011011100",
  63387=>"010010001",
  63388=>"000110100",
  63389=>"111111111",
  63390=>"001011111",
  63391=>"001100011",
  63392=>"110000100",
  63393=>"001000010",
  63394=>"110000000",
  63395=>"000110110",
  63396=>"000011010",
  63397=>"010000111",
  63398=>"100001100",
  63399=>"100000010",
  63400=>"001010001",
  63401=>"111001110",
  63402=>"010000111",
  63403=>"111111100",
  63404=>"111101110",
  63405=>"000001110",
  63406=>"011011100",
  63407=>"010111010",
  63408=>"110001000",
  63409=>"010011001",
  63410=>"111001001",
  63411=>"000001111",
  63412=>"101100110",
  63413=>"000011100",
  63414=>"110101110",
  63415=>"111101110",
  63416=>"100010110",
  63417=>"110010000",
  63418=>"101001111",
  63419=>"100111000",
  63420=>"000110011",
  63421=>"000000000",
  63422=>"100010010",
  63423=>"011000010",
  63424=>"100000101",
  63425=>"011010000",
  63426=>"001001011",
  63427=>"000001011",
  63428=>"101000011",
  63429=>"001010001",
  63430=>"111110000",
  63431=>"010101010",
  63432=>"101110011",
  63433=>"100101010",
  63434=>"110011010",
  63435=>"100110101",
  63436=>"101101111",
  63437=>"011000111",
  63438=>"110011010",
  63439=>"111000100",
  63440=>"101101010",
  63441=>"110101001",
  63442=>"011000101",
  63443=>"100100111",
  63444=>"010101101",
  63445=>"101101111",
  63446=>"100001000",
  63447=>"011100101",
  63448=>"100110010",
  63449=>"001110100",
  63450=>"111110101",
  63451=>"001011001",
  63452=>"000111101",
  63453=>"010000100",
  63454=>"110010000",
  63455=>"000111010",
  63456=>"001110011",
  63457=>"011111101",
  63458=>"001000100",
  63459=>"011010010",
  63460=>"000111111",
  63461=>"000101111",
  63462=>"100111110",
  63463=>"010001000",
  63464=>"011100001",
  63465=>"110101111",
  63466=>"000110111",
  63467=>"000111100",
  63468=>"011110010",
  63469=>"000101100",
  63470=>"111100101",
  63471=>"100000011",
  63472=>"110100110",
  63473=>"001101100",
  63474=>"111101000",
  63475=>"000111110",
  63476=>"011110011",
  63477=>"101110011",
  63478=>"011101100",
  63479=>"001100010",
  63480=>"111010110",
  63481=>"011011101",
  63482=>"101111101",
  63483=>"001111000",
  63484=>"101101111",
  63485=>"110100000",
  63486=>"011111111",
  63487=>"111010101",
  63488=>"010010000",
  63489=>"110110110",
  63490=>"000000100",
  63491=>"010010111",
  63492=>"110011011",
  63493=>"000111011",
  63494=>"111101000",
  63495=>"001001000",
  63496=>"110001111",
  63497=>"010110110",
  63498=>"010001010",
  63499=>"000110010",
  63500=>"101001110",
  63501=>"101111000",
  63502=>"110111010",
  63503=>"000000011",
  63504=>"001010011",
  63505=>"010111011",
  63506=>"110001011",
  63507=>"101001101",
  63508=>"011000010",
  63509=>"101111111",
  63510=>"001011101",
  63511=>"000000000",
  63512=>"110000110",
  63513=>"001001101",
  63514=>"001011000",
  63515=>"100011010",
  63516=>"110100011",
  63517=>"010000101",
  63518=>"111100001",
  63519=>"111001001",
  63520=>"001011011",
  63521=>"110000011",
  63522=>"000011000",
  63523=>"100111011",
  63524=>"101110000",
  63525=>"000000110",
  63526=>"100011000",
  63527=>"010100000",
  63528=>"011010101",
  63529=>"001011010",
  63530=>"000001100",
  63531=>"100011101",
  63532=>"010110000",
  63533=>"011000001",
  63534=>"111110000",
  63535=>"101101111",
  63536=>"011001001",
  63537=>"010000101",
  63538=>"110010110",
  63539=>"010011001",
  63540=>"100011010",
  63541=>"111000000",
  63542=>"001101111",
  63543=>"011110111",
  63544=>"100101110",
  63545=>"100111100",
  63546=>"001101011",
  63547=>"000000100",
  63548=>"110101010",
  63549=>"101011111",
  63550=>"101010000",
  63551=>"011110001",
  63552=>"111110110",
  63553=>"011000011",
  63554=>"000110101",
  63555=>"000101101",
  63556=>"111100111",
  63557=>"110101100",
  63558=>"101100100",
  63559=>"110000100",
  63560=>"011111000",
  63561=>"101011001",
  63562=>"100011000",
  63563=>"001101110",
  63564=>"001101111",
  63565=>"011001000",
  63566=>"011111001",
  63567=>"011001111",
  63568=>"010101010",
  63569=>"001101000",
  63570=>"101111011",
  63571=>"011100111",
  63572=>"101011000",
  63573=>"110010101",
  63574=>"101100001",
  63575=>"000001100",
  63576=>"001100101",
  63577=>"010011100",
  63578=>"010101011",
  63579=>"011000010",
  63580=>"110110111",
  63581=>"000001110",
  63582=>"001001111",
  63583=>"111000010",
  63584=>"000011001",
  63585=>"001011010",
  63586=>"001001000",
  63587=>"010101100",
  63588=>"111111010",
  63589=>"010000010",
  63590=>"111001011",
  63591=>"010100110",
  63592=>"000110001",
  63593=>"100000111",
  63594=>"010100011",
  63595=>"001110001",
  63596=>"101010110",
  63597=>"111111001",
  63598=>"110001101",
  63599=>"100000000",
  63600=>"000101111",
  63601=>"010101000",
  63602=>"000101011",
  63603=>"010100101",
  63604=>"010110110",
  63605=>"101111100",
  63606=>"111101110",
  63607=>"000111010",
  63608=>"000000101",
  63609=>"101011101",
  63610=>"011100111",
  63611=>"010111000",
  63612=>"100000100",
  63613=>"100110000",
  63614=>"011001011",
  63615=>"001110100",
  63616=>"001011110",
  63617=>"000100111",
  63618=>"000000010",
  63619=>"010110100",
  63620=>"111101010",
  63621=>"110000101",
  63622=>"101011000",
  63623=>"100110000",
  63624=>"000100100",
  63625=>"010111010",
  63626=>"110000100",
  63627=>"111001111",
  63628=>"101100001",
  63629=>"110010111",
  63630=>"011001111",
  63631=>"111110111",
  63632=>"101100001",
  63633=>"001001010",
  63634=>"100111001",
  63635=>"110110001",
  63636=>"001011100",
  63637=>"000011011",
  63638=>"001011111",
  63639=>"111000000",
  63640=>"000111001",
  63641=>"010100100",
  63642=>"111111011",
  63643=>"101010001",
  63644=>"100011101",
  63645=>"101011000",
  63646=>"100010010",
  63647=>"100100111",
  63648=>"000010010",
  63649=>"110110100",
  63650=>"010011100",
  63651=>"111101101",
  63652=>"011001101",
  63653=>"011101010",
  63654=>"100000110",
  63655=>"111111001",
  63656=>"110000010",
  63657=>"101111000",
  63658=>"111111100",
  63659=>"000110000",
  63660=>"000010110",
  63661=>"110110001",
  63662=>"011011111",
  63663=>"101100101",
  63664=>"000000010",
  63665=>"000000110",
  63666=>"100010010",
  63667=>"111010010",
  63668=>"000001110",
  63669=>"001000100",
  63670=>"011101010",
  63671=>"011101100",
  63672=>"001100110",
  63673=>"111111100",
  63674=>"010000000",
  63675=>"011111100",
  63676=>"011111110",
  63677=>"001101111",
  63678=>"101001100",
  63679=>"010010001",
  63680=>"100000101",
  63681=>"011011110",
  63682=>"000110010",
  63683=>"011011010",
  63684=>"110110010",
  63685=>"011000111",
  63686=>"001001100",
  63687=>"111100010",
  63688=>"001000001",
  63689=>"101101000",
  63690=>"101110010",
  63691=>"110100110",
  63692=>"011101011",
  63693=>"010000100",
  63694=>"010011011",
  63695=>"110010111",
  63696=>"011010000",
  63697=>"101000010",
  63698=>"000000001",
  63699=>"111000100",
  63700=>"010001111",
  63701=>"011000000",
  63702=>"001100001",
  63703=>"011001100",
  63704=>"011011001",
  63705=>"011110010",
  63706=>"110000011",
  63707=>"101011101",
  63708=>"111010000",
  63709=>"110100010",
  63710=>"110011011",
  63711=>"110011001",
  63712=>"110101100",
  63713=>"101101111",
  63714=>"101010111",
  63715=>"010111011",
  63716=>"101010000",
  63717=>"000110000",
  63718=>"111101100",
  63719=>"001001111",
  63720=>"110010110",
  63721=>"110110001",
  63722=>"101010111",
  63723=>"100101110",
  63724=>"100000001",
  63725=>"100001010",
  63726=>"111000011",
  63727=>"111001101",
  63728=>"110001110",
  63729=>"001110111",
  63730=>"100011000",
  63731=>"011000110",
  63732=>"110110110",
  63733=>"100000110",
  63734=>"101011111",
  63735=>"001100110",
  63736=>"101001010",
  63737=>"111011110",
  63738=>"011100111",
  63739=>"010011011",
  63740=>"100110110",
  63741=>"001001000",
  63742=>"100001100",
  63743=>"000010110",
  63744=>"101100111",
  63745=>"101111011",
  63746=>"100101000",
  63747=>"111001000",
  63748=>"100100011",
  63749=>"111110110",
  63750=>"010111100",
  63751=>"001101111",
  63752=>"101101010",
  63753=>"101100000",
  63754=>"011110000",
  63755=>"000010110",
  63756=>"100011010",
  63757=>"111000111",
  63758=>"010000100",
  63759=>"001011110",
  63760=>"010011011",
  63761=>"010000110",
  63762=>"111011110",
  63763=>"100010101",
  63764=>"001011101",
  63765=>"001000101",
  63766=>"000110001",
  63767=>"001010000",
  63768=>"011001111",
  63769=>"101011111",
  63770=>"111100110",
  63771=>"110100001",
  63772=>"011110100",
  63773=>"100100110",
  63774=>"100000100",
  63775=>"010110001",
  63776=>"001010100",
  63777=>"110010101",
  63778=>"110101101",
  63779=>"111110111",
  63780=>"100101111",
  63781=>"000010011",
  63782=>"001101101",
  63783=>"110101101",
  63784=>"001001111",
  63785=>"000010011",
  63786=>"101010001",
  63787=>"000010110",
  63788=>"110011100",
  63789=>"100011000",
  63790=>"111011111",
  63791=>"111000100",
  63792=>"000000100",
  63793=>"010001011",
  63794=>"001100110",
  63795=>"111011010",
  63796=>"111110011",
  63797=>"000001100",
  63798=>"101010101",
  63799=>"111100001",
  63800=>"001000001",
  63801=>"100000101",
  63802=>"000010000",
  63803=>"011011111",
  63804=>"011001010",
  63805=>"010000000",
  63806=>"001011100",
  63807=>"111110110",
  63808=>"101101101",
  63809=>"000010110",
  63810=>"000001001",
  63811=>"011000011",
  63812=>"011000000",
  63813=>"000011101",
  63814=>"111111001",
  63815=>"111100101",
  63816=>"101000001",
  63817=>"110101110",
  63818=>"001001011",
  63819=>"011010011",
  63820=>"011010010",
  63821=>"010001001",
  63822=>"101000001",
  63823=>"001101011",
  63824=>"100000000",
  63825=>"011000100",
  63826=>"010011100",
  63827=>"010101011",
  63828=>"001100000",
  63829=>"001100000",
  63830=>"000000001",
  63831=>"000011000",
  63832=>"010101110",
  63833=>"010011100",
  63834=>"000001111",
  63835=>"100111000",
  63836=>"000000111",
  63837=>"001010111",
  63838=>"110010001",
  63839=>"010000001",
  63840=>"110001000",
  63841=>"010000000",
  63842=>"001001111",
  63843=>"001011001",
  63844=>"000111110",
  63845=>"100011000",
  63846=>"011100101",
  63847=>"000010000",
  63848=>"000000111",
  63849=>"011000010",
  63850=>"001110001",
  63851=>"000111101",
  63852=>"110000000",
  63853=>"100001101",
  63854=>"101110100",
  63855=>"000000010",
  63856=>"110011011",
  63857=>"110010000",
  63858=>"111011111",
  63859=>"100100001",
  63860=>"101100110",
  63861=>"011010001",
  63862=>"011100000",
  63863=>"000001111",
  63864=>"000011101",
  63865=>"011111111",
  63866=>"110100011",
  63867=>"100110100",
  63868=>"100000001",
  63869=>"110100100",
  63870=>"001101010",
  63871=>"011001010",
  63872=>"010001010",
  63873=>"001101101",
  63874=>"001110101",
  63875=>"100101000",
  63876=>"011100011",
  63877=>"101110001",
  63878=>"101011010",
  63879=>"011010101",
  63880=>"010100101",
  63881=>"011000011",
  63882=>"011011111",
  63883=>"011110001",
  63884=>"010101100",
  63885=>"111100000",
  63886=>"000100100",
  63887=>"000100010",
  63888=>"110011111",
  63889=>"011101110",
  63890=>"010010110",
  63891=>"110011111",
  63892=>"010110010",
  63893=>"111111110",
  63894=>"001000010",
  63895=>"101010000",
  63896=>"000101001",
  63897=>"100000111",
  63898=>"000011010",
  63899=>"100001010",
  63900=>"001101000",
  63901=>"011101100",
  63902=>"100100000",
  63903=>"010001101",
  63904=>"000100000",
  63905=>"101010010",
  63906=>"010011110",
  63907=>"010001010",
  63908=>"011001111",
  63909=>"011001000",
  63910=>"110111011",
  63911=>"101100001",
  63912=>"000111111",
  63913=>"000010010",
  63914=>"000010110",
  63915=>"001101010",
  63916=>"001101011",
  63917=>"011101100",
  63918=>"000000001",
  63919=>"100111100",
  63920=>"001011101",
  63921=>"000010010",
  63922=>"101111001",
  63923=>"101100000",
  63924=>"001111000",
  63925=>"000100000",
  63926=>"101101000",
  63927=>"111101001",
  63928=>"001000101",
  63929=>"011010100",
  63930=>"011001000",
  63931=>"111011100",
  63932=>"101100100",
  63933=>"101110001",
  63934=>"100100010",
  63935=>"001001101",
  63936=>"010110001",
  63937=>"101000110",
  63938=>"001000101",
  63939=>"001011001",
  63940=>"101110000",
  63941=>"001000010",
  63942=>"100110000",
  63943=>"011101011",
  63944=>"011101111",
  63945=>"110111011",
  63946=>"101000000",
  63947=>"101011011",
  63948=>"000011110",
  63949=>"010010011",
  63950=>"100001110",
  63951=>"101001001",
  63952=>"110000010",
  63953=>"010100010",
  63954=>"000110110",
  63955=>"101011100",
  63956=>"001010100",
  63957=>"011000110",
  63958=>"010100111",
  63959=>"000001011",
  63960=>"101110000",
  63961=>"111100111",
  63962=>"101101110",
  63963=>"001100101",
  63964=>"011101011",
  63965=>"111001010",
  63966=>"110010011",
  63967=>"101000011",
  63968=>"100111011",
  63969=>"010010001",
  63970=>"101001111",
  63971=>"111111110",
  63972=>"011001101",
  63973=>"111101000",
  63974=>"111111100",
  63975=>"011101011",
  63976=>"000101111",
  63977=>"001101010",
  63978=>"101011000",
  63979=>"101111001",
  63980=>"111101111",
  63981=>"011110111",
  63982=>"110111000",
  63983=>"000000110",
  63984=>"111011110",
  63985=>"001111000",
  63986=>"111100000",
  63987=>"000011001",
  63988=>"100101101",
  63989=>"000110000",
  63990=>"101011111",
  63991=>"101011100",
  63992=>"100100001",
  63993=>"110000110",
  63994=>"100100111",
  63995=>"001101101",
  63996=>"001001100",
  63997=>"001000111",
  63998=>"000010111",
  63999=>"001110110",
  64000=>"100101011",
  64001=>"110000011",
  64002=>"111011111",
  64003=>"100101001",
  64004=>"111001111",
  64005=>"111100001",
  64006=>"000100000",
  64007=>"000000101",
  64008=>"010001111",
  64009=>"010110011",
  64010=>"000101011",
  64011=>"000101100",
  64012=>"100000101",
  64013=>"011000011",
  64014=>"110110011",
  64015=>"110011001",
  64016=>"110101001",
  64017=>"000000000",
  64018=>"100000111",
  64019=>"011101011",
  64020=>"101110011",
  64021=>"111000000",
  64022=>"111011110",
  64023=>"000010111",
  64024=>"100100111",
  64025=>"011111111",
  64026=>"011101001",
  64027=>"111011100",
  64028=>"001111111",
  64029=>"000010110",
  64030=>"110000111",
  64031=>"111110010",
  64032=>"001010110",
  64033=>"111001010",
  64034=>"001011111",
  64035=>"011111110",
  64036=>"110010110",
  64037=>"110100100",
  64038=>"000000000",
  64039=>"011010110",
  64040=>"111000001",
  64041=>"100110111",
  64042=>"000000111",
  64043=>"011001110",
  64044=>"001011011",
  64045=>"110111000",
  64046=>"011011111",
  64047=>"111101000",
  64048=>"010101001",
  64049=>"111111111",
  64050=>"000000110",
  64051=>"000100101",
  64052=>"110011010",
  64053=>"100010100",
  64054=>"001011111",
  64055=>"110101100",
  64056=>"100001011",
  64057=>"001000111",
  64058=>"110011100",
  64059=>"000111110",
  64060=>"111110011",
  64061=>"000001100",
  64062=>"101111011",
  64063=>"001001100",
  64064=>"011100010",
  64065=>"000101011",
  64066=>"000101101",
  64067=>"000101010",
  64068=>"011100010",
  64069=>"010100100",
  64070=>"010001011",
  64071=>"010100100",
  64072=>"100010000",
  64073=>"000110000",
  64074=>"111111110",
  64075=>"010111100",
  64076=>"000011111",
  64077=>"101110100",
  64078=>"001010000",
  64079=>"100000110",
  64080=>"000000010",
  64081=>"111111001",
  64082=>"001001110",
  64083=>"000010010",
  64084=>"100110001",
  64085=>"000010001",
  64086=>"000000101",
  64087=>"101001100",
  64088=>"101101010",
  64089=>"100000111",
  64090=>"101110101",
  64091=>"101010101",
  64092=>"011011011",
  64093=>"000000110",
  64094=>"000111001",
  64095=>"111111010",
  64096=>"101110011",
  64097=>"010110000",
  64098=>"110000010",
  64099=>"011110011",
  64100=>"011101110",
  64101=>"001101000",
  64102=>"111111101",
  64103=>"100001000",
  64104=>"101000110",
  64105=>"001100110",
  64106=>"001011000",
  64107=>"011001011",
  64108=>"000110000",
  64109=>"100101010",
  64110=>"011100001",
  64111=>"110101011",
  64112=>"000100101",
  64113=>"000111001",
  64114=>"100101110",
  64115=>"110001111",
  64116=>"011110101",
  64117=>"111110100",
  64118=>"111111011",
  64119=>"100011001",
  64120=>"000000111",
  64121=>"010000001",
  64122=>"101010101",
  64123=>"000010010",
  64124=>"010010011",
  64125=>"100010100",
  64126=>"110101101",
  64127=>"010100111",
  64128=>"011001011",
  64129=>"111110110",
  64130=>"001011101",
  64131=>"101000011",
  64132=>"001111010",
  64133=>"001100011",
  64134=>"001100111",
  64135=>"100100110",
  64136=>"001111100",
  64137=>"100001001",
  64138=>"011011010",
  64139=>"110111010",
  64140=>"001110110",
  64141=>"101111011",
  64142=>"001111101",
  64143=>"010000010",
  64144=>"011101001",
  64145=>"100111100",
  64146=>"111001011",
  64147=>"110010000",
  64148=>"010111001",
  64149=>"111111110",
  64150=>"001110000",
  64151=>"000101001",
  64152=>"101110010",
  64153=>"001011111",
  64154=>"001110100",
  64155=>"001011111",
  64156=>"000001101",
  64157=>"100001001",
  64158=>"011100001",
  64159=>"011000000",
  64160=>"001001000",
  64161=>"110111000",
  64162=>"111100101",
  64163=>"110000100",
  64164=>"101000010",
  64165=>"001010010",
  64166=>"101000100",
  64167=>"101001001",
  64168=>"000100010",
  64169=>"100100011",
  64170=>"100000110",
  64171=>"001011110",
  64172=>"100000001",
  64173=>"111010010",
  64174=>"100010100",
  64175=>"110010000",
  64176=>"100001000",
  64177=>"010110110",
  64178=>"010100111",
  64179=>"100010011",
  64180=>"001101100",
  64181=>"110111011",
  64182=>"100100101",
  64183=>"110011010",
  64184=>"010111111",
  64185=>"110000011",
  64186=>"101101100",
  64187=>"110111101",
  64188=>"100100011",
  64189=>"111011000",
  64190=>"001100100",
  64191=>"101010110",
  64192=>"111001110",
  64193=>"100100101",
  64194=>"010110111",
  64195=>"111100111",
  64196=>"000101101",
  64197=>"111011011",
  64198=>"101010110",
  64199=>"101110110",
  64200=>"000010000",
  64201=>"011000111",
  64202=>"101111111",
  64203=>"111001110",
  64204=>"101110110",
  64205=>"100100101",
  64206=>"111011000",
  64207=>"110011111",
  64208=>"010101100",
  64209=>"010010010",
  64210=>"100010000",
  64211=>"101011001",
  64212=>"100111100",
  64213=>"000000000",
  64214=>"101111100",
  64215=>"011000001",
  64216=>"001000100",
  64217=>"110000101",
  64218=>"011100001",
  64219=>"111011000",
  64220=>"000000111",
  64221=>"001111011",
  64222=>"111000010",
  64223=>"010001100",
  64224=>"110011110",
  64225=>"011101110",
  64226=>"011111111",
  64227=>"100110000",
  64228=>"101001101",
  64229=>"000010001",
  64230=>"001010110",
  64231=>"110010011",
  64232=>"000011100",
  64233=>"111111101",
  64234=>"010010101",
  64235=>"000011000",
  64236=>"110011111",
  64237=>"001011111",
  64238=>"111111110",
  64239=>"000100100",
  64240=>"111101110",
  64241=>"000001011",
  64242=>"100011101",
  64243=>"010001010",
  64244=>"100101100",
  64245=>"101100110",
  64246=>"101100110",
  64247=>"110100001",
  64248=>"001010100",
  64249=>"001110111",
  64250=>"100111110",
  64251=>"010010010",
  64252=>"010101101",
  64253=>"110000000",
  64254=>"101101010",
  64255=>"000110001",
  64256=>"011100011",
  64257=>"111101100",
  64258=>"001110001",
  64259=>"011010111",
  64260=>"000111111",
  64261=>"011010010",
  64262=>"011101100",
  64263=>"010100011",
  64264=>"001010000",
  64265=>"110001001",
  64266=>"111001011",
  64267=>"001000100",
  64268=>"001110101",
  64269=>"101001001",
  64270=>"101001011",
  64271=>"000011011",
  64272=>"111000010",
  64273=>"100001011",
  64274=>"000001101",
  64275=>"001100100",
  64276=>"111100001",
  64277=>"000101010",
  64278=>"100110000",
  64279=>"011000001",
  64280=>"011000011",
  64281=>"010010001",
  64282=>"000100011",
  64283=>"101100010",
  64284=>"001101000",
  64285=>"011000101",
  64286=>"111011001",
  64287=>"110110111",
  64288=>"110101010",
  64289=>"000111100",
  64290=>"101110010",
  64291=>"100010110",
  64292=>"111101101",
  64293=>"011111111",
  64294=>"011100101",
  64295=>"111011001",
  64296=>"110000001",
  64297=>"011001100",
  64298=>"100110001",
  64299=>"101101010",
  64300=>"010000100",
  64301=>"011001101",
  64302=>"001100100",
  64303=>"100110000",
  64304=>"010101110",
  64305=>"100011001",
  64306=>"001010000",
  64307=>"010011010",
  64308=>"011000011",
  64309=>"010101100",
  64310=>"001010010",
  64311=>"000001011",
  64312=>"010000101",
  64313=>"011100110",
  64314=>"010000100",
  64315=>"010001001",
  64316=>"100001000",
  64317=>"111001001",
  64318=>"110001000",
  64319=>"000011000",
  64320=>"001001001",
  64321=>"101001100",
  64322=>"101101000",
  64323=>"100001110",
  64324=>"011110101",
  64325=>"101111010",
  64326=>"101010101",
  64327=>"011100010",
  64328=>"111101111",
  64329=>"000110101",
  64330=>"110110000",
  64331=>"110011101",
  64332=>"011101001",
  64333=>"101101010",
  64334=>"001101100",
  64335=>"011001100",
  64336=>"111111101",
  64337=>"110001011",
  64338=>"100010110",
  64339=>"100101001",
  64340=>"000110010",
  64341=>"011110101",
  64342=>"001011010",
  64343=>"000100000",
  64344=>"010010111",
  64345=>"100110001",
  64346=>"000101100",
  64347=>"000100111",
  64348=>"111101100",
  64349=>"101111110",
  64350=>"000011101",
  64351=>"110101010",
  64352=>"010111000",
  64353=>"011010011",
  64354=>"010010011",
  64355=>"111101011",
  64356=>"011010000",
  64357=>"000001011",
  64358=>"000010110",
  64359=>"011001111",
  64360=>"000010101",
  64361=>"110110000",
  64362=>"011001001",
  64363=>"000110000",
  64364=>"010001000",
  64365=>"101110001",
  64366=>"110111100",
  64367=>"111111111",
  64368=>"001111011",
  64369=>"001000010",
  64370=>"111001111",
  64371=>"111101001",
  64372=>"000111110",
  64373=>"000101110",
  64374=>"110111001",
  64375=>"110000100",
  64376=>"111001110",
  64377=>"011101111",
  64378=>"100111110",
  64379=>"110110100",
  64380=>"000110000",
  64381=>"001110111",
  64382=>"000101111",
  64383=>"111000000",
  64384=>"111110101",
  64385=>"111111000",
  64386=>"010111110",
  64387=>"000000011",
  64388=>"010111010",
  64389=>"010010001",
  64390=>"101001101",
  64391=>"111111100",
  64392=>"111110101",
  64393=>"110100011",
  64394=>"001010100",
  64395=>"101110010",
  64396=>"101010001",
  64397=>"110011111",
  64398=>"010100001",
  64399=>"101011111",
  64400=>"000011100",
  64401=>"111100111",
  64402=>"001100000",
  64403=>"001000000",
  64404=>"100011110",
  64405=>"010111101",
  64406=>"101111000",
  64407=>"001000011",
  64408=>"000101101",
  64409=>"111100111",
  64410=>"010101111",
  64411=>"110001111",
  64412=>"011000111",
  64413=>"010100100",
  64414=>"011001110",
  64415=>"001011010",
  64416=>"110010110",
  64417=>"101110111",
  64418=>"000000100",
  64419=>"111100010",
  64420=>"001111010",
  64421=>"111100010",
  64422=>"110001010",
  64423=>"001110001",
  64424=>"001110010",
  64425=>"010111010",
  64426=>"010000011",
  64427=>"001000110",
  64428=>"111001000",
  64429=>"011111111",
  64430=>"101101000",
  64431=>"101101111",
  64432=>"000011000",
  64433=>"110111000",
  64434=>"011010101",
  64435=>"010010101",
  64436=>"100010111",
  64437=>"011010101",
  64438=>"111101111",
  64439=>"101110111",
  64440=>"101100010",
  64441=>"000000010",
  64442=>"100011010",
  64443=>"000001100",
  64444=>"101010011",
  64445=>"000101001",
  64446=>"011111101",
  64447=>"011010110",
  64448=>"000110010",
  64449=>"111111001",
  64450=>"111101100",
  64451=>"100001001",
  64452=>"000100110",
  64453=>"001100111",
  64454=>"001100001",
  64455=>"011111110",
  64456=>"001010010",
  64457=>"101010000",
  64458=>"011010101",
  64459=>"100101100",
  64460=>"100111110",
  64461=>"100000001",
  64462=>"110000101",
  64463=>"010100100",
  64464=>"010010100",
  64465=>"110100111",
  64466=>"001000001",
  64467=>"111101001",
  64468=>"010011100",
  64469=>"101001000",
  64470=>"110100100",
  64471=>"000001010",
  64472=>"100001110",
  64473=>"101001101",
  64474=>"011101011",
  64475=>"110110111",
  64476=>"011110101",
  64477=>"111000000",
  64478=>"110101101",
  64479=>"011001111",
  64480=>"000100010",
  64481=>"000110001",
  64482=>"101100010",
  64483=>"011110001",
  64484=>"100010010",
  64485=>"110110010",
  64486=>"101000110",
  64487=>"100111001",
  64488=>"011011000",
  64489=>"110100010",
  64490=>"100110001",
  64491=>"101111001",
  64492=>"100011100",
  64493=>"101001111",
  64494=>"000100110",
  64495=>"100011000",
  64496=>"010011001",
  64497=>"001111111",
  64498=>"000110000",
  64499=>"101111001",
  64500=>"101111010",
  64501=>"111000010",
  64502=>"110011011",
  64503=>"111010000",
  64504=>"001100101",
  64505=>"110110111",
  64506=>"110010001",
  64507=>"100110101",
  64508=>"111011000",
  64509=>"101011100",
  64510=>"011000001",
  64511=>"010111010",
  64512=>"000001011",
  64513=>"101011010",
  64514=>"000101010",
  64515=>"100001001",
  64516=>"010111100",
  64517=>"000001101",
  64518=>"001100011",
  64519=>"100011110",
  64520=>"111011101",
  64521=>"000011010",
  64522=>"001000011",
  64523=>"000001101",
  64524=>"010000000",
  64525=>"000010011",
  64526=>"100101011",
  64527=>"001101111",
  64528=>"000010100",
  64529=>"010110000",
  64530=>"001100101",
  64531=>"000001011",
  64532=>"111111110",
  64533=>"100001000",
  64534=>"010111011",
  64535=>"001110110",
  64536=>"011000010",
  64537=>"011011110",
  64538=>"011110011",
  64539=>"101101110",
  64540=>"110011111",
  64541=>"100101101",
  64542=>"110001000",
  64543=>"011010100",
  64544=>"001110000",
  64545=>"000111000",
  64546=>"001001010",
  64547=>"111010011",
  64548=>"010100000",
  64549=>"001000001",
  64550=>"001100100",
  64551=>"101010000",
  64552=>"111010100",
  64553=>"010011111",
  64554=>"110001100",
  64555=>"000111101",
  64556=>"101101001",
  64557=>"101100001",
  64558=>"111001011",
  64559=>"000110000",
  64560=>"001001110",
  64561=>"010101110",
  64562=>"001001101",
  64563=>"111010111",
  64564=>"100111000",
  64565=>"111001110",
  64566=>"101001001",
  64567=>"100011010",
  64568=>"000110100",
  64569=>"010111101",
  64570=>"000011101",
  64571=>"001100100",
  64572=>"101110111",
  64573=>"010110111",
  64574=>"111100000",
  64575=>"110110101",
  64576=>"001010011",
  64577=>"001100000",
  64578=>"010010000",
  64579=>"001001100",
  64580=>"000000011",
  64581=>"100000110",
  64582=>"011000110",
  64583=>"001110000",
  64584=>"010000110",
  64585=>"001101010",
  64586=>"001101011",
  64587=>"100001110",
  64588=>"000001100",
  64589=>"111111011",
  64590=>"001101011",
  64591=>"101000100",
  64592=>"100011101",
  64593=>"111100111",
  64594=>"101111100",
  64595=>"000010010",
  64596=>"111000000",
  64597=>"110001101",
  64598=>"111101001",
  64599=>"111100011",
  64600=>"101011110",
  64601=>"000100011",
  64602=>"011110010",
  64603=>"110110100",
  64604=>"010001110",
  64605=>"010110101",
  64606=>"110110000",
  64607=>"110100100",
  64608=>"111001100",
  64609=>"111011110",
  64610=>"011001111",
  64611=>"111110111",
  64612=>"000010001",
  64613=>"100011110",
  64614=>"101010011",
  64615=>"000011000",
  64616=>"011100011",
  64617=>"000001101",
  64618=>"000011001",
  64619=>"000111010",
  64620=>"111110000",
  64621=>"011100010",
  64622=>"000001010",
  64623=>"101111111",
  64624=>"100100001",
  64625=>"100100101",
  64626=>"111110011",
  64627=>"100011111",
  64628=>"001110011",
  64629=>"100110011",
  64630=>"010010110",
  64631=>"111010010",
  64632=>"111110001",
  64633=>"010100001",
  64634=>"001101110",
  64635=>"001101010",
  64636=>"111011101",
  64637=>"110101000",
  64638=>"101101111",
  64639=>"010000100",
  64640=>"100100000",
  64641=>"111100010",
  64642=>"000111001",
  64643=>"000011000",
  64644=>"010110111",
  64645=>"101000101",
  64646=>"001011001",
  64647=>"111100110",
  64648=>"101001110",
  64649=>"110101000",
  64650=>"100011101",
  64651=>"010011111",
  64652=>"110110000",
  64653=>"111000011",
  64654=>"001101010",
  64655=>"110111000",
  64656=>"011000011",
  64657=>"000001111",
  64658=>"100100111",
  64659=>"110111111",
  64660=>"100100001",
  64661=>"011101001",
  64662=>"000100010",
  64663=>"000110100",
  64664=>"000010111",
  64665=>"111010110",
  64666=>"111101011",
  64667=>"001011101",
  64668=>"000111110",
  64669=>"100110100",
  64670=>"100111000",
  64671=>"101001111",
  64672=>"000100010",
  64673=>"010101001",
  64674=>"001001111",
  64675=>"111010110",
  64676=>"001011110",
  64677=>"111011000",
  64678=>"101100111",
  64679=>"101111110",
  64680=>"001010100",
  64681=>"100011111",
  64682=>"101100011",
  64683=>"000011001",
  64684=>"101111001",
  64685=>"110111110",
  64686=>"111000010",
  64687=>"100111010",
  64688=>"000110011",
  64689=>"111100101",
  64690=>"100100010",
  64691=>"100010010",
  64692=>"001011101",
  64693=>"111000111",
  64694=>"110110110",
  64695=>"001001101",
  64696=>"011010011",
  64697=>"000011110",
  64698=>"011011011",
  64699=>"101101100",
  64700=>"101100111",
  64701=>"000000010",
  64702=>"001111001",
  64703=>"101000110",
  64704=>"101110000",
  64705=>"110011010",
  64706=>"110011010",
  64707=>"010111111",
  64708=>"110001000",
  64709=>"101001001",
  64710=>"001111111",
  64711=>"110011011",
  64712=>"100001001",
  64713=>"011000110",
  64714=>"111001100",
  64715=>"000100110",
  64716=>"000111110",
  64717=>"111100010",
  64718=>"001000001",
  64719=>"101011011",
  64720=>"000011010",
  64721=>"101001100",
  64722=>"100000001",
  64723=>"110011100",
  64724=>"001011001",
  64725=>"010011001",
  64726=>"000100111",
  64727=>"000110000",
  64728=>"000010011",
  64729=>"010101000",
  64730=>"010000010",
  64731=>"111111110",
  64732=>"000000100",
  64733=>"000110101",
  64734=>"001001100",
  64735=>"100101001",
  64736=>"001000100",
  64737=>"011100111",
  64738=>"001100000",
  64739=>"000000011",
  64740=>"101111001",
  64741=>"000001111",
  64742=>"111011011",
  64743=>"011101100",
  64744=>"001011001",
  64745=>"001110011",
  64746=>"010000101",
  64747=>"110000000",
  64748=>"110110010",
  64749=>"001011111",
  64750=>"111101101",
  64751=>"011011010",
  64752=>"000110011",
  64753=>"000101100",
  64754=>"001110110",
  64755=>"110011000",
  64756=>"111010011",
  64757=>"111010110",
  64758=>"110001001",
  64759=>"110101101",
  64760=>"101110111",
  64761=>"111010101",
  64762=>"100010111",
  64763=>"001000111",
  64764=>"111100011",
  64765=>"110101011",
  64766=>"110110111",
  64767=>"001000011",
  64768=>"001001100",
  64769=>"001100000",
  64770=>"110111011",
  64771=>"111100101",
  64772=>"000011001",
  64773=>"101100000",
  64774=>"000001000",
  64775=>"111001110",
  64776=>"111000101",
  64777=>"000011011",
  64778=>"011011001",
  64779=>"100110011",
  64780=>"111111011",
  64781=>"011101011",
  64782=>"110110001",
  64783=>"000111010",
  64784=>"010110100",
  64785=>"011010001",
  64786=>"111010101",
  64787=>"111101110",
  64788=>"100111101",
  64789=>"100101110",
  64790=>"111111111",
  64791=>"100111011",
  64792=>"001100100",
  64793=>"000111011",
  64794=>"000010110",
  64795=>"010110011",
  64796=>"000110110",
  64797=>"000100100",
  64798=>"011001101",
  64799=>"010101111",
  64800=>"110000001",
  64801=>"110100110",
  64802=>"110011001",
  64803=>"011000011",
  64804=>"111001001",
  64805=>"111001010",
  64806=>"000000000",
  64807=>"111111001",
  64808=>"111111100",
  64809=>"000111010",
  64810=>"001010100",
  64811=>"111010011",
  64812=>"010111111",
  64813=>"011011101",
  64814=>"000001111",
  64815=>"000101111",
  64816=>"110111111",
  64817=>"011010001",
  64818=>"010001010",
  64819=>"001000000",
  64820=>"011101101",
  64821=>"111001001",
  64822=>"101111100",
  64823=>"101100110",
  64824=>"111010101",
  64825=>"001010111",
  64826=>"101001001",
  64827=>"001111100",
  64828=>"110001010",
  64829=>"000100101",
  64830=>"011000011",
  64831=>"001011100",
  64832=>"000100101",
  64833=>"011010000",
  64834=>"010110101",
  64835=>"011101100",
  64836=>"000111111",
  64837=>"100001011",
  64838=>"001001011",
  64839=>"011001100",
  64840=>"110010111",
  64841=>"101011111",
  64842=>"101000010",
  64843=>"101001110",
  64844=>"111000111",
  64845=>"000001110",
  64846=>"101000010",
  64847=>"100010000",
  64848=>"000111010",
  64849=>"011011000",
  64850=>"000000010",
  64851=>"010111011",
  64852=>"000010011",
  64853=>"111100101",
  64854=>"011000100",
  64855=>"001100101",
  64856=>"110100001",
  64857=>"101001011",
  64858=>"100000001",
  64859=>"011111000",
  64860=>"111001010",
  64861=>"010111110",
  64862=>"010100100",
  64863=>"000100111",
  64864=>"000000000",
  64865=>"101011101",
  64866=>"111100001",
  64867=>"010001011",
  64868=>"001100000",
  64869=>"011101100",
  64870=>"111100000",
  64871=>"010010000",
  64872=>"100011100",
  64873=>"111011001",
  64874=>"110100110",
  64875=>"000010010",
  64876=>"110001101",
  64877=>"110111111",
  64878=>"110010110",
  64879=>"101010110",
  64880=>"110001111",
  64881=>"111010110",
  64882=>"101100101",
  64883=>"011111110",
  64884=>"100101010",
  64885=>"000101000",
  64886=>"110000001",
  64887=>"001010100",
  64888=>"000000011",
  64889=>"111101011",
  64890=>"010100011",
  64891=>"110001000",
  64892=>"111000001",
  64893=>"101111110",
  64894=>"100111000",
  64895=>"001001000",
  64896=>"111011000",
  64897=>"001011011",
  64898=>"011000100",
  64899=>"011100001",
  64900=>"101011111",
  64901=>"101100000",
  64902=>"101000000",
  64903=>"001010111",
  64904=>"111111000",
  64905=>"111011111",
  64906=>"011000000",
  64907=>"101001111",
  64908=>"111000100",
  64909=>"111011000",
  64910=>"111101101",
  64911=>"000100100",
  64912=>"001000010",
  64913=>"011000101",
  64914=>"011110011",
  64915=>"110111100",
  64916=>"001111010",
  64917=>"010010010",
  64918=>"101111110",
  64919=>"101001011",
  64920=>"101010111",
  64921=>"110010011",
  64922=>"111101011",
  64923=>"111101101",
  64924=>"110010010",
  64925=>"010001101",
  64926=>"000011111",
  64927=>"100001001",
  64928=>"101101110",
  64929=>"110111111",
  64930=>"001100100",
  64931=>"100111010",
  64932=>"010001111",
  64933=>"000001100",
  64934=>"110111011",
  64935=>"011111111",
  64936=>"011110101",
  64937=>"111101001",
  64938=>"001001011",
  64939=>"000111001",
  64940=>"100010111",
  64941=>"111000001",
  64942=>"100011000",
  64943=>"010100010",
  64944=>"011101111",
  64945=>"010011100",
  64946=>"001100011",
  64947=>"110101111",
  64948=>"101110001",
  64949=>"111111110",
  64950=>"010110011",
  64951=>"110001000",
  64952=>"110100001",
  64953=>"010010011",
  64954=>"010100010",
  64955=>"101011110",
  64956=>"010100000",
  64957=>"111101000",
  64958=>"000010111",
  64959=>"100000011",
  64960=>"001011000",
  64961=>"000000010",
  64962=>"110010111",
  64963=>"001110101",
  64964=>"000111010",
  64965=>"100011001",
  64966=>"111101010",
  64967=>"111000101",
  64968=>"001101101",
  64969=>"110001100",
  64970=>"111011000",
  64971=>"110001111",
  64972=>"101111101",
  64973=>"100111101",
  64974=>"111001111",
  64975=>"010100100",
  64976=>"001011010",
  64977=>"011000111",
  64978=>"010110011",
  64979=>"111110010",
  64980=>"101011011",
  64981=>"110011111",
  64982=>"000011011",
  64983=>"011011000",
  64984=>"110011001",
  64985=>"001101000",
  64986=>"001011101",
  64987=>"000111010",
  64988=>"100000100",
  64989=>"111111110",
  64990=>"111011010",
  64991=>"110000111",
  64992=>"011000001",
  64993=>"011110010",
  64994=>"001101110",
  64995=>"010101000",
  64996=>"100100111",
  64997=>"101111111",
  64998=>"010111110",
  64999=>"001110011",
  65000=>"000010010",
  65001=>"000010000",
  65002=>"101111111",
  65003=>"000101011",
  65004=>"000001001",
  65005=>"000000010",
  65006=>"111000101",
  65007=>"000111000",
  65008=>"011101010",
  65009=>"110111000",
  65010=>"010101001",
  65011=>"000110110",
  65012=>"110000001",
  65013=>"011011111",
  65014=>"111111111",
  65015=>"111110110",
  65016=>"111000010",
  65017=>"001110110",
  65018=>"001010000",
  65019=>"000100010",
  65020=>"101000000",
  65021=>"010010011",
  65022=>"010001111",
  65023=>"100000001",
  65024=>"000110100",
  65025=>"000111011",
  65026=>"101000000",
  65027=>"111000011",
  65028=>"110110011",
  65029=>"101111101",
  65030=>"011110101",
  65031=>"100110110",
  65032=>"111000001",
  65033=>"011001100",
  65034=>"000100011",
  65035=>"000011000",
  65036=>"011111101",
  65037=>"001011111",
  65038=>"110110100",
  65039=>"101000000",
  65040=>"100111100",
  65041=>"011110100",
  65042=>"000000011",
  65043=>"111100001",
  65044=>"010001010",
  65045=>"110111111",
  65046=>"011101100",
  65047=>"010110100",
  65048=>"100010000",
  65049=>"000010111",
  65050=>"000001100",
  65051=>"001000011",
  65052=>"001010010",
  65053=>"111100111",
  65054=>"001000110",
  65055=>"101100111",
  65056=>"011110101",
  65057=>"110000001",
  65058=>"101110101",
  65059=>"011101000",
  65060=>"111001110",
  65061=>"011001111",
  65062=>"110011000",
  65063=>"110010100",
  65064=>"101100000",
  65065=>"000101111",
  65066=>"111111000",
  65067=>"000011011",
  65068=>"110001111",
  65069=>"111001000",
  65070=>"101101111",
  65071=>"110010111",
  65072=>"000000100",
  65073=>"001101000",
  65074=>"000000001",
  65075=>"110000100",
  65076=>"110000001",
  65077=>"110011011",
  65078=>"011001101",
  65079=>"100111100",
  65080=>"010111110",
  65081=>"010101101",
  65082=>"110110100",
  65083=>"010100111",
  65084=>"010000101",
  65085=>"011010101",
  65086=>"010101000",
  65087=>"101011010",
  65088=>"100100111",
  65089=>"010000000",
  65090=>"011000001",
  65091=>"010001000",
  65092=>"101111110",
  65093=>"111101011",
  65094=>"111010100",
  65095=>"011001010",
  65096=>"011111011",
  65097=>"100110110",
  65098=>"100011000",
  65099=>"111011110",
  65100=>"011010100",
  65101=>"101110001",
  65102=>"100001001",
  65103=>"100110101",
  65104=>"110000110",
  65105=>"010011010",
  65106=>"111011100",
  65107=>"010111011",
  65108=>"010011110",
  65109=>"100101110",
  65110=>"110110111",
  65111=>"011010001",
  65112=>"111001011",
  65113=>"010001111",
  65114=>"101101000",
  65115=>"000000100",
  65116=>"110110000",
  65117=>"100001011",
  65118=>"110100001",
  65119=>"011100110",
  65120=>"111010100",
  65121=>"000000000",
  65122=>"101000101",
  65123=>"011010100",
  65124=>"011101100",
  65125=>"000001100",
  65126=>"010100000",
  65127=>"100011101",
  65128=>"100101011",
  65129=>"010011110",
  65130=>"001001000",
  65131=>"001011011",
  65132=>"000101111",
  65133=>"100001101",
  65134=>"110010010",
  65135=>"001101000",
  65136=>"001100000",
  65137=>"000010110",
  65138=>"100110111",
  65139=>"000100001",
  65140=>"010100000",
  65141=>"110001011",
  65142=>"100000111",
  65143=>"101110110",
  65144=>"001000100",
  65145=>"000001111",
  65146=>"111010001",
  65147=>"100100010",
  65148=>"111111001",
  65149=>"000000010",
  65150=>"011101001",
  65151=>"011100001",
  65152=>"010011101",
  65153=>"001001101",
  65154=>"001011111",
  65155=>"010001001",
  65156=>"101000000",
  65157=>"101111010",
  65158=>"111111111",
  65159=>"010011000",
  65160=>"100011111",
  65161=>"011111100",
  65162=>"000001100",
  65163=>"111101000",
  65164=>"001111000",
  65165=>"111100110",
  65166=>"111001100",
  65167=>"000110111",
  65168=>"010010010",
  65169=>"010111010",
  65170=>"010001100",
  65171=>"010001011",
  65172=>"010111100",
  65173=>"110100000",
  65174=>"110010011",
  65175=>"000101001",
  65176=>"111011001",
  65177=>"111100000",
  65178=>"100010111",
  65179=>"101101000",
  65180=>"101011000",
  65181=>"111100011",
  65182=>"110001001",
  65183=>"000100010",
  65184=>"011000101",
  65185=>"111100101",
  65186=>"110001110",
  65187=>"001001110",
  65188=>"011101010",
  65189=>"110011101",
  65190=>"010001111",
  65191=>"111001100",
  65192=>"111111000",
  65193=>"110110001",
  65194=>"110001001",
  65195=>"101010010",
  65196=>"100100010",
  65197=>"110110011",
  65198=>"011111001",
  65199=>"101111001",
  65200=>"011000001",
  65201=>"110010001",
  65202=>"111100011",
  65203=>"001001111",
  65204=>"100101110",
  65205=>"100101110",
  65206=>"000010111",
  65207=>"001000010",
  65208=>"011011101",
  65209=>"001000000",
  65210=>"100000010",
  65211=>"010111000",
  65212=>"111001110",
  65213=>"100000011",
  65214=>"010100010",
  65215=>"100111011",
  65216=>"101011111",
  65217=>"111001100",
  65218=>"101111011",
  65219=>"000011110",
  65220=>"101101111",
  65221=>"000100010",
  65222=>"101000101",
  65223=>"010101101",
  65224=>"000000000",
  65225=>"111101011",
  65226=>"111001110",
  65227=>"110110101",
  65228=>"011011100",
  65229=>"010111100",
  65230=>"100111101",
  65231=>"101000000",
  65232=>"001001111",
  65233=>"101111101",
  65234=>"111111100",
  65235=>"111111000",
  65236=>"110010100",
  65237=>"000111010",
  65238=>"000001111",
  65239=>"100100111",
  65240=>"111110111",
  65241=>"100000101",
  65242=>"000001001",
  65243=>"010100101",
  65244=>"110011111",
  65245=>"111111011",
  65246=>"110010111",
  65247=>"101011000",
  65248=>"110111111",
  65249=>"100101111",
  65250=>"000101011",
  65251=>"101100011",
  65252=>"110111101",
  65253=>"100101011",
  65254=>"000011010",
  65255=>"010010111",
  65256=>"110111101",
  65257=>"011011011",
  65258=>"000010100",
  65259=>"101110111",
  65260=>"000011111",
  65261=>"100011000",
  65262=>"101111011",
  65263=>"110000100",
  65264=>"000000110",
  65265=>"111101101",
  65266=>"110101111",
  65267=>"010000110",
  65268=>"010101000",
  65269=>"111010000",
  65270=>"010010000",
  65271=>"010101110",
  65272=>"100100011",
  65273=>"001101000",
  65274=>"111111111",
  65275=>"111100000",
  65276=>"101111010",
  65277=>"111001111",
  65278=>"010111011",
  65279=>"011100111",
  65280=>"100101111",
  65281=>"001010100",
  65282=>"011101100",
  65283=>"010100001",
  65284=>"010101111",
  65285=>"000111000",
  65286=>"000100100",
  65287=>"001000001",
  65288=>"100111100",
  65289=>"011100001",
  65290=>"011100001",
  65291=>"110010111",
  65292=>"000011010",
  65293=>"110000011",
  65294=>"000111100",
  65295=>"010101110",
  65296=>"101010110",
  65297=>"010100101",
  65298=>"001001000",
  65299=>"000110100",
  65300=>"000000100",
  65301=>"110101100",
  65302=>"010010000",
  65303=>"011011101",
  65304=>"101101111",
  65305=>"010000000",
  65306=>"101100000",
  65307=>"010110100",
  65308=>"101000111",
  65309=>"111111110",
  65310=>"011101011",
  65311=>"011101010",
  65312=>"001001100",
  65313=>"111001101",
  65314=>"001011010",
  65315=>"001010110",
  65316=>"011010010",
  65317=>"101101111",
  65318=>"100101100",
  65319=>"100111100",
  65320=>"110010101",
  65321=>"001001000",
  65322=>"001001000",
  65323=>"001000011",
  65324=>"111000101",
  65325=>"100001111",
  65326=>"111101101",
  65327=>"101011111",
  65328=>"010000010",
  65329=>"000011001",
  65330=>"111000010",
  65331=>"111011010",
  65332=>"000011111",
  65333=>"001001000",
  65334=>"100011100",
  65335=>"110010000",
  65336=>"010110001",
  65337=>"011111111",
  65338=>"010101110",
  65339=>"001000010",
  65340=>"010100110",
  65341=>"110100011",
  65342=>"100010010",
  65343=>"001111111",
  65344=>"001010110",
  65345=>"111000000",
  65346=>"001111100",
  65347=>"001101111",
  65348=>"110001100",
  65349=>"011001000",
  65350=>"111111110",
  65351=>"000010001",
  65352=>"011000111",
  65353=>"111101011",
  65354=>"000111111",
  65355=>"111001001",
  65356=>"001000001",
  65357=>"111011101",
  65358=>"010100111",
  65359=>"111111010",
  65360=>"110000010",
  65361=>"110011001",
  65362=>"111111000",
  65363=>"111001111",
  65364=>"011010111",
  65365=>"000001110",
  65366=>"111100111",
  65367=>"000100010",
  65368=>"101010110",
  65369=>"010101011",
  65370=>"000111010",
  65371=>"101100110",
  65372=>"000101110",
  65373=>"001001100",
  65374=>"010100101",
  65375=>"001100111",
  65376=>"000010001",
  65377=>"010101101",
  65378=>"101001100",
  65379=>"111100110",
  65380=>"000111100",
  65381=>"100000110",
  65382=>"101100011",
  65383=>"111111010",
  65384=>"111000110",
  65385=>"110010011",
  65386=>"100111001",
  65387=>"010101010",
  65388=>"100001110",
  65389=>"100000111",
  65390=>"101000110",
  65391=>"000110101",
  65392=>"111111101",
  65393=>"110000010",
  65394=>"100010010",
  65395=>"101010101",
  65396=>"010111011",
  65397=>"010010000",
  65398=>"001001110",
  65399=>"001010010",
  65400=>"111001000",
  65401=>"000011101",
  65402=>"100001101",
  65403=>"000101010",
  65404=>"011110001",
  65405=>"110110011",
  65406=>"010111000",
  65407=>"010011110",
  65408=>"011000000",
  65409=>"111111110",
  65410=>"010111101",
  65411=>"000101100",
  65412=>"000000011",
  65413=>"111111100",
  65414=>"110111001",
  65415=>"100001110",
  65416=>"101110001",
  65417=>"111001010",
  65418=>"101010101",
  65419=>"000011011",
  65420=>"000000010",
  65421=>"000010100",
  65422=>"101101101",
  65423=>"100011000",
  65424=>"111010110",
  65425=>"110010101",
  65426=>"101010101",
  65427=>"100100000",
  65428=>"100111011",
  65429=>"111101010",
  65430=>"001100001",
  65431=>"001100110",
  65432=>"110101110",
  65433=>"000001001",
  65434=>"100111100",
  65435=>"101001000",
  65436=>"010111101",
  65437=>"101111011",
  65438=>"001000101",
  65439=>"111110000",
  65440=>"101011010",
  65441=>"101001001",
  65442=>"001010111",
  65443=>"010011011",
  65444=>"010010001",
  65445=>"100110110",
  65446=>"111111010",
  65447=>"100010110",
  65448=>"000011011",
  65449=>"010111111",
  65450=>"010101111",
  65451=>"001010110",
  65452=>"111001011",
  65453=>"000011100",
  65454=>"001010111",
  65455=>"101011101",
  65456=>"111000000",
  65457=>"111001001",
  65458=>"000000110",
  65459=>"010010010",
  65460=>"010010010",
  65461=>"111000000",
  65462=>"101111000",
  65463=>"000010101",
  65464=>"101001011",
  65465=>"000011011",
  65466=>"001100110",
  65467=>"110111010",
  65468=>"011000110",
  65469=>"000100101",
  65470=>"100001110",
  65471=>"110101110",
  65472=>"110000010",
  65473=>"010111111",
  65474=>"100110100",
  65475=>"111001011",
  65476=>"111111000",
  65477=>"000110100",
  65478=>"100000001",
  65479=>"100101111",
  65480=>"001101101",
  65481=>"110010011",
  65482=>"010010111",
  65483=>"111001000",
  65484=>"110110000",
  65485=>"110100111",
  65486=>"000100110",
  65487=>"011111001",
  65488=>"111000001",
  65489=>"011011111",
  65490=>"101010010",
  65491=>"101000101",
  65492=>"111111111",
  65493=>"010011001",
  65494=>"001011101",
  65495=>"010111111",
  65496=>"010111110",
  65497=>"111111011",
  65498=>"111110111",
  65499=>"000001000",
  65500=>"100010001",
  65501=>"101000101",
  65502=>"100001100",
  65503=>"000100010",
  65504=>"101100001",
  65505=>"110010001",
  65506=>"000011000",
  65507=>"111010101",
  65508=>"010101011",
  65509=>"000000011",
  65510=>"100110111",
  65511=>"110111111",
  65512=>"111101000",
  65513=>"011011101",
  65514=>"100100110",
  65515=>"111011001",
  65516=>"110000101",
  65517=>"000000110",
  65518=>"110100000",
  65519=>"001001001",
  65520=>"100000111",
  65521=>"001111110",
  65522=>"000000001",
  65523=>"110000111",
  65524=>"000001110",
  65525=>"010010000",
  65526=>"101110100",
  65527=>"001001100",
  65528=>"011100100",
  65529=>"010000110",
  65530=>"000011000",
  65531=>"100110000",
  65532=>"001000111",
  65533=>"111110101",
  65534=>"100110111",
  65535=>"001100011");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;