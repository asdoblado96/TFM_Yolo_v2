LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L2_1_BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(3 DOWNTO 0));
END L2_1_BNROM;

ARCHITECTURE RTL OF L2_1_BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"1110110001011111"&"0001011110011100",
    1=>"0010011001101010"&"0000110100010011",
    2=>"0000100100001100"&"0010001111001000",
    3=>"0000011101010100"&"0001110101010100",
    4=>"0000100010010100"&"0010001011101001",
    5=>"0000001110010111"&"0000111100000101",
    6=>"0011111111101001"&"0001001010011001",
    7=>"0010010111001110"&"0000111011011001",
    8=>"1111111010001110"&"0001101001100010",
    9=>"0001100101111010"&"0001000101100101",
    10=>"0000110111010110"&"0001110010100111",
    11=>"1111111100001001"&"0000110001010000",
    12=>"1110000100100000"&"0000011111101101",
    13=>"0000111001100101"&"0010000000001110",
    14=>"0010000101110101"&"0001100100011110",
    15=>"0001110011011000"&"0001110101101011");
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;