LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_9_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_9_BNROM;

ARCHITECTURE RTL OF L8_9_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0001011010001000"&"0001111101101101",
  1=>"0001111101000101"&"0010000110011000",
  2=>"0010110011111100"&"0010010010011000",
  3=>"0010101100111001"&"0010001010100100",
  4=>"0001000000001110"&"0010011111000011",
  5=>"1100110110001101"&"0001010011000100",
  6=>"0000111011110110"&"0010011100110011",
  7=>"0001000000110011"&"0001111111110000",
  8=>"0000111000001110"&"0001111010111000",
  9=>"0001101111001011"&"0010011001010101",
  10=>"0000100001100111"&"0001111100100101",
  11=>"0010101110111011"&"0001111110101100",
  12=>"0010000001001000"&"0010011010100010",
  13=>"0001110100111010"&"0010000011001010",
  14=>"0000110010111010"&"0010100000001100",
  15=>"0000101111000000"&"0010011111110011",
  16=>"0000101111111001"&"0010011000100001",
  17=>"0001100110100100"&"0010011110111001",
  18=>"0000111100101101"&"0010010010011110",
  19=>"0001100100000011"&"0010000100110100",
  20=>"0001001010100011"&"0010010100011000",
  21=>"0000101100001100"&"0001101010011011",
  22=>"0001011001000110"&"0010001010101011",
  23=>"0000101011000101"&"0010001010001010",
  24=>"1111011011101000"&"0010001101100101",
  25=>"0001000000001001"&"0010101000101011",
  26=>"1111010010111011"&"0001110110101000",
  27=>"0000101011011110"&"0001100010100011",
  28=>"0001010011000001"&"0001110101000000",
  29=>"0001011101110101"&"0010010111101001",
  30=>"0001001100010010"&"0010001000110011",
  31=>"1111111110110000"&"0010011000101111",
  32=>"0001000010001011"&"0010010000111000",
  33=>"1111111000110011"&"0001111010000001",
  34=>"0010100111010101"&"0010010001111011",
  35=>"0001111001001001"&"0010011011000010",
  36=>"0000101101010101"&"0010000100000110",
  37=>"0001010111111100"&"0010011101000100",
  38=>"0000101111101001"&"0001101010110111",
  39=>"0001101100110111"&"0010011010011011",
  40=>"0000010011110011"&"0010011001111110",
  41=>"0010111101000011"&"0010000100000001",
  42=>"0000001001110010"&"0010010110010000",
  43=>"0000010110100101"&"0010010000100101",
  44=>"0001010000111011"&"0010010111100001",
  45=>"0001101011010110"&"0010100000000110",
  46=>"0000101100100101"&"0010001101110011",
  47=>"0010100000010100"&"0010000110111110",
  48=>"0001000110110000"&"0010010111101110",
  49=>"0000101110000100"&"0010001010110011",
  50=>"0001110111010011"&"0001101101100101",
  51=>"0010111111011101"&"0001111010101100",
  52=>"0000111100101010"&"0010101001101011",
  53=>"0000100101010100"&"0010011010101110",
  54=>"0010000101010010"&"0010000100101101",
  55=>"0001110101101010"&"0010001100011110",
  56=>"0001011001011010"&"0010010001111010",
  57=>"0000100100100001"&"0001110100001101",
  58=>"0001110110100110"&"0001111101000101",
  59=>"0010000011011111"&"0010010001001010",
  60=>"0000011110110111"&"0001110001110010",
  61=>"0000111110011111"&"0010001101110001",
  62=>"0000001101100010"&"0001111110010101",
  63=>"1111001101110110"&"0001101001011001");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;