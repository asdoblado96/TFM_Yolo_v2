LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_3_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(6 DOWNTO 0));
END L7_3_BNROM;

ARCHITECTURE RTL OF L7_3_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"1111000110110111"&"0010110000111000",
  1=>"1111010010111010"&"0010010111100011",
  2=>"1111001111100011"&"0010011000000011",
  3=>"1111001101000100"&"0010110000001000",
  4=>"1111110010100111"&"0010001100100110",
  5=>"1111000101011101"&"0010011110110010",
  6=>"1111011100001011"&"0010011111111011",
  7=>"1111001110100000"&"0010001100011111",
  8=>"1111101000111110"&"0010001110011000",
  9=>"1110110111111100"&"0010011001000100",
  10=>"1110111010110011"&"0010110010111111",
  11=>"1110101000111011"&"0010011000011001",
  12=>"1111001110101110"&"0010001110100100",
  13=>"1110111010110010"&"0010010001110010",
  14=>"1111010001010001"&"0010011010010001",
  15=>"1110010101010111"&"0010010010111000",
  16=>"1111001100011100"&"0010010110110111",
  17=>"1111011110110010"&"0010000111111111",
  18=>"1110011111001110"&"0010100011110000",
  19=>"1110010110100111"&"0010011111011110",
  20=>"1111001001110010"&"0010011001001010",
  21=>"1111000110000100"&"0010001001011110",
  22=>"1111110010111001"&"0010001000011111",
  23=>"1110011000000000"&"0010100100011010",
  24=>"1110001011111110"&"0010011011100110",
  25=>"1110001111110111"&"0010101100101010",
  26=>"1110111010110000"&"0010001011100111",
  27=>"1110101011001111"&"0010011000001111",
  28=>"1111011111111101"&"0010001100010001",
  29=>"1110100011001111"&"0010100101010000",
  30=>"1111100110010001"&"0010010010011101",
  31=>"1111010001111111"&"0010010100110001",
  32=>"1110000001001111"&"0010101110000110",
  33=>"1110111001110000"&"0010001100100111",
  34=>"1110110000100100"&"0010011111100101",
  35=>"1111101101110010"&"0010010011100011",
  36=>"1111000010101011"&"0010001111001010",
  37=>"1111110100110011"&"0010001111110110",
  38=>"0000100001100111"&"0010000111011011",
  39=>"1111001110001110"&"0010010101101111",
  40=>"1110101011110111"&"0010101001110101",
  41=>"1110110001000111"&"0010011010011000",
  42=>"1111011010111000"&"0010001101111111",
  43=>"1111000101000100"&"0010000001110100",
  44=>"1111010111100111"&"0010011000101001",
  45=>"1111001100101010"&"0010011001111110",
  46=>"1110011001000001"&"0010010111011100",
  47=>"0000000011000111"&"0010010111011011",
  48=>"1111111010001101"&"0010010100101110",
  49=>"1110011011000110"&"0010011000011010",
  50=>"1110110100000111"&"0010001010111000",
  51=>"1110110100101010"&"0010011101010110",
  52=>"1111001010010110"&"0010001011100101",
  53=>"1110110100100011"&"0010100011110010",
  54=>"1111011000001001"&"0010100010100001",
  55=>"1110100011101111"&"0010001111011001",
  56=>"1110100010010101"&"0010000101000100",
  57=>"1111010011001000"&"0010011011000100",
  58=>"1111011101100111"&"0010001001110110",
  59=>"1111111011111010"&"0010100101001100",
  60=>"1111010111110110"&"0010010001110001",
  61=>"1111010111000101"&"0010100101010111",
  62=>"1111010010011010"&"0010010100000000",
  63=>"1111011111111001"&"0010001101101000",
  64=>"1111101011011011"&"0010000111100011",
  65=>"1110011111000100"&"0010011110100100",
  66=>"1111110001111000"&"0010010111100110",
  67=>"1110010100111110"&"0010000101101101",
  68=>"1111101001101111"&"0010000100011010",
  69=>"1110110110011101"&"0010101100010100",
  70=>"1110100100000101"&"0010011100111111",
  71=>"1111010110000001"&"0010011001100110",
  72=>"1110111110000111"&"0010100001110110",
  73=>"1110001111101110"&"0001111110001110",
  74=>"1111010011010101"&"0010001110001011",
  75=>"1110011011010001"&"0010001011000111",
  76=>"1110110011100110"&"0010100100000111",
  77=>"1110010000001011"&"0010111101101000",
  78=>"1111000101001110"&"0001111111111011",
  79=>"1110011010000101"&"0001111110100110",
  80=>"1110100011101010"&"0010010000100001",
  81=>"1110001111110001"&"0010111010100001",
  82=>"1111010101110010"&"0010010101010101",
  83=>"1111111111001110"&"0010010110010011",
  84=>"1111000111100011"&"0010110010101110",
  85=>"1110110111100000"&"0010000000111111",
  86=>"1110011110100100"&"0010011001010111",
  87=>"1111001001101110"&"0010011010010111",
  88=>"1111101010101001"&"0010010011100100",
  89=>"1110100011111000"&"0010000001001001",
  90=>"1110100010000101"&"0010001010010111",
  91=>"1111000001110000"&"0010010011100110",
  92=>"1110100000001111"&"0010001010000010",
  93=>"1111001000001001"&"0010101010001011",
  94=>"1110110110011001"&"0010011100000011",
  95=>"1111001011101100"&"0010100011100001",
  96=>"1111000110110000"&"0010000101101100",
  97=>"0000000100001001"&"0010011000001001",
  98=>"1110111010001011"&"0010101100100111",
  99=>"1110100111111010"&"0010011001111000",
  100=>"1111011100100100"&"0010100110100010",
  101=>"1111001000111110"&"0010011110100011",
  102=>"1110111100010011"&"0010101010110111",
  103=>"1110101101101100"&"0010010011000110",
  104=>"1111101000111010"&"0010001110011000",
  105=>"1110101101011101"&"0010010000001110",
  106=>"1111011100001111"&"0010010100111011",
  107=>"1110110110101001"&"0010101101111011",
  108=>"1110110000110010"&"0010001011001111",
  109=>"1110001000101001"&"0011000010000000",
  110=>"1110001000110111"&"0010100010110100",
  111=>"1111001100111110"&"0010011110011111",
  112=>"1110110100011011"&"0010010101111000",
  113=>"1110001011111011"&"0010101001010000",
  114=>"1111001000110011"&"0010100001010010",
  115=>"0000000010001111"&"0010001110000011",
  116=>"1110101100101001"&"0010111100011000",
  117=>"1110000111011010"&"0010001101110000",
  118=>"1101111111010100"&"0010011101001111",
  119=>"1111001100011010"&"0010010110100111",
  120=>"1111001101001000"&"0010011101100101",
  121=>"1110011011010000"&"0010001010011010",
  122=>"1111010001110010"&"0010101000110001",
  123=>"1110101111100111"&"0010011001111100",
  124=>"1110011111001110"&"0010001001100000",
  125=>"1111100001010100"&"0010011101001100",
  126=>"1111100000100010"&"0010110101011000",
  127=>"1110010010101101"&"0010001011000011");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;