LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_3_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8) - 1 DOWNTO 0));
END L8_3_WROM;

ARCHITECTURE RTL OF L8_3_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"100001000",
  1=>"001001100",
  2=>"000010111",
  3=>"001111010",
  4=>"110001101",
  5=>"111100001",
  6=>"011011001",
  7=>"110101010",
  8=>"011101101",
  9=>"100100000",
  10=>"001110110",
  11=>"101000101",
  12=>"111000101",
  13=>"011010110",
  14=>"011110011",
  15=>"111001110",
  16=>"000000111",
  17=>"011010001",
  18=>"010101101",
  19=>"000110111",
  20=>"000011101",
  21=>"100011101",
  22=>"100111110",
  23=>"011111011",
  24=>"101001010",
  25=>"011011000",
  26=>"111000010",
  27=>"111010101",
  28=>"111000001",
  29=>"101001101",
  30=>"111101101",
  31=>"000001101",
  32=>"000000011",
  33=>"100101101",
  34=>"100001111",
  35=>"011000001",
  36=>"100101100",
  37=>"111011011",
  38=>"100101111",
  39=>"110110101",
  40=>"111101111",
  41=>"010010100",
  42=>"101011000",
  43=>"101111011",
  44=>"000100111",
  45=>"010000110",
  46=>"101001111",
  47=>"000010001",
  48=>"011000101",
  49=>"100011000",
  50=>"000100001",
  51=>"110011101",
  52=>"000000110",
  53=>"011100011",
  54=>"100011011",
  55=>"011000001",
  56=>"111001101",
  57=>"011011100",
  58=>"100010111",
  59=>"001011000",
  60=>"000111101",
  61=>"101010010",
  62=>"110000000",
  63=>"000011111",
  64=>"001011001",
  65=>"110110100",
  66=>"111010101",
  67=>"100111111",
  68=>"011101010",
  69=>"010011011",
  70=>"000110001",
  71=>"111000001",
  72=>"101100111",
  73=>"110101010",
  74=>"101101110",
  75=>"010101010",
  76=>"111011101",
  77=>"111011001",
  78=>"000100111",
  79=>"101110111",
  80=>"001101110",
  81=>"111101111",
  82=>"011101111",
  83=>"000101101",
  84=>"000010001",
  85=>"111100011",
  86=>"000000001",
  87=>"101101011",
  88=>"011011101",
  89=>"100001100",
  90=>"011011110",
  91=>"101000000",
  92=>"100101010",
  93=>"000110001",
  94=>"010011010",
  95=>"100011111",
  96=>"010011101",
  97=>"011011010",
  98=>"000000000",
  99=>"101100110",
  100=>"110000001",
  101=>"001011001",
  102=>"010100001",
  103=>"101111001",
  104=>"011010110",
  105=>"101101111",
  106=>"000010111",
  107=>"100000111",
  108=>"000111000",
  109=>"100110110",
  110=>"110110001",
  111=>"000000101",
  112=>"000000100",
  113=>"101011010",
  114=>"110001100",
  115=>"010111101",
  116=>"010010010",
  117=>"101001011",
  118=>"100011001",
  119=>"100111101",
  120=>"000000100",
  121=>"101100101",
  122=>"000000001",
  123=>"011100100",
  124=>"100011101",
  125=>"001110110",
  126=>"010010010",
  127=>"000100100",
  128=>"011001010",
  129=>"001100000",
  130=>"100010100",
  131=>"000110000",
  132=>"001010111",
  133=>"110111111",
  134=>"111010001",
  135=>"010110000",
  136=>"111101101",
  137=>"110011010",
  138=>"001011000",
  139=>"000010011",
  140=>"011101111",
  141=>"110001100",
  142=>"110111000",
  143=>"010011111",
  144=>"010000000",
  145=>"101111100",
  146=>"101010010",
  147=>"001110111",
  148=>"101100001",
  149=>"101000111",
  150=>"000001001",
  151=>"111001000",
  152=>"001100111",
  153=>"111011100",
  154=>"000011100",
  155=>"110111110",
  156=>"001000100",
  157=>"000111110",
  158=>"001110111",
  159=>"001111000",
  160=>"100100001",
  161=>"110001110",
  162=>"111101011",
  163=>"000101100",
  164=>"000000101",
  165=>"011010101",
  166=>"101110100",
  167=>"001100010",
  168=>"010001000",
  169=>"011111011",
  170=>"101101100",
  171=>"100110010",
  172=>"001001000",
  173=>"111010111",
  174=>"001101001",
  175=>"010111010",
  176=>"100010010",
  177=>"011100011",
  178=>"011010000",
  179=>"010011011",
  180=>"010100100",
  181=>"010000000",
  182=>"010100001",
  183=>"100000110",
  184=>"011110110",
  185=>"110100000",
  186=>"001100010",
  187=>"110111101",
  188=>"110110001",
  189=>"100111001",
  190=>"010000101",
  191=>"010000100",
  192=>"001110111",
  193=>"111000111",
  194=>"101111000",
  195=>"110010010",
  196=>"011000001",
  197=>"111001011",
  198=>"000001001",
  199=>"101100111",
  200=>"111011110",
  201=>"100101101",
  202=>"101100011",
  203=>"100010111",
  204=>"101101111",
  205=>"110001011",
  206=>"010001000",
  207=>"110101001",
  208=>"000010100",
  209=>"001111000",
  210=>"010111001",
  211=>"001010011",
  212=>"101111110",
  213=>"110010011",
  214=>"111111110",
  215=>"100011010",
  216=>"110100010",
  217=>"011001011",
  218=>"101101011",
  219=>"111000001",
  220=>"110101001",
  221=>"111000100",
  222=>"101101101",
  223=>"110101111",
  224=>"000010001",
  225=>"001110010",
  226=>"101110111",
  227=>"101011011",
  228=>"111010001",
  229=>"111101010",
  230=>"110100011",
  231=>"111110100",
  232=>"111100000",
  233=>"010110000",
  234=>"000000111",
  235=>"100001010",
  236=>"100011000",
  237=>"000111111",
  238=>"101100111",
  239=>"101111111",
  240=>"101000101",
  241=>"011000101",
  242=>"010100000",
  243=>"001000000",
  244=>"000010101",
  245=>"001100100",
  246=>"011011001",
  247=>"000100001",
  248=>"100000000",
  249=>"010001100",
  250=>"011111110",
  251=>"000000011",
  252=>"000110110",
  253=>"110100000",
  254=>"001000001",
  255=>"100111111",
  256=>"100101000",
  257=>"000000010",
  258=>"101000110",
  259=>"110000001",
  260=>"011000011",
  261=>"000111001",
  262=>"100000010",
  263=>"101101011",
  264=>"000001101",
  265=>"001001011",
  266=>"000010001",
  267=>"110111000",
  268=>"000111010",
  269=>"100010010",
  270=>"110111000",
  271=>"101110001",
  272=>"101011011",
  273=>"000000110",
  274=>"000000101",
  275=>"000111111",
  276=>"111001101",
  277=>"111100000",
  278=>"101000000",
  279=>"100110010",
  280=>"000100001",
  281=>"011100000",
  282=>"010110000",
  283=>"010111010",
  284=>"000000010",
  285=>"000110011",
  286=>"110100111",
  287=>"000010110",
  288=>"110010101",
  289=>"110100010",
  290=>"000010011",
  291=>"011010011",
  292=>"100000100",
  293=>"101010001",
  294=>"101000111",
  295=>"100111000",
  296=>"000111100",
  297=>"110101110",
  298=>"111110111",
  299=>"010000010",
  300=>"100001111",
  301=>"000100001",
  302=>"110000100",
  303=>"111110000",
  304=>"110111101",
  305=>"110101011",
  306=>"010000001",
  307=>"001101110",
  308=>"011011000",
  309=>"100111101",
  310=>"100010000",
  311=>"100001001",
  312=>"000001111",
  313=>"001001011",
  314=>"011111111",
  315=>"100101011",
  316=>"000010101",
  317=>"101001111",
  318=>"111111101",
  319=>"011100101",
  320=>"011100110",
  321=>"010000101",
  322=>"010001100",
  323=>"100100101",
  324=>"011100011",
  325=>"001001010",
  326=>"000000100",
  327=>"000000101",
  328=>"000100111",
  329=>"010101110",
  330=>"000110111",
  331=>"001101001",
  332=>"000000010",
  333=>"111100011",
  334=>"011011111",
  335=>"110110111",
  336=>"101011011",
  337=>"111000101",
  338=>"100000011",
  339=>"101000100",
  340=>"001000101",
  341=>"100100111",
  342=>"110110110",
  343=>"111110010",
  344=>"101000110",
  345=>"101011100",
  346=>"111001100",
  347=>"100001000",
  348=>"000000000",
  349=>"110010010",
  350=>"111110010",
  351=>"011110100",
  352=>"001101110",
  353=>"100111010",
  354=>"011011010",
  355=>"000110000",
  356=>"111011101",
  357=>"010110000",
  358=>"101010110",
  359=>"110011101",
  360=>"011110001",
  361=>"001100000",
  362=>"101101101",
  363=>"001000000",
  364=>"000011011",
  365=>"010101001",
  366=>"001111101",
  367=>"101010011",
  368=>"001011000",
  369=>"010110100",
  370=>"011011100",
  371=>"110101011",
  372=>"100101010",
  373=>"001111011",
  374=>"100001001",
  375=>"101101110",
  376=>"110000010",
  377=>"010111110",
  378=>"000001011",
  379=>"011110101",
  380=>"011111110",
  381=>"010000001",
  382=>"111011110",
  383=>"011100110",
  384=>"000010001",
  385=>"110111001",
  386=>"111000100",
  387=>"010111000",
  388=>"010111101",
  389=>"110111010",
  390=>"000101101",
  391=>"000100100",
  392=>"101110101",
  393=>"110010011",
  394=>"110100111",
  395=>"111010001",
  396=>"100001001",
  397=>"100111110",
  398=>"101101000",
  399=>"111101111",
  400=>"101010110",
  401=>"001000010",
  402=>"101111100",
  403=>"001010010",
  404=>"000111101",
  405=>"110001101",
  406=>"101101111",
  407=>"000010100",
  408=>"110011110",
  409=>"011001000",
  410=>"100000001",
  411=>"100110001",
  412=>"011001011",
  413=>"010110010",
  414=>"101001111",
  415=>"100000000",
  416=>"101110101",
  417=>"101010100",
  418=>"110000000",
  419=>"101000010",
  420=>"101101110",
  421=>"111100101",
  422=>"111110000",
  423=>"100001100",
  424=>"111100010",
  425=>"100100111",
  426=>"101000000",
  427=>"001010010",
  428=>"000010110",
  429=>"000101100",
  430=>"011100101",
  431=>"000110100",
  432=>"000000100",
  433=>"111101111",
  434=>"111110110",
  435=>"101101110",
  436=>"010010010",
  437=>"100110101",
  438=>"101111010",
  439=>"010000101",
  440=>"010101011",
  441=>"010111011",
  442=>"000000010",
  443=>"011010011",
  444=>"010010001",
  445=>"010010101",
  446=>"101010110",
  447=>"001100010",
  448=>"011111011",
  449=>"111000010",
  450=>"011010010",
  451=>"111101000",
  452=>"100000101",
  453=>"010011001",
  454=>"000100011",
  455=>"011110010",
  456=>"011110001",
  457=>"001110100",
  458=>"001111000",
  459=>"100111111",
  460=>"010110011",
  461=>"100011000",
  462=>"100000001",
  463=>"010000010",
  464=>"000011000",
  465=>"100101000",
  466=>"000010110",
  467=>"100000000",
  468=>"110100011",
  469=>"101010010",
  470=>"101111110",
  471=>"001010110",
  472=>"010110010",
  473=>"101111111",
  474=>"110011110",
  475=>"000101001",
  476=>"101001001",
  477=>"110010111",
  478=>"010100111",
  479=>"111001111",
  480=>"101011100",
  481=>"100011001",
  482=>"111010000",
  483=>"110011010",
  484=>"111101000",
  485=>"111111100",
  486=>"100000100",
  487=>"010101001",
  488=>"000101011",
  489=>"101110110",
  490=>"111000110",
  491=>"101010101",
  492=>"010110111",
  493=>"001110001",
  494=>"100010011",
  495=>"000111111",
  496=>"000010000",
  497=>"111001110",
  498=>"100100011",
  499=>"111011000",
  500=>"101010100",
  501=>"111111111",
  502=>"110100110",
  503=>"000110010",
  504=>"000110101",
  505=>"010111010",
  506=>"001001001",
  507=>"111010010",
  508=>"100010101",
  509=>"110101100",
  510=>"100101001",
  511=>"111101001",
  512=>"000011111",
  513=>"000010100",
  514=>"111000100",
  515=>"111111110",
  516=>"001010101",
  517=>"010000001",
  518=>"001001100",
  519=>"000111100",
  520=>"000110101",
  521=>"001010000",
  522=>"001011101",
  523=>"001110010",
  524=>"101001001",
  525=>"111111101",
  526=>"110000000",
  527=>"111110001",
  528=>"011100001",
  529=>"011011011",
  530=>"101111000",
  531=>"000011101",
  532=>"001011000",
  533=>"110110110",
  534=>"010001100",
  535=>"001000101",
  536=>"110001111",
  537=>"000001111",
  538=>"001101100",
  539=>"100011000",
  540=>"110001100",
  541=>"011101100",
  542=>"111111011",
  543=>"001001111",
  544=>"000100100",
  545=>"100110011",
  546=>"110010100",
  547=>"000011010",
  548=>"001010110",
  549=>"101000000",
  550=>"110000000",
  551=>"100111000",
  552=>"011110010",
  553=>"000100000",
  554=>"110101000",
  555=>"110000111",
  556=>"010001101",
  557=>"000011100",
  558=>"111100000",
  559=>"001101010",
  560=>"110111100",
  561=>"011100101",
  562=>"011011010",
  563=>"100011101",
  564=>"001011110",
  565=>"000111011",
  566=>"001000100",
  567=>"011110101",
  568=>"000000110",
  569=>"001000110",
  570=>"000110111",
  571=>"100000110",
  572=>"000010000",
  573=>"010011000",
  574=>"100110101",
  575=>"110111110",
  576=>"110010100",
  577=>"111001011",
  578=>"101100111",
  579=>"111010100",
  580=>"000110000",
  581=>"010001101",
  582=>"000010100",
  583=>"001111011",
  584=>"001110111",
  585=>"001100001",
  586=>"000001100",
  587=>"101000011",
  588=>"100111010",
  589=>"001101000",
  590=>"100010001",
  591=>"010110001",
  592=>"100100100",
  593=>"011110000",
  594=>"100101101",
  595=>"000101000",
  596=>"001101110",
  597=>"110000001",
  598=>"010000000",
  599=>"100010110",
  600=>"011111011",
  601=>"111101110",
  602=>"010111011",
  603=>"000011010",
  604=>"011001100",
  605=>"111100000",
  606=>"101001110",
  607=>"101101100",
  608=>"110100000",
  609=>"000000011",
  610=>"101111110",
  611=>"111100101",
  612=>"100011110",
  613=>"111000000",
  614=>"000011010",
  615=>"110001000",
  616=>"000000011",
  617=>"101000010",
  618=>"010011011",
  619=>"010010001",
  620=>"011111100",
  621=>"001001010",
  622=>"100100111",
  623=>"000010101",
  624=>"111110101",
  625=>"001100010",
  626=>"010000101",
  627=>"110111100",
  628=>"111101100",
  629=>"110101001",
  630=>"011100010",
  631=>"010000100",
  632=>"111000000",
  633=>"101111011",
  634=>"011010000",
  635=>"101001001",
  636=>"000101010",
  637=>"101100010",
  638=>"101000010",
  639=>"101110110",
  640=>"000001010",
  641=>"001110010",
  642=>"001110001",
  643=>"000100010",
  644=>"110000100",
  645=>"001001011",
  646=>"101111000",
  647=>"000100101",
  648=>"001001001",
  649=>"001111110",
  650=>"110101010",
  651=>"011110101",
  652=>"101000100",
  653=>"011001101",
  654=>"001101001",
  655=>"101110110",
  656=>"111110101",
  657=>"110001000",
  658=>"000101110",
  659=>"100001101",
  660=>"011101000",
  661=>"111111011",
  662=>"101000100",
  663=>"000000111",
  664=>"101010110",
  665=>"111110101",
  666=>"111100001",
  667=>"101111010",
  668=>"011111001",
  669=>"110000000",
  670=>"011111001",
  671=>"100000011",
  672=>"001001011",
  673=>"000111010",
  674=>"000101101",
  675=>"111100000",
  676=>"111100010",
  677=>"011111111",
  678=>"100000010",
  679=>"010110110",
  680=>"110010100",
  681=>"000000011",
  682=>"110100011",
  683=>"001001010",
  684=>"010000100",
  685=>"001101101",
  686=>"111000010",
  687=>"101001111",
  688=>"100001110",
  689=>"110100000",
  690=>"101001101",
  691=>"110011010",
  692=>"010011100",
  693=>"110101111",
  694=>"000000110",
  695=>"100110001",
  696=>"110011000",
  697=>"111011000",
  698=>"101010110",
  699=>"110110111",
  700=>"101101011",
  701=>"111001001",
  702=>"001110110",
  703=>"110001011",
  704=>"101110011",
  705=>"000000110",
  706=>"101000011",
  707=>"010111100",
  708=>"110110111",
  709=>"001000011",
  710=>"100000101",
  711=>"110011000",
  712=>"100101100",
  713=>"011101010",
  714=>"000001111",
  715=>"011110011",
  716=>"001001000",
  717=>"000010000",
  718=>"111001111",
  719=>"110001100",
  720=>"110111101",
  721=>"011001100",
  722=>"000010000",
  723=>"001011011",
  724=>"001111101",
  725=>"010000100",
  726=>"010011000",
  727=>"110010100",
  728=>"010000011",
  729=>"001001111",
  730=>"001100100",
  731=>"101001010",
  732=>"001110110",
  733=>"101111001",
  734=>"100010001",
  735=>"010001001",
  736=>"011010100",
  737=>"100100110",
  738=>"001101110",
  739=>"010110101",
  740=>"011010101",
  741=>"100001110",
  742=>"001100100",
  743=>"101100000",
  744=>"101001001",
  745=>"101110101",
  746=>"000101010",
  747=>"001101110",
  748=>"010011100",
  749=>"111010100",
  750=>"010101011",
  751=>"000011110",
  752=>"010111001",
  753=>"000010100",
  754=>"001010010",
  755=>"010011100",
  756=>"101011101",
  757=>"100111110",
  758=>"010101110",
  759=>"000111011",
  760=>"011000101",
  761=>"100011101",
  762=>"010110101",
  763=>"101010011",
  764=>"111010111",
  765=>"000110001",
  766=>"001010101",
  767=>"101110000",
  768=>"011000110",
  769=>"101111011",
  770=>"111111000",
  771=>"011010110",
  772=>"100000011",
  773=>"100110011",
  774=>"101100100",
  775=>"100011001",
  776=>"000001111",
  777=>"100110100",
  778=>"100000100",
  779=>"011010101",
  780=>"010010000",
  781=>"111110010",
  782=>"111010100",
  783=>"100010111",
  784=>"100001101",
  785=>"000000100",
  786=>"010011110",
  787=>"100101101",
  788=>"111000100",
  789=>"000000111",
  790=>"010011101",
  791=>"000010101",
  792=>"001000101",
  793=>"010110000",
  794=>"010101000",
  795=>"101001011",
  796=>"001001101",
  797=>"110110000",
  798=>"110001011",
  799=>"010100001",
  800=>"010010011",
  801=>"010101110",
  802=>"101001110",
  803=>"011010010",
  804=>"101000010",
  805=>"011001010",
  806=>"101100000",
  807=>"110100001",
  808=>"011111100",
  809=>"001000001",
  810=>"111010011",
  811=>"111010001",
  812=>"101000000",
  813=>"110100111",
  814=>"101011100",
  815=>"101001010",
  816=>"010101101",
  817=>"110001011",
  818=>"100111000",
  819=>"001010001",
  820=>"001000011",
  821=>"010101100",
  822=>"001010010",
  823=>"111010010",
  824=>"100001000",
  825=>"110101100",
  826=>"010001011",
  827=>"100111110",
  828=>"100011110",
  829=>"001100011",
  830=>"101011111",
  831=>"100110100",
  832=>"100010111",
  833=>"101101010",
  834=>"011001101",
  835=>"000000000",
  836=>"111110100",
  837=>"110111100",
  838=>"111101101",
  839=>"111010110",
  840=>"001011110",
  841=>"100000111",
  842=>"011111101",
  843=>"000100011",
  844=>"111001100",
  845=>"011100000",
  846=>"000000010",
  847=>"000001001",
  848=>"001010100",
  849=>"111000111",
  850=>"000110111",
  851=>"000000101",
  852=>"010111110",
  853=>"000111101",
  854=>"010101110",
  855=>"000011000",
  856=>"100111000",
  857=>"001000101",
  858=>"000001100",
  859=>"101101000",
  860=>"110010011",
  861=>"100100011",
  862=>"111100001",
  863=>"000001101",
  864=>"110101100",
  865=>"101000010",
  866=>"111110100",
  867=>"001011100",
  868=>"100101011",
  869=>"101000101",
  870=>"001110000",
  871=>"001010110",
  872=>"000011001",
  873=>"100000010",
  874=>"010100110",
  875=>"001110111",
  876=>"010000010",
  877=>"111111011",
  878=>"000000011",
  879=>"011000011",
  880=>"000100011",
  881=>"010100011",
  882=>"101101011",
  883=>"101111101",
  884=>"101111101",
  885=>"010101110",
  886=>"001011100",
  887=>"010011000",
  888=>"101100001",
  889=>"011000001",
  890=>"110000111",
  891=>"010101111",
  892=>"001101101",
  893=>"110111110",
  894=>"001000111",
  895=>"001100100",
  896=>"001010111",
  897=>"010110011",
  898=>"101101101",
  899=>"100010100",
  900=>"010101010",
  901=>"000000000",
  902=>"010111010",
  903=>"110010010",
  904=>"111001001",
  905=>"111011111",
  906=>"000111011",
  907=>"000101010",
  908=>"011111111",
  909=>"010110100",
  910=>"000010101",
  911=>"110110111",
  912=>"111000110",
  913=>"001110100",
  914=>"011111100",
  915=>"011111101",
  916=>"110111100",
  917=>"111110111",
  918=>"110010101",
  919=>"111011110",
  920=>"101000111",
  921=>"111101100",
  922=>"001011000",
  923=>"001000100",
  924=>"010011000",
  925=>"010001001",
  926=>"100000010",
  927=>"011010010",
  928=>"100110001",
  929=>"010110110",
  930=>"010011000",
  931=>"100000010",
  932=>"101000101",
  933=>"101001011",
  934=>"101010100",
  935=>"110100011",
  936=>"001010010",
  937=>"001000001",
  938=>"110011010",
  939=>"101111001",
  940=>"000111111",
  941=>"100100101",
  942=>"101101111",
  943=>"000010111",
  944=>"001000000",
  945=>"010001101",
  946=>"010001011",
  947=>"100011010",
  948=>"001010111",
  949=>"101110011",
  950=>"001011101",
  951=>"101101010",
  952=>"011111110",
  953=>"110100000",
  954=>"001110011",
  955=>"010000111",
  956=>"001001011",
  957=>"000100000",
  958=>"001001001",
  959=>"011000000",
  960=>"000000101",
  961=>"111000100",
  962=>"011011111",
  963=>"010101111",
  964=>"001111111",
  965=>"110001010",
  966=>"100110110",
  967=>"010010010",
  968=>"100111100",
  969=>"001110011",
  970=>"101010010",
  971=>"000110100",
  972=>"101011111",
  973=>"000101110",
  974=>"000010000",
  975=>"101010111",
  976=>"011111100",
  977=>"000000011",
  978=>"011111011",
  979=>"000100001",
  980=>"010110010",
  981=>"001101100",
  982=>"110010111",
  983=>"111001111",
  984=>"110000000",
  985=>"110001111",
  986=>"100110101",
  987=>"010010000",
  988=>"100000001",
  989=>"010110100",
  990=>"010010010",
  991=>"101101111",
  992=>"111011111",
  993=>"101011100",
  994=>"011101001",
  995=>"100000001",
  996=>"111001001",
  997=>"111000100",
  998=>"101100111",
  999=>"111110000",
  1000=>"101101011",
  1001=>"111100010",
  1002=>"111100001",
  1003=>"100010101",
  1004=>"110100111",
  1005=>"110000001",
  1006=>"000001101",
  1007=>"110111100",
  1008=>"000001100",
  1009=>"101010011",
  1010=>"110010101",
  1011=>"100100011",
  1012=>"101000010",
  1013=>"011100100",
  1014=>"010111011",
  1015=>"100000010",
  1016=>"101001101",
  1017=>"000001110",
  1018=>"100101010",
  1019=>"010010010",
  1020=>"111111111",
  1021=>"111001010",
  1022=>"111001010",
  1023=>"010110110",
  1024=>"110011111",
  1025=>"100100100",
  1026=>"001100110",
  1027=>"010001010",
  1028=>"000100110",
  1029=>"000010011",
  1030=>"110010011",
  1031=>"111010000",
  1032=>"000000101",
  1033=>"001100101",
  1034=>"001010011",
  1035=>"110101110",
  1036=>"000001000",
  1037=>"001000011",
  1038=>"011000001",
  1039=>"010111100",
  1040=>"000110000",
  1041=>"101011000",
  1042=>"100000010",
  1043=>"000010000",
  1044=>"000110110",
  1045=>"110001110",
  1046=>"100001111",
  1047=>"011001001",
  1048=>"100000111",
  1049=>"101111000",
  1050=>"011111110",
  1051=>"101000110",
  1052=>"101111011",
  1053=>"001001110",
  1054=>"001110110",
  1055=>"101000011",
  1056=>"001001001",
  1057=>"101110101",
  1058=>"110011110",
  1059=>"100100100",
  1060=>"000111010",
  1061=>"000100000",
  1062=>"101100111",
  1063=>"111010100",
  1064=>"011010000",
  1065=>"111101101",
  1066=>"011110110",
  1067=>"001100101",
  1068=>"110010111",
  1069=>"111011100",
  1070=>"000010111",
  1071=>"100100010",
  1072=>"101000001",
  1073=>"110000000",
  1074=>"100000100",
  1075=>"001011100",
  1076=>"000000000",
  1077=>"110010010",
  1078=>"010101010",
  1079=>"011110011",
  1080=>"101000011",
  1081=>"011000100",
  1082=>"111010110",
  1083=>"010010011",
  1084=>"000010011",
  1085=>"111100101",
  1086=>"001000001",
  1087=>"111000110",
  1088=>"000111111",
  1089=>"110000100",
  1090=>"011111001",
  1091=>"101001000",
  1092=>"001101111",
  1093=>"000010101",
  1094=>"001011110",
  1095=>"101000100",
  1096=>"001000001",
  1097=>"110010010",
  1098=>"010000001",
  1099=>"011011010",
  1100=>"101100101",
  1101=>"011001110",
  1102=>"111010101",
  1103=>"111100010",
  1104=>"011101111",
  1105=>"111100010",
  1106=>"011000110",
  1107=>"110010110",
  1108=>"000011000",
  1109=>"010111001",
  1110=>"010101110",
  1111=>"000011100",
  1112=>"100010010",
  1113=>"010101011",
  1114=>"010101111",
  1115=>"011000101",
  1116=>"011011001",
  1117=>"011100001",
  1118=>"000101110",
  1119=>"010110011",
  1120=>"100111010",
  1121=>"110011110",
  1122=>"101100100",
  1123=>"011011000",
  1124=>"101111101",
  1125=>"000011110",
  1126=>"000010010",
  1127=>"000000010",
  1128=>"111011111",
  1129=>"110100111",
  1130=>"000111100",
  1131=>"100100010",
  1132=>"001110100",
  1133=>"001001100",
  1134=>"010111001",
  1135=>"111101111",
  1136=>"001101110",
  1137=>"010000011",
  1138=>"000101101",
  1139=>"011000111",
  1140=>"111111101",
  1141=>"011110110",
  1142=>"101111011",
  1143=>"110000000",
  1144=>"100101001",
  1145=>"000111010",
  1146=>"100010000",
  1147=>"100111001",
  1148=>"010100010",
  1149=>"110110011",
  1150=>"010111111",
  1151=>"111110110",
  1152=>"010000101",
  1153=>"111110101",
  1154=>"111011101",
  1155=>"011010001",
  1156=>"111100111",
  1157=>"001001010",
  1158=>"000101011",
  1159=>"101111101",
  1160=>"101000101",
  1161=>"110111111",
  1162=>"100011010",
  1163=>"101101100",
  1164=>"001110000",
  1165=>"100001111",
  1166=>"110111111",
  1167=>"010111011",
  1168=>"110101011",
  1169=>"010100100",
  1170=>"111101110",
  1171=>"111000000",
  1172=>"011111001",
  1173=>"001011011",
  1174=>"100110001",
  1175=>"111111110",
  1176=>"011000110",
  1177=>"000011011",
  1178=>"100011111",
  1179=>"000000111",
  1180=>"000110100",
  1181=>"100101100",
  1182=>"100010111",
  1183=>"010110100",
  1184=>"101100010",
  1185=>"110010011",
  1186=>"011010000",
  1187=>"110000100",
  1188=>"000011100",
  1189=>"101110001",
  1190=>"000010010",
  1191=>"100111000",
  1192=>"101110110",
  1193=>"000010001",
  1194=>"011000101",
  1195=>"000100000",
  1196=>"011010010",
  1197=>"101100111",
  1198=>"110011111",
  1199=>"011001010",
  1200=>"000100111",
  1201=>"000111000",
  1202=>"111101100",
  1203=>"000100000",
  1204=>"110110110",
  1205=>"111110110",
  1206=>"001000000",
  1207=>"110110100",
  1208=>"011001111",
  1209=>"000011000",
  1210=>"011111000",
  1211=>"100100110",
  1212=>"000111000",
  1213=>"101011010",
  1214=>"001011001",
  1215=>"100001001",
  1216=>"111101001",
  1217=>"100000010",
  1218=>"001010110",
  1219=>"000001110",
  1220=>"011011101",
  1221=>"111011111",
  1222=>"101110100",
  1223=>"111000100",
  1224=>"011000111",
  1225=>"100111001",
  1226=>"101100101",
  1227=>"011001110",
  1228=>"100000100",
  1229=>"001001110",
  1230=>"000000010",
  1231=>"111110001",
  1232=>"011111001",
  1233=>"001010101",
  1234=>"000100100",
  1235=>"000000001",
  1236=>"110010010",
  1237=>"000111111",
  1238=>"111011000",
  1239=>"000011000",
  1240=>"000010010",
  1241=>"000101101",
  1242=>"001100000",
  1243=>"111010001",
  1244=>"011110111",
  1245=>"101100110",
  1246=>"111110000",
  1247=>"011000000",
  1248=>"011111010",
  1249=>"100010101",
  1250=>"011001100",
  1251=>"000011000",
  1252=>"110000101",
  1253=>"000000000",
  1254=>"101100000",
  1255=>"001000010",
  1256=>"101111001",
  1257=>"010100000",
  1258=>"001010011",
  1259=>"001101110",
  1260=>"110101111",
  1261=>"010000010",
  1262=>"101000000",
  1263=>"110100010",
  1264=>"111111000",
  1265=>"110100000",
  1266=>"000000001",
  1267=>"000100101",
  1268=>"100101011",
  1269=>"111110010",
  1270=>"101000111",
  1271=>"110111111",
  1272=>"011111010",
  1273=>"110011111",
  1274=>"001000111",
  1275=>"100101001",
  1276=>"110000011",
  1277=>"111001101",
  1278=>"010101010",
  1279=>"111000101",
  1280=>"101000101",
  1281=>"101001110",
  1282=>"100111000",
  1283=>"010111111",
  1284=>"110110100",
  1285=>"111110000",
  1286=>"110110011",
  1287=>"000101001",
  1288=>"010010110",
  1289=>"111111100",
  1290=>"001100010",
  1291=>"010110011",
  1292=>"010101110",
  1293=>"010010011",
  1294=>"010010011",
  1295=>"011000101",
  1296=>"010010000",
  1297=>"001001011",
  1298=>"110110111",
  1299=>"101010100",
  1300=>"011101100",
  1301=>"001111000",
  1302=>"001100000",
  1303=>"101110000",
  1304=>"110010110",
  1305=>"010000011",
  1306=>"100111000",
  1307=>"000101111",
  1308=>"000000110",
  1309=>"001011101",
  1310=>"011010001",
  1311=>"010110100",
  1312=>"111010110",
  1313=>"110000010",
  1314=>"101100100",
  1315=>"010010010",
  1316=>"110111111",
  1317=>"001001110",
  1318=>"000011001",
  1319=>"111011000",
  1320=>"100100011",
  1321=>"010011010",
  1322=>"000011110",
  1323=>"001111111",
  1324=>"000101100",
  1325=>"011111001",
  1326=>"111001001",
  1327=>"010011111",
  1328=>"100111101",
  1329=>"101101000",
  1330=>"010101111",
  1331=>"000111010",
  1332=>"101101011",
  1333=>"111100111",
  1334=>"100100000",
  1335=>"110001111",
  1336=>"010010010",
  1337=>"000001111",
  1338=>"110011010",
  1339=>"101111110",
  1340=>"110100101",
  1341=>"001001000",
  1342=>"110110100",
  1343=>"110010011",
  1344=>"111110001",
  1345=>"101011100",
  1346=>"000010001",
  1347=>"100000010",
  1348=>"010010101",
  1349=>"010001111",
  1350=>"001001110",
  1351=>"101101010",
  1352=>"001010101",
  1353=>"001001110",
  1354=>"101101101",
  1355=>"000111101",
  1356=>"011000101",
  1357=>"100011110",
  1358=>"100110111",
  1359=>"000111100",
  1360=>"001100000",
  1361=>"001000111",
  1362=>"110101101",
  1363=>"101001000",
  1364=>"110111000",
  1365=>"001111010",
  1366=>"000100011",
  1367=>"001110100",
  1368=>"001001001",
  1369=>"010010111",
  1370=>"110000111",
  1371=>"001000001",
  1372=>"000101001",
  1373=>"010100011",
  1374=>"111010001",
  1375=>"001010000",
  1376=>"011110111",
  1377=>"010100111",
  1378=>"010001000",
  1379=>"001000000",
  1380=>"000001100",
  1381=>"111101111",
  1382=>"010111001",
  1383=>"101101110",
  1384=>"100000010",
  1385=>"000011001",
  1386=>"101001010",
  1387=>"011010101",
  1388=>"010100110",
  1389=>"010101010",
  1390=>"010001111",
  1391=>"001100011",
  1392=>"000111100",
  1393=>"111111101",
  1394=>"100011010",
  1395=>"100111000",
  1396=>"011010000",
  1397=>"100111001",
  1398=>"011011000",
  1399=>"000010011",
  1400=>"000010111",
  1401=>"100000111",
  1402=>"100111001",
  1403=>"000100100",
  1404=>"010000011",
  1405=>"011000011",
  1406=>"011101000",
  1407=>"110000001",
  1408=>"111111111",
  1409=>"001110110",
  1410=>"111011101",
  1411=>"101110111",
  1412=>"011110001",
  1413=>"100000101",
  1414=>"011110100",
  1415=>"110101110",
  1416=>"000000000",
  1417=>"100110101",
  1418=>"100001011",
  1419=>"111100100",
  1420=>"110111000",
  1421=>"011011011",
  1422=>"101100100",
  1423=>"111110001",
  1424=>"000011110",
  1425=>"010010010",
  1426=>"001000101",
  1427=>"010011010",
  1428=>"111001111",
  1429=>"011010111",
  1430=>"000110111",
  1431=>"001010011",
  1432=>"001110010",
  1433=>"010000001",
  1434=>"001011111",
  1435=>"000101110",
  1436=>"001010001",
  1437=>"110101100",
  1438=>"001000010",
  1439=>"100110110",
  1440=>"100110100",
  1441=>"001011001",
  1442=>"111100111",
  1443=>"001001011",
  1444=>"110001010",
  1445=>"001011110",
  1446=>"000001101",
  1447=>"101000101",
  1448=>"111110100",
  1449=>"001000000",
  1450=>"000000110",
  1451=>"001010010",
  1452=>"010000011",
  1453=>"110011101",
  1454=>"110100000",
  1455=>"000111001",
  1456=>"001001101",
  1457=>"001110000",
  1458=>"001110101",
  1459=>"010001011",
  1460=>"000111110",
  1461=>"110000010",
  1462=>"011000110",
  1463=>"100000100",
  1464=>"111011001",
  1465=>"011001011",
  1466=>"000110000",
  1467=>"111111110",
  1468=>"001110111",
  1469=>"010101110",
  1470=>"111001001",
  1471=>"111111110",
  1472=>"111101101",
  1473=>"011011010",
  1474=>"111011001",
  1475=>"110001001",
  1476=>"111111010",
  1477=>"010010001",
  1478=>"000000000",
  1479=>"110111000",
  1480=>"010010100",
  1481=>"010111000",
  1482=>"011111111",
  1483=>"101000010",
  1484=>"010001001",
  1485=>"110010101",
  1486=>"001001000",
  1487=>"100101011",
  1488=>"010010011",
  1489=>"110110001",
  1490=>"011000100",
  1491=>"011011011",
  1492=>"011000000",
  1493=>"111111010",
  1494=>"110111111",
  1495=>"000011110",
  1496=>"001000111",
  1497=>"101110000",
  1498=>"110000101",
  1499=>"111110010",
  1500=>"010011111",
  1501=>"011001011",
  1502=>"001100011",
  1503=>"001011111",
  1504=>"010111100",
  1505=>"001111001",
  1506=>"010100000",
  1507=>"010001101",
  1508=>"010000010",
  1509=>"111010011",
  1510=>"111001011",
  1511=>"010101000",
  1512=>"010100010",
  1513=>"101001000",
  1514=>"000101101",
  1515=>"110001110",
  1516=>"101100110",
  1517=>"100101110",
  1518=>"011100100",
  1519=>"110100100",
  1520=>"100000000",
  1521=>"010100011",
  1522=>"111010001",
  1523=>"101101100",
  1524=>"010000110",
  1525=>"111001000",
  1526=>"110111101",
  1527=>"010011001",
  1528=>"011010000",
  1529=>"001000010",
  1530=>"110110100",
  1531=>"110100111",
  1532=>"000101111",
  1533=>"111010000",
  1534=>"000010000",
  1535=>"111111000",
  1536=>"110110011",
  1537=>"110001100",
  1538=>"101101111",
  1539=>"000111100",
  1540=>"010100000",
  1541=>"111001101",
  1542=>"111001000",
  1543=>"001101100",
  1544=>"100001100",
  1545=>"111011101",
  1546=>"001000110",
  1547=>"100101110",
  1548=>"101011101",
  1549=>"001110100",
  1550=>"100001110",
  1551=>"011000100",
  1552=>"100101101",
  1553=>"111010011",
  1554=>"010010000",
  1555=>"100110010",
  1556=>"100010010",
  1557=>"000101010",
  1558=>"001111110",
  1559=>"111010001",
  1560=>"101110100",
  1561=>"000011101",
  1562=>"010001001",
  1563=>"010001001",
  1564=>"010011000",
  1565=>"000110100",
  1566=>"101110101",
  1567=>"101101101",
  1568=>"010001100",
  1569=>"110010000",
  1570=>"000001011",
  1571=>"000001000",
  1572=>"110110101",
  1573=>"100101011",
  1574=>"101110110",
  1575=>"110010111",
  1576=>"111110110",
  1577=>"111010011",
  1578=>"010000011",
  1579=>"001000010",
  1580=>"011001010",
  1581=>"011110000",
  1582=>"011000111",
  1583=>"000011010",
  1584=>"111001111",
  1585=>"011000000",
  1586=>"001100110",
  1587=>"101111111",
  1588=>"011001111",
  1589=>"010101000",
  1590=>"101010111",
  1591=>"101111001",
  1592=>"010101011",
  1593=>"100100100",
  1594=>"101100011",
  1595=>"101101001",
  1596=>"101110111",
  1597=>"111000110",
  1598=>"100110110",
  1599=>"111101000",
  1600=>"110010111",
  1601=>"010000000",
  1602=>"101011000",
  1603=>"110000110",
  1604=>"010111000",
  1605=>"010110100",
  1606=>"001101000",
  1607=>"101100111",
  1608=>"010101001",
  1609=>"111101101",
  1610=>"001100001",
  1611=>"001011010",
  1612=>"100101011",
  1613=>"101100010",
  1614=>"110001000",
  1615=>"111110110",
  1616=>"010000001",
  1617=>"011000010",
  1618=>"011011010",
  1619=>"001011000",
  1620=>"111100001",
  1621=>"010100001",
  1622=>"000001011",
  1623=>"000011110",
  1624=>"110100001",
  1625=>"010000100",
  1626=>"011001001",
  1627=>"000111111",
  1628=>"001111100",
  1629=>"111011010",
  1630=>"110000010",
  1631=>"101111000",
  1632=>"000000101",
  1633=>"001000001",
  1634=>"000101111",
  1635=>"001000000",
  1636=>"101000011",
  1637=>"101001110",
  1638=>"100000111",
  1639=>"010101111",
  1640=>"101110010",
  1641=>"001011000",
  1642=>"010101101",
  1643=>"110110000",
  1644=>"000101011",
  1645=>"001011010",
  1646=>"000111111",
  1647=>"011001110",
  1648=>"010100101",
  1649=>"010010100",
  1650=>"101011111",
  1651=>"110000000",
  1652=>"000000010",
  1653=>"111100101",
  1654=>"000110000",
  1655=>"100011010",
  1656=>"000111111",
  1657=>"100010100",
  1658=>"010101001",
  1659=>"110100110",
  1660=>"111000101",
  1661=>"010001110",
  1662=>"101100000",
  1663=>"100111101",
  1664=>"101000000",
  1665=>"001011100",
  1666=>"010000100",
  1667=>"010111101",
  1668=>"000110010",
  1669=>"011011100",
  1670=>"110110011",
  1671=>"010010010",
  1672=>"001101110",
  1673=>"100100110",
  1674=>"001001001",
  1675=>"110101101",
  1676=>"010101011",
  1677=>"011000100",
  1678=>"111100100",
  1679=>"010000111",
  1680=>"110100001",
  1681=>"001100001",
  1682=>"001111111",
  1683=>"111001011",
  1684=>"001101101",
  1685=>"001000011",
  1686=>"111111011",
  1687=>"101011000",
  1688=>"001011010",
  1689=>"011000101",
  1690=>"011011101",
  1691=>"101000111",
  1692=>"011100000",
  1693=>"100110111",
  1694=>"101010000",
  1695=>"011001110",
  1696=>"101101000",
  1697=>"011110110",
  1698=>"110000100",
  1699=>"100010001",
  1700=>"001111001",
  1701=>"000011111",
  1702=>"110010010",
  1703=>"000011000",
  1704=>"011011000",
  1705=>"010010011",
  1706=>"111000001",
  1707=>"000101010",
  1708=>"101101111",
  1709=>"000000100",
  1710=>"011101010",
  1711=>"110010001",
  1712=>"111011010",
  1713=>"010010110",
  1714=>"111101110",
  1715=>"010011101",
  1716=>"100100001",
  1717=>"011100101",
  1718=>"000100101",
  1719=>"001010100",
  1720=>"110100111",
  1721=>"111101110",
  1722=>"000111110",
  1723=>"111010111",
  1724=>"101100000",
  1725=>"110111010",
  1726=>"000001001",
  1727=>"110011111",
  1728=>"100111010",
  1729=>"010110100",
  1730=>"111101101",
  1731=>"100110010",
  1732=>"111011001",
  1733=>"101100110",
  1734=>"111010111",
  1735=>"111011110",
  1736=>"111111111",
  1737=>"000101011",
  1738=>"100100001",
  1739=>"011100000",
  1740=>"010100011",
  1741=>"010101011",
  1742=>"000011000",
  1743=>"000100101",
  1744=>"001110011",
  1745=>"110010101",
  1746=>"001111100",
  1747=>"100001000",
  1748=>"101110100",
  1749=>"010101011",
  1750=>"110110111",
  1751=>"110001100",
  1752=>"000001111",
  1753=>"101000001",
  1754=>"110011010",
  1755=>"010010100",
  1756=>"010000001",
  1757=>"111001001",
  1758=>"101100110",
  1759=>"011010101",
  1760=>"000110111",
  1761=>"001011000",
  1762=>"110000101",
  1763=>"001101000",
  1764=>"010101100",
  1765=>"111011001",
  1766=>"111110110",
  1767=>"010101100",
  1768=>"111111111",
  1769=>"101011000",
  1770=>"000110100",
  1771=>"000110110",
  1772=>"011110111",
  1773=>"100010111",
  1774=>"111000001",
  1775=>"110010001",
  1776=>"011000011",
  1777=>"100010010",
  1778=>"111000101",
  1779=>"010001101",
  1780=>"111111111",
  1781=>"100010100",
  1782=>"110111111",
  1783=>"110110001",
  1784=>"100001110",
  1785=>"100000111",
  1786=>"011001111",
  1787=>"110011111",
  1788=>"010010001",
  1789=>"110110101",
  1790=>"010011110",
  1791=>"100111111",
  1792=>"001100010",
  1793=>"001111111",
  1794=>"101100011",
  1795=>"011100000",
  1796=>"110011110",
  1797=>"000100001",
  1798=>"101111001",
  1799=>"110111010",
  1800=>"000100101",
  1801=>"011110101",
  1802=>"001010010",
  1803=>"111011001",
  1804=>"111001010",
  1805=>"010111110",
  1806=>"000010111",
  1807=>"111011011",
  1808=>"010000111",
  1809=>"001001101",
  1810=>"111000011",
  1811=>"001001101",
  1812=>"111111101",
  1813=>"110010100",
  1814=>"110101101",
  1815=>"010011111",
  1816=>"010000011",
  1817=>"000010110",
  1818=>"000100110",
  1819=>"111100110",
  1820=>"100000100",
  1821=>"111001011",
  1822=>"010110101",
  1823=>"101000010",
  1824=>"111100100",
  1825=>"010000010",
  1826=>"001001111",
  1827=>"101100010",
  1828=>"110001110",
  1829=>"110100011",
  1830=>"001100100",
  1831=>"110001010",
  1832=>"001000101",
  1833=>"010110111",
  1834=>"101111010",
  1835=>"101000111",
  1836=>"111001010",
  1837=>"100001001",
  1838=>"011011001",
  1839=>"010110100",
  1840=>"010001000",
  1841=>"000111010",
  1842=>"000000000",
  1843=>"000110011",
  1844=>"101100001",
  1845=>"001011110",
  1846=>"001011101",
  1847=>"110111101",
  1848=>"111010100",
  1849=>"011111000",
  1850=>"001100011",
  1851=>"101111000",
  1852=>"110100110",
  1853=>"000110110",
  1854=>"000110101",
  1855=>"010111011",
  1856=>"011000101",
  1857=>"011101111",
  1858=>"010111111",
  1859=>"111100011",
  1860=>"111111001",
  1861=>"001100101",
  1862=>"101110000",
  1863=>"110111001",
  1864=>"110110011",
  1865=>"101100111",
  1866=>"000110101",
  1867=>"100001101",
  1868=>"000011001",
  1869=>"000100000",
  1870=>"001000111",
  1871=>"101010110",
  1872=>"010111010",
  1873=>"100010100",
  1874=>"011110110",
  1875=>"101101001",
  1876=>"000011000",
  1877=>"101101100",
  1878=>"010001000",
  1879=>"110010110",
  1880=>"100010011",
  1881=>"101010111",
  1882=>"000001010",
  1883=>"110010010",
  1884=>"111110010",
  1885=>"101000011",
  1886=>"011110110",
  1887=>"100101010",
  1888=>"010101110",
  1889=>"001001101",
  1890=>"100001010",
  1891=>"101010111",
  1892=>"001010010",
  1893=>"000110001",
  1894=>"001001110",
  1895=>"001100110",
  1896=>"100101001",
  1897=>"111010010",
  1898=>"010000010",
  1899=>"110101101",
  1900=>"000000011",
  1901=>"001101011",
  1902=>"010101001",
  1903=>"001010111",
  1904=>"010001101",
  1905=>"001100001",
  1906=>"100110000",
  1907=>"101001000",
  1908=>"000010111",
  1909=>"011011011",
  1910=>"101111100",
  1911=>"111110101",
  1912=>"011100000",
  1913=>"010000100",
  1914=>"101100110",
  1915=>"111110011",
  1916=>"101010100",
  1917=>"010011010",
  1918=>"000100000",
  1919=>"111010100",
  1920=>"010110101",
  1921=>"100011001",
  1922=>"111100101",
  1923=>"000011101",
  1924=>"101111001",
  1925=>"110111100",
  1926=>"111001011",
  1927=>"001000000",
  1928=>"100001010",
  1929=>"010101011",
  1930=>"111010001",
  1931=>"101100111",
  1932=>"100010100",
  1933=>"011001110",
  1934=>"111001000",
  1935=>"100000100",
  1936=>"011101100",
  1937=>"000100010",
  1938=>"010001111",
  1939=>"000000110",
  1940=>"101111000",
  1941=>"111101010",
  1942=>"101101000",
  1943=>"011100010",
  1944=>"001011101",
  1945=>"010001000",
  1946=>"111110100",
  1947=>"001101101",
  1948=>"000111000",
  1949=>"001000100",
  1950=>"110100110",
  1951=>"100000001",
  1952=>"000110010",
  1953=>"100000001",
  1954=>"010011011",
  1955=>"000011100",
  1956=>"100001100",
  1957=>"001100000",
  1958=>"001110101",
  1959=>"110010000",
  1960=>"100000000",
  1961=>"101101111",
  1962=>"010111011",
  1963=>"101100011",
  1964=>"111000000",
  1965=>"100100101",
  1966=>"110001101",
  1967=>"000100111",
  1968=>"110011001",
  1969=>"010111111",
  1970=>"101110111",
  1971=>"000100001",
  1972=>"100110001",
  1973=>"100111000",
  1974=>"101101000",
  1975=>"010111000",
  1976=>"001000010",
  1977=>"100111110",
  1978=>"111100101",
  1979=>"100101110",
  1980=>"111101011",
  1981=>"100011000",
  1982=>"110100000",
  1983=>"010010010",
  1984=>"000100101",
  1985=>"110111110",
  1986=>"000010001",
  1987=>"101001000",
  1988=>"111110111",
  1989=>"101100110",
  1990=>"000110101",
  1991=>"101111000",
  1992=>"101010110",
  1993=>"110011011",
  1994=>"101100111",
  1995=>"001110111",
  1996=>"111010010",
  1997=>"011100101",
  1998=>"111011010",
  1999=>"000011010",
  2000=>"001101100",
  2001=>"110101111",
  2002=>"110101010",
  2003=>"010110011",
  2004=>"100000000",
  2005=>"000110011",
  2006=>"001100110",
  2007=>"000000000",
  2008=>"010010110",
  2009=>"110110000",
  2010=>"100000000",
  2011=>"111100110",
  2012=>"000000010",
  2013=>"001101100",
  2014=>"000001010",
  2015=>"110000000",
  2016=>"011111101",
  2017=>"101100010",
  2018=>"000110111",
  2019=>"000001001",
  2020=>"011101000",
  2021=>"110000100",
  2022=>"010100000",
  2023=>"010110101",
  2024=>"010010100",
  2025=>"000000101",
  2026=>"101001010",
  2027=>"101111111",
  2028=>"011111001",
  2029=>"110100101",
  2030=>"011110001",
  2031=>"000011011",
  2032=>"101100100",
  2033=>"011101110",
  2034=>"101100010",
  2035=>"110010001",
  2036=>"001101101",
  2037=>"111001111",
  2038=>"101010000",
  2039=>"110011001",
  2040=>"111111111",
  2041=>"111111011",
  2042=>"110101010",
  2043=>"001000000",
  2044=>"100101110",
  2045=>"010000101",
  2046=>"001111111",
  2047=>"011011001",
  2048=>"011110101",
  2049=>"110100001",
  2050=>"011001000",
  2051=>"010011101",
  2052=>"010111000",
  2053=>"010010010",
  2054=>"000000100",
  2055=>"100100101",
  2056=>"100111011",
  2057=>"100101010",
  2058=>"111101000",
  2059=>"010001000",
  2060=>"010000000",
  2061=>"010000101",
  2062=>"001110100",
  2063=>"000110110",
  2064=>"000110011",
  2065=>"011100110",
  2066=>"010011111",
  2067=>"101000101",
  2068=>"101010001",
  2069=>"110011111",
  2070=>"010011010",
  2071=>"000001100",
  2072=>"010100011",
  2073=>"001010100",
  2074=>"001110010",
  2075=>"011101011",
  2076=>"001001011",
  2077=>"101110101",
  2078=>"110110100",
  2079=>"000110001",
  2080=>"000000101",
  2081=>"110111110",
  2082=>"001100100",
  2083=>"010001000",
  2084=>"100111111",
  2085=>"000000010",
  2086=>"000110010",
  2087=>"100110010",
  2088=>"001111100",
  2089=>"101010101",
  2090=>"101001111",
  2091=>"101000110",
  2092=>"111101100",
  2093=>"000011010",
  2094=>"000000101",
  2095=>"000011110",
  2096=>"001111110",
  2097=>"100101111",
  2098=>"001101010",
  2099=>"010000001",
  2100=>"010110111",
  2101=>"111010001",
  2102=>"000100110",
  2103=>"001010101",
  2104=>"101000010",
  2105=>"011110111",
  2106=>"101100111",
  2107=>"111101110",
  2108=>"111010000",
  2109=>"001100100",
  2110=>"111010101",
  2111=>"000110001",
  2112=>"000101111",
  2113=>"000011001",
  2114=>"000110011",
  2115=>"000000100",
  2116=>"010010010",
  2117=>"001111101",
  2118=>"010011000",
  2119=>"110111011",
  2120=>"101001100",
  2121=>"110101001",
  2122=>"101110110",
  2123=>"110000110",
  2124=>"000000110",
  2125=>"111101101",
  2126=>"010010111",
  2127=>"110000010",
  2128=>"110000101",
  2129=>"111111000",
  2130=>"010101100",
  2131=>"011111010",
  2132=>"010110000",
  2133=>"000110100",
  2134=>"111011110",
  2135=>"100111111",
  2136=>"010011001",
  2137=>"000110110",
  2138=>"011100110",
  2139=>"111111101",
  2140=>"111111011",
  2141=>"011011011",
  2142=>"001001011",
  2143=>"111100000",
  2144=>"011111001",
  2145=>"101111011",
  2146=>"111111111",
  2147=>"010010010",
  2148=>"100001010",
  2149=>"110010000",
  2150=>"001100110",
  2151=>"000010010",
  2152=>"110001111",
  2153=>"110011010",
  2154=>"110000010",
  2155=>"011101110",
  2156=>"101101001",
  2157=>"101110010",
  2158=>"000111010",
  2159=>"111100110",
  2160=>"111101001",
  2161=>"011101101",
  2162=>"100110111",
  2163=>"100011100",
  2164=>"111110110",
  2165=>"111001100",
  2166=>"101100101",
  2167=>"100001110",
  2168=>"010001010",
  2169=>"101011011",
  2170=>"111001001",
  2171=>"111010101",
  2172=>"100100010",
  2173=>"011000100",
  2174=>"111011111",
  2175=>"111000110",
  2176=>"001101111",
  2177=>"100001110",
  2178=>"010111101",
  2179=>"111101110",
  2180=>"001101100",
  2181=>"100110011",
  2182=>"000110110",
  2183=>"011111010",
  2184=>"000101000",
  2185=>"001000000",
  2186=>"111000011",
  2187=>"001011000",
  2188=>"000110001",
  2189=>"011001011",
  2190=>"110001000",
  2191=>"001000010",
  2192=>"100010101",
  2193=>"100110110",
  2194=>"011111110",
  2195=>"111110011",
  2196=>"111110110",
  2197=>"001010100",
  2198=>"111111100",
  2199=>"110001011",
  2200=>"011011101",
  2201=>"010010001",
  2202=>"011111111",
  2203=>"100000010",
  2204=>"010101100",
  2205=>"011101110",
  2206=>"000100001",
  2207=>"011010000",
  2208=>"100001100",
  2209=>"011010110",
  2210=>"111100011",
  2211=>"110111111",
  2212=>"110111100",
  2213=>"010011000",
  2214=>"100011100",
  2215=>"000001000",
  2216=>"111001100",
  2217=>"110111110",
  2218=>"001010000",
  2219=>"001100010",
  2220=>"000101010",
  2221=>"010001010",
  2222=>"101110111",
  2223=>"110000100",
  2224=>"011111101",
  2225=>"011101100",
  2226=>"111010101",
  2227=>"011001010",
  2228=>"111111110",
  2229=>"100111111",
  2230=>"100100110",
  2231=>"011000101",
  2232=>"100100110",
  2233=>"111100000",
  2234=>"011010000",
  2235=>"011110001",
  2236=>"100011110",
  2237=>"100001011",
  2238=>"111111110",
  2239=>"000111101",
  2240=>"110110001",
  2241=>"000100100",
  2242=>"010010100",
  2243=>"100000011",
  2244=>"110001111",
  2245=>"101111101",
  2246=>"000010011",
  2247=>"000010100",
  2248=>"000011010",
  2249=>"110000000",
  2250=>"011101011",
  2251=>"100110010",
  2252=>"100011101",
  2253=>"010011010",
  2254=>"011101001",
  2255=>"110101110",
  2256=>"101111011",
  2257=>"110001110",
  2258=>"000011100",
  2259=>"101001010",
  2260=>"110010100",
  2261=>"110100101",
  2262=>"110111001",
  2263=>"001111111",
  2264=>"011010101",
  2265=>"100111001",
  2266=>"101111000",
  2267=>"100101011",
  2268=>"101001000",
  2269=>"011100011",
  2270=>"000000111",
  2271=>"000111110",
  2272=>"000101010",
  2273=>"000000011",
  2274=>"101011010",
  2275=>"000010000",
  2276=>"010101101",
  2277=>"011101001",
  2278=>"110011010",
  2279=>"001111001",
  2280=>"110111000",
  2281=>"110111010",
  2282=>"100011010",
  2283=>"111011110",
  2284=>"000100101",
  2285=>"101010101",
  2286=>"101011000",
  2287=>"011000111",
  2288=>"011001001",
  2289=>"001011101",
  2290=>"001110000",
  2291=>"000011111",
  2292=>"110000000",
  2293=>"100111000",
  2294=>"101010011",
  2295=>"110000000",
  2296=>"000101011",
  2297=>"100111001",
  2298=>"000111011",
  2299=>"000010001",
  2300=>"011110110",
  2301=>"000110111",
  2302=>"011001101",
  2303=>"111110011",
  2304=>"111100111",
  2305=>"111001011",
  2306=>"000100101",
  2307=>"011101111",
  2308=>"110000000",
  2309=>"100111111",
  2310=>"100100000",
  2311=>"110101110",
  2312=>"110001000",
  2313=>"101000111",
  2314=>"101010110",
  2315=>"011001000",
  2316=>"000100000",
  2317=>"100001100",
  2318=>"110010001",
  2319=>"111110001",
  2320=>"011100010",
  2321=>"100001011",
  2322=>"011001000",
  2323=>"111111111",
  2324=>"110011010",
  2325=>"001011010",
  2326=>"110001000",
  2327=>"100101001",
  2328=>"000111110",
  2329=>"010010101",
  2330=>"001111111",
  2331=>"111000110",
  2332=>"110110001",
  2333=>"001111001",
  2334=>"101110000",
  2335=>"110000001",
  2336=>"001110110",
  2337=>"101011101",
  2338=>"111001110",
  2339=>"110011010",
  2340=>"001101101",
  2341=>"001000010",
  2342=>"001010000",
  2343=>"000111011",
  2344=>"001110100",
  2345=>"001000110",
  2346=>"000011001",
  2347=>"100010010",
  2348=>"000101010",
  2349=>"001100001",
  2350=>"111000010",
  2351=>"101110000",
  2352=>"100010000",
  2353=>"000001000",
  2354=>"000010001",
  2355=>"011100100",
  2356=>"001010111",
  2357=>"011100011",
  2358=>"110001010",
  2359=>"111101011",
  2360=>"000000010",
  2361=>"001011000",
  2362=>"000011101",
  2363=>"000011001",
  2364=>"001111010",
  2365=>"011011000",
  2366=>"011000011",
  2367=>"010000111",
  2368=>"101000110",
  2369=>"110010111",
  2370=>"100100110",
  2371=>"010000111",
  2372=>"111000100",
  2373=>"101100111",
  2374=>"111010111",
  2375=>"000101000",
  2376=>"101101111",
  2377=>"111110011",
  2378=>"111011110",
  2379=>"111100000",
  2380=>"010101001",
  2381=>"011000111",
  2382=>"100110011",
  2383=>"111010110",
  2384=>"110101001",
  2385=>"101011000",
  2386=>"110001011",
  2387=>"101111110",
  2388=>"010001000",
  2389=>"011100111",
  2390=>"110100001",
  2391=>"001010101",
  2392=>"010001010",
  2393=>"001010001",
  2394=>"110100000",
  2395=>"111011001",
  2396=>"010001101",
  2397=>"010110110",
  2398=>"010110011",
  2399=>"000101110",
  2400=>"000110011",
  2401=>"010110101",
  2402=>"111110001",
  2403=>"100111010",
  2404=>"010001110",
  2405=>"101101010",
  2406=>"110010110",
  2407=>"100011010",
  2408=>"001000110",
  2409=>"001001111",
  2410=>"000110101",
  2411=>"111011110",
  2412=>"011100001",
  2413=>"101110010",
  2414=>"010101000",
  2415=>"001011001",
  2416=>"101000110",
  2417=>"111000001",
  2418=>"110101100",
  2419=>"011110110",
  2420=>"110100110",
  2421=>"111111011",
  2422=>"100011010",
  2423=>"010101101",
  2424=>"000100011",
  2425=>"110001011",
  2426=>"010001010",
  2427=>"000111100",
  2428=>"100100011",
  2429=>"101110011",
  2430=>"110101010",
  2431=>"110011101",
  2432=>"101001100",
  2433=>"001101011",
  2434=>"101000011",
  2435=>"001000101",
  2436=>"011111110",
  2437=>"011110010",
  2438=>"000010110",
  2439=>"101010010",
  2440=>"001011001",
  2441=>"111111101",
  2442=>"010001001",
  2443=>"101101101",
  2444=>"010100010",
  2445=>"010100010",
  2446=>"000110011",
  2447=>"100011001",
  2448=>"111101001",
  2449=>"111111111",
  2450=>"010001010",
  2451=>"011111100",
  2452=>"001100010",
  2453=>"011000101",
  2454=>"010011011",
  2455=>"101010100",
  2456=>"110110010",
  2457=>"001000011",
  2458=>"101010001",
  2459=>"110011001",
  2460=>"101110110",
  2461=>"110110000",
  2462=>"011011110",
  2463=>"101011011",
  2464=>"000101011",
  2465=>"111110011",
  2466=>"110101111",
  2467=>"010111101",
  2468=>"011100101",
  2469=>"111110100",
  2470=>"011100010",
  2471=>"101100110",
  2472=>"110101010",
  2473=>"010110000",
  2474=>"100011111",
  2475=>"001000011",
  2476=>"010110001",
  2477=>"110001000",
  2478=>"001101001",
  2479=>"101110000",
  2480=>"010000000",
  2481=>"001111101",
  2482=>"010010101",
  2483=>"000011111",
  2484=>"101010111",
  2485=>"110001110",
  2486=>"101110110",
  2487=>"101110010",
  2488=>"111001001",
  2489=>"010111000",
  2490=>"101110100",
  2491=>"010001110",
  2492=>"111111111",
  2493=>"101111101",
  2494=>"001101111",
  2495=>"101110000",
  2496=>"100011100",
  2497=>"011011000",
  2498=>"101111001",
  2499=>"110110010",
  2500=>"001111101",
  2501=>"001001110",
  2502=>"101111110",
  2503=>"111111000",
  2504=>"011011010",
  2505=>"111001111",
  2506=>"010010110",
  2507=>"101000011",
  2508=>"010010111",
  2509=>"100011100",
  2510=>"011110001",
  2511=>"100100001",
  2512=>"000111011",
  2513=>"001011000",
  2514=>"010100111",
  2515=>"111100101",
  2516=>"100001110",
  2517=>"010101111",
  2518=>"000100110",
  2519=>"110101111",
  2520=>"111111101",
  2521=>"110101110",
  2522=>"100001010",
  2523=>"100100010",
  2524=>"110010100",
  2525=>"010110100",
  2526=>"100001001",
  2527=>"000100011",
  2528=>"100110001",
  2529=>"111011111",
  2530=>"011110100",
  2531=>"111101100",
  2532=>"101101100",
  2533=>"000000001",
  2534=>"110111100",
  2535=>"000011111",
  2536=>"100001101",
  2537=>"001011110",
  2538=>"100110010",
  2539=>"011000010",
  2540=>"000110101",
  2541=>"101011111",
  2542=>"101111010",
  2543=>"101010000",
  2544=>"000000010",
  2545=>"011110101",
  2546=>"010000001",
  2547=>"011001110",
  2548=>"101001000",
  2549=>"010011100",
  2550=>"100100111",
  2551=>"010010000",
  2552=>"101101011",
  2553=>"001001110",
  2554=>"101001010",
  2555=>"010011101",
  2556=>"010011111",
  2557=>"110000101",
  2558=>"101110001",
  2559=>"010011100",
  2560=>"000111101",
  2561=>"001101011",
  2562=>"000001011",
  2563=>"001111101",
  2564=>"000100111",
  2565=>"101010100",
  2566=>"011010000",
  2567=>"100110111",
  2568=>"000110110",
  2569=>"001010010",
  2570=>"111111010",
  2571=>"110010110",
  2572=>"011110001",
  2573=>"001010110",
  2574=>"111000010",
  2575=>"001000011",
  2576=>"111100110",
  2577=>"101101100",
  2578=>"001110000",
  2579=>"010000010",
  2580=>"001000000",
  2581=>"001101110",
  2582=>"000101110",
  2583=>"010111101",
  2584=>"101001110",
  2585=>"100010000",
  2586=>"010010001",
  2587=>"110011000",
  2588=>"000110111",
  2589=>"100001111",
  2590=>"111111100",
  2591=>"000111110",
  2592=>"000110001",
  2593=>"010010100",
  2594=>"000110011",
  2595=>"100001100",
  2596=>"011101100",
  2597=>"000111110",
  2598=>"001101010",
  2599=>"100101100",
  2600=>"011011101",
  2601=>"000000001",
  2602=>"101011010",
  2603=>"000111011",
  2604=>"100010101",
  2605=>"000100100",
  2606=>"010100110",
  2607=>"111100110",
  2608=>"100111100",
  2609=>"010100110",
  2610=>"010011000",
  2611=>"100111000",
  2612=>"000001111",
  2613=>"001010100",
  2614=>"000101011",
  2615=>"100100101",
  2616=>"010011000",
  2617=>"001011111",
  2618=>"111001100",
  2619=>"111010010",
  2620=>"011001110",
  2621=>"110001110",
  2622=>"000100101",
  2623=>"010000101",
  2624=>"110000000",
  2625=>"011110000",
  2626=>"101000111",
  2627=>"011101000",
  2628=>"110000111",
  2629=>"110011110",
  2630=>"001111111",
  2631=>"110000100",
  2632=>"110110011",
  2633=>"111111111",
  2634=>"000101000",
  2635=>"010110101",
  2636=>"001101011",
  2637=>"000111101",
  2638=>"100010101",
  2639=>"101100110",
  2640=>"100001100",
  2641=>"000001000",
  2642=>"111101101",
  2643=>"110000011",
  2644=>"110110000",
  2645=>"010011100",
  2646=>"010111010",
  2647=>"100111111",
  2648=>"010111100",
  2649=>"100101000",
  2650=>"000000100",
  2651=>"111001101",
  2652=>"000010010",
  2653=>"001001000",
  2654=>"100110110",
  2655=>"101101101",
  2656=>"100000101",
  2657=>"000111111",
  2658=>"110000111",
  2659=>"100100000",
  2660=>"111000101",
  2661=>"001111101",
  2662=>"010011001",
  2663=>"101001010",
  2664=>"000000001",
  2665=>"101000000",
  2666=>"111011010",
  2667=>"001001110",
  2668=>"000000001",
  2669=>"100010100",
  2670=>"101100010",
  2671=>"010111100",
  2672=>"000001001",
  2673=>"111100100",
  2674=>"110011100",
  2675=>"101000010",
  2676=>"110110001",
  2677=>"001110100",
  2678=>"010001011",
  2679=>"010000100",
  2680=>"100100010",
  2681=>"111010101",
  2682=>"000001111",
  2683=>"000001101",
  2684=>"011110010",
  2685=>"111000000",
  2686=>"000001110",
  2687=>"001010000",
  2688=>"110001001",
  2689=>"010010100",
  2690=>"100100010",
  2691=>"001010001",
  2692=>"010111101",
  2693=>"010100101",
  2694=>"010011010",
  2695=>"001101100",
  2696=>"110101111",
  2697=>"110011000",
  2698=>"100010101",
  2699=>"100100110",
  2700=>"110111101",
  2701=>"000100000",
  2702=>"101111000",
  2703=>"101000010",
  2704=>"110111111",
  2705=>"001011111",
  2706=>"111111011",
  2707=>"101111000",
  2708=>"100011011",
  2709=>"000100010",
  2710=>"001000101",
  2711=>"101101010",
  2712=>"000001101",
  2713=>"001011010",
  2714=>"010101100",
  2715=>"000110111",
  2716=>"001000111",
  2717=>"000101000",
  2718=>"110001010",
  2719=>"111010101",
  2720=>"111101101",
  2721=>"100001110",
  2722=>"010001000",
  2723=>"000000111",
  2724=>"111110110",
  2725=>"101100101",
  2726=>"010100101",
  2727=>"001111000",
  2728=>"110110001",
  2729=>"100111101",
  2730=>"100100001",
  2731=>"101011010",
  2732=>"101000111",
  2733=>"010110111",
  2734=>"111010010",
  2735=>"001110010",
  2736=>"011110110",
  2737=>"010011101",
  2738=>"011011001",
  2739=>"010000100",
  2740=>"100001001",
  2741=>"001101001",
  2742=>"010111001",
  2743=>"101111010",
  2744=>"011111010",
  2745=>"000000100",
  2746=>"100011011",
  2747=>"010111011",
  2748=>"100000111",
  2749=>"100110000",
  2750=>"000110000",
  2751=>"101011101",
  2752=>"011110110",
  2753=>"110111011",
  2754=>"001000100",
  2755=>"101001101",
  2756=>"000010010",
  2757=>"001110110",
  2758=>"111101010",
  2759=>"000011011",
  2760=>"101100100",
  2761=>"111111001",
  2762=>"011000101",
  2763=>"110000011",
  2764=>"011001000",
  2765=>"010110000",
  2766=>"100101000",
  2767=>"100111100",
  2768=>"011000010",
  2769=>"101111000",
  2770=>"010001011",
  2771=>"001000100",
  2772=>"010110010",
  2773=>"011010101",
  2774=>"000011100",
  2775=>"010101011",
  2776=>"000100010",
  2777=>"100010111",
  2778=>"011001101",
  2779=>"011111000",
  2780=>"000000110",
  2781=>"110011000",
  2782=>"110111011",
  2783=>"110101101",
  2784=>"000000100",
  2785=>"110100000",
  2786=>"111000000",
  2787=>"000100000",
  2788=>"101111001",
  2789=>"000001011",
  2790=>"101111010",
  2791=>"001111110",
  2792=>"011101110",
  2793=>"110000000",
  2794=>"101010101",
  2795=>"011111011",
  2796=>"010000011",
  2797=>"110110100",
  2798=>"110100011",
  2799=>"110111000",
  2800=>"011000000",
  2801=>"100010110",
  2802=>"110011001",
  2803=>"101110011",
  2804=>"000000011",
  2805=>"100111101",
  2806=>"111101101",
  2807=>"010111110",
  2808=>"111101001",
  2809=>"001111010",
  2810=>"000111111",
  2811=>"001110000",
  2812=>"000100100",
  2813=>"001010101",
  2814=>"110001110",
  2815=>"001011111",
  2816=>"101111101",
  2817=>"010000110",
  2818=>"010111000",
  2819=>"011100000",
  2820=>"101101010",
  2821=>"000100110",
  2822=>"110011110",
  2823=>"000111110",
  2824=>"011111001",
  2825=>"001000100",
  2826=>"001000100",
  2827=>"011001010",
  2828=>"101000010",
  2829=>"001011010",
  2830=>"000010010",
  2831=>"100000011",
  2832=>"010111011",
  2833=>"001100111",
  2834=>"111011010",
  2835=>"001011000",
  2836=>"110100111",
  2837=>"111011110",
  2838=>"110100101",
  2839=>"010110000",
  2840=>"000011100",
  2841=>"000111110",
  2842=>"111000010",
  2843=>"111111010",
  2844=>"111001011",
  2845=>"011100000",
  2846=>"111101000",
  2847=>"100001000",
  2848=>"111000100",
  2849=>"111101111",
  2850=>"110011000",
  2851=>"001000100",
  2852=>"000101101",
  2853=>"011000000",
  2854=>"110101100",
  2855=>"000101100",
  2856=>"010001001",
  2857=>"110000100",
  2858=>"110110001",
  2859=>"000010010",
  2860=>"110110011",
  2861=>"001001100",
  2862=>"111001100",
  2863=>"110101000",
  2864=>"000001010",
  2865=>"100010100",
  2866=>"100100101",
  2867=>"101111110",
  2868=>"111010111",
  2869=>"100001111",
  2870=>"111010000",
  2871=>"011001001",
  2872=>"010011111",
  2873=>"001101111",
  2874=>"010010000",
  2875=>"111000101",
  2876=>"011011111",
  2877=>"000010010",
  2878=>"010010100",
  2879=>"011001100",
  2880=>"100011111",
  2881=>"010010110",
  2882=>"110010101",
  2883=>"001110101",
  2884=>"110000100",
  2885=>"001010000",
  2886=>"110101010",
  2887=>"110100010",
  2888=>"100100000",
  2889=>"110110000",
  2890=>"110011011",
  2891=>"011001101",
  2892=>"010000000",
  2893=>"010110001",
  2894=>"111110001",
  2895=>"110101101",
  2896=>"011010111",
  2897=>"000101111",
  2898=>"000010000",
  2899=>"111110000",
  2900=>"010100100",
  2901=>"100110110",
  2902=>"011010100",
  2903=>"000010100",
  2904=>"110011011",
  2905=>"101100111",
  2906=>"110011000",
  2907=>"100100000",
  2908=>"010101000",
  2909=>"011010111",
  2910=>"001010111",
  2911=>"001001111",
  2912=>"001001111",
  2913=>"111111101",
  2914=>"100001001",
  2915=>"110100100",
  2916=>"111001110",
  2917=>"010100010",
  2918=>"111100110",
  2919=>"011001000",
  2920=>"110111110",
  2921=>"010110000",
  2922=>"010101110",
  2923=>"100101011",
  2924=>"110000011",
  2925=>"011111000",
  2926=>"000011010",
  2927=>"010110010",
  2928=>"010110100",
  2929=>"011000000",
  2930=>"111001101",
  2931=>"000001100",
  2932=>"100010000",
  2933=>"011011001",
  2934=>"000000110",
  2935=>"101101111",
  2936=>"111011100",
  2937=>"110101101",
  2938=>"001010100",
  2939=>"101000000",
  2940=>"101010110",
  2941=>"000100010",
  2942=>"010111001",
  2943=>"111011111",
  2944=>"100100001",
  2945=>"101111000",
  2946=>"000010011",
  2947=>"110101100",
  2948=>"010011111",
  2949=>"110100110",
  2950=>"111001000",
  2951=>"010011110",
  2952=>"111100101",
  2953=>"000001101",
  2954=>"110111001",
  2955=>"101110101",
  2956=>"100111101",
  2957=>"000001010",
  2958=>"100101011",
  2959=>"001000111",
  2960=>"110110100",
  2961=>"001101011",
  2962=>"000111110",
  2963=>"101001010",
  2964=>"110011111",
  2965=>"011101000",
  2966=>"001010011",
  2967=>"100001011",
  2968=>"100110011",
  2969=>"011101101",
  2970=>"001000100",
  2971=>"111010011",
  2972=>"101000001",
  2973=>"011110101",
  2974=>"011101100",
  2975=>"101101000",
  2976=>"100011001",
  2977=>"101001011",
  2978=>"001100000",
  2979=>"011000010",
  2980=>"101111000",
  2981=>"010101110",
  2982=>"010100110",
  2983=>"110000111",
  2984=>"011111011",
  2985=>"000110011",
  2986=>"000111110",
  2987=>"010100100",
  2988=>"110111101",
  2989=>"000100000",
  2990=>"010001010",
  2991=>"010100111",
  2992=>"010011111",
  2993=>"101111101",
  2994=>"101001101",
  2995=>"101110110",
  2996=>"001110111",
  2997=>"110110111",
  2998=>"000010111",
  2999=>"000010000",
  3000=>"000001010",
  3001=>"101010011",
  3002=>"111010101",
  3003=>"000011000",
  3004=>"000011000",
  3005=>"001001111",
  3006=>"001100110",
  3007=>"100000010",
  3008=>"100110110",
  3009=>"111011010",
  3010=>"001111110",
  3011=>"101100001",
  3012=>"111101110",
  3013=>"111100110",
  3014=>"110111111",
  3015=>"101011100",
  3016=>"011101111",
  3017=>"010001011",
  3018=>"100011101",
  3019=>"110111010",
  3020=>"100001111",
  3021=>"111001111",
  3022=>"011100000",
  3023=>"111000010",
  3024=>"111101000",
  3025=>"100101000",
  3026=>"000011000",
  3027=>"100101110",
  3028=>"100101001",
  3029=>"011001101",
  3030=>"111100000",
  3031=>"100110110",
  3032=>"011111111",
  3033=>"110001000",
  3034=>"000111110",
  3035=>"011110011",
  3036=>"001100111",
  3037=>"101101011",
  3038=>"111110001",
  3039=>"111010000",
  3040=>"001111100",
  3041=>"001011110",
  3042=>"010011101",
  3043=>"110010100",
  3044=>"111001001",
  3045=>"000100011",
  3046=>"001100100",
  3047=>"000000101",
  3048=>"100010110",
  3049=>"011110101",
  3050=>"000000110",
  3051=>"010110100",
  3052=>"011001001",
  3053=>"111000011",
  3054=>"111111111",
  3055=>"100010000",
  3056=>"110000111",
  3057=>"100111001",
  3058=>"100101111",
  3059=>"111101001",
  3060=>"001001111",
  3061=>"011000101",
  3062=>"000000000",
  3063=>"011000000",
  3064=>"111011010",
  3065=>"110011000",
  3066=>"101010000",
  3067=>"011111010",
  3068=>"110101001",
  3069=>"011001011",
  3070=>"011110000",
  3071=>"100101100",
  3072=>"000000011",
  3073=>"110000010",
  3074=>"000111011",
  3075=>"010000101",
  3076=>"111110010",
  3077=>"000001100",
  3078=>"111110111",
  3079=>"110001001",
  3080=>"001101110",
  3081=>"000010011",
  3082=>"001010001",
  3083=>"111111110",
  3084=>"101000111",
  3085=>"101110100",
  3086=>"101000101",
  3087=>"010000010",
  3088=>"100100000",
  3089=>"010001101",
  3090=>"111111010",
  3091=>"100010001",
  3092=>"001100000",
  3093=>"101001100",
  3094=>"000111100",
  3095=>"011010010",
  3096=>"111000011",
  3097=>"111000011",
  3098=>"110101110",
  3099=>"101110100",
  3100=>"111001111",
  3101=>"111101100",
  3102=>"111100000",
  3103=>"110101110",
  3104=>"010011010",
  3105=>"100110101",
  3106=>"111000001",
  3107=>"101110101",
  3108=>"100110010",
  3109=>"110000001",
  3110=>"010000001",
  3111=>"001100001",
  3112=>"000010100",
  3113=>"001111101",
  3114=>"010011011",
  3115=>"010011100",
  3116=>"100001001",
  3117=>"100101000",
  3118=>"011110010",
  3119=>"100111001",
  3120=>"001101000",
  3121=>"101111110",
  3122=>"110110010",
  3123=>"110011011",
  3124=>"110101001",
  3125=>"000111111",
  3126=>"111000110",
  3127=>"001001100",
  3128=>"101101001",
  3129=>"010111010",
  3130=>"111100111",
  3131=>"001100110",
  3132=>"000100000",
  3133=>"000000010",
  3134=>"011001001",
  3135=>"101110110",
  3136=>"110110000",
  3137=>"100010010",
  3138=>"000011011",
  3139=>"000111011",
  3140=>"011100101",
  3141=>"111010001",
  3142=>"101011101",
  3143=>"111011000",
  3144=>"000101101",
  3145=>"110111111",
  3146=>"010010001",
  3147=>"100001111",
  3148=>"000001101",
  3149=>"111001100",
  3150=>"100001101",
  3151=>"111100110",
  3152=>"001110110",
  3153=>"001000010",
  3154=>"111100111",
  3155=>"101001000",
  3156=>"001101000",
  3157=>"010010001",
  3158=>"101101110",
  3159=>"011011010",
  3160=>"110110101",
  3161=>"000001111",
  3162=>"010100110",
  3163=>"000010011",
  3164=>"100000111",
  3165=>"100101001",
  3166=>"011110100",
  3167=>"001101111",
  3168=>"010100111",
  3169=>"111011000",
  3170=>"000001000",
  3171=>"011100000",
  3172=>"001110100",
  3173=>"111001110",
  3174=>"010100100",
  3175=>"100000110",
  3176=>"000100010",
  3177=>"011101110",
  3178=>"100001100",
  3179=>"001100000",
  3180=>"111000111",
  3181=>"110111011",
  3182=>"111001000",
  3183=>"111101101",
  3184=>"001001110",
  3185=>"010110100",
  3186=>"011111110",
  3187=>"100101100",
  3188=>"110010010",
  3189=>"000010001",
  3190=>"110110010",
  3191=>"111000001",
  3192=>"011001100",
  3193=>"111011000",
  3194=>"001101101",
  3195=>"100101010",
  3196=>"011000011",
  3197=>"101010010",
  3198=>"100001010",
  3199=>"001001111",
  3200=>"101101011",
  3201=>"110010001",
  3202=>"000011010",
  3203=>"001100000",
  3204=>"001111000",
  3205=>"110001100",
  3206=>"111100011",
  3207=>"011110111",
  3208=>"010000000",
  3209=>"001010100",
  3210=>"100010010",
  3211=>"101111111",
  3212=>"011111000",
  3213=>"001001111",
  3214=>"010101111",
  3215=>"100000011",
  3216=>"110011001",
  3217=>"100111010",
  3218=>"000001111",
  3219=>"100100110",
  3220=>"110010011",
  3221=>"011101100",
  3222=>"010001000",
  3223=>"111101111",
  3224=>"010101011",
  3225=>"000011101",
  3226=>"001101111",
  3227=>"000111101",
  3228=>"110011011",
  3229=>"010111011",
  3230=>"100101000",
  3231=>"010001100",
  3232=>"111110110",
  3233=>"011101000",
  3234=>"100110001",
  3235=>"111100110",
  3236=>"111010111",
  3237=>"110111010",
  3238=>"010100100",
  3239=>"010011010",
  3240=>"111011000",
  3241=>"111010111",
  3242=>"101001011",
  3243=>"011000010",
  3244=>"001000000",
  3245=>"011000011",
  3246=>"100000100",
  3247=>"001000110",
  3248=>"011001010",
  3249=>"000100010",
  3250=>"011011000",
  3251=>"011000001",
  3252=>"101010011",
  3253=>"010000010",
  3254=>"010000000",
  3255=>"100001001",
  3256=>"000001110",
  3257=>"101101011",
  3258=>"101110000",
  3259=>"000110111",
  3260=>"111101100",
  3261=>"010000010",
  3262=>"000001101",
  3263=>"010111010",
  3264=>"001000000",
  3265=>"101010110",
  3266=>"001010110",
  3267=>"101101010",
  3268=>"001010011",
  3269=>"011100100",
  3270=>"111001110",
  3271=>"101011111",
  3272=>"100011101",
  3273=>"010011111",
  3274=>"111111100",
  3275=>"011110001",
  3276=>"001001010",
  3277=>"100100001",
  3278=>"011111111",
  3279=>"110010011",
  3280=>"101010000",
  3281=>"000001001",
  3282=>"100010101",
  3283=>"001001101",
  3284=>"100000001",
  3285=>"011010110",
  3286=>"110100110",
  3287=>"101000000",
  3288=>"100111010",
  3289=>"110110100",
  3290=>"001100001",
  3291=>"110000110",
  3292=>"000111001",
  3293=>"001101101",
  3294=>"000100001",
  3295=>"111001000",
  3296=>"000000001",
  3297=>"111010011",
  3298=>"000111100",
  3299=>"000000111",
  3300=>"010010101",
  3301=>"000011011",
  3302=>"001000011",
  3303=>"100111110",
  3304=>"111110011",
  3305=>"001101101",
  3306=>"110000111",
  3307=>"111010101",
  3308=>"111111011",
  3309=>"110101010",
  3310=>"001101100",
  3311=>"101010101",
  3312=>"110111111",
  3313=>"110100010",
  3314=>"010110010",
  3315=>"001010001",
  3316=>"001111111",
  3317=>"001010001",
  3318=>"100110010",
  3319=>"111100110",
  3320=>"011010101",
  3321=>"100110110",
  3322=>"001001011",
  3323=>"011010010",
  3324=>"010001100",
  3325=>"000000010",
  3326=>"100111001",
  3327=>"011000011",
  3328=>"100000000",
  3329=>"000100010",
  3330=>"010101101",
  3331=>"110000110",
  3332=>"101110110",
  3333=>"000001001",
  3334=>"010011000",
  3335=>"100010100",
  3336=>"100001111",
  3337=>"000111011",
  3338=>"101110011",
  3339=>"110110011",
  3340=>"101001100",
  3341=>"001010111",
  3342=>"011001010",
  3343=>"100110000",
  3344=>"010000100",
  3345=>"101001001",
  3346=>"111111100",
  3347=>"111010000",
  3348=>"101101110",
  3349=>"010111000",
  3350=>"000010111",
  3351=>"001110011",
  3352=>"000010100",
  3353=>"111010100",
  3354=>"100100100",
  3355=>"000101110",
  3356=>"111101100",
  3357=>"011010001",
  3358=>"111010001",
  3359=>"110011010",
  3360=>"000010011",
  3361=>"101010010",
  3362=>"000100010",
  3363=>"010001010",
  3364=>"000111110",
  3365=>"000101011",
  3366=>"000100101",
  3367=>"111111010",
  3368=>"110100000",
  3369=>"100111011",
  3370=>"001111010",
  3371=>"111001101",
  3372=>"101001110",
  3373=>"010111110",
  3374=>"111111111",
  3375=>"000100000",
  3376=>"110101010",
  3377=>"111001010",
  3378=>"110111101",
  3379=>"011001011",
  3380=>"001011000",
  3381=>"001110010",
  3382=>"100001001",
  3383=>"001101011",
  3384=>"001001001",
  3385=>"101001011",
  3386=>"100101011",
  3387=>"010110001",
  3388=>"001000100",
  3389=>"001001110",
  3390=>"001001101",
  3391=>"011001110",
  3392=>"001111000",
  3393=>"101110100",
  3394=>"010100100",
  3395=>"001001011",
  3396=>"000010010",
  3397=>"000100001",
  3398=>"011001010",
  3399=>"000101011",
  3400=>"010000111",
  3401=>"000000010",
  3402=>"010100101",
  3403=>"100000010",
  3404=>"110110111",
  3405=>"000110100",
  3406=>"000110000",
  3407=>"010101101",
  3408=>"101000001",
  3409=>"000000000",
  3410=>"010010011",
  3411=>"101110111",
  3412=>"001101010",
  3413=>"010000110",
  3414=>"110011000",
  3415=>"101000100",
  3416=>"100100010",
  3417=>"110111000",
  3418=>"101011111",
  3419=>"001101110",
  3420=>"101011000",
  3421=>"000001111",
  3422=>"000001111",
  3423=>"101101101",
  3424=>"011110100",
  3425=>"001111111",
  3426=>"111000110",
  3427=>"111011001",
  3428=>"011101101",
  3429=>"010001111",
  3430=>"101000111",
  3431=>"100110110",
  3432=>"000110010",
  3433=>"110001011",
  3434=>"111000001",
  3435=>"110101000",
  3436=>"111000000",
  3437=>"101101111",
  3438=>"001010011",
  3439=>"101110011",
  3440=>"011100110",
  3441=>"011101110",
  3442=>"010110100",
  3443=>"000111000",
  3444=>"110011011",
  3445=>"100001101",
  3446=>"001000011",
  3447=>"001111110",
  3448=>"001000110",
  3449=>"001101101",
  3450=>"111100011",
  3451=>"011100100",
  3452=>"111010111",
  3453=>"011100100",
  3454=>"110111111",
  3455=>"100111111",
  3456=>"000010001",
  3457=>"100011111",
  3458=>"010000100",
  3459=>"000101010",
  3460=>"101000011",
  3461=>"000110101",
  3462=>"010010000",
  3463=>"000001100",
  3464=>"111110010",
  3465=>"100011001",
  3466=>"110011011",
  3467=>"010011110",
  3468=>"111010011",
  3469=>"001000001",
  3470=>"111011010",
  3471=>"010110010",
  3472=>"101010010",
  3473=>"000010010",
  3474=>"110000110",
  3475=>"000010010",
  3476=>"100110000",
  3477=>"011011011",
  3478=>"000111100",
  3479=>"000111010",
  3480=>"111001110",
  3481=>"110100010",
  3482=>"011101100",
  3483=>"101111111",
  3484=>"010110100",
  3485=>"100100011",
  3486=>"111000001",
  3487=>"111101010",
  3488=>"010100000",
  3489=>"100011110",
  3490=>"110110100",
  3491=>"000110110",
  3492=>"001010110",
  3493=>"111111011",
  3494=>"001110110",
  3495=>"010000010",
  3496=>"010100011",
  3497=>"101001111",
  3498=>"010010101",
  3499=>"111110100",
  3500=>"000000101",
  3501=>"110010100",
  3502=>"101110001",
  3503=>"000001101",
  3504=>"011101000",
  3505=>"101011010",
  3506=>"010010011",
  3507=>"111111110",
  3508=>"011111100",
  3509=>"101110010",
  3510=>"000010111",
  3511=>"100010111",
  3512=>"110111010",
  3513=>"111000100",
  3514=>"101110110",
  3515=>"001100011",
  3516=>"101100110",
  3517=>"111111111",
  3518=>"100101000",
  3519=>"111100010",
  3520=>"001010010",
  3521=>"101110111",
  3522=>"100101111",
  3523=>"110111110",
  3524=>"011000001",
  3525=>"001010110",
  3526=>"000011111",
  3527=>"000100111",
  3528=>"110110111",
  3529=>"100111100",
  3530=>"111110011",
  3531=>"000010010",
  3532=>"011000111",
  3533=>"100000011",
  3534=>"010110110",
  3535=>"100000011",
  3536=>"001000000",
  3537=>"001111001",
  3538=>"101101010",
  3539=>"111011001",
  3540=>"001110000",
  3541=>"001100000",
  3542=>"101111001",
  3543=>"001111100",
  3544=>"111111001",
  3545=>"001101001",
  3546=>"001110111",
  3547=>"111100111",
  3548=>"010001110",
  3549=>"100001001",
  3550=>"111000001",
  3551=>"000000100",
  3552=>"100000111",
  3553=>"010001100",
  3554=>"010101011",
  3555=>"110101111",
  3556=>"000111010",
  3557=>"111001001",
  3558=>"101111111",
  3559=>"000111110",
  3560=>"110010110",
  3561=>"000011111",
  3562=>"000011111",
  3563=>"110111010",
  3564=>"010000000",
  3565=>"001110000",
  3566=>"101111111",
  3567=>"000110110",
  3568=>"111111100",
  3569=>"110110100",
  3570=>"011100000",
  3571=>"000110011",
  3572=>"110000011",
  3573=>"110110011",
  3574=>"001111011",
  3575=>"111100100",
  3576=>"010101101",
  3577=>"111010111",
  3578=>"010101010",
  3579=>"011110011",
  3580=>"111110111",
  3581=>"011000001",
  3582=>"111001110",
  3583=>"010011000",
  3584=>"011000000",
  3585=>"010011011",
  3586=>"101101101",
  3587=>"001011101",
  3588=>"000011100",
  3589=>"101001100",
  3590=>"010111111",
  3591=>"010010100",
  3592=>"010000011",
  3593=>"001001101",
  3594=>"010001001",
  3595=>"111111101",
  3596=>"010011011",
  3597=>"111010101",
  3598=>"000011111",
  3599=>"000010010",
  3600=>"111010110",
  3601=>"010111000",
  3602=>"101001001",
  3603=>"011000001",
  3604=>"011011111",
  3605=>"010010101",
  3606=>"110011110",
  3607=>"111000110",
  3608=>"110111100",
  3609=>"001011100",
  3610=>"010010010",
  3611=>"110001011",
  3612=>"101001001",
  3613=>"100011111",
  3614=>"111010111",
  3615=>"111010001",
  3616=>"110011110",
  3617=>"101101001",
  3618=>"010000100",
  3619=>"001100000",
  3620=>"110010000",
  3621=>"001110011",
  3622=>"110111011",
  3623=>"100011000",
  3624=>"001101110",
  3625=>"100101101",
  3626=>"011111111",
  3627=>"111001000",
  3628=>"110010001",
  3629=>"111011010",
  3630=>"111000110",
  3631=>"111010011",
  3632=>"010011001",
  3633=>"110100011",
  3634=>"100001110",
  3635=>"010000000",
  3636=>"010100010",
  3637=>"000111100",
  3638=>"101001100",
  3639=>"111110001",
  3640=>"000111100",
  3641=>"111011011",
  3642=>"100001101",
  3643=>"001100101",
  3644=>"110111111",
  3645=>"010001110",
  3646=>"000000001",
  3647=>"010000101",
  3648=>"010111001",
  3649=>"001100101",
  3650=>"001011110",
  3651=>"100011111",
  3652=>"010111111",
  3653=>"111101110",
  3654=>"000000110",
  3655=>"101001000",
  3656=>"011111010",
  3657=>"001011111",
  3658=>"111111100",
  3659=>"010000010",
  3660=>"001001110",
  3661=>"100001101",
  3662=>"011001111",
  3663=>"001010111",
  3664=>"110011011",
  3665=>"111001011",
  3666=>"111111110",
  3667=>"111000111",
  3668=>"011010011",
  3669=>"101100111",
  3670=>"111100111",
  3671=>"010010011",
  3672=>"101110010",
  3673=>"010011110",
  3674=>"101100100",
  3675=>"001110111",
  3676=>"010001011",
  3677=>"101101110",
  3678=>"011011011",
  3679=>"000100000",
  3680=>"011101101",
  3681=>"000001100",
  3682=>"111010010",
  3683=>"011101000",
  3684=>"010001110",
  3685=>"111100001",
  3686=>"010100111",
  3687=>"001000100",
  3688=>"000101000",
  3689=>"001010110",
  3690=>"100110011",
  3691=>"100000011",
  3692=>"011000000",
  3693=>"111110101",
  3694=>"010101001",
  3695=>"001001111",
  3696=>"010000010",
  3697=>"010111011",
  3698=>"000011111",
  3699=>"000010100",
  3700=>"010011011",
  3701=>"001001010",
  3702=>"111100000",
  3703=>"001000000",
  3704=>"110100001",
  3705=>"010010010",
  3706=>"101001000",
  3707=>"111001011",
  3708=>"110111000",
  3709=>"011000111",
  3710=>"011110011",
  3711=>"110010000",
  3712=>"000100011",
  3713=>"000100111",
  3714=>"100000111",
  3715=>"000000101",
  3716=>"001110010",
  3717=>"000100110",
  3718=>"011110101",
  3719=>"011011100",
  3720=>"101110101",
  3721=>"011010110",
  3722=>"111101000",
  3723=>"100111110",
  3724=>"110000110",
  3725=>"000011101",
  3726=>"110010010",
  3727=>"100000110",
  3728=>"111010000",
  3729=>"000000001",
  3730=>"111001110",
  3731=>"100001011",
  3732=>"011010000",
  3733=>"110101010",
  3734=>"001000001",
  3735=>"001101111",
  3736=>"101110010",
  3737=>"110000101",
  3738=>"001000001",
  3739=>"010100000",
  3740=>"011100111",
  3741=>"111011000",
  3742=>"000110111",
  3743=>"010001100",
  3744=>"100011010",
  3745=>"110111011",
  3746=>"110010010",
  3747=>"011011110",
  3748=>"101111011",
  3749=>"001111111",
  3750=>"001011010",
  3751=>"110000100",
  3752=>"100010101",
  3753=>"001000010",
  3754=>"111001010",
  3755=>"110101100",
  3756=>"011000111",
  3757=>"010010011",
  3758=>"111001000",
  3759=>"001110111",
  3760=>"100011000",
  3761=>"101101101",
  3762=>"110110001",
  3763=>"110011111",
  3764=>"001101000",
  3765=>"011110011",
  3766=>"110100010",
  3767=>"001100000",
  3768=>"001110010",
  3769=>"000000101",
  3770=>"000000011",
  3771=>"000011000",
  3772=>"011011000",
  3773=>"010000001",
  3774=>"111010001",
  3775=>"000001000",
  3776=>"111010010",
  3777=>"101111001",
  3778=>"001111100",
  3779=>"000101001",
  3780=>"011101010",
  3781=>"000101100",
  3782=>"000101101",
  3783=>"100011111",
  3784=>"111101000",
  3785=>"110000011",
  3786=>"011000000",
  3787=>"100100101",
  3788=>"001100101",
  3789=>"110101100",
  3790=>"100100111",
  3791=>"101110010",
  3792=>"011010111",
  3793=>"111111011",
  3794=>"001100011",
  3795=>"110110010",
  3796=>"100010100",
  3797=>"100000000",
  3798=>"000000001",
  3799=>"000101000",
  3800=>"101011000",
  3801=>"101000110",
  3802=>"010001101",
  3803=>"000100011",
  3804=>"011100001",
  3805=>"010101000",
  3806=>"101110100",
  3807=>"001000011",
  3808=>"011101110",
  3809=>"111001001",
  3810=>"001011011",
  3811=>"011110111",
  3812=>"110110001",
  3813=>"100000111",
  3814=>"011111011",
  3815=>"111110100",
  3816=>"010100100",
  3817=>"000101001",
  3818=>"011010101",
  3819=>"000001010",
  3820=>"110010111",
  3821=>"001101010",
  3822=>"100100101",
  3823=>"111101101",
  3824=>"110011000",
  3825=>"101100010",
  3826=>"111100010",
  3827=>"111001100",
  3828=>"000011111",
  3829=>"100010000",
  3830=>"011100010",
  3831=>"100000000",
  3832=>"001001111",
  3833=>"100111100",
  3834=>"010000001",
  3835=>"010000001",
  3836=>"110111100",
  3837=>"001000111",
  3838=>"110010000",
  3839=>"000000011",
  3840=>"111001010",
  3841=>"001010000",
  3842=>"110101010",
  3843=>"011110101",
  3844=>"100111000",
  3845=>"101100010",
  3846=>"001011010",
  3847=>"111111101",
  3848=>"011100000",
  3849=>"110111110",
  3850=>"011100011",
  3851=>"010011111",
  3852=>"001011110",
  3853=>"100101000",
  3854=>"000011011",
  3855=>"011111100",
  3856=>"011111100",
  3857=>"100011000",
  3858=>"010011000",
  3859=>"110000110",
  3860=>"100000111",
  3861=>"000100001",
  3862=>"110111100",
  3863=>"001010001",
  3864=>"010000011",
  3865=>"000010001",
  3866=>"000000110",
  3867=>"110011101",
  3868=>"101101101",
  3869=>"110110111",
  3870=>"010100100",
  3871=>"110000001",
  3872=>"010100001",
  3873=>"111101101",
  3874=>"101011100",
  3875=>"000000111",
  3876=>"111101010",
  3877=>"110001010",
  3878=>"101010001",
  3879=>"010011101",
  3880=>"000011110",
  3881=>"111010110",
  3882=>"000010101",
  3883=>"011000101",
  3884=>"101011010",
  3885=>"110111010",
  3886=>"000010001",
  3887=>"001011101",
  3888=>"000111100",
  3889=>"011000101",
  3890=>"101110001",
  3891=>"010100111",
  3892=>"000011011",
  3893=>"010011001",
  3894=>"001010000",
  3895=>"000100010",
  3896=>"100101100",
  3897=>"011010110",
  3898=>"011111010",
  3899=>"110110111",
  3900=>"001110000",
  3901=>"011000100",
  3902=>"101111100",
  3903=>"000110100",
  3904=>"100010101",
  3905=>"011000000",
  3906=>"001101111",
  3907=>"100001001",
  3908=>"011001000",
  3909=>"111011101",
  3910=>"010011010",
  3911=>"000000110",
  3912=>"100100001",
  3913=>"110101111",
  3914=>"001111110",
  3915=>"111000100",
  3916=>"100001000",
  3917=>"011010001",
  3918=>"001000101",
  3919=>"111010010",
  3920=>"011011000",
  3921=>"101001101",
  3922=>"000101000",
  3923=>"011011111",
  3924=>"101110011",
  3925=>"011110100",
  3926=>"110000111",
  3927=>"100010111",
  3928=>"011010010",
  3929=>"010100011",
  3930=>"000011000",
  3931=>"101101011",
  3932=>"100100101",
  3933=>"000001001",
  3934=>"010000111",
  3935=>"010010101",
  3936=>"001100001",
  3937=>"010000110",
  3938=>"100100011",
  3939=>"110011011",
  3940=>"110001011",
  3941=>"001101110",
  3942=>"101110011",
  3943=>"100110100",
  3944=>"110111010",
  3945=>"111000101",
  3946=>"001011111",
  3947=>"101010100",
  3948=>"001000001",
  3949=>"001111011",
  3950=>"000110110",
  3951=>"101110111",
  3952=>"101000001",
  3953=>"001001001",
  3954=>"111010101",
  3955=>"111011000",
  3956=>"100000000",
  3957=>"111010111",
  3958=>"110010011",
  3959=>"101111110",
  3960=>"111100100",
  3961=>"010011110",
  3962=>"100011010",
  3963=>"101011101",
  3964=>"000001010",
  3965=>"011000100",
  3966=>"011111110",
  3967=>"001001010",
  3968=>"000101011",
  3969=>"100000101",
  3970=>"000010001",
  3971=>"100011111",
  3972=>"000011011",
  3973=>"110111100",
  3974=>"011000110",
  3975=>"001010101",
  3976=>"000000100",
  3977=>"001000011",
  3978=>"110101111",
  3979=>"111111001",
  3980=>"000110000",
  3981=>"111100101",
  3982=>"001001110",
  3983=>"110101101",
  3984=>"010101110",
  3985=>"010111100",
  3986=>"000001111",
  3987=>"010111010",
  3988=>"000001101",
  3989=>"111110001",
  3990=>"000010110",
  3991=>"000001110",
  3992=>"000001101",
  3993=>"001100011",
  3994=>"111001000",
  3995=>"011101100",
  3996=>"100010001",
  3997=>"010001101",
  3998=>"000111000",
  3999=>"010001010",
  4000=>"011110001",
  4001=>"101010101",
  4002=>"011010111",
  4003=>"110110110",
  4004=>"110101010",
  4005=>"010000111",
  4006=>"001010011",
  4007=>"101101111",
  4008=>"001010000",
  4009=>"011100000",
  4010=>"111100010",
  4011=>"110000110",
  4012=>"110010111",
  4013=>"101111101",
  4014=>"111001001",
  4015=>"111010110",
  4016=>"001101100",
  4017=>"010111110",
  4018=>"000000101",
  4019=>"101010111",
  4020=>"101011000",
  4021=>"101101101",
  4022=>"100111000",
  4023=>"010101001",
  4024=>"110100101",
  4025=>"111101101",
  4026=>"000011110",
  4027=>"001011110",
  4028=>"010101110",
  4029=>"100001000",
  4030=>"110110000",
  4031=>"000001011",
  4032=>"111111010",
  4033=>"100010110",
  4034=>"010111111",
  4035=>"001010110",
  4036=>"010111101",
  4037=>"000010101",
  4038=>"011010101",
  4039=>"101001001",
  4040=>"010000001",
  4041=>"000011111",
  4042=>"101101100",
  4043=>"010000001",
  4044=>"110100100",
  4045=>"001100100",
  4046=>"110100000",
  4047=>"100010000",
  4048=>"010110011",
  4049=>"001101000",
  4050=>"000001111",
  4051=>"111111001",
  4052=>"100111100",
  4053=>"000011101",
  4054=>"001000100",
  4055=>"111001101",
  4056=>"111101010",
  4057=>"110101001",
  4058=>"100011101",
  4059=>"110101101",
  4060=>"000000110",
  4061=>"100111111",
  4062=>"011001010",
  4063=>"111111100",
  4064=>"101010001",
  4065=>"011101101",
  4066=>"001010010",
  4067=>"000010010",
  4068=>"000010000",
  4069=>"100000110",
  4070=>"010000001",
  4071=>"100111010",
  4072=>"111001111",
  4073=>"010110110",
  4074=>"000001100",
  4075=>"001101111",
  4076=>"101011011",
  4077=>"000110000",
  4078=>"100010110",
  4079=>"101100001",
  4080=>"010101110",
  4081=>"010111010",
  4082=>"011100110",
  4083=>"110010100",
  4084=>"000100111",
  4085=>"111100111",
  4086=>"111110010",
  4087=>"111111000",
  4088=>"000010010",
  4089=>"001001110",
  4090=>"010101011",
  4091=>"010000110",
  4092=>"110101101",
  4093=>"001100111",
  4094=>"110100111",
  4095=>"000100011",
  4096=>"110101011",
  4097=>"101001011",
  4098=>"110011111",
  4099=>"101100110",
  4100=>"010101011",
  4101=>"100110011",
  4102=>"101001011",
  4103=>"011110111",
  4104=>"101011000",
  4105=>"000101010",
  4106=>"010001100",
  4107=>"000010010",
  4108=>"101010100",
  4109=>"110110000",
  4110=>"101000011",
  4111=>"110101101",
  4112=>"111111011",
  4113=>"011111100",
  4114=>"110101000",
  4115=>"011111100",
  4116=>"110111101",
  4117=>"101000001",
  4118=>"101110001",
  4119=>"110110111",
  4120=>"100010111",
  4121=>"001110010",
  4122=>"111100100",
  4123=>"001000000",
  4124=>"000100100",
  4125=>"111001010",
  4126=>"010001000",
  4127=>"001010011",
  4128=>"101001011",
  4129=>"111111001",
  4130=>"101010010",
  4131=>"001001000",
  4132=>"101100111",
  4133=>"000010000",
  4134=>"101110011",
  4135=>"011010000",
  4136=>"010000001",
  4137=>"111101110",
  4138=>"000110100",
  4139=>"101101011",
  4140=>"000111111",
  4141=>"001011010",
  4142=>"000001101",
  4143=>"001101100",
  4144=>"000011101",
  4145=>"110001101",
  4146=>"011000110",
  4147=>"011101101",
  4148=>"101010111",
  4149=>"001101101",
  4150=>"111000011",
  4151=>"111100001",
  4152=>"010111110",
  4153=>"110110011",
  4154=>"010011000",
  4155=>"000110010",
  4156=>"001000011",
  4157=>"111000110",
  4158=>"111111000",
  4159=>"110111011",
  4160=>"100111000",
  4161=>"101000101",
  4162=>"010001010",
  4163=>"100000010",
  4164=>"010110010",
  4165=>"101110111",
  4166=>"101011001",
  4167=>"010000111",
  4168=>"000001011",
  4169=>"111111001",
  4170=>"101010100",
  4171=>"100100000",
  4172=>"000101101",
  4173=>"010101010",
  4174=>"100000001",
  4175=>"101010001",
  4176=>"010001011",
  4177=>"101001100",
  4178=>"010001000",
  4179=>"011111011",
  4180=>"110011001",
  4181=>"111000001",
  4182=>"011111010",
  4183=>"111001101",
  4184=>"001011101",
  4185=>"111111111",
  4186=>"000110001",
  4187=>"011101001",
  4188=>"001000001",
  4189=>"001101010",
  4190=>"001000011",
  4191=>"011111110",
  4192=>"010110110",
  4193=>"111011110",
  4194=>"001110111",
  4195=>"001000101",
  4196=>"110000011",
  4197=>"011000011",
  4198=>"010000011",
  4199=>"101101100",
  4200=>"001001001",
  4201=>"001010000",
  4202=>"001110100",
  4203=>"000001011",
  4204=>"010100000",
  4205=>"000110010",
  4206=>"111111000",
  4207=>"110111100",
  4208=>"010001101",
  4209=>"010101011",
  4210=>"000001011",
  4211=>"010000111",
  4212=>"101110111",
  4213=>"010110110",
  4214=>"101100111",
  4215=>"010001100",
  4216=>"011100011",
  4217=>"110011110",
  4218=>"010101100",
  4219=>"001110000",
  4220=>"000100011",
  4221=>"000000000",
  4222=>"010101011",
  4223=>"100101001",
  4224=>"010111010",
  4225=>"111110101",
  4226=>"000011001",
  4227=>"110111011",
  4228=>"101101010",
  4229=>"011011110",
  4230=>"011011011",
  4231=>"010100001",
  4232=>"110000101",
  4233=>"101001110",
  4234=>"010101010",
  4235=>"111111110",
  4236=>"110110011",
  4237=>"100010011",
  4238=>"100001000",
  4239=>"000000001",
  4240=>"110111111",
  4241=>"001101101",
  4242=>"010011110",
  4243=>"100011100",
  4244=>"100000110",
  4245=>"100001111",
  4246=>"000100000",
  4247=>"001111110",
  4248=>"110000111",
  4249=>"011011010",
  4250=>"111111110",
  4251=>"100100100",
  4252=>"010101001",
  4253=>"100010110",
  4254=>"101000000",
  4255=>"101101001",
  4256=>"110101011",
  4257=>"000001000",
  4258=>"110110010",
  4259=>"111010101",
  4260=>"000111001",
  4261=>"010010010",
  4262=>"010100111",
  4263=>"100000100",
  4264=>"010011111",
  4265=>"100010111",
  4266=>"100100111",
  4267=>"010001001",
  4268=>"011111101",
  4269=>"010100000",
  4270=>"110001101",
  4271=>"110011101",
  4272=>"101110111",
  4273=>"010111101",
  4274=>"110001111",
  4275=>"110010111",
  4276=>"010010001",
  4277=>"001011110",
  4278=>"000111000",
  4279=>"100101010",
  4280=>"010001101",
  4281=>"011100101",
  4282=>"100110000",
  4283=>"100010110",
  4284=>"111001001",
  4285=>"001010010",
  4286=>"011110001",
  4287=>"011100111",
  4288=>"010110101",
  4289=>"100010100",
  4290=>"110110000",
  4291=>"110111111",
  4292=>"001001101",
  4293=>"100111010",
  4294=>"101001011",
  4295=>"110100001",
  4296=>"010100100",
  4297=>"001111111",
  4298=>"001101111",
  4299=>"001101100",
  4300=>"010001101",
  4301=>"111010010",
  4302=>"111010000",
  4303=>"000000101",
  4304=>"101110100",
  4305=>"100101100",
  4306=>"100010101",
  4307=>"101011111",
  4308=>"001110100",
  4309=>"001000100",
  4310=>"000100110",
  4311=>"101011001",
  4312=>"001011101",
  4313=>"011000111",
  4314=>"111000000",
  4315=>"000111010",
  4316=>"011110111",
  4317=>"100001001",
  4318=>"001100001",
  4319=>"011111010",
  4320=>"000100100",
  4321=>"010011011",
  4322=>"110001000",
  4323=>"101010000",
  4324=>"101110011",
  4325=>"100010000",
  4326=>"111011011",
  4327=>"001100110",
  4328=>"010000001",
  4329=>"010101010",
  4330=>"001101011",
  4331=>"111100001",
  4332=>"011000011",
  4333=>"100100011",
  4334=>"011001101",
  4335=>"101111110",
  4336=>"110000101",
  4337=>"011100001",
  4338=>"101010001",
  4339=>"000111100",
  4340=>"101001011",
  4341=>"100010001",
  4342=>"000110000",
  4343=>"000111001",
  4344=>"001010110",
  4345=>"110101100",
  4346=>"101001101",
  4347=>"011010011",
  4348=>"001101111",
  4349=>"111110011",
  4350=>"001101111",
  4351=>"111101011",
  4352=>"111110111",
  4353=>"110101111",
  4354=>"011101011",
  4355=>"100100010",
  4356=>"100001111",
  4357=>"001111111",
  4358=>"011101101",
  4359=>"001110100",
  4360=>"110110111",
  4361=>"000001100",
  4362=>"100111111",
  4363=>"000000001",
  4364=>"110000101",
  4365=>"100100001",
  4366=>"010111011",
  4367=>"101011100",
  4368=>"111001000",
  4369=>"110110000",
  4370=>"110000011",
  4371=>"110011000",
  4372=>"111000001",
  4373=>"001110100",
  4374=>"000011001",
  4375=>"001101101",
  4376=>"110100100",
  4377=>"100001011",
  4378=>"111000000",
  4379=>"001001001",
  4380=>"100110010",
  4381=>"100001111",
  4382=>"111001000",
  4383=>"111101101",
  4384=>"000001011",
  4385=>"000000000",
  4386=>"101100011",
  4387=>"101100001",
  4388=>"111110110",
  4389=>"000011110",
  4390=>"010111101",
  4391=>"100101001",
  4392=>"001000101",
  4393=>"001111100",
  4394=>"101000001",
  4395=>"111011101",
  4396=>"110111011",
  4397=>"100010000",
  4398=>"111011111",
  4399=>"111101111",
  4400=>"100011001",
  4401=>"100111110",
  4402=>"110001011",
  4403=>"111111101",
  4404=>"001000000",
  4405=>"011101111",
  4406=>"011111010",
  4407=>"011101100",
  4408=>"100011100",
  4409=>"011010011",
  4410=>"011011111",
  4411=>"100100100",
  4412=>"100011001",
  4413=>"110110100",
  4414=>"010110001",
  4415=>"100101110",
  4416=>"110010101",
  4417=>"011101100",
  4418=>"001110101",
  4419=>"000010101",
  4420=>"100010000",
  4421=>"010100110",
  4422=>"111111000",
  4423=>"001010000",
  4424=>"101101111",
  4425=>"001000100",
  4426=>"001111010",
  4427=>"000110100",
  4428=>"101110001",
  4429=>"110111000",
  4430=>"100000001",
  4431=>"010111000",
  4432=>"100000011",
  4433=>"100000001",
  4434=>"011011100",
  4435=>"010110010",
  4436=>"010011011",
  4437=>"111000100",
  4438=>"001010001",
  4439=>"101000000",
  4440=>"111001000",
  4441=>"001101010",
  4442=>"000111011",
  4443=>"101010001",
  4444=>"100010101",
  4445=>"100110000",
  4446=>"111111101",
  4447=>"101100101",
  4448=>"010011000",
  4449=>"011010010",
  4450=>"000101111",
  4451=>"110100000",
  4452=>"011111000",
  4453=>"000000101",
  4454=>"010110010",
  4455=>"010001111",
  4456=>"011101100",
  4457=>"010100010",
  4458=>"101101111",
  4459=>"101011111",
  4460=>"111010111",
  4461=>"100101110",
  4462=>"111000000",
  4463=>"101100000",
  4464=>"011101000",
  4465=>"111101011",
  4466=>"110111001",
  4467=>"010011011",
  4468=>"010001000",
  4469=>"101001111",
  4470=>"010100110",
  4471=>"110110111",
  4472=>"101100110",
  4473=>"110010000",
  4474=>"101001111",
  4475=>"001111110",
  4476=>"000111110",
  4477=>"101010000",
  4478=>"101100010",
  4479=>"101011101",
  4480=>"101101101",
  4481=>"101000000",
  4482=>"010011010",
  4483=>"101001101",
  4484=>"111010010",
  4485=>"011000110",
  4486=>"010110001",
  4487=>"000011010",
  4488=>"000000010",
  4489=>"100111101",
  4490=>"011011010",
  4491=>"010100111",
  4492=>"100001010",
  4493=>"011100100",
  4494=>"010111001",
  4495=>"100101001",
  4496=>"111001001",
  4497=>"000001111",
  4498=>"100011111",
  4499=>"011011001",
  4500=>"101010101",
  4501=>"110001111",
  4502=>"000100111",
  4503=>"010000101",
  4504=>"011101011",
  4505=>"010111111",
  4506=>"001010011",
  4507=>"011010101",
  4508=>"111000111",
  4509=>"000010111",
  4510=>"001110111",
  4511=>"100110010",
  4512=>"100001110",
  4513=>"000010100",
  4514=>"101100110",
  4515=>"000011001",
  4516=>"000011000",
  4517=>"011110100",
  4518=>"111110100",
  4519=>"011110101",
  4520=>"001111101",
  4521=>"100101100",
  4522=>"010001010",
  4523=>"000011001",
  4524=>"110101001",
  4525=>"100100010",
  4526=>"111010110",
  4527=>"100010110",
  4528=>"010111011",
  4529=>"010110011",
  4530=>"111101001",
  4531=>"011100011",
  4532=>"100110101",
  4533=>"111001010",
  4534=>"000110000",
  4535=>"110110011",
  4536=>"111100101",
  4537=>"010011110",
  4538=>"000111111",
  4539=>"101110000",
  4540=>"001010010",
  4541=>"011011001",
  4542=>"011001010",
  4543=>"011100011",
  4544=>"001101110",
  4545=>"010110101",
  4546=>"011111011",
  4547=>"100111110",
  4548=>"011100010",
  4549=>"010000111",
  4550=>"001001111",
  4551=>"000011110",
  4552=>"110101011",
  4553=>"001010010",
  4554=>"100001111",
  4555=>"000100101",
  4556=>"110110001",
  4557=>"001001100",
  4558=>"000010101",
  4559=>"111000010",
  4560=>"100101001",
  4561=>"010111110",
  4562=>"100110001",
  4563=>"110101110",
  4564=>"111010101",
  4565=>"110100000",
  4566=>"001110000",
  4567=>"000011010",
  4568=>"100011011",
  4569=>"111000000",
  4570=>"010111010",
  4571=>"101011011",
  4572=>"000101111",
  4573=>"100011100",
  4574=>"010010010",
  4575=>"001110010",
  4576=>"111111110",
  4577=>"101011000",
  4578=>"100011000",
  4579=>"010111000",
  4580=>"001000001",
  4581=>"110011010",
  4582=>"011101110",
  4583=>"001100110",
  4584=>"010010011",
  4585=>"100000110",
  4586=>"101110110",
  4587=>"111011010",
  4588=>"101000100",
  4589=>"101110111",
  4590=>"111101101",
  4591=>"000100100",
  4592=>"101110110",
  4593=>"101100001",
  4594=>"011101001",
  4595=>"010010010",
  4596=>"001000010",
  4597=>"010100111",
  4598=>"001011101",
  4599=>"000101011",
  4600=>"111101001",
  4601=>"011101111",
  4602=>"001010010",
  4603=>"101010111",
  4604=>"011101110",
  4605=>"011101001",
  4606=>"101100101",
  4607=>"001111000",
  4608=>"000000110",
  4609=>"100111111",
  4610=>"101111010",
  4611=>"101000110",
  4612=>"100000100",
  4613=>"010111101",
  4614=>"001100111",
  4615=>"010011110",
  4616=>"000100100",
  4617=>"000011010",
  4618=>"010111001",
  4619=>"111000110",
  4620=>"011011101",
  4621=>"001010010",
  4622=>"010110010",
  4623=>"011110010",
  4624=>"000100110",
  4625=>"011110110",
  4626=>"010001011",
  4627=>"100101000",
  4628=>"011100000",
  4629=>"100000010",
  4630=>"000111011",
  4631=>"101001111",
  4632=>"000101101",
  4633=>"011111110",
  4634=>"011010011",
  4635=>"110100010",
  4636=>"001010000",
  4637=>"100010011",
  4638=>"101000010",
  4639=>"110010111",
  4640=>"000110100",
  4641=>"100110100",
  4642=>"010100011",
  4643=>"011011011",
  4644=>"101001101",
  4645=>"111011110",
  4646=>"011101101",
  4647=>"110011111",
  4648=>"100001011",
  4649=>"100110110",
  4650=>"000010101",
  4651=>"001011000",
  4652=>"101000100",
  4653=>"001011101",
  4654=>"100010110",
  4655=>"100101110",
  4656=>"010010110",
  4657=>"100101111",
  4658=>"100110001",
  4659=>"100101001",
  4660=>"100111000",
  4661=>"101111111",
  4662=>"000110110",
  4663=>"111001001",
  4664=>"001110000",
  4665=>"111001111",
  4666=>"110000011",
  4667=>"101101111",
  4668=>"110110100",
  4669=>"010011110",
  4670=>"101001000",
  4671=>"000110000",
  4672=>"010110010",
  4673=>"000100110",
  4674=>"011111010",
  4675=>"100100010",
  4676=>"110110101",
  4677=>"100100100",
  4678=>"001001010",
  4679=>"010111000",
  4680=>"000000100",
  4681=>"111100111",
  4682=>"010100100",
  4683=>"001110001",
  4684=>"011101101",
  4685=>"010100001",
  4686=>"010100000",
  4687=>"000111100",
  4688=>"000000101",
  4689=>"001101110",
  4690=>"010100100",
  4691=>"111000110",
  4692=>"000010000",
  4693=>"100011100",
  4694=>"100001110",
  4695=>"101010001",
  4696=>"101001011",
  4697=>"001000000",
  4698=>"001010110",
  4699=>"010101110",
  4700=>"100000000",
  4701=>"000011010",
  4702=>"001111010",
  4703=>"010100010",
  4704=>"011011000",
  4705=>"100011010",
  4706=>"100001011",
  4707=>"100101010",
  4708=>"111011011",
  4709=>"010000101",
  4710=>"011001011",
  4711=>"010000100",
  4712=>"100011101",
  4713=>"100110010",
  4714=>"110110011",
  4715=>"100101100",
  4716=>"110110101",
  4717=>"111001100",
  4718=>"101100000",
  4719=>"001011100",
  4720=>"011010101",
  4721=>"001000010",
  4722=>"001001111",
  4723=>"001001001",
  4724=>"011110100",
  4725=>"100111010",
  4726=>"111111000",
  4727=>"010010110",
  4728=>"100100111",
  4729=>"001010000",
  4730=>"011000101",
  4731=>"011010001",
  4732=>"011101011",
  4733=>"110101000",
  4734=>"100000011",
  4735=>"110000110",
  4736=>"100011000",
  4737=>"110111101",
  4738=>"111101101",
  4739=>"100000001",
  4740=>"000010100",
  4741=>"000010101",
  4742=>"001100000",
  4743=>"111100001",
  4744=>"000110111",
  4745=>"000110110",
  4746=>"001110100",
  4747=>"101111110",
  4748=>"101100010",
  4749=>"001111101",
  4750=>"111000100",
  4751=>"111011010",
  4752=>"111000011",
  4753=>"001101100",
  4754=>"001010000",
  4755=>"000000010",
  4756=>"010000010",
  4757=>"101001111",
  4758=>"111111000",
  4759=>"001111101",
  4760=>"001010000",
  4761=>"010101101",
  4762=>"001100010",
  4763=>"110010000",
  4764=>"000111100",
  4765=>"010000110",
  4766=>"001011000",
  4767=>"100001010",
  4768=>"000110010",
  4769=>"010001010",
  4770=>"110011011",
  4771=>"001000111",
  4772=>"101001011",
  4773=>"000101111",
  4774=>"000000111",
  4775=>"011001101",
  4776=>"110011000",
  4777=>"100110110",
  4778=>"010110011",
  4779=>"011100001",
  4780=>"000000111",
  4781=>"101001000",
  4782=>"110010010",
  4783=>"011011101",
  4784=>"010001100",
  4785=>"110001111",
  4786=>"010101000",
  4787=>"100100000",
  4788=>"111000010",
  4789=>"101001011",
  4790=>"100010110",
  4791=>"111010101",
  4792=>"011101000",
  4793=>"100000110",
  4794=>"011010111",
  4795=>"010110100",
  4796=>"001100110",
  4797=>"010010101",
  4798=>"011110010",
  4799=>"010011011",
  4800=>"011011110",
  4801=>"111100000",
  4802=>"101111110",
  4803=>"010011001",
  4804=>"000000011",
  4805=>"011001110",
  4806=>"110001111",
  4807=>"000101011",
  4808=>"110010111",
  4809=>"101110011",
  4810=>"000110010",
  4811=>"111111110",
  4812=>"010100010",
  4813=>"110011111",
  4814=>"111111100",
  4815=>"110010011",
  4816=>"000011110",
  4817=>"001100111",
  4818=>"011111011",
  4819=>"110001010",
  4820=>"100001101",
  4821=>"000010111",
  4822=>"100000010",
  4823=>"101000000",
  4824=>"011100000",
  4825=>"100110001",
  4826=>"010000000",
  4827=>"011111011",
  4828=>"001011111",
  4829=>"110111100",
  4830=>"001001111",
  4831=>"101111001",
  4832=>"010011001",
  4833=>"001111010",
  4834=>"010000011",
  4835=>"010100101",
  4836=>"000111001",
  4837=>"001110110",
  4838=>"111111001",
  4839=>"011000010",
  4840=>"011111000",
  4841=>"011111111",
  4842=>"010010010",
  4843=>"000111000",
  4844=>"000000001",
  4845=>"000010011",
  4846=>"111001010",
  4847=>"110100001",
  4848=>"011001000",
  4849=>"111001001",
  4850=>"011101001",
  4851=>"000011011",
  4852=>"100001011",
  4853=>"100110101",
  4854=>"010110110",
  4855=>"100101101",
  4856=>"000000101",
  4857=>"100110110",
  4858=>"001100110",
  4859=>"000110001",
  4860=>"010010100",
  4861=>"001110100",
  4862=>"011010110",
  4863=>"001011110",
  4864=>"101110001",
  4865=>"011110100",
  4866=>"111001000",
  4867=>"010101000",
  4868=>"101111101",
  4869=>"101100111",
  4870=>"000100010",
  4871=>"101011111",
  4872=>"001100101",
  4873=>"011000111",
  4874=>"111001101",
  4875=>"100000100",
  4876=>"010000111",
  4877=>"000101101",
  4878=>"000100101",
  4879=>"001001110",
  4880=>"100101000",
  4881=>"010000010",
  4882=>"111111000",
  4883=>"111110100",
  4884=>"011010000",
  4885=>"100000111",
  4886=>"111111111",
  4887=>"101011011",
  4888=>"101110101",
  4889=>"110000001",
  4890=>"000001000",
  4891=>"001111011",
  4892=>"101011110",
  4893=>"001101011",
  4894=>"001110001",
  4895=>"101011000",
  4896=>"000000100",
  4897=>"110111110",
  4898=>"101111001",
  4899=>"011011110",
  4900=>"100011011",
  4901=>"111101001",
  4902=>"101000010",
  4903=>"011000100",
  4904=>"010011100",
  4905=>"010011010",
  4906=>"000001000",
  4907=>"111100001",
  4908=>"110101000",
  4909=>"100110100",
  4910=>"111100001",
  4911=>"000001100",
  4912=>"001100110",
  4913=>"111010101",
  4914=>"001100111",
  4915=>"101010100",
  4916=>"100110011",
  4917=>"110011000",
  4918=>"100001101",
  4919=>"110110001",
  4920=>"011110011",
  4921=>"110001011",
  4922=>"111000100",
  4923=>"101101000",
  4924=>"001001000",
  4925=>"111110001",
  4926=>"010000001",
  4927=>"100100111",
  4928=>"100110111",
  4929=>"000000001",
  4930=>"111010001",
  4931=>"101111011",
  4932=>"010010110",
  4933=>"111101000",
  4934=>"111010101",
  4935=>"011110101",
  4936=>"111010001",
  4937=>"111001110",
  4938=>"111111011",
  4939=>"001001100",
  4940=>"011100111",
  4941=>"010111101",
  4942=>"100011011",
  4943=>"100010001",
  4944=>"101111101",
  4945=>"000011001",
  4946=>"000001000",
  4947=>"011010011",
  4948=>"001001101",
  4949=>"101000101",
  4950=>"011101100",
  4951=>"111110010",
  4952=>"011111100",
  4953=>"110000010",
  4954=>"011011100",
  4955=>"110001011",
  4956=>"101100010",
  4957=>"111111000",
  4958=>"100000010",
  4959=>"010101101",
  4960=>"011101111",
  4961=>"111010111",
  4962=>"100001100",
  4963=>"011011101",
  4964=>"101110100",
  4965=>"010110110",
  4966=>"110011111",
  4967=>"011111011",
  4968=>"111111100",
  4969=>"100001000",
  4970=>"010110110",
  4971=>"001010001",
  4972=>"000001001",
  4973=>"110110110",
  4974=>"001011101",
  4975=>"011010011",
  4976=>"101101110",
  4977=>"100101110",
  4978=>"111010000",
  4979=>"010110101",
  4980=>"000001000",
  4981=>"111000000",
  4982=>"000110010",
  4983=>"110111111",
  4984=>"011011010",
  4985=>"011000100",
  4986=>"110000010",
  4987=>"100100111",
  4988=>"011101000",
  4989=>"111010011",
  4990=>"000100010",
  4991=>"011100001",
  4992=>"000101001",
  4993=>"111000000",
  4994=>"000101101",
  4995=>"010011011",
  4996=>"010001100",
  4997=>"110010010",
  4998=>"000110010",
  4999=>"001100000",
  5000=>"101110111",
  5001=>"000101000",
  5002=>"010010010",
  5003=>"111011111",
  5004=>"101110000",
  5005=>"111010110",
  5006=>"011001010",
  5007=>"011011001",
  5008=>"000001001",
  5009=>"100101010",
  5010=>"000111100",
  5011=>"000001001",
  5012=>"111111100",
  5013=>"011100100",
  5014=>"110110010",
  5015=>"101100010",
  5016=>"001001101",
  5017=>"001000000",
  5018=>"100110011",
  5019=>"110110011",
  5020=>"010100100",
  5021=>"011101011",
  5022=>"110011001",
  5023=>"010010010",
  5024=>"011101001",
  5025=>"000110111",
  5026=>"101001100",
  5027=>"001100101",
  5028=>"011111101",
  5029=>"001111100",
  5030=>"100000110",
  5031=>"011111101",
  5032=>"001001100",
  5033=>"101111100",
  5034=>"110001110",
  5035=>"101001110",
  5036=>"101011011",
  5037=>"101001011",
  5038=>"101111000",
  5039=>"000110000",
  5040=>"001000101",
  5041=>"110000110",
  5042=>"100010000",
  5043=>"111000001",
  5044=>"110001011",
  5045=>"111010111",
  5046=>"000101001",
  5047=>"001111110",
  5048=>"010011011",
  5049=>"010111101",
  5050=>"101010001",
  5051=>"101011000",
  5052=>"101101111",
  5053=>"010001010",
  5054=>"010011111",
  5055=>"010011011",
  5056=>"001011111",
  5057=>"110100101",
  5058=>"011011101",
  5059=>"011110101",
  5060=>"001011111",
  5061=>"111101001",
  5062=>"101011000",
  5063=>"011101001",
  5064=>"110011000",
  5065=>"101101111",
  5066=>"010111010",
  5067=>"011110100",
  5068=>"100001110",
  5069=>"111011000",
  5070=>"010000111",
  5071=>"011010110",
  5072=>"100111111",
  5073=>"010100000",
  5074=>"000001000",
  5075=>"011000111",
  5076=>"111101101",
  5077=>"101110010",
  5078=>"010011011",
  5079=>"011011111",
  5080=>"011001000",
  5081=>"010011011",
  5082=>"000011110",
  5083=>"000000100",
  5084=>"001100001",
  5085=>"111110011",
  5086=>"011100000",
  5087=>"011101001",
  5088=>"000001001",
  5089=>"011110010",
  5090=>"111010111",
  5091=>"110000110",
  5092=>"010001111",
  5093=>"100100010",
  5094=>"001011001",
  5095=>"101101011",
  5096=>"001100001",
  5097=>"110101101",
  5098=>"100100101",
  5099=>"001000101",
  5100=>"011000100",
  5101=>"001000001",
  5102=>"001011110",
  5103=>"010110100",
  5104=>"000111010",
  5105=>"111001001",
  5106=>"100001010",
  5107=>"001101000",
  5108=>"001001011",
  5109=>"010110010",
  5110=>"000101101",
  5111=>"001100111",
  5112=>"110000011",
  5113=>"101000011",
  5114=>"111110111",
  5115=>"001110000",
  5116=>"010110010",
  5117=>"011010001",
  5118=>"010011101",
  5119=>"101001100",
  5120=>"101010100",
  5121=>"100111000",
  5122=>"011111000",
  5123=>"111100110",
  5124=>"000000000",
  5125=>"000000101",
  5126=>"101100100",
  5127=>"111100001",
  5128=>"001100000",
  5129=>"000111110",
  5130=>"000000000",
  5131=>"101011000",
  5132=>"010110010",
  5133=>"011000100",
  5134=>"110001010",
  5135=>"011010000",
  5136=>"010011001",
  5137=>"010111010",
  5138=>"011110010",
  5139=>"100000011",
  5140=>"000011000",
  5141=>"011011100",
  5142=>"010001000",
  5143=>"100100101",
  5144=>"110001011",
  5145=>"101000011",
  5146=>"101010010",
  5147=>"011001101",
  5148=>"110001000",
  5149=>"100001001",
  5150=>"011100001",
  5151=>"000011100",
  5152=>"010001111",
  5153=>"100011101",
  5154=>"010100000",
  5155=>"111000011",
  5156=>"110100011",
  5157=>"110010110",
  5158=>"010010011",
  5159=>"100101010",
  5160=>"001010000",
  5161=>"001001111",
  5162=>"010110100",
  5163=>"110110100",
  5164=>"100110100",
  5165=>"000101111",
  5166=>"010000111",
  5167=>"100010110",
  5168=>"100011001",
  5169=>"001010101",
  5170=>"010011111",
  5171=>"101000001",
  5172=>"010101000",
  5173=>"010100011",
  5174=>"001101011",
  5175=>"110101100",
  5176=>"101011100",
  5177=>"110110000",
  5178=>"010100110",
  5179=>"110001011",
  5180=>"100000011",
  5181=>"000000001",
  5182=>"011010100",
  5183=>"001111111",
  5184=>"001101001",
  5185=>"001101001",
  5186=>"111100100",
  5187=>"101001100",
  5188=>"110111110",
  5189=>"011011000",
  5190=>"000000011",
  5191=>"011101110",
  5192=>"101110001",
  5193=>"000010001",
  5194=>"111111111",
  5195=>"100011101",
  5196=>"110101000",
  5197=>"111100101",
  5198=>"110011110",
  5199=>"000000000",
  5200=>"001110011",
  5201=>"000010110",
  5202=>"101111010",
  5203=>"100000111",
  5204=>"101101110",
  5205=>"010010010",
  5206=>"011010111",
  5207=>"100101001",
  5208=>"000110101",
  5209=>"100100111",
  5210=>"010101101",
  5211=>"000010000",
  5212=>"110011010",
  5213=>"000011110",
  5214=>"000000011",
  5215=>"111000110",
  5216=>"011000000",
  5217=>"010010100",
  5218=>"111111011",
  5219=>"100001010",
  5220=>"000100110",
  5221=>"001001110",
  5222=>"101001110",
  5223=>"001111000",
  5224=>"101101010",
  5225=>"010111001",
  5226=>"000010010",
  5227=>"101111010",
  5228=>"001100101",
  5229=>"010011010",
  5230=>"010110011",
  5231=>"000011111",
  5232=>"110100000",
  5233=>"101011001",
  5234=>"111111101",
  5235=>"110110100",
  5236=>"010111010",
  5237=>"011001100",
  5238=>"100100101",
  5239=>"001000111",
  5240=>"011011011",
  5241=>"101110000",
  5242=>"000001110",
  5243=>"000000010",
  5244=>"111000000",
  5245=>"010101110",
  5246=>"010011000",
  5247=>"001001000",
  5248=>"011000101",
  5249=>"011100010",
  5250=>"010011001",
  5251=>"000001011",
  5252=>"101010100",
  5253=>"100111001",
  5254=>"001101010",
  5255=>"111101111",
  5256=>"101000100",
  5257=>"000100001",
  5258=>"100100000",
  5259=>"100010011",
  5260=>"001000111",
  5261=>"011110010",
  5262=>"101111100",
  5263=>"000110101",
  5264=>"010000111",
  5265=>"111000001",
  5266=>"111100111",
  5267=>"100010110",
  5268=>"111111010",
  5269=>"010010000",
  5270=>"001010001",
  5271=>"011000001",
  5272=>"101011001",
  5273=>"000010000",
  5274=>"000011000",
  5275=>"100101000",
  5276=>"010010001",
  5277=>"011100000",
  5278=>"100010001",
  5279=>"010101001",
  5280=>"100110101",
  5281=>"110110110",
  5282=>"000000000",
  5283=>"000010000",
  5284=>"010100000",
  5285=>"101110111",
  5286=>"100010011",
  5287=>"101010101",
  5288=>"001011000",
  5289=>"010011000",
  5290=>"101101100",
  5291=>"001100101",
  5292=>"110000001",
  5293=>"111110111",
  5294=>"100000100",
  5295=>"101111111",
  5296=>"101101100",
  5297=>"010100101",
  5298=>"000000001",
  5299=>"011010010",
  5300=>"011011110",
  5301=>"000011010",
  5302=>"010010000",
  5303=>"001011110",
  5304=>"010010011",
  5305=>"111000111",
  5306=>"111100101",
  5307=>"001100011",
  5308=>"011110111",
  5309=>"000111001",
  5310=>"000001101",
  5311=>"011011110",
  5312=>"000101101",
  5313=>"010001100",
  5314=>"000101100",
  5315=>"000101010",
  5316=>"110001111",
  5317=>"000001110",
  5318=>"001100110",
  5319=>"010111000",
  5320=>"001110011",
  5321=>"010010001",
  5322=>"011101110",
  5323=>"100100000",
  5324=>"100001011",
  5325=>"001101001",
  5326=>"111111001",
  5327=>"111000001",
  5328=>"100001000",
  5329=>"010011110",
  5330=>"001100000",
  5331=>"101011110",
  5332=>"011000110",
  5333=>"101011111",
  5334=>"001000111",
  5335=>"001110011",
  5336=>"100111110",
  5337=>"111010000",
  5338=>"000010100",
  5339=>"010110001",
  5340=>"001011010",
  5341=>"100100110",
  5342=>"000100100",
  5343=>"011011101",
  5344=>"000011110",
  5345=>"011111000",
  5346=>"100100001",
  5347=>"001110000",
  5348=>"100110101",
  5349=>"001110011",
  5350=>"000001111",
  5351=>"000110110",
  5352=>"100011001",
  5353=>"110010110",
  5354=>"000010000",
  5355=>"100001011",
  5356=>"101010001",
  5357=>"011100001",
  5358=>"010011110",
  5359=>"001110111",
  5360=>"110101010",
  5361=>"000010110",
  5362=>"001001001",
  5363=>"110100101",
  5364=>"101111011",
  5365=>"100110101",
  5366=>"101011100",
  5367=>"110001111",
  5368=>"000100010",
  5369=>"011001010",
  5370=>"110000101",
  5371=>"101000000",
  5372=>"111001100",
  5373=>"100001110",
  5374=>"000110001",
  5375=>"000100101",
  5376=>"001010001",
  5377=>"010011111",
  5378=>"001010010",
  5379=>"101010011",
  5380=>"000000111",
  5381=>"111010001",
  5382=>"011001110",
  5383=>"011001011",
  5384=>"001000000",
  5385=>"001000101",
  5386=>"100001000",
  5387=>"011000111",
  5388=>"011111001",
  5389=>"010000000",
  5390=>"001000101",
  5391=>"000011001",
  5392=>"111001000",
  5393=>"101011010",
  5394=>"010100111",
  5395=>"110101101",
  5396=>"001100000",
  5397=>"000000001",
  5398=>"000101111",
  5399=>"010001010",
  5400=>"111011000",
  5401=>"101111100",
  5402=>"000010000",
  5403=>"111111010",
  5404=>"001111000",
  5405=>"111000000",
  5406=>"101101010",
  5407=>"101000110",
  5408=>"110000010",
  5409=>"000011101",
  5410=>"111000110",
  5411=>"010000111",
  5412=>"110000111",
  5413=>"010101000",
  5414=>"100101110",
  5415=>"000111110",
  5416=>"001011001",
  5417=>"010000101",
  5418=>"100100111",
  5419=>"111011010",
  5420=>"101000001",
  5421=>"001010000",
  5422=>"000011111",
  5423=>"111011111",
  5424=>"000110111",
  5425=>"010000001",
  5426=>"111101000",
  5427=>"101000001",
  5428=>"000000000",
  5429=>"010000001",
  5430=>"110000011",
  5431=>"011101001",
  5432=>"110110001",
  5433=>"001000010",
  5434=>"011100011",
  5435=>"000111001",
  5436=>"010101110",
  5437=>"001111001",
  5438=>"011111011",
  5439=>"110100110",
  5440=>"001110010",
  5441=>"001000100",
  5442=>"101110111",
  5443=>"100011101",
  5444=>"000010111",
  5445=>"110110110",
  5446=>"111001100",
  5447=>"001001001",
  5448=>"010100101",
  5449=>"011010000",
  5450=>"101011110",
  5451=>"000000100",
  5452=>"001111110",
  5453=>"111011000",
  5454=>"000001010",
  5455=>"010111110",
  5456=>"101110000",
  5457=>"011111111",
  5458=>"100111101",
  5459=>"000110000",
  5460=>"010111010",
  5461=>"101000101",
  5462=>"110100100",
  5463=>"001011001",
  5464=>"000101010",
  5465=>"010000000",
  5466=>"100101100",
  5467=>"010100100",
  5468=>"110101001",
  5469=>"001001100",
  5470=>"010000001",
  5471=>"100010000",
  5472=>"111010110",
  5473=>"111010100",
  5474=>"011111110",
  5475=>"001100011",
  5476=>"111110010",
  5477=>"100001110",
  5478=>"001101000",
  5479=>"110001100",
  5480=>"011000111",
  5481=>"000001011",
  5482=>"101000001",
  5483=>"101000011",
  5484=>"000101111",
  5485=>"110001011",
  5486=>"100111000",
  5487=>"101001010",
  5488=>"111001110",
  5489=>"001001011",
  5490=>"101110110",
  5491=>"100110101",
  5492=>"010001001",
  5493=>"010000100",
  5494=>"010000000",
  5495=>"000000110",
  5496=>"001000001",
  5497=>"101101010",
  5498=>"111101101",
  5499=>"011101000",
  5500=>"110001101",
  5501=>"111111011",
  5502=>"110111000",
  5503=>"011000001",
  5504=>"001110010",
  5505=>"111010111",
  5506=>"100110110",
  5507=>"011110010",
  5508=>"111111011",
  5509=>"000010000",
  5510=>"101001100",
  5511=>"111101111",
  5512=>"011100001",
  5513=>"100111111",
  5514=>"010011011",
  5515=>"101010011",
  5516=>"010010001",
  5517=>"001100110",
  5518=>"101010100",
  5519=>"001011000",
  5520=>"001000000",
  5521=>"100010000",
  5522=>"011100100",
  5523=>"000111100",
  5524=>"100001000",
  5525=>"111111111",
  5526=>"001000000",
  5527=>"101000000",
  5528=>"011110100",
  5529=>"010110101",
  5530=>"000100000",
  5531=>"010100110",
  5532=>"110000010",
  5533=>"000011101",
  5534=>"000110100",
  5535=>"011001111",
  5536=>"011110101",
  5537=>"010001000",
  5538=>"010110100",
  5539=>"000010101",
  5540=>"111100101",
  5541=>"110001010",
  5542=>"001010010",
  5543=>"001000011",
  5544=>"100100110",
  5545=>"110011011",
  5546=>"000110111",
  5547=>"111110011",
  5548=>"010100101",
  5549=>"101011111",
  5550=>"000100001",
  5551=>"110011000",
  5552=>"101011110",
  5553=>"110000111",
  5554=>"000101001",
  5555=>"010000111",
  5556=>"111110100",
  5557=>"100101010",
  5558=>"000100111",
  5559=>"110100011",
  5560=>"111001100",
  5561=>"101000101",
  5562=>"100001110",
  5563=>"100011110",
  5564=>"100111100",
  5565=>"011110100",
  5566=>"010100110",
  5567=>"111100001",
  5568=>"001001011",
  5569=>"001011110",
  5570=>"010001000",
  5571=>"011010000",
  5572=>"100000000",
  5573=>"001100101",
  5574=>"011110010",
  5575=>"010010100",
  5576=>"011101110",
  5577=>"101110000",
  5578=>"110111001",
  5579=>"100100110",
  5580=>"000100010",
  5581=>"100111110",
  5582=>"111001101",
  5583=>"111000011",
  5584=>"101111010",
  5585=>"100000111",
  5586=>"101100000",
  5587=>"110110010",
  5588=>"000001001",
  5589=>"000001110",
  5590=>"101101110",
  5591=>"010100110",
  5592=>"001000110",
  5593=>"001010010",
  5594=>"110110011",
  5595=>"111101001",
  5596=>"111101010",
  5597=>"001100100",
  5598=>"100011101",
  5599=>"000011100",
  5600=>"010100000",
  5601=>"100010001",
  5602=>"100100110",
  5603=>"101110000",
  5604=>"011000110",
  5605=>"111101111",
  5606=>"000111000",
  5607=>"010111110",
  5608=>"011000101",
  5609=>"010001111",
  5610=>"010001001",
  5611=>"001100010",
  5612=>"111010100",
  5613=>"100010111",
  5614=>"110111001",
  5615=>"011100010",
  5616=>"111001111",
  5617=>"110111101",
  5618=>"000011100",
  5619=>"010001100",
  5620=>"110010101",
  5621=>"100111110",
  5622=>"011111101",
  5623=>"100010100",
  5624=>"100010100",
  5625=>"000111101",
  5626=>"010010110",
  5627=>"101011110",
  5628=>"111111110",
  5629=>"000010011",
  5630=>"011001111",
  5631=>"100101100",
  5632=>"111100010",
  5633=>"010001110",
  5634=>"110000010",
  5635=>"100000001",
  5636=>"000010000",
  5637=>"010001111",
  5638=>"110010110",
  5639=>"010100000",
  5640=>"010110101",
  5641=>"010110011",
  5642=>"110111110",
  5643=>"000010100",
  5644=>"001001100",
  5645=>"110001111",
  5646=>"111110111",
  5647=>"101111110",
  5648=>"001100110",
  5649=>"110101101",
  5650=>"101110111",
  5651=>"111111100",
  5652=>"101110101",
  5653=>"101010010",
  5654=>"001110000",
  5655=>"010110010",
  5656=>"110000010",
  5657=>"011000000",
  5658=>"101111000",
  5659=>"111101011",
  5660=>"100100110",
  5661=>"000011011",
  5662=>"000111110",
  5663=>"011010000",
  5664=>"010010000",
  5665=>"100001111",
  5666=>"011011011",
  5667=>"000100001",
  5668=>"110111101",
  5669=>"001011010",
  5670=>"000101001",
  5671=>"001000010",
  5672=>"011000001",
  5673=>"111011111",
  5674=>"111100001",
  5675=>"100010100",
  5676=>"101101010",
  5677=>"100110100",
  5678=>"100001001",
  5679=>"111010000",
  5680=>"101010100",
  5681=>"110111011",
  5682=>"000111100",
  5683=>"100000100",
  5684=>"011011001",
  5685=>"011111111",
  5686=>"101000101",
  5687=>"000001001",
  5688=>"010110011",
  5689=>"111101111",
  5690=>"100100111",
  5691=>"101010010",
  5692=>"011010101",
  5693=>"100100110",
  5694=>"100011011",
  5695=>"100111010",
  5696=>"110000000",
  5697=>"010111011",
  5698=>"010101100",
  5699=>"000100000",
  5700=>"011100000",
  5701=>"100000100",
  5702=>"110101000",
  5703=>"010100011",
  5704=>"101100101",
  5705=>"101011110",
  5706=>"100101100",
  5707=>"100100000",
  5708=>"101001001",
  5709=>"100100001",
  5710=>"101100101",
  5711=>"011000110",
  5712=>"111010101",
  5713=>"001100111",
  5714=>"111100111",
  5715=>"101000011",
  5716=>"001101011",
  5717=>"001001001",
  5718=>"111110110",
  5719=>"111101000",
  5720=>"000000000",
  5721=>"100111001",
  5722=>"111111111",
  5723=>"001001110",
  5724=>"010011000",
  5725=>"100010111",
  5726=>"000010101",
  5727=>"111001010",
  5728=>"001001001",
  5729=>"100000001",
  5730=>"100011000",
  5731=>"100111011",
  5732=>"100010110",
  5733=>"001110101",
  5734=>"100000000",
  5735=>"100010101",
  5736=>"101001011",
  5737=>"010011010",
  5738=>"100101110",
  5739=>"101101001",
  5740=>"001111101",
  5741=>"111101011",
  5742=>"111010100",
  5743=>"111110110",
  5744=>"010001101",
  5745=>"001011110",
  5746=>"011001101",
  5747=>"010001100",
  5748=>"110111101",
  5749=>"100100111",
  5750=>"101110010",
  5751=>"010000100",
  5752=>"010100001",
  5753=>"101000101",
  5754=>"111011110",
  5755=>"101110001",
  5756=>"111001010",
  5757=>"011010011",
  5758=>"110101001",
  5759=>"100011000",
  5760=>"000010011",
  5761=>"011100000",
  5762=>"010001000",
  5763=>"000001110",
  5764=>"110101010",
  5765=>"001100000",
  5766=>"011110001",
  5767=>"111000111",
  5768=>"000101000",
  5769=>"111101101",
  5770=>"101010111",
  5771=>"000100011",
  5772=>"100001000",
  5773=>"000101101",
  5774=>"010111011",
  5775=>"010010000",
  5776=>"001001001",
  5777=>"100001101",
  5778=>"000000100",
  5779=>"000101010",
  5780=>"000110001",
  5781=>"011100011",
  5782=>"101110000",
  5783=>"010111100",
  5784=>"111110111",
  5785=>"100011000",
  5786=>"001110001",
  5787=>"110111001",
  5788=>"110001101",
  5789=>"010101000",
  5790=>"101000001",
  5791=>"001000000",
  5792=>"110010000",
  5793=>"010001001",
  5794=>"011000000",
  5795=>"100000110",
  5796=>"100100010",
  5797=>"111101000",
  5798=>"001000100",
  5799=>"100100000",
  5800=>"010110100",
  5801=>"111010101",
  5802=>"001000001",
  5803=>"011000000",
  5804=>"111101011",
  5805=>"010010000",
  5806=>"001111110",
  5807=>"100110011",
  5808=>"101110110",
  5809=>"010000110",
  5810=>"100110110",
  5811=>"011011101",
  5812=>"000000000",
  5813=>"100110100",
  5814=>"011000111",
  5815=>"110010100",
  5816=>"001011110",
  5817=>"000010011",
  5818=>"110111100",
  5819=>"101001111",
  5820=>"001000111",
  5821=>"101011110",
  5822=>"000101011",
  5823=>"000011100",
  5824=>"100101011",
  5825=>"000101001",
  5826=>"111011110",
  5827=>"100001010",
  5828=>"101001010",
  5829=>"000111000",
  5830=>"101010111",
  5831=>"000001110",
  5832=>"100100110",
  5833=>"100100100",
  5834=>"001101011",
  5835=>"010000101",
  5836=>"100111001",
  5837=>"100110111",
  5838=>"111010101",
  5839=>"011110011",
  5840=>"110001010",
  5841=>"101110000",
  5842=>"110000010",
  5843=>"111111100",
  5844=>"111010101",
  5845=>"011101011",
  5846=>"101111100",
  5847=>"000011010",
  5848=>"011000011",
  5849=>"001010101",
  5850=>"011010001",
  5851=>"001111111",
  5852=>"110110010",
  5853=>"000010000",
  5854=>"100111000",
  5855=>"111010000",
  5856=>"100111001",
  5857=>"011000100",
  5858=>"011100011",
  5859=>"110100000",
  5860=>"000111100",
  5861=>"111100000",
  5862=>"110100000",
  5863=>"000011111",
  5864=>"001101001",
  5865=>"110010101",
  5866=>"101011110",
  5867=>"101100011",
  5868=>"001101110",
  5869=>"000111001",
  5870=>"110010000",
  5871=>"000001001",
  5872=>"100001111",
  5873=>"101001110",
  5874=>"111000111",
  5875=>"001001010",
  5876=>"000011101",
  5877=>"010011100",
  5878=>"110000001",
  5879=>"000010000",
  5880=>"101110010",
  5881=>"100000100",
  5882=>"111011011",
  5883=>"000100010",
  5884=>"100101001",
  5885=>"010001110",
  5886=>"010000101",
  5887=>"001101100",
  5888=>"101110101",
  5889=>"100000111",
  5890=>"010111100",
  5891=>"000111000",
  5892=>"011001110",
  5893=>"010010011",
  5894=>"000001101",
  5895=>"010101000",
  5896=>"000101011",
  5897=>"010010111",
  5898=>"000010000",
  5899=>"101101101",
  5900=>"010010000",
  5901=>"101111100",
  5902=>"111000101",
  5903=>"011000000",
  5904=>"111101111",
  5905=>"001101100",
  5906=>"110000011",
  5907=>"100000100",
  5908=>"100001001",
  5909=>"000111000",
  5910=>"011001100",
  5911=>"100110101",
  5912=>"111001100",
  5913=>"110101000",
  5914=>"000000110",
  5915=>"111100110",
  5916=>"001010101",
  5917=>"010111001",
  5918=>"010110001",
  5919=>"000001001",
  5920=>"110001101",
  5921=>"000011000",
  5922=>"101001111",
  5923=>"100011101",
  5924=>"110110110",
  5925=>"000000111",
  5926=>"011011000",
  5927=>"000010100",
  5928=>"000011100",
  5929=>"101011010",
  5930=>"101010010",
  5931=>"111111100",
  5932=>"011010001",
  5933=>"011010111",
  5934=>"000010110",
  5935=>"000110101",
  5936=>"100111010",
  5937=>"000000100",
  5938=>"010000000",
  5939=>"110001110",
  5940=>"001110010",
  5941=>"010111110",
  5942=>"000010000",
  5943=>"000010111",
  5944=>"001000010",
  5945=>"010011101",
  5946=>"011110110",
  5947=>"110111111",
  5948=>"001100010",
  5949=>"110011100",
  5950=>"110111110",
  5951=>"010011110",
  5952=>"011101111",
  5953=>"101001001",
  5954=>"011110010",
  5955=>"111100101",
  5956=>"000111110",
  5957=>"100000010",
  5958=>"110110111",
  5959=>"001011110",
  5960=>"100101011",
  5961=>"000010000",
  5962=>"101110001",
  5963=>"010110100",
  5964=>"010110001",
  5965=>"110101101",
  5966=>"011010101",
  5967=>"100011011",
  5968=>"011000000",
  5969=>"011100110",
  5970=>"010011100",
  5971=>"011000110",
  5972=>"101001110",
  5973=>"010001111",
  5974=>"001100100",
  5975=>"110010111",
  5976=>"010110010",
  5977=>"111011010",
  5978=>"101101001",
  5979=>"110000111",
  5980=>"101000100",
  5981=>"111000100",
  5982=>"111011101",
  5983=>"101000111",
  5984=>"101010111",
  5985=>"010111011",
  5986=>"000000001",
  5987=>"011101111",
  5988=>"010010000",
  5989=>"001100001",
  5990=>"001010110",
  5991=>"001000110",
  5992=>"011010100",
  5993=>"010111101",
  5994=>"010101110",
  5995=>"110010110",
  5996=>"111001000",
  5997=>"000000111",
  5998=>"001001111",
  5999=>"001001001",
  6000=>"001101010",
  6001=>"000111100",
  6002=>"111110000",
  6003=>"111111101",
  6004=>"000000100",
  6005=>"001000011",
  6006=>"001111110",
  6007=>"100010000",
  6008=>"101100010",
  6009=>"010000010",
  6010=>"111100101",
  6011=>"100000011",
  6012=>"000000000",
  6013=>"010000000",
  6014=>"000001111",
  6015=>"101110011",
  6016=>"000001110",
  6017=>"111110000",
  6018=>"000000100",
  6019=>"100000000",
  6020=>"011100100",
  6021=>"110010011",
  6022=>"111111101",
  6023=>"101010001",
  6024=>"110110011",
  6025=>"011100100",
  6026=>"010110001",
  6027=>"000010011",
  6028=>"100100100",
  6029=>"100100011",
  6030=>"010100110",
  6031=>"000100010",
  6032=>"001011100",
  6033=>"011011011",
  6034=>"100000101",
  6035=>"101000011",
  6036=>"110111111",
  6037=>"001111110",
  6038=>"000010111",
  6039=>"110110011",
  6040=>"001001100",
  6041=>"100100011",
  6042=>"011011111",
  6043=>"110111010",
  6044=>"010110111",
  6045=>"111101100",
  6046=>"010111001",
  6047=>"100000011",
  6048=>"100001001",
  6049=>"110001000",
  6050=>"101100001",
  6051=>"111000101",
  6052=>"000000000",
  6053=>"000111000",
  6054=>"011100100",
  6055=>"110000010",
  6056=>"100100011",
  6057=>"000001101",
  6058=>"111111111",
  6059=>"000100011",
  6060=>"000001010",
  6061=>"100000011",
  6062=>"001110010",
  6063=>"010111011",
  6064=>"000001001",
  6065=>"101110010",
  6066=>"111000011",
  6067=>"010100001",
  6068=>"000000010",
  6069=>"101111001",
  6070=>"010010111",
  6071=>"000111001",
  6072=>"110101111",
  6073=>"101000110",
  6074=>"001001001",
  6075=>"101110011",
  6076=>"100010010",
  6077=>"011010011",
  6078=>"101100110",
  6079=>"001101000",
  6080=>"100100110",
  6081=>"110010011",
  6082=>"000111011",
  6083=>"000101001",
  6084=>"000000110",
  6085=>"111000110",
  6086=>"000000010",
  6087=>"011010111",
  6088=>"100100110",
  6089=>"001100000",
  6090=>"001101010",
  6091=>"110001001",
  6092=>"100110111",
  6093=>"110000010",
  6094=>"101000011",
  6095=>"010011111",
  6096=>"000100000",
  6097=>"100000000",
  6098=>"000010111",
  6099=>"010000000",
  6100=>"011100101",
  6101=>"110001100",
  6102=>"110101000",
  6103=>"011101111",
  6104=>"100000000",
  6105=>"010010101",
  6106=>"011101010",
  6107=>"000001010",
  6108=>"000001100",
  6109=>"001100101",
  6110=>"011010000",
  6111=>"000000110",
  6112=>"011110111",
  6113=>"001011101",
  6114=>"100011101",
  6115=>"110000110",
  6116=>"100010010",
  6117=>"000001111",
  6118=>"111001101",
  6119=>"001000100",
  6120=>"110001000",
  6121=>"111011110",
  6122=>"110011011",
  6123=>"010110111",
  6124=>"111000101",
  6125=>"001010101",
  6126=>"001011100",
  6127=>"111011011",
  6128=>"010000110",
  6129=>"100010011",
  6130=>"101111110",
  6131=>"111111100",
  6132=>"011000111",
  6133=>"101111111",
  6134=>"010101110",
  6135=>"111100001",
  6136=>"111111001",
  6137=>"111000001",
  6138=>"000111011",
  6139=>"101110111",
  6140=>"000000011",
  6141=>"110000111",
  6142=>"000011000",
  6143=>"111000100",
  6144=>"111011111",
  6145=>"111111001",
  6146=>"110011000",
  6147=>"010101110",
  6148=>"100111001",
  6149=>"110101110",
  6150=>"000100111",
  6151=>"110101110",
  6152=>"111010011",
  6153=>"100110000",
  6154=>"010101010",
  6155=>"111011000",
  6156=>"010000001",
  6157=>"110111110",
  6158=>"111110100",
  6159=>"000110111",
  6160=>"011010010",
  6161=>"010000001",
  6162=>"001111101",
  6163=>"000101111",
  6164=>"110001110",
  6165=>"110011001",
  6166=>"000111000",
  6167=>"101101011",
  6168=>"010011111",
  6169=>"101001010",
  6170=>"000001110",
  6171=>"010011000",
  6172=>"100010011",
  6173=>"111011011",
  6174=>"000010100",
  6175=>"001101001",
  6176=>"100000111",
  6177=>"000011111",
  6178=>"001000000",
  6179=>"011100111",
  6180=>"010100000",
  6181=>"100101110",
  6182=>"100100011",
  6183=>"111000010",
  6184=>"011010111",
  6185=>"000111000",
  6186=>"010000100",
  6187=>"010100110",
  6188=>"101010001",
  6189=>"011101100",
  6190=>"111011011",
  6191=>"000000000",
  6192=>"000000110",
  6193=>"001011110",
  6194=>"001011000",
  6195=>"100111001",
  6196=>"010101111",
  6197=>"010001100",
  6198=>"101100001",
  6199=>"110101000",
  6200=>"111110001",
  6201=>"011010000",
  6202=>"001001001",
  6203=>"001000010",
  6204=>"110010001",
  6205=>"110011110",
  6206=>"100001010",
  6207=>"010010000",
  6208=>"111110011",
  6209=>"000001111",
  6210=>"110000000",
  6211=>"000000111",
  6212=>"101011101",
  6213=>"101110001",
  6214=>"100110010",
  6215=>"110100000",
  6216=>"001111011",
  6217=>"101010111",
  6218=>"001111111",
  6219=>"001100010",
  6220=>"101011000",
  6221=>"100000110",
  6222=>"111001011",
  6223=>"011010000",
  6224=>"111001100",
  6225=>"110101100",
  6226=>"101101010",
  6227=>"111111101",
  6228=>"010000000",
  6229=>"111110001",
  6230=>"010110011",
  6231=>"000111000",
  6232=>"111000011",
  6233=>"010001011",
  6234=>"100000011",
  6235=>"001100110",
  6236=>"111101101",
  6237=>"000001010",
  6238=>"001010010",
  6239=>"001100101",
  6240=>"011000111",
  6241=>"101111100",
  6242=>"001110001",
  6243=>"111001001",
  6244=>"101101011",
  6245=>"101001011",
  6246=>"101010001",
  6247=>"000101001",
  6248=>"001100100",
  6249=>"110100001",
  6250=>"100000101",
  6251=>"001010010",
  6252=>"101110100",
  6253=>"111101110",
  6254=>"000011010",
  6255=>"011100101",
  6256=>"111001110",
  6257=>"001110001",
  6258=>"001111001",
  6259=>"011010010",
  6260=>"111100100",
  6261=>"010111001",
  6262=>"110100101",
  6263=>"001100101",
  6264=>"011010111",
  6265=>"100001001",
  6266=>"010001111",
  6267=>"011011011",
  6268=>"001011000",
  6269=>"100101001",
  6270=>"101000010",
  6271=>"001000110",
  6272=>"111111110",
  6273=>"101100111",
  6274=>"010000001",
  6275=>"000100001",
  6276=>"000010000",
  6277=>"111001101",
  6278=>"100111010",
  6279=>"001111100",
  6280=>"011101101",
  6281=>"111000100",
  6282=>"100001100",
  6283=>"001110010",
  6284=>"000100110",
  6285=>"001010101",
  6286=>"010110000",
  6287=>"111111011",
  6288=>"001001011",
  6289=>"001001011",
  6290=>"001011010",
  6291=>"111111000",
  6292=>"010111001",
  6293=>"011000010",
  6294=>"111010110",
  6295=>"101011001",
  6296=>"101000001",
  6297=>"001000000",
  6298=>"001111100",
  6299=>"101001011",
  6300=>"100101011",
  6301=>"011000001",
  6302=>"001100001",
  6303=>"110101101",
  6304=>"111111110",
  6305=>"111111111",
  6306=>"010111100",
  6307=>"001011011",
  6308=>"110101001",
  6309=>"100100011",
  6310=>"011101010",
  6311=>"011110011",
  6312=>"111010000",
  6313=>"110011100",
  6314=>"001001000",
  6315=>"111010001",
  6316=>"010101110",
  6317=>"110000010",
  6318=>"100111100",
  6319=>"111011010",
  6320=>"101101011",
  6321=>"000000100",
  6322=>"110101011",
  6323=>"011010011",
  6324=>"111011001",
  6325=>"111010111",
  6326=>"000000111",
  6327=>"110001010",
  6328=>"101000100",
  6329=>"101010011",
  6330=>"001000001",
  6331=>"101010110",
  6332=>"001001100",
  6333=>"010001101",
  6334=>"001100110",
  6335=>"111111111",
  6336=>"000011011",
  6337=>"010011011",
  6338=>"000011010",
  6339=>"101000110",
  6340=>"000010111",
  6341=>"000110000",
  6342=>"111000010",
  6343=>"111000011",
  6344=>"100001101",
  6345=>"100101100",
  6346=>"110001011",
  6347=>"010100011",
  6348=>"011000100",
  6349=>"011110011",
  6350=>"011101010",
  6351=>"100001011",
  6352=>"010100101",
  6353=>"101000010",
  6354=>"000011001",
  6355=>"110100101",
  6356=>"110110000",
  6357=>"110111010",
  6358=>"101000100",
  6359=>"011110011",
  6360=>"100011010",
  6361=>"111000110",
  6362=>"010000001",
  6363=>"110000001",
  6364=>"001000001",
  6365=>"101000101",
  6366=>"011101100",
  6367=>"010000100",
  6368=>"011101111",
  6369=>"000100111",
  6370=>"011101011",
  6371=>"000000000",
  6372=>"101101001",
  6373=>"101001000",
  6374=>"001010001",
  6375=>"100101011",
  6376=>"001000010",
  6377=>"000001000",
  6378=>"100011111",
  6379=>"101100111",
  6380=>"110000001",
  6381=>"110000111",
  6382=>"000000011",
  6383=>"010100000",
  6384=>"011111111",
  6385=>"001111111",
  6386=>"000101001",
  6387=>"000001010",
  6388=>"011110101",
  6389=>"111101110",
  6390=>"111111100",
  6391=>"010010010",
  6392=>"001001111",
  6393=>"010100000",
  6394=>"101110000",
  6395=>"100010011",
  6396=>"111000110",
  6397=>"010001101",
  6398=>"010101011",
  6399=>"101110000",
  6400=>"111111010",
  6401=>"010000001",
  6402=>"101011101",
  6403=>"000111010",
  6404=>"100101000",
  6405=>"110001111",
  6406=>"011010100",
  6407=>"011101100",
  6408=>"001101010",
  6409=>"101011001",
  6410=>"010001010",
  6411=>"100001011",
  6412=>"110111100",
  6413=>"001001011",
  6414=>"101100010",
  6415=>"001011111",
  6416=>"011001011",
  6417=>"110011010",
  6418=>"011001001",
  6419=>"011111100",
  6420=>"001001110",
  6421=>"000001010",
  6422=>"010000111",
  6423=>"110110101",
  6424=>"110100011",
  6425=>"000001001",
  6426=>"001010110",
  6427=>"110000111",
  6428=>"010000001",
  6429=>"011000111",
  6430=>"111110111",
  6431=>"000110100",
  6432=>"000100100",
  6433=>"100111000",
  6434=>"100100100",
  6435=>"100000001",
  6436=>"100110110",
  6437=>"000100111",
  6438=>"011000111",
  6439=>"011001011",
  6440=>"111111111",
  6441=>"100001011",
  6442=>"000001010",
  6443=>"011110000",
  6444=>"101010110",
  6445=>"000000110",
  6446=>"101001000",
  6447=>"101011000",
  6448=>"010000011",
  6449=>"100110111",
  6450=>"011111001",
  6451=>"001101000",
  6452=>"111000101",
  6453=>"000010000",
  6454=>"010111101",
  6455=>"100100111",
  6456=>"000000110",
  6457=>"011010111",
  6458=>"100110110",
  6459=>"001111000",
  6460=>"001101001",
  6461=>"010011001",
  6462=>"111011010",
  6463=>"001011000",
  6464=>"111101010",
  6465=>"100110000",
  6466=>"101001001",
  6467=>"110011101",
  6468=>"001111000",
  6469=>"010100110",
  6470=>"001000000",
  6471=>"000110100",
  6472=>"001011001",
  6473=>"011100111",
  6474=>"100110101",
  6475=>"101001010",
  6476=>"100110101",
  6477=>"101111110",
  6478=>"111000111",
  6479=>"111011100",
  6480=>"010001100",
  6481=>"101100101",
  6482=>"111101000",
  6483=>"000101000",
  6484=>"000011010",
  6485=>"001000010",
  6486=>"110010111",
  6487=>"110111100",
  6488=>"101110001",
  6489=>"000001000",
  6490=>"101011111",
  6491=>"001000001",
  6492=>"110010111",
  6493=>"001110101",
  6494=>"111011000",
  6495=>"000010001",
  6496=>"111000010",
  6497=>"010011101",
  6498=>"000111010",
  6499=>"000001110",
  6500=>"010000000",
  6501=>"011000001",
  6502=>"110100111",
  6503=>"101110111",
  6504=>"000111111",
  6505=>"001011111",
  6506=>"101100011",
  6507=>"111101111",
  6508=>"101011111",
  6509=>"100001011",
  6510=>"001001111",
  6511=>"111000101",
  6512=>"001110101",
  6513=>"101011010",
  6514=>"011100011",
  6515=>"111100111",
  6516=>"010101110",
  6517=>"001000001",
  6518=>"110001010",
  6519=>"001011001",
  6520=>"111000101",
  6521=>"111110111",
  6522=>"010001101",
  6523=>"010000010",
  6524=>"111000111",
  6525=>"111001111",
  6526=>"000111010",
  6527=>"010001101",
  6528=>"000011010",
  6529=>"100100001",
  6530=>"001100011",
  6531=>"101000101",
  6532=>"100100101",
  6533=>"001010001",
  6534=>"101010010",
  6535=>"111001100",
  6536=>"100001110",
  6537=>"101110011",
  6538=>"011001100",
  6539=>"110100000",
  6540=>"011010001",
  6541=>"001010111",
  6542=>"010100101",
  6543=>"111011010",
  6544=>"001010101",
  6545=>"111100111",
  6546=>"111100111",
  6547=>"000111111",
  6548=>"001101110",
  6549=>"111011000",
  6550=>"011100011",
  6551=>"111111111",
  6552=>"001001011",
  6553=>"011001011",
  6554=>"011010100",
  6555=>"011000001",
  6556=>"110010010",
  6557=>"101010010",
  6558=>"000110100",
  6559=>"001101100",
  6560=>"000000010",
  6561=>"001110010",
  6562=>"010111111",
  6563=>"101000011",
  6564=>"111000101",
  6565=>"000000011",
  6566=>"010001110",
  6567=>"100101101",
  6568=>"101110011",
  6569=>"011010101",
  6570=>"000100100",
  6571=>"010011000",
  6572=>"000011010",
  6573=>"100111011",
  6574=>"100110001",
  6575=>"010000011",
  6576=>"101100110",
  6577=>"011000000",
  6578=>"100100111",
  6579=>"000010110",
  6580=>"010001011",
  6581=>"110111000",
  6582=>"000000000",
  6583=>"000011000",
  6584=>"000001000",
  6585=>"101000000",
  6586=>"000110101",
  6587=>"111010001",
  6588=>"001100000",
  6589=>"011110110",
  6590=>"101001000",
  6591=>"010011111",
  6592=>"110010010",
  6593=>"101010101",
  6594=>"000110001",
  6595=>"010011101",
  6596=>"100000000",
  6597=>"000001101",
  6598=>"111101101",
  6599=>"111000010",
  6600=>"110101011",
  6601=>"100001110",
  6602=>"010110010",
  6603=>"110011110",
  6604=>"011110010",
  6605=>"010000100",
  6606=>"011000010",
  6607=>"001000101",
  6608=>"011110011",
  6609=>"001000000",
  6610=>"110010101",
  6611=>"000001110",
  6612=>"000111010",
  6613=>"011111111",
  6614=>"111011110",
  6615=>"000000100",
  6616=>"111011010",
  6617=>"111110101",
  6618=>"111110001",
  6619=>"001000000",
  6620=>"110001100",
  6621=>"110111000",
  6622=>"101011001",
  6623=>"000100101",
  6624=>"001100110",
  6625=>"111000111",
  6626=>"111110010",
  6627=>"111111001",
  6628=>"101110010",
  6629=>"011111110",
  6630=>"001000010",
  6631=>"010101110",
  6632=>"000100101",
  6633=>"110011100",
  6634=>"000010110",
  6635=>"100000100",
  6636=>"010100011",
  6637=>"111110101",
  6638=>"010000010",
  6639=>"111110101",
  6640=>"110111000",
  6641=>"001001110",
  6642=>"000111011",
  6643=>"000001010",
  6644=>"001100011",
  6645=>"111000111",
  6646=>"110001001",
  6647=>"100011000",
  6648=>"001100000",
  6649=>"110100100",
  6650=>"111110111",
  6651=>"000000101",
  6652=>"001010000",
  6653=>"101100101",
  6654=>"111101100",
  6655=>"010110111",
  6656=>"101011110",
  6657=>"001001010",
  6658=>"111011001",
  6659=>"101011010",
  6660=>"010111101",
  6661=>"101100000",
  6662=>"011101110",
  6663=>"110110000",
  6664=>"110100111",
  6665=>"001001101",
  6666=>"000101011",
  6667=>"001101101",
  6668=>"011011001",
  6669=>"110110000",
  6670=>"111101010",
  6671=>"110100011",
  6672=>"011011001",
  6673=>"110110011",
  6674=>"011001110",
  6675=>"111111100",
  6676=>"001101011",
  6677=>"100001010",
  6678=>"110000110",
  6679=>"100011011",
  6680=>"101010101",
  6681=>"110101001",
  6682=>"000101100",
  6683=>"011011001",
  6684=>"110011010",
  6685=>"010100000",
  6686=>"101110100",
  6687=>"110101100",
  6688=>"011011101",
  6689=>"000011010",
  6690=>"000100001",
  6691=>"111100111",
  6692=>"111111001",
  6693=>"100010011",
  6694=>"111001100",
  6695=>"111000010",
  6696=>"010010100",
  6697=>"111101011",
  6698=>"010001010",
  6699=>"101111011",
  6700=>"100111010",
  6701=>"101100110",
  6702=>"110101100",
  6703=>"000011001",
  6704=>"110000101",
  6705=>"110001000",
  6706=>"110100011",
  6707=>"011110010",
  6708=>"000101100",
  6709=>"010110110",
  6710=>"000101101",
  6711=>"000000010",
  6712=>"100000001",
  6713=>"110110111",
  6714=>"101111000",
  6715=>"000100001",
  6716=>"011100010",
  6717=>"110111101",
  6718=>"101010000",
  6719=>"111000010",
  6720=>"100000101",
  6721=>"000111000",
  6722=>"100101111",
  6723=>"111001110",
  6724=>"001000001",
  6725=>"100110100",
  6726=>"011011001",
  6727=>"001101000",
  6728=>"010011010",
  6729=>"101001010",
  6730=>"101001010",
  6731=>"101011000",
  6732=>"111001010",
  6733=>"100000111",
  6734=>"110110101",
  6735=>"010111011",
  6736=>"010110010",
  6737=>"111010011",
  6738=>"001010100",
  6739=>"011001101",
  6740=>"100110100",
  6741=>"000010101",
  6742=>"011001101",
  6743=>"110001100",
  6744=>"011001001",
  6745=>"110010000",
  6746=>"110111100",
  6747=>"000101001",
  6748=>"000010010",
  6749=>"010110001",
  6750=>"010000011",
  6751=>"001010011",
  6752=>"101011110",
  6753=>"110110110",
  6754=>"100111010",
  6755=>"000010010",
  6756=>"101001110",
  6757=>"010101000",
  6758=>"011100110",
  6759=>"011011110",
  6760=>"000000001",
  6761=>"001011101",
  6762=>"000010111",
  6763=>"101101010",
  6764=>"000001110",
  6765=>"100100001",
  6766=>"000011010",
  6767=>"101010001",
  6768=>"110100000",
  6769=>"100110010",
  6770=>"101100111",
  6771=>"110111110",
  6772=>"111010111",
  6773=>"110011001",
  6774=>"000100010",
  6775=>"101001011",
  6776=>"000000101",
  6777=>"000000100",
  6778=>"011111001",
  6779=>"001110011",
  6780=>"000111110",
  6781=>"001100100",
  6782=>"110110010",
  6783=>"111000011",
  6784=>"111011111",
  6785=>"011001011",
  6786=>"101110000",
  6787=>"100001111",
  6788=>"100010000",
  6789=>"010101000",
  6790=>"010111100",
  6791=>"100111111",
  6792=>"001000100",
  6793=>"101010111",
  6794=>"001111011",
  6795=>"110011000",
  6796=>"011110000",
  6797=>"111001000",
  6798=>"100110001",
  6799=>"000010000",
  6800=>"010001110",
  6801=>"010100100",
  6802=>"111111000",
  6803=>"011010100",
  6804=>"000100110",
  6805=>"010011000",
  6806=>"111010100",
  6807=>"000100111",
  6808=>"111000011",
  6809=>"110011011",
  6810=>"111010010",
  6811=>"100000110",
  6812=>"011110001",
  6813=>"011100101",
  6814=>"110011110",
  6815=>"111101000",
  6816=>"011001100",
  6817=>"010100111",
  6818=>"100001111",
  6819=>"110110010",
  6820=>"000010111",
  6821=>"000100001",
  6822=>"000111111",
  6823=>"110000010",
  6824=>"000111001",
  6825=>"110010100",
  6826=>"101001001",
  6827=>"010001010",
  6828=>"011010010",
  6829=>"111001000",
  6830=>"010111101",
  6831=>"111011100",
  6832=>"000001010",
  6833=>"010010010",
  6834=>"000010100",
  6835=>"010101010",
  6836=>"111111001",
  6837=>"101111111",
  6838=>"001011010",
  6839=>"111111111",
  6840=>"001010100",
  6841=>"100101110",
  6842=>"000000001",
  6843=>"111000001",
  6844=>"011111000",
  6845=>"000011001",
  6846=>"001100011",
  6847=>"010000111",
  6848=>"111010011",
  6849=>"101110000",
  6850=>"001011001",
  6851=>"010111010",
  6852=>"011010111",
  6853=>"111000010",
  6854=>"110010111",
  6855=>"001101110",
  6856=>"110110000",
  6857=>"111101111",
  6858=>"110100011",
  6859=>"100000010",
  6860=>"001110101",
  6861=>"000000010",
  6862=>"110011010",
  6863=>"100111111",
  6864=>"100110110",
  6865=>"100011110",
  6866=>"100101010",
  6867=>"011010000",
  6868=>"000101100",
  6869=>"010000110",
  6870=>"110111100",
  6871=>"001101100",
  6872=>"000000111",
  6873=>"111001010",
  6874=>"000111001",
  6875=>"111000111",
  6876=>"001101101",
  6877=>"010100011",
  6878=>"001011000",
  6879=>"011100010",
  6880=>"001000110",
  6881=>"100100100",
  6882=>"100100100",
  6883=>"111010001",
  6884=>"101101000",
  6885=>"111101000",
  6886=>"010010001",
  6887=>"001000100",
  6888=>"101110110",
  6889=>"111101100",
  6890=>"010101001",
  6891=>"101001001",
  6892=>"010010111",
  6893=>"101100110",
  6894=>"001000110",
  6895=>"100110001",
  6896=>"111001101",
  6897=>"011101101",
  6898=>"100001111",
  6899=>"011101000",
  6900=>"100010100",
  6901=>"111011101",
  6902=>"010110011",
  6903=>"001000111",
  6904=>"110011001",
  6905=>"011111000",
  6906=>"110100111",
  6907=>"101000100",
  6908=>"000110100",
  6909=>"111011001",
  6910=>"100000000",
  6911=>"100011111",
  6912=>"110010011",
  6913=>"100000000",
  6914=>"110011011",
  6915=>"001000011",
  6916=>"001000010",
  6917=>"101101001",
  6918=>"011000101",
  6919=>"011111101",
  6920=>"100001001",
  6921=>"100100001",
  6922=>"110111011",
  6923=>"001010111",
  6924=>"010011111",
  6925=>"110011100",
  6926=>"010010000",
  6927=>"010000011",
  6928=>"100001110",
  6929=>"001110110",
  6930=>"110001000",
  6931=>"001010100",
  6932=>"011001110",
  6933=>"010001001",
  6934=>"011010010",
  6935=>"110110100",
  6936=>"010010111",
  6937=>"000100111",
  6938=>"101111111",
  6939=>"010100100",
  6940=>"110010100",
  6941=>"000000100",
  6942=>"000110100",
  6943=>"000011000",
  6944=>"101000000",
  6945=>"000111000",
  6946=>"101010011",
  6947=>"000110011",
  6948=>"001100101",
  6949=>"100101000",
  6950=>"010000010",
  6951=>"011000111",
  6952=>"111100110",
  6953=>"111100101",
  6954=>"010000101",
  6955=>"001100010",
  6956=>"010100010",
  6957=>"101100011",
  6958=>"001111001",
  6959=>"000110000",
  6960=>"000010000",
  6961=>"100000000",
  6962=>"111100001",
  6963=>"100100011",
  6964=>"110111110",
  6965=>"111010111",
  6966=>"111100010",
  6967=>"010101110",
  6968=>"100110000",
  6969=>"011111000",
  6970=>"111110100",
  6971=>"100001011",
  6972=>"011001000",
  6973=>"011000111",
  6974=>"010100011",
  6975=>"110100011",
  6976=>"100010011",
  6977=>"110110111",
  6978=>"001101010",
  6979=>"001001001",
  6980=>"011001010",
  6981=>"101101111",
  6982=>"011011011",
  6983=>"000010110",
  6984=>"111111011",
  6985=>"101110100",
  6986=>"000110111",
  6987=>"110000011",
  6988=>"100101000",
  6989=>"110110000",
  6990=>"001001101",
  6991=>"101101110",
  6992=>"100110110",
  6993=>"011001001",
  6994=>"010100000",
  6995=>"011001000",
  6996=>"100010000",
  6997=>"110110111",
  6998=>"001101010",
  6999=>"010111000",
  7000=>"001011111",
  7001=>"100101001",
  7002=>"110010101",
  7003=>"000110100",
  7004=>"101011110",
  7005=>"010110011",
  7006=>"100011000",
  7007=>"000100000",
  7008=>"000101101",
  7009=>"010001000",
  7010=>"100011111",
  7011=>"010100111",
  7012=>"111000100",
  7013=>"011110001",
  7014=>"110100001",
  7015=>"011110111",
  7016=>"001111111",
  7017=>"111010111",
  7018=>"101101000",
  7019=>"010111101",
  7020=>"100010101",
  7021=>"111011000",
  7022=>"100011111",
  7023=>"111001111",
  7024=>"101101000",
  7025=>"001000011",
  7026=>"111110110",
  7027=>"111011001",
  7028=>"011110001",
  7029=>"110100001",
  7030=>"011101110",
  7031=>"010110100",
  7032=>"110110000",
  7033=>"101010001",
  7034=>"100101011",
  7035=>"000010101",
  7036=>"000000000",
  7037=>"100010010",
  7038=>"100000111",
  7039=>"110001011",
  7040=>"001011100",
  7041=>"000000001",
  7042=>"010001010",
  7043=>"000010110",
  7044=>"010111101",
  7045=>"110100111",
  7046=>"100100100",
  7047=>"011000110",
  7048=>"110000111",
  7049=>"110000101",
  7050=>"000001001",
  7051=>"001010110",
  7052=>"010100000",
  7053=>"010100101",
  7054=>"100011100",
  7055=>"010101011",
  7056=>"010001100",
  7057=>"011101011",
  7058=>"100100000",
  7059=>"101001010",
  7060=>"010110011",
  7061=>"100111111",
  7062=>"111110111",
  7063=>"101110000",
  7064=>"010100001",
  7065=>"111111010",
  7066=>"000111010",
  7067=>"100111010",
  7068=>"010010111",
  7069=>"111111111",
  7070=>"101111011",
  7071=>"010000100",
  7072=>"100110001",
  7073=>"101110110",
  7074=>"111101011",
  7075=>"010000101",
  7076=>"100100000",
  7077=>"101101111",
  7078=>"011100111",
  7079=>"000101110",
  7080=>"011011101",
  7081=>"010000100",
  7082=>"011010011",
  7083=>"011010110",
  7084=>"110010110",
  7085=>"110010110",
  7086=>"101001110",
  7087=>"000000001",
  7088=>"101101101",
  7089=>"010011011",
  7090=>"111010110",
  7091=>"010000000",
  7092=>"101001100",
  7093=>"010000101",
  7094=>"100101010",
  7095=>"100000100",
  7096=>"101001010",
  7097=>"001000110",
  7098=>"101011111",
  7099=>"110000001",
  7100=>"110101001",
  7101=>"101101100",
  7102=>"110111010",
  7103=>"111000000",
  7104=>"110101001",
  7105=>"010101000",
  7106=>"101111000",
  7107=>"110110101",
  7108=>"001011000",
  7109=>"100001111",
  7110=>"100111110",
  7111=>"011001000",
  7112=>"100001100",
  7113=>"000110100",
  7114=>"101011011",
  7115=>"100011111",
  7116=>"110101110",
  7117=>"001000011",
  7118=>"111111011",
  7119=>"111100000",
  7120=>"100011010",
  7121=>"001000011",
  7122=>"101110001",
  7123=>"111000001",
  7124=>"001000110",
  7125=>"010110111",
  7126=>"110001011",
  7127=>"000100010",
  7128=>"001001101",
  7129=>"110100011",
  7130=>"110111100",
  7131=>"011011000",
  7132=>"001000101",
  7133=>"110100001",
  7134=>"011000110",
  7135=>"111001100",
  7136=>"000001000",
  7137=>"100010011",
  7138=>"011111011",
  7139=>"110001010",
  7140=>"000011000",
  7141=>"100111000",
  7142=>"100100100",
  7143=>"010010110",
  7144=>"000111110",
  7145=>"100000011",
  7146=>"000111101",
  7147=>"010111000",
  7148=>"100101011",
  7149=>"110011010",
  7150=>"000100011",
  7151=>"010000100",
  7152=>"001011100",
  7153=>"011100001",
  7154=>"000111100",
  7155=>"000000000",
  7156=>"111000010",
  7157=>"111000011",
  7158=>"000000010",
  7159=>"000111100",
  7160=>"001011111",
  7161=>"100100000",
  7162=>"010110100",
  7163=>"100010110",
  7164=>"001000101",
  7165=>"101000101",
  7166=>"001110101",
  7167=>"001010000",
  7168=>"101001100",
  7169=>"100000011",
  7170=>"010011101",
  7171=>"101010110",
  7172=>"111011110",
  7173=>"110111011",
  7174=>"111111011",
  7175=>"110010001",
  7176=>"010110101",
  7177=>"100010101",
  7178=>"011111000",
  7179=>"001011110",
  7180=>"101110010",
  7181=>"001011111",
  7182=>"000011110",
  7183=>"001000010",
  7184=>"101000110",
  7185=>"100110110",
  7186=>"011110000",
  7187=>"101111100",
  7188=>"001110111",
  7189=>"001000110",
  7190=>"011101001",
  7191=>"111101011",
  7192=>"111001011",
  7193=>"111110001",
  7194=>"111101000",
  7195=>"111000111",
  7196=>"100010001",
  7197=>"110010000",
  7198=>"011010001",
  7199=>"000010001",
  7200=>"111111111",
  7201=>"110001111",
  7202=>"010000100",
  7203=>"110001010",
  7204=>"001001110",
  7205=>"011111111",
  7206=>"000001110",
  7207=>"101110101",
  7208=>"010111011",
  7209=>"000110010",
  7210=>"110001101",
  7211=>"010101111",
  7212=>"100001001",
  7213=>"000101001",
  7214=>"111111111",
  7215=>"101001010",
  7216=>"010010100",
  7217=>"000000000",
  7218=>"111100010",
  7219=>"010000100",
  7220=>"001100100",
  7221=>"001001100",
  7222=>"001001111",
  7223=>"010110001",
  7224=>"000000111",
  7225=>"011011100",
  7226=>"011001011",
  7227=>"101010011",
  7228=>"101001011",
  7229=>"111101100",
  7230=>"001110111",
  7231=>"101111111",
  7232=>"011000111",
  7233=>"101010111",
  7234=>"001000011",
  7235=>"100001100",
  7236=>"000101101",
  7237=>"100101101",
  7238=>"100111010",
  7239=>"011101100",
  7240=>"010011010",
  7241=>"111101101",
  7242=>"111110011",
  7243=>"001010101",
  7244=>"111110000",
  7245=>"001110011",
  7246=>"010110001",
  7247=>"010000101",
  7248=>"110001110",
  7249=>"110101010",
  7250=>"111001110",
  7251=>"110100110",
  7252=>"001101110",
  7253=>"101111010",
  7254=>"101100011",
  7255=>"010101000",
  7256=>"100000011",
  7257=>"010001100",
  7258=>"011111000",
  7259=>"111100110",
  7260=>"011110101",
  7261=>"001011111",
  7262=>"001101100",
  7263=>"101101111",
  7264=>"000100100",
  7265=>"011100001",
  7266=>"110101110",
  7267=>"000001110",
  7268=>"010111111",
  7269=>"001111010",
  7270=>"001011001",
  7271=>"101010001",
  7272=>"011011011",
  7273=>"100100001",
  7274=>"100101010",
  7275=>"111010101",
  7276=>"100010001",
  7277=>"111110000",
  7278=>"110001101",
  7279=>"111101011",
  7280=>"010010001",
  7281=>"001111101",
  7282=>"110101111",
  7283=>"010001111",
  7284=>"001011011",
  7285=>"111000000",
  7286=>"010101000",
  7287=>"011100000",
  7288=>"111000101",
  7289=>"000001001",
  7290=>"000110000",
  7291=>"111100000",
  7292=>"101111111",
  7293=>"010011110",
  7294=>"111001111",
  7295=>"100101010",
  7296=>"000001101",
  7297=>"000110011",
  7298=>"110101011",
  7299=>"101100100",
  7300=>"010011000",
  7301=>"100000100",
  7302=>"100011111",
  7303=>"100000100",
  7304=>"000111000",
  7305=>"110000100",
  7306=>"001010110",
  7307=>"001111001",
  7308=>"010010110",
  7309=>"011000000",
  7310=>"011011111",
  7311=>"011111000",
  7312=>"000101011",
  7313=>"110010100",
  7314=>"111000000",
  7315=>"111001010",
  7316=>"111010011",
  7317=>"101111001",
  7318=>"111001011",
  7319=>"110000110",
  7320=>"111100100",
  7321=>"110001110",
  7322=>"011111011",
  7323=>"100100001",
  7324=>"100110011",
  7325=>"110110010",
  7326=>"100101100",
  7327=>"011101100",
  7328=>"000001111",
  7329=>"101111110",
  7330=>"100101101",
  7331=>"001100110",
  7332=>"110001110",
  7333=>"110111101",
  7334=>"110001111",
  7335=>"001110111",
  7336=>"001110101",
  7337=>"000000010",
  7338=>"111011000",
  7339=>"000010111",
  7340=>"110110111",
  7341=>"101101010",
  7342=>"011000001",
  7343=>"110111100",
  7344=>"010000100",
  7345=>"100101010",
  7346=>"101001111",
  7347=>"011011000",
  7348=>"110001000",
  7349=>"101010100",
  7350=>"111101110",
  7351=>"010000000",
  7352=>"011000010",
  7353=>"000010010",
  7354=>"101001110",
  7355=>"101100011",
  7356=>"111111100",
  7357=>"001011000",
  7358=>"011011000",
  7359=>"010001100",
  7360=>"001111000",
  7361=>"010000001",
  7362=>"000001011",
  7363=>"111011101",
  7364=>"110111001",
  7365=>"000110010",
  7366=>"100111010",
  7367=>"011000000",
  7368=>"001100001",
  7369=>"110001001",
  7370=>"110010110",
  7371=>"001101001",
  7372=>"110001101",
  7373=>"110001110",
  7374=>"111101111",
  7375=>"100111111",
  7376=>"011001000",
  7377=>"010110000",
  7378=>"100110000",
  7379=>"111111100",
  7380=>"000100000",
  7381=>"001101000",
  7382=>"101100000",
  7383=>"000011111",
  7384=>"001100010",
  7385=>"011101000",
  7386=>"001011101",
  7387=>"010101101",
  7388=>"011110101",
  7389=>"001110110",
  7390=>"000000001",
  7391=>"001010100",
  7392=>"011101111",
  7393=>"111111110",
  7394=>"011100001",
  7395=>"110010000",
  7396=>"000111000",
  7397=>"111111000",
  7398=>"101011111",
  7399=>"110110001",
  7400=>"111001101",
  7401=>"110010110",
  7402=>"101111110",
  7403=>"111010000",
  7404=>"001011101",
  7405=>"111101101",
  7406=>"000000110",
  7407=>"001000011",
  7408=>"111101000",
  7409=>"011111100",
  7410=>"100000100",
  7411=>"110101110",
  7412=>"100110000",
  7413=>"010001111",
  7414=>"110111100",
  7415=>"100011110",
  7416=>"111100001",
  7417=>"110011110",
  7418=>"100101010",
  7419=>"100010000",
  7420=>"101001010",
  7421=>"101011111",
  7422=>"010111110",
  7423=>"101000001",
  7424=>"110010010",
  7425=>"101111001",
  7426=>"101101101",
  7427=>"000111010",
  7428=>"001111100",
  7429=>"111101001",
  7430=>"011110011",
  7431=>"111001101",
  7432=>"111111000",
  7433=>"100100100",
  7434=>"001001001",
  7435=>"100110001",
  7436=>"101100010",
  7437=>"011000000",
  7438=>"101111101",
  7439=>"001100100",
  7440=>"100010100",
  7441=>"001100001",
  7442=>"001100101",
  7443=>"111010111",
  7444=>"111110001",
  7445=>"100000001",
  7446=>"101011000",
  7447=>"011100100",
  7448=>"010011100",
  7449=>"011001011",
  7450=>"111101100",
  7451=>"000000010",
  7452=>"000110111",
  7453=>"011111101",
  7454=>"100100101",
  7455=>"011010111",
  7456=>"000000101",
  7457=>"100110100",
  7458=>"101110110",
  7459=>"101111010",
  7460=>"110000111",
  7461=>"000000001",
  7462=>"000101010",
  7463=>"011011011",
  7464=>"110101101",
  7465=>"100110010",
  7466=>"000100101",
  7467=>"111100011",
  7468=>"101101100",
  7469=>"000100010",
  7470=>"001000110",
  7471=>"111110011",
  7472=>"000010000",
  7473=>"111011110",
  7474=>"101001111",
  7475=>"101101111",
  7476=>"100111010",
  7477=>"100000010",
  7478=>"011111010",
  7479=>"001100010",
  7480=>"101010110",
  7481=>"011101010",
  7482=>"101011000",
  7483=>"011000010",
  7484=>"110010100",
  7485=>"010100011",
  7486=>"010011000",
  7487=>"100101001",
  7488=>"000110101",
  7489=>"010101001",
  7490=>"101100011",
  7491=>"000100000",
  7492=>"111011111",
  7493=>"010011011",
  7494=>"011011110",
  7495=>"110000111",
  7496=>"101010010",
  7497=>"101010111",
  7498=>"100100111",
  7499=>"100101000",
  7500=>"000010101",
  7501=>"000100000",
  7502=>"000001111",
  7503=>"001110010",
  7504=>"000001000",
  7505=>"001111111",
  7506=>"101110111",
  7507=>"110100001",
  7508=>"110010101",
  7509=>"001010111",
  7510=>"000010000",
  7511=>"111101100",
  7512=>"000001111",
  7513=>"110110000",
  7514=>"111110101",
  7515=>"000100010",
  7516=>"001101000",
  7517=>"101001110",
  7518=>"001110011",
  7519=>"010101011",
  7520=>"000101000",
  7521=>"011110111",
  7522=>"101111111",
  7523=>"000001001",
  7524=>"101010100",
  7525=>"100101001",
  7526=>"100001110",
  7527=>"000011100",
  7528=>"010111011",
  7529=>"110110111",
  7530=>"001011111",
  7531=>"001111011",
  7532=>"100101111",
  7533=>"000011100",
  7534=>"111010100",
  7535=>"110010000",
  7536=>"001110111",
  7537=>"011100110",
  7538=>"111000001",
  7539=>"010010001",
  7540=>"011101110",
  7541=>"101001100",
  7542=>"001010000",
  7543=>"100100000",
  7544=>"010010010",
  7545=>"110111101",
  7546=>"101110111",
  7547=>"001101111",
  7548=>"010011111",
  7549=>"101100001",
  7550=>"000110001",
  7551=>"000100111",
  7552=>"111111001",
  7553=>"111100100",
  7554=>"111000011",
  7555=>"011011100",
  7556=>"001111101",
  7557=>"000010111",
  7558=>"111000001",
  7559=>"110001111",
  7560=>"111111111",
  7561=>"111100110",
  7562=>"010111011",
  7563=>"111101011",
  7564=>"100100001",
  7565=>"111010011",
  7566=>"010001001",
  7567=>"101100111",
  7568=>"011111011",
  7569=>"100100011",
  7570=>"101100110",
  7571=>"110110011",
  7572=>"101011111",
  7573=>"110001001",
  7574=>"010100000",
  7575=>"111001101",
  7576=>"110010111",
  7577=>"011000111",
  7578=>"111000111",
  7579=>"111101000",
  7580=>"011101000",
  7581=>"110011110",
  7582=>"010001000",
  7583=>"001101111",
  7584=>"111100000",
  7585=>"100011010",
  7586=>"010010101",
  7587=>"000110010",
  7588=>"110011111",
  7589=>"010100000",
  7590=>"011011000",
  7591=>"011111111",
  7592=>"000010100",
  7593=>"001000100",
  7594=>"001110001",
  7595=>"101011111",
  7596=>"000001011",
  7597=>"100110111",
  7598=>"000010111",
  7599=>"101010000",
  7600=>"000010010",
  7601=>"010010000",
  7602=>"100101010",
  7603=>"000101111",
  7604=>"001110101",
  7605=>"001000010",
  7606=>"111001110",
  7607=>"001001101",
  7608=>"011010101",
  7609=>"101001111",
  7610=>"101111000",
  7611=>"011000100",
  7612=>"010101110",
  7613=>"011000100",
  7614=>"100010110",
  7615=>"010000110",
  7616=>"010101111",
  7617=>"101111010",
  7618=>"010010000",
  7619=>"110101110",
  7620=>"101111111",
  7621=>"011000100",
  7622=>"110100010",
  7623=>"011001011",
  7624=>"011100010",
  7625=>"101001001",
  7626=>"101101111",
  7627=>"111011101",
  7628=>"111010000",
  7629=>"100010001",
  7630=>"000001100",
  7631=>"101101001",
  7632=>"111100010",
  7633=>"101111111",
  7634=>"110010000",
  7635=>"111001010",
  7636=>"000110011",
  7637=>"111000011",
  7638=>"000111111",
  7639=>"111001011",
  7640=>"011100001",
  7641=>"110000011",
  7642=>"011010110",
  7643=>"111001001",
  7644=>"010100110",
  7645=>"000000101",
  7646=>"001110011",
  7647=>"011100010",
  7648=>"010101111",
  7649=>"110110000",
  7650=>"111011101",
  7651=>"001111000",
  7652=>"011010001",
  7653=>"101111100",
  7654=>"100001000",
  7655=>"001000110",
  7656=>"100101011",
  7657=>"001101110",
  7658=>"010110010",
  7659=>"111110010",
  7660=>"000101001",
  7661=>"010000111",
  7662=>"101111110",
  7663=>"101000001",
  7664=>"011110011",
  7665=>"011001011",
  7666=>"000101100",
  7667=>"110011010",
  7668=>"110011110",
  7669=>"010011000",
  7670=>"001100110",
  7671=>"101011110",
  7672=>"100110101",
  7673=>"010111011",
  7674=>"110000000",
  7675=>"101110010",
  7676=>"110011001",
  7677=>"110000110",
  7678=>"010011010",
  7679=>"011000101",
  7680=>"110111001",
  7681=>"001111110",
  7682=>"001111001",
  7683=>"100101010",
  7684=>"100100001",
  7685=>"100011001",
  7686=>"010010011",
  7687=>"011011110",
  7688=>"010111010",
  7689=>"100110100",
  7690=>"011100110",
  7691=>"001001101",
  7692=>"001001010",
  7693=>"101101101",
  7694=>"100011101",
  7695=>"100000111",
  7696=>"100010110",
  7697=>"000011011",
  7698=>"011101110",
  7699=>"001101101",
  7700=>"110000110",
  7701=>"000001100",
  7702=>"101000100",
  7703=>"110110110",
  7704=>"000110110",
  7705=>"111111000",
  7706=>"100100101",
  7707=>"101010111",
  7708=>"111000001",
  7709=>"110000101",
  7710=>"010011110",
  7711=>"100111100",
  7712=>"001001110",
  7713=>"010100111",
  7714=>"001000001",
  7715=>"100000101",
  7716=>"011011110",
  7717=>"101100001",
  7718=>"100101111",
  7719=>"100101101",
  7720=>"000011000",
  7721=>"100111100",
  7722=>"101001011",
  7723=>"001001111",
  7724=>"000001001",
  7725=>"101111111",
  7726=>"000001111",
  7727=>"001010010",
  7728=>"000000100",
  7729=>"011000101",
  7730=>"000000001",
  7731=>"010011100",
  7732=>"011101001",
  7733=>"101010011",
  7734=>"010100110",
  7735=>"110100111",
  7736=>"000011000",
  7737=>"000110010",
  7738=>"010001100",
  7739=>"011100000",
  7740=>"100011010",
  7741=>"010011100",
  7742=>"110110111",
  7743=>"101110011",
  7744=>"101000110",
  7745=>"000010111",
  7746=>"011101101",
  7747=>"000000001",
  7748=>"010001101",
  7749=>"101101100",
  7750=>"000100011",
  7751=>"110001101",
  7752=>"100111011",
  7753=>"110100000",
  7754=>"000001011",
  7755=>"010011000",
  7756=>"100000100",
  7757=>"100011010",
  7758=>"001101000",
  7759=>"011001111",
  7760=>"100000110",
  7761=>"100100111",
  7762=>"001101001",
  7763=>"001011001",
  7764=>"111100110",
  7765=>"110000011",
  7766=>"101100001",
  7767=>"010101110",
  7768=>"100111101",
  7769=>"001101110",
  7770=>"101100110",
  7771=>"001010110",
  7772=>"100010001",
  7773=>"110000111",
  7774=>"100111101",
  7775=>"110101010",
  7776=>"110010000",
  7777=>"111001100",
  7778=>"001000101",
  7779=>"001111011",
  7780=>"001010000",
  7781=>"110001110",
  7782=>"000110100",
  7783=>"001010101",
  7784=>"000011100",
  7785=>"111111110",
  7786=>"001010011",
  7787=>"001001011",
  7788=>"100001110",
  7789=>"010101001",
  7790=>"010010010",
  7791=>"011010010",
  7792=>"111110110",
  7793=>"101110111",
  7794=>"001011010",
  7795=>"000110011",
  7796=>"101111110",
  7797=>"110110101",
  7798=>"001111101",
  7799=>"000001111",
  7800=>"110100101",
  7801=>"011001110",
  7802=>"000000010",
  7803=>"010101010",
  7804=>"011010111",
  7805=>"110001100",
  7806=>"011010110",
  7807=>"101110111",
  7808=>"111101011",
  7809=>"110101011",
  7810=>"101010101",
  7811=>"100001110",
  7812=>"010001000",
  7813=>"000001001",
  7814=>"000110111",
  7815=>"100100111",
  7816=>"011100100",
  7817=>"001111001",
  7818=>"000010111",
  7819=>"111100011",
  7820=>"111000001",
  7821=>"100010111",
  7822=>"000001101",
  7823=>"011111111",
  7824=>"001110001",
  7825=>"001100011",
  7826=>"000111101",
  7827=>"010011010",
  7828=>"010000101",
  7829=>"001001001",
  7830=>"001101011",
  7831=>"011101101",
  7832=>"001000111",
  7833=>"010010000",
  7834=>"110101011",
  7835=>"000100111",
  7836=>"000000001",
  7837=>"011101101",
  7838=>"110111010",
  7839=>"100010100",
  7840=>"010000111",
  7841=>"010101100",
  7842=>"001110101",
  7843=>"001110110",
  7844=>"100111101",
  7845=>"111101101",
  7846=>"000001100",
  7847=>"101000000",
  7848=>"010000001",
  7849=>"000000000",
  7850=>"001110001",
  7851=>"110010101",
  7852=>"011011010",
  7853=>"001101101",
  7854=>"001101101",
  7855=>"000101001",
  7856=>"001101000",
  7857=>"011110000",
  7858=>"000101011",
  7859=>"111101010",
  7860=>"001101110",
  7861=>"000110011",
  7862=>"111110101",
  7863=>"100110011",
  7864=>"100101001",
  7865=>"111111111",
  7866=>"110000010",
  7867=>"101001110",
  7868=>"001101110",
  7869=>"001000000",
  7870=>"000111101",
  7871=>"110111111",
  7872=>"011010100",
  7873=>"000111110",
  7874=>"111110010",
  7875=>"001100000",
  7876=>"101111001",
  7877=>"101101001",
  7878=>"000001001",
  7879=>"011111001",
  7880=>"111000110",
  7881=>"110001100",
  7882=>"100110001",
  7883=>"110101100",
  7884=>"110010100",
  7885=>"011001101",
  7886=>"000101011",
  7887=>"101001000",
  7888=>"010100011",
  7889=>"101101111",
  7890=>"101001110",
  7891=>"001010101",
  7892=>"100011000",
  7893=>"111101010",
  7894=>"011001111",
  7895=>"110011000",
  7896=>"100100011",
  7897=>"110000000",
  7898=>"001110111",
  7899=>"000010100",
  7900=>"101011110",
  7901=>"110010110",
  7902=>"000110110",
  7903=>"011000010",
  7904=>"001011101",
  7905=>"010001110",
  7906=>"010001010",
  7907=>"011000000",
  7908=>"000100010",
  7909=>"010110100",
  7910=>"101111101",
  7911=>"100110000",
  7912=>"010110000",
  7913=>"010101110",
  7914=>"001000000",
  7915=>"100101001",
  7916=>"001111101",
  7917=>"111100111",
  7918=>"111001000",
  7919=>"100001110",
  7920=>"010100000",
  7921=>"110001101",
  7922=>"001101001",
  7923=>"110011011",
  7924=>"101001001",
  7925=>"001110011",
  7926=>"110011011",
  7927=>"000010010",
  7928=>"001110100",
  7929=>"001001000",
  7930=>"101010001",
  7931=>"011010101",
  7932=>"001111011",
  7933=>"110010011",
  7934=>"011101110",
  7935=>"101010101",
  7936=>"101100101",
  7937=>"100110001",
  7938=>"100010000",
  7939=>"000010000",
  7940=>"101010000",
  7941=>"000000010",
  7942=>"101001011",
  7943=>"100010000",
  7944=>"000100001",
  7945=>"011011010",
  7946=>"101101111",
  7947=>"011000111",
  7948=>"100101011",
  7949=>"010011011",
  7950=>"000110110",
  7951=>"000100100",
  7952=>"110010001",
  7953=>"101101000",
  7954=>"000101000",
  7955=>"000101011",
  7956=>"011100001",
  7957=>"000110111",
  7958=>"111100100",
  7959=>"101100101",
  7960=>"001001101",
  7961=>"011111101",
  7962=>"001000010",
  7963=>"000001011",
  7964=>"110110110",
  7965=>"111111111",
  7966=>"110111110",
  7967=>"111011011",
  7968=>"100111011",
  7969=>"000100001",
  7970=>"010000011",
  7971=>"110101111",
  7972=>"100000100",
  7973=>"100010110",
  7974=>"111110001",
  7975=>"100101111",
  7976=>"001000010",
  7977=>"001110100",
  7978=>"101001001",
  7979=>"010011010",
  7980=>"010101011",
  7981=>"101100001",
  7982=>"000001100",
  7983=>"000110100",
  7984=>"100001101",
  7985=>"010010100",
  7986=>"011000010",
  7987=>"110101010",
  7988=>"100000110",
  7989=>"110011001",
  7990=>"011010111",
  7991=>"010000101",
  7992=>"011010010",
  7993=>"100100010",
  7994=>"101001010",
  7995=>"110110011",
  7996=>"011011100",
  7997=>"011110000",
  7998=>"001001110",
  7999=>"011001011",
  8000=>"110100011",
  8001=>"101000011",
  8002=>"000110100",
  8003=>"010000000",
  8004=>"010110111",
  8005=>"110011111",
  8006=>"001110111",
  8007=>"111010011",
  8008=>"101000111",
  8009=>"010111100",
  8010=>"001111001",
  8011=>"100101010",
  8012=>"001011110",
  8013=>"000000000",
  8014=>"110001101",
  8015=>"100111100",
  8016=>"000000001",
  8017=>"110001010",
  8018=>"010000010",
  8019=>"011111101",
  8020=>"010111010",
  8021=>"000101101",
  8022=>"011100010",
  8023=>"111111110",
  8024=>"111010000",
  8025=>"101101011",
  8026=>"001010001",
  8027=>"101100111",
  8028=>"010010101",
  8029=>"110111101",
  8030=>"100010111",
  8031=>"100111110",
  8032=>"011111010",
  8033=>"101110100",
  8034=>"001001011",
  8035=>"111011100",
  8036=>"011100001",
  8037=>"111101001",
  8038=>"011010110",
  8039=>"111010000",
  8040=>"011001011",
  8041=>"010100101",
  8042=>"001010110",
  8043=>"110110011",
  8044=>"000100110",
  8045=>"001001101",
  8046=>"001000110",
  8047=>"000100111",
  8048=>"010100000",
  8049=>"001101001",
  8050=>"000100111",
  8051=>"011110010",
  8052=>"010101010",
  8053=>"101011111",
  8054=>"100101001",
  8055=>"110110000",
  8056=>"000000110",
  8057=>"101101011",
  8058=>"110100000",
  8059=>"111010101",
  8060=>"110010010",
  8061=>"010111010",
  8062=>"111110011",
  8063=>"101001001",
  8064=>"110100001",
  8065=>"000010110",
  8066=>"000000011",
  8067=>"100010010",
  8068=>"010110001",
  8069=>"101101100",
  8070=>"111000001",
  8071=>"000000000",
  8072=>"110001000",
  8073=>"000011010",
  8074=>"010100011",
  8075=>"101110001",
  8076=>"000010111",
  8077=>"101001101",
  8078=>"011101001",
  8079=>"110101100",
  8080=>"100101101",
  8081=>"011000110",
  8082=>"101111000",
  8083=>"001000100",
  8084=>"000111101",
  8085=>"110000011",
  8086=>"110010101",
  8087=>"001000100",
  8088=>"010100010",
  8089=>"011001001",
  8090=>"100000010",
  8091=>"111101010",
  8092=>"011100101",
  8093=>"010001110",
  8094=>"010001101",
  8095=>"011111011",
  8096=>"000011100",
  8097=>"011111110",
  8098=>"001010100",
  8099=>"001011101",
  8100=>"000010101",
  8101=>"111011110",
  8102=>"000011011",
  8103=>"001101111",
  8104=>"101001100",
  8105=>"101101011",
  8106=>"111111100",
  8107=>"010101111",
  8108=>"001111000",
  8109=>"001000110",
  8110=>"000110011",
  8111=>"110001111",
  8112=>"101000000",
  8113=>"100111011",
  8114=>"111000010",
  8115=>"100000010",
  8116=>"000111100",
  8117=>"101100000",
  8118=>"011101100",
  8119=>"000010100",
  8120=>"000101111",
  8121=>"110001110",
  8122=>"100000000",
  8123=>"111110000",
  8124=>"101011111",
  8125=>"011011101",
  8126=>"111001001",
  8127=>"001101100",
  8128=>"001100010",
  8129=>"010111000",
  8130=>"100001011",
  8131=>"000110001",
  8132=>"010100011",
  8133=>"101111010",
  8134=>"010011010",
  8135=>"111100100",
  8136=>"100100000",
  8137=>"000001000",
  8138=>"000010100",
  8139=>"001101111",
  8140=>"000011110",
  8141=>"000110010",
  8142=>"010111001",
  8143=>"000001000",
  8144=>"111110011",
  8145=>"111011000",
  8146=>"100001011",
  8147=>"110101111",
  8148=>"100111000",
  8149=>"111110110",
  8150=>"101011011",
  8151=>"101001000",
  8152=>"010001010",
  8153=>"110100000",
  8154=>"101000011",
  8155=>"101000111",
  8156=>"111010101",
  8157=>"111010001",
  8158=>"010010101",
  8159=>"100100101",
  8160=>"010110101",
  8161=>"100000011",
  8162=>"100000100",
  8163=>"011011110",
  8164=>"010011100",
  8165=>"001000111",
  8166=>"100101001",
  8167=>"110100011",
  8168=>"000011000",
  8169=>"011000001",
  8170=>"010100000",
  8171=>"001001100",
  8172=>"101110111",
  8173=>"001000001",
  8174=>"100111110",
  8175=>"111001101",
  8176=>"011101000",
  8177=>"000001010",
  8178=>"000001010",
  8179=>"000100000",
  8180=>"011010010",
  8181=>"001100101",
  8182=>"110110100",
  8183=>"001000100",
  8184=>"010000001",
  8185=>"100001111",
  8186=>"110010101",
  8187=>"011011001",
  8188=>"101111101",
  8189=>"101000101",
  8190=>"001101111",
  8191=>"111110011",
  8192=>"000010100",
  8193=>"011101000",
  8194=>"101111000",
  8195=>"100100000",
  8196=>"011101011",
  8197=>"001010100",
  8198=>"000000101",
  8199=>"100001100",
  8200=>"111100000",
  8201=>"001000001",
  8202=>"000100000",
  8203=>"111111001",
  8204=>"100010000",
  8205=>"001100000",
  8206=>"100100111",
  8207=>"010011111",
  8208=>"000001000",
  8209=>"001011111",
  8210=>"101011110",
  8211=>"100110100",
  8212=>"000010110",
  8213=>"110011001",
  8214=>"011011101",
  8215=>"011100001",
  8216=>"101111000",
  8217=>"000100011",
  8218=>"011001001",
  8219=>"001001010",
  8220=>"010100101",
  8221=>"100100011",
  8222=>"100010100",
  8223=>"000010000",
  8224=>"100001110",
  8225=>"110111110",
  8226=>"010101110",
  8227=>"111011000",
  8228=>"011111101",
  8229=>"110111001",
  8230=>"000000100",
  8231=>"110101110",
  8232=>"000111011",
  8233=>"010100001",
  8234=>"001111110",
  8235=>"101110010",
  8236=>"001101110",
  8237=>"001111110",
  8238=>"001100101",
  8239=>"101110100",
  8240=>"000010110",
  8241=>"010100111",
  8242=>"101101110",
  8243=>"011101000",
  8244=>"001000000",
  8245=>"111011001",
  8246=>"111000100",
  8247=>"111010000",
  8248=>"000100000",
  8249=>"000000111",
  8250=>"010101111",
  8251=>"110111001",
  8252=>"111011000",
  8253=>"011000001",
  8254=>"110100101",
  8255=>"100101010",
  8256=>"011000011",
  8257=>"001000100",
  8258=>"100101011",
  8259=>"110100111",
  8260=>"110001000",
  8261=>"101101010",
  8262=>"011111011",
  8263=>"011000011",
  8264=>"010100000",
  8265=>"000000001",
  8266=>"110100000",
  8267=>"101000111",
  8268=>"010111010",
  8269=>"010011100",
  8270=>"011011101",
  8271=>"111100110",
  8272=>"111011011",
  8273=>"010000011",
  8274=>"100111000",
  8275=>"101111110",
  8276=>"101100110",
  8277=>"010000000",
  8278=>"111011101",
  8279=>"001101101",
  8280=>"010001000",
  8281=>"001101000",
  8282=>"000110110",
  8283=>"011010000",
  8284=>"011101011",
  8285=>"100010010",
  8286=>"001000111",
  8287=>"001011101",
  8288=>"011000011",
  8289=>"100100011",
  8290=>"111101000",
  8291=>"010000011",
  8292=>"000011001",
  8293=>"111110000",
  8294=>"111001100",
  8295=>"111000101",
  8296=>"000010001",
  8297=>"110001100",
  8298=>"001010011",
  8299=>"100110110",
  8300=>"001000101",
  8301=>"010100010",
  8302=>"101010111",
  8303=>"101000000",
  8304=>"111000001",
  8305=>"110101011",
  8306=>"110001101",
  8307=>"110011001",
  8308=>"000101010",
  8309=>"011110000",
  8310=>"101101100",
  8311=>"100111110",
  8312=>"000100110",
  8313=>"010100110",
  8314=>"111000011",
  8315=>"010000101",
  8316=>"110000100",
  8317=>"110111010",
  8318=>"000101010",
  8319=>"100000000",
  8320=>"000101101",
  8321=>"111111110",
  8322=>"100011000",
  8323=>"101000010",
  8324=>"001110000",
  8325=>"010010000",
  8326=>"011000000",
  8327=>"111110000",
  8328=>"000001000",
  8329=>"101010101",
  8330=>"100001100",
  8331=>"010100100",
  8332=>"011000011",
  8333=>"000100000",
  8334=>"101011101",
  8335=>"111001101",
  8336=>"110110101",
  8337=>"010001000",
  8338=>"010010010",
  8339=>"111010101",
  8340=>"111011101",
  8341=>"100100000",
  8342=>"001100010",
  8343=>"101010001",
  8344=>"110011011",
  8345=>"110110011",
  8346=>"001010110",
  8347=>"110111000",
  8348=>"101111110",
  8349=>"100000110",
  8350=>"101000000",
  8351=>"000100110",
  8352=>"010101100",
  8353=>"011110010",
  8354=>"100101010",
  8355=>"100111001",
  8356=>"001001101",
  8357=>"101001100",
  8358=>"110110111",
  8359=>"010010111",
  8360=>"111000101",
  8361=>"010001001",
  8362=>"000110000",
  8363=>"011000100",
  8364=>"000100101",
  8365=>"000010011",
  8366=>"010000000",
  8367=>"101001111",
  8368=>"111100101",
  8369=>"101110100",
  8370=>"010000110",
  8371=>"000101111",
  8372=>"101000110",
  8373=>"110101011",
  8374=>"001101011",
  8375=>"001100101",
  8376=>"000011111",
  8377=>"111100110",
  8378=>"000111101",
  8379=>"000100010",
  8380=>"111001101",
  8381=>"011011110",
  8382=>"001001001",
  8383=>"000101100",
  8384=>"001000110",
  8385=>"100111110",
  8386=>"000001111",
  8387=>"101100000",
  8388=>"011010000",
  8389=>"111001110",
  8390=>"000110100",
  8391=>"100001010",
  8392=>"010010011",
  8393=>"000100110",
  8394=>"111001011",
  8395=>"011000110",
  8396=>"000110001",
  8397=>"111100110",
  8398=>"010000000",
  8399=>"111111111",
  8400=>"000011111",
  8401=>"100010110",
  8402=>"100000101",
  8403=>"100110110",
  8404=>"111110111",
  8405=>"011110001",
  8406=>"101011010",
  8407=>"100111100",
  8408=>"000100001",
  8409=>"101111111",
  8410=>"000110010",
  8411=>"111010101",
  8412=>"111100110",
  8413=>"100010100",
  8414=>"000101000",
  8415=>"100111111",
  8416=>"111111100",
  8417=>"000011010",
  8418=>"001101110",
  8419=>"100011110",
  8420=>"010111001",
  8421=>"011011110",
  8422=>"111000011",
  8423=>"101101111",
  8424=>"101001100",
  8425=>"100100001",
  8426=>"000011001",
  8427=>"111011000",
  8428=>"111100010",
  8429=>"000011001",
  8430=>"000000001",
  8431=>"101111101",
  8432=>"111011110",
  8433=>"111111111",
  8434=>"100000010",
  8435=>"100111111",
  8436=>"000011100",
  8437=>"001010101",
  8438=>"010000110",
  8439=>"011010001",
  8440=>"000010010",
  8441=>"110011111",
  8442=>"101010110",
  8443=>"100110101",
  8444=>"011100110",
  8445=>"111000101",
  8446=>"001000100",
  8447=>"101100110",
  8448=>"010001101",
  8449=>"000100101",
  8450=>"101101010",
  8451=>"110111010",
  8452=>"111011111",
  8453=>"000111111",
  8454=>"011100100",
  8455=>"000111001",
  8456=>"101100101",
  8457=>"010001110",
  8458=>"101101111",
  8459=>"101110110",
  8460=>"001110100",
  8461=>"110010100",
  8462=>"000000000",
  8463=>"010010110",
  8464=>"010101000",
  8465=>"001110110",
  8466=>"011101011",
  8467=>"111111100",
  8468=>"001000011",
  8469=>"010110000",
  8470=>"111110100",
  8471=>"111001110",
  8472=>"110111000",
  8473=>"000101111",
  8474=>"010000100",
  8475=>"101101111",
  8476=>"111000101",
  8477=>"000110010",
  8478=>"011010001",
  8479=>"111000100",
  8480=>"001100100",
  8481=>"000101000",
  8482=>"010011110",
  8483=>"011111010",
  8484=>"101110101",
  8485=>"100100011",
  8486=>"111000000",
  8487=>"111001001",
  8488=>"011100000",
  8489=>"010010101",
  8490=>"001110011",
  8491=>"010010011",
  8492=>"011000010",
  8493=>"000100111",
  8494=>"111010101",
  8495=>"100100001",
  8496=>"101000101",
  8497=>"111000011",
  8498=>"001000000",
  8499=>"011101010",
  8500=>"100001000",
  8501=>"000000000",
  8502=>"101111010",
  8503=>"011111111",
  8504=>"001000000",
  8505=>"110011000",
  8506=>"110100111",
  8507=>"001001111",
  8508=>"111010010",
  8509=>"111000111",
  8510=>"100000110",
  8511=>"000010110",
  8512=>"001100011",
  8513=>"100110011",
  8514=>"110001101",
  8515=>"101001110",
  8516=>"111101001",
  8517=>"101000101",
  8518=>"101010000",
  8519=>"000001000",
  8520=>"100011000",
  8521=>"010100110",
  8522=>"111111001",
  8523=>"000000110",
  8524=>"010000000",
  8525=>"100001101",
  8526=>"111010000",
  8527=>"110101010",
  8528=>"001111111",
  8529=>"110111101",
  8530=>"101101001",
  8531=>"101010101",
  8532=>"011100000",
  8533=>"010101100",
  8534=>"010010011",
  8535=>"001110000",
  8536=>"111110001",
  8537=>"000001010",
  8538=>"000010011",
  8539=>"101000011",
  8540=>"000100001",
  8541=>"011101111",
  8542=>"001001101",
  8543=>"111111010",
  8544=>"000001000",
  8545=>"011001101",
  8546=>"100111111",
  8547=>"000001001",
  8548=>"111111001",
  8549=>"010010010",
  8550=>"101111000",
  8551=>"100100101",
  8552=>"110110101",
  8553=>"000011011",
  8554=>"101110010",
  8555=>"010001110",
  8556=>"001000011",
  8557=>"101101101",
  8558=>"100111001",
  8559=>"111001010",
  8560=>"000000111",
  8561=>"000101011",
  8562=>"100100010",
  8563=>"111001101",
  8564=>"010010001",
  8565=>"011001001",
  8566=>"101101001",
  8567=>"101001100",
  8568=>"000010100",
  8569=>"111100010",
  8570=>"100001011",
  8571=>"110001111",
  8572=>"111000010",
  8573=>"000001111",
  8574=>"010011010",
  8575=>"100001000",
  8576=>"000110111",
  8577=>"000011000",
  8578=>"000111001",
  8579=>"010111101",
  8580=>"100011001",
  8581=>"010100010",
  8582=>"100001100",
  8583=>"110010011",
  8584=>"100011000",
  8585=>"100110110",
  8586=>"011101100",
  8587=>"010110101",
  8588=>"110100110",
  8589=>"111000010",
  8590=>"100101101",
  8591=>"010011000",
  8592=>"100101100",
  8593=>"001000111",
  8594=>"101101110",
  8595=>"111101111",
  8596=>"100111110",
  8597=>"010110100",
  8598=>"101110000",
  8599=>"100111110",
  8600=>"110110011",
  8601=>"000010111",
  8602=>"010001101",
  8603=>"111010110",
  8604=>"011110100",
  8605=>"011011100",
  8606=>"010100111",
  8607=>"100101001",
  8608=>"101101111",
  8609=>"001001001",
  8610=>"010011101",
  8611=>"001110011",
  8612=>"000010011",
  8613=>"100010001",
  8614=>"000111100",
  8615=>"100101101",
  8616=>"010001010",
  8617=>"111001100",
  8618=>"001001001",
  8619=>"000110010",
  8620=>"111001110",
  8621=>"100111100",
  8622=>"101110011",
  8623=>"000100100",
  8624=>"001000000",
  8625=>"101001111",
  8626=>"101010000",
  8627=>"001001010",
  8628=>"010101101",
  8629=>"100001111",
  8630=>"100001111",
  8631=>"011100100",
  8632=>"010110101",
  8633=>"110101011",
  8634=>"000000000",
  8635=>"010000110",
  8636=>"110111101",
  8637=>"000011111",
  8638=>"111111101",
  8639=>"111011000",
  8640=>"010101010",
  8641=>"110100101",
  8642=>"111111000",
  8643=>"110111010",
  8644=>"000110100",
  8645=>"001110100",
  8646=>"010001101",
  8647=>"111101000",
  8648=>"000001101",
  8649=>"100101010",
  8650=>"001111000",
  8651=>"110100100",
  8652=>"101011011",
  8653=>"011011111",
  8654=>"010011111",
  8655=>"100011010",
  8656=>"111111001",
  8657=>"010100100",
  8658=>"110111100",
  8659=>"010011101",
  8660=>"101011100",
  8661=>"000001000",
  8662=>"100110111",
  8663=>"010011110",
  8664=>"001001100",
  8665=>"101010011",
  8666=>"001011000",
  8667=>"010101110",
  8668=>"110001101",
  8669=>"100101111",
  8670=>"101111010",
  8671=>"100011101",
  8672=>"101101010",
  8673=>"110000001",
  8674=>"100011000",
  8675=>"011001101",
  8676=>"101001011",
  8677=>"111011110",
  8678=>"111011011",
  8679=>"010000101",
  8680=>"011000100",
  8681=>"101010101",
  8682=>"000000111",
  8683=>"000011111",
  8684=>"010100001",
  8685=>"001010100",
  8686=>"100011110",
  8687=>"000001000",
  8688=>"001110110",
  8689=>"011101110",
  8690=>"001101000",
  8691=>"000001111",
  8692=>"100000101",
  8693=>"000000011",
  8694=>"111011101",
  8695=>"110011110",
  8696=>"000000001",
  8697=>"100011110",
  8698=>"011100000",
  8699=>"010110111",
  8700=>"100010110",
  8701=>"000101001",
  8702=>"110011001",
  8703=>"111111100",
  8704=>"011001000",
  8705=>"111100010",
  8706=>"001000100",
  8707=>"000100101",
  8708=>"011111111",
  8709=>"111101100",
  8710=>"000110111",
  8711=>"101001010",
  8712=>"101001010",
  8713=>"011000001",
  8714=>"100100110",
  8715=>"011011000",
  8716=>"000110101",
  8717=>"101000110",
  8718=>"101001010",
  8719=>"111011101",
  8720=>"101010001",
  8721=>"000001010",
  8722=>"110111010",
  8723=>"001110011",
  8724=>"110000110",
  8725=>"111001010",
  8726=>"010111111",
  8727=>"100010110",
  8728=>"010100001",
  8729=>"010110110",
  8730=>"001001111",
  8731=>"100001111",
  8732=>"110111001",
  8733=>"000001111",
  8734=>"110000011",
  8735=>"001100010",
  8736=>"101011101",
  8737=>"010110111",
  8738=>"010011010",
  8739=>"000000010",
  8740=>"000110101",
  8741=>"001011100",
  8742=>"100100111",
  8743=>"111000111",
  8744=>"101110011",
  8745=>"100100011",
  8746=>"010110000",
  8747=>"010111101",
  8748=>"111100111",
  8749=>"000111001",
  8750=>"001010110",
  8751=>"011011000",
  8752=>"000111011",
  8753=>"011101110",
  8754=>"100110001",
  8755=>"000011000",
  8756=>"111010111",
  8757=>"100111001",
  8758=>"111000001",
  8759=>"110110111",
  8760=>"110011111",
  8761=>"100010110",
  8762=>"001111010",
  8763=>"011011011",
  8764=>"100111110",
  8765=>"010010011",
  8766=>"101101001",
  8767=>"111001101",
  8768=>"001101111",
  8769=>"001111110",
  8770=>"000000010",
  8771=>"111001010",
  8772=>"011110001",
  8773=>"101110011",
  8774=>"001110000",
  8775=>"000111011",
  8776=>"100000000",
  8777=>"100000001",
  8778=>"101110101",
  8779=>"111011000",
  8780=>"000100011",
  8781=>"010000011",
  8782=>"001011110",
  8783=>"000011110",
  8784=>"011011011",
  8785=>"011000010",
  8786=>"100010101",
  8787=>"000101001",
  8788=>"011001111",
  8789=>"110011011",
  8790=>"111111000",
  8791=>"100000000",
  8792=>"110111011",
  8793=>"010110011",
  8794=>"010010101",
  8795=>"110111101",
  8796=>"001110111",
  8797=>"001101100",
  8798=>"000101100",
  8799=>"010001110",
  8800=>"110100101",
  8801=>"000001001",
  8802=>"011001111",
  8803=>"101001001",
  8804=>"100000111",
  8805=>"100000000",
  8806=>"100101100",
  8807=>"011001110",
  8808=>"000010010",
  8809=>"001110110",
  8810=>"100111101",
  8811=>"010011110",
  8812=>"111111000",
  8813=>"000101100",
  8814=>"010011000",
  8815=>"010111101",
  8816=>"110010001",
  8817=>"000001010",
  8818=>"000111100",
  8819=>"010001011",
  8820=>"000011111",
  8821=>"000000010",
  8822=>"011100001",
  8823=>"011001111",
  8824=>"101111011",
  8825=>"011101011",
  8826=>"101100001",
  8827=>"100000111",
  8828=>"111100011",
  8829=>"001001111",
  8830=>"111010100",
  8831=>"100111001",
  8832=>"001000100",
  8833=>"110010001",
  8834=>"111001101",
  8835=>"100110001",
  8836=>"101011001",
  8837=>"011000110",
  8838=>"111011101",
  8839=>"100110101",
  8840=>"001110100",
  8841=>"010000111",
  8842=>"000000100",
  8843=>"100011011",
  8844=>"111011111",
  8845=>"111101111",
  8846=>"011010011",
  8847=>"000110011",
  8848=>"101010100",
  8849=>"101001100",
  8850=>"100100000",
  8851=>"011001101",
  8852=>"001010100",
  8853=>"111111100",
  8854=>"011001100",
  8855=>"101001001",
  8856=>"001111010",
  8857=>"000010100",
  8858=>"100010100",
  8859=>"111111001",
  8860=>"100011101",
  8861=>"111110110",
  8862=>"000001011",
  8863=>"110111011",
  8864=>"101110100",
  8865=>"100101011",
  8866=>"010010001",
  8867=>"101000101",
  8868=>"011111111",
  8869=>"110111000",
  8870=>"001010000",
  8871=>"010010001",
  8872=>"110111101",
  8873=>"001110001",
  8874=>"101100010",
  8875=>"001111100",
  8876=>"110001011",
  8877=>"001010011",
  8878=>"100000100",
  8879=>"110100001",
  8880=>"010001011",
  8881=>"011101001",
  8882=>"000101011",
  8883=>"000101000",
  8884=>"011011111",
  8885=>"100111101",
  8886=>"100011010",
  8887=>"001000111",
  8888=>"001001111",
  8889=>"000111010",
  8890=>"000010111",
  8891=>"100111001",
  8892=>"010010010",
  8893=>"000100011",
  8894=>"000011101",
  8895=>"011001101",
  8896=>"000111110",
  8897=>"011101000",
  8898=>"101110111",
  8899=>"110101110",
  8900=>"100111000",
  8901=>"001011010",
  8902=>"000111111",
  8903=>"101000010",
  8904=>"011001001",
  8905=>"101010001",
  8906=>"111111001",
  8907=>"101110011",
  8908=>"001011001",
  8909=>"000000101",
  8910=>"000010000",
  8911=>"010000110",
  8912=>"100000011",
  8913=>"001010100",
  8914=>"000010010",
  8915=>"000101010",
  8916=>"100010000",
  8917=>"111110000",
  8918=>"000101100",
  8919=>"101011001",
  8920=>"101010110",
  8921=>"010101110",
  8922=>"000110010",
  8923=>"000110010",
  8924=>"010010100",
  8925=>"101110100",
  8926=>"110110011",
  8927=>"101001111",
  8928=>"000001111",
  8929=>"000000000",
  8930=>"011010001",
  8931=>"111100001",
  8932=>"101101110",
  8933=>"101110110",
  8934=>"110111001",
  8935=>"000000010",
  8936=>"000101001",
  8937=>"101110100",
  8938=>"101000000",
  8939=>"010100001",
  8940=>"000010010",
  8941=>"101100111",
  8942=>"000110011",
  8943=>"100110011",
  8944=>"000111110",
  8945=>"101000100",
  8946=>"110000000",
  8947=>"101011110",
  8948=>"100111100",
  8949=>"000011000",
  8950=>"111100001",
  8951=>"000010111",
  8952=>"011011101",
  8953=>"001010111",
  8954=>"100110010",
  8955=>"010001101",
  8956=>"001011101",
  8957=>"010110111",
  8958=>"110000011",
  8959=>"010100100",
  8960=>"100000110",
  8961=>"001000100",
  8962=>"011000011",
  8963=>"000101100",
  8964=>"010010101",
  8965=>"100110000",
  8966=>"110101010",
  8967=>"011000010",
  8968=>"100110101",
  8969=>"010010010",
  8970=>"010001101",
  8971=>"000001111",
  8972=>"001011010",
  8973=>"000100010",
  8974=>"100101011",
  8975=>"100001100",
  8976=>"110111000",
  8977=>"000000001",
  8978=>"000101000",
  8979=>"001111010",
  8980=>"101001100",
  8981=>"110011110",
  8982=>"101001101",
  8983=>"101011011",
  8984=>"101100001",
  8985=>"001001100",
  8986=>"100001000",
  8987=>"010001011",
  8988=>"100101101",
  8989=>"000000110",
  8990=>"100111101",
  8991=>"111011001",
  8992=>"110110111",
  8993=>"111011000",
  8994=>"000010101",
  8995=>"000101011",
  8996=>"011011111",
  8997=>"100001111",
  8998=>"011010110",
  8999=>"001110011",
  9000=>"001001110",
  9001=>"000001100",
  9002=>"111011111",
  9003=>"101011110",
  9004=>"101000011",
  9005=>"000001111",
  9006=>"101011111",
  9007=>"110111110",
  9008=>"001101000",
  9009=>"000110111",
  9010=>"101001011",
  9011=>"010000110",
  9012=>"111111010",
  9013=>"110101001",
  9014=>"000110010",
  9015=>"010110100",
  9016=>"100000111",
  9017=>"111101101",
  9018=>"001000011",
  9019=>"000101100",
  9020=>"011000111",
  9021=>"010011101",
  9022=>"001000110",
  9023=>"111111100",
  9024=>"011001001",
  9025=>"101100011",
  9026=>"111111011",
  9027=>"100100100",
  9028=>"111001000",
  9029=>"100110001",
  9030=>"000101001",
  9031=>"111001101",
  9032=>"011100110",
  9033=>"001100000",
  9034=>"100000000",
  9035=>"011000010",
  9036=>"110111010",
  9037=>"000000101",
  9038=>"101000000",
  9039=>"010110000",
  9040=>"111110011",
  9041=>"101000100",
  9042=>"001100000",
  9043=>"001000010",
  9044=>"010001111",
  9045=>"000000100",
  9046=>"100101111",
  9047=>"100100011",
  9048=>"010111010",
  9049=>"010010111",
  9050=>"000101000",
  9051=>"101111111",
  9052=>"110110101",
  9053=>"111001110",
  9054=>"110100110",
  9055=>"000111011",
  9056=>"011011101",
  9057=>"000000101",
  9058=>"000001110",
  9059=>"111001000",
  9060=>"011001111",
  9061=>"000110111",
  9062=>"100000001",
  9063=>"111001011",
  9064=>"000101101",
  9065=>"010110111",
  9066=>"000111101",
  9067=>"000011110",
  9068=>"000001001",
  9069=>"101111100",
  9070=>"101100000",
  9071=>"101101011",
  9072=>"010101000",
  9073=>"100000111",
  9074=>"100101010",
  9075=>"100011100",
  9076=>"011100110",
  9077=>"000110010",
  9078=>"000111000",
  9079=>"111001111",
  9080=>"100011110",
  9081=>"011100001",
  9082=>"000011011",
  9083=>"111000011",
  9084=>"000001110",
  9085=>"110111100",
  9086=>"100010011",
  9087=>"001000001",
  9088=>"010010001",
  9089=>"011110111",
  9090=>"111110001",
  9091=>"001000110",
  9092=>"100100001",
  9093=>"111001011",
  9094=>"100100010",
  9095=>"010111100",
  9096=>"111010001",
  9097=>"101111100",
  9098=>"000001100",
  9099=>"111110111",
  9100=>"100000010",
  9101=>"101000111",
  9102=>"110000110",
  9103=>"100110100",
  9104=>"100101100",
  9105=>"111010110",
  9106=>"000000101",
  9107=>"101000001",
  9108=>"010000000",
  9109=>"100111111",
  9110=>"000101101",
  9111=>"111100101",
  9112=>"110001001",
  9113=>"000110100",
  9114=>"111011101",
  9115=>"000101100",
  9116=>"110011100",
  9117=>"000011011",
  9118=>"100100000",
  9119=>"111010001",
  9120=>"101111001",
  9121=>"011111100",
  9122=>"000100000",
  9123=>"000000111",
  9124=>"110011110",
  9125=>"011100001",
  9126=>"110100001",
  9127=>"000010000",
  9128=>"001011111",
  9129=>"111111101",
  9130=>"011111011",
  9131=>"010100100",
  9132=>"001001011",
  9133=>"011010011",
  9134=>"001111011",
  9135=>"100010011",
  9136=>"111000010",
  9137=>"110110011",
  9138=>"100010101",
  9139=>"001101010",
  9140=>"101111100",
  9141=>"010110010",
  9142=>"110111001",
  9143=>"011000000",
  9144=>"111000110",
  9145=>"101110001",
  9146=>"110111000",
  9147=>"100100010",
  9148=>"100100000",
  9149=>"001000001",
  9150=>"111100011",
  9151=>"000000100",
  9152=>"011001101",
  9153=>"001010010",
  9154=>"000110001",
  9155=>"100001101",
  9156=>"111011100",
  9157=>"100010010",
  9158=>"110000000",
  9159=>"010001111",
  9160=>"001000000",
  9161=>"011101111",
  9162=>"110010011",
  9163=>"111111000",
  9164=>"001011000",
  9165=>"101000011",
  9166=>"111110101",
  9167=>"100100110",
  9168=>"010010001",
  9169=>"000000001",
  9170=>"111111101",
  9171=>"110100011",
  9172=>"010001111",
  9173=>"111001011",
  9174=>"000010110",
  9175=>"010100010",
  9176=>"100000111",
  9177=>"110111101",
  9178=>"101000011",
  9179=>"000100000",
  9180=>"101111110",
  9181=>"110111111",
  9182=>"001111100",
  9183=>"111001001",
  9184=>"111110000",
  9185=>"101000001",
  9186=>"110010101",
  9187=>"101101100",
  9188=>"011101010",
  9189=>"010001001",
  9190=>"001000000",
  9191=>"010100010",
  9192=>"000000111",
  9193=>"011011011",
  9194=>"001001010",
  9195=>"001101110",
  9196=>"001111010",
  9197=>"010100111",
  9198=>"000101111",
  9199=>"010111110",
  9200=>"100100000",
  9201=>"010100000",
  9202=>"110000000",
  9203=>"100100001",
  9204=>"000010101",
  9205=>"100000101",
  9206=>"101000010",
  9207=>"011000000",
  9208=>"101000001",
  9209=>"001001001",
  9210=>"000110100",
  9211=>"010010110",
  9212=>"111001010",
  9213=>"010101000",
  9214=>"110001000",
  9215=>"001011000",
  9216=>"010100100",
  9217=>"001000001",
  9218=>"011001011",
  9219=>"000010000",
  9220=>"111011110",
  9221=>"100101010",
  9222=>"111111001",
  9223=>"011100000",
  9224=>"011010000",
  9225=>"000001011",
  9226=>"011101011",
  9227=>"100001000",
  9228=>"011101100",
  9229=>"011011010",
  9230=>"101100100",
  9231=>"100000100",
  9232=>"111100110",
  9233=>"101101110",
  9234=>"110100011",
  9235=>"011101001",
  9236=>"101111010",
  9237=>"000110111",
  9238=>"010100111",
  9239=>"001010001",
  9240=>"010001110",
  9241=>"100100101",
  9242=>"100011010",
  9243=>"001001110",
  9244=>"111000111",
  9245=>"111010001",
  9246=>"000001001",
  9247=>"100101100",
  9248=>"110011001",
  9249=>"001010100",
  9250=>"001110010",
  9251=>"001101000",
  9252=>"110100000",
  9253=>"110001111",
  9254=>"101110110",
  9255=>"011011101",
  9256=>"111011001",
  9257=>"111100101",
  9258=>"011110001",
  9259=>"100001011",
  9260=>"110001000",
  9261=>"110011001",
  9262=>"011000011",
  9263=>"101000110",
  9264=>"101110001",
  9265=>"001111111",
  9266=>"011111010",
  9267=>"110110110",
  9268=>"110111010",
  9269=>"000000101",
  9270=>"000100111",
  9271=>"011110000",
  9272=>"100101111",
  9273=>"110011101",
  9274=>"101001101",
  9275=>"000110111",
  9276=>"001010100",
  9277=>"000000011",
  9278=>"101111111",
  9279=>"000010000",
  9280=>"100110110",
  9281=>"110001011",
  9282=>"010101001",
  9283=>"000010101",
  9284=>"101010110",
  9285=>"000001001",
  9286=>"000111000",
  9287=>"011000111",
  9288=>"110011011",
  9289=>"101110001",
  9290=>"001011000",
  9291=>"010011111",
  9292=>"001001100",
  9293=>"101001011",
  9294=>"101011011",
  9295=>"101011111",
  9296=>"111100001",
  9297=>"000001100",
  9298=>"010001111",
  9299=>"010000001",
  9300=>"000011110",
  9301=>"111001100",
  9302=>"000111000",
  9303=>"001010001",
  9304=>"001110100",
  9305=>"011000001",
  9306=>"011001111",
  9307=>"100000000",
  9308=>"111011000",
  9309=>"011110010",
  9310=>"010000101",
  9311=>"010000000",
  9312=>"000111000",
  9313=>"010100111",
  9314=>"001100011",
  9315=>"010001000",
  9316=>"011101011",
  9317=>"010110010",
  9318=>"111101100",
  9319=>"011100001",
  9320=>"000100011",
  9321=>"001100111",
  9322=>"110010110",
  9323=>"000101001",
  9324=>"001001100",
  9325=>"011011010",
  9326=>"010110001",
  9327=>"100110001",
  9328=>"100111000",
  9329=>"010001110",
  9330=>"000000010",
  9331=>"100110100",
  9332=>"110001010",
  9333=>"111010100",
  9334=>"110111000",
  9335=>"000110001",
  9336=>"000001001",
  9337=>"000011011",
  9338=>"111000000",
  9339=>"000101011",
  9340=>"010010000",
  9341=>"111101001",
  9342=>"110111111",
  9343=>"011010011",
  9344=>"001010001",
  9345=>"110101101",
  9346=>"000000001",
  9347=>"111100101",
  9348=>"011111100",
  9349=>"101001110",
  9350=>"001000101",
  9351=>"001111110",
  9352=>"101000111",
  9353=>"000000100",
  9354=>"000100001",
  9355=>"000011011",
  9356=>"000100010",
  9357=>"011111001",
  9358=>"011011000",
  9359=>"100101100",
  9360=>"010001110",
  9361=>"101001011",
  9362=>"111010100",
  9363=>"000010000",
  9364=>"000100101",
  9365=>"100000010",
  9366=>"001101011",
  9367=>"001011011",
  9368=>"110001101",
  9369=>"110010111",
  9370=>"111000100",
  9371=>"111010010",
  9372=>"011101011",
  9373=>"000011011",
  9374=>"000000001",
  9375=>"101000001",
  9376=>"100011101",
  9377=>"101001111",
  9378=>"100110010",
  9379=>"010001111",
  9380=>"101111000",
  9381=>"110010111",
  9382=>"101010001",
  9383=>"011110111",
  9384=>"000000010",
  9385=>"100001111",
  9386=>"111101000",
  9387=>"111111101",
  9388=>"110100000",
  9389=>"101001010",
  9390=>"000010100",
  9391=>"011110011",
  9392=>"100011011",
  9393=>"000100010",
  9394=>"000100000",
  9395=>"101000101",
  9396=>"001101100",
  9397=>"001011100",
  9398=>"100101111",
  9399=>"100001101",
  9400=>"101110011",
  9401=>"011001110",
  9402=>"101000101",
  9403=>"100010000",
  9404=>"110011101",
  9405=>"101000110",
  9406=>"011001000",
  9407=>"111101110",
  9408=>"000001010",
  9409=>"000111010",
  9410=>"111011101",
  9411=>"011100101",
  9412=>"110101010",
  9413=>"101000101",
  9414=>"000111000",
  9415=>"010001101",
  9416=>"001000100",
  9417=>"000111001",
  9418=>"101001011",
  9419=>"000111110",
  9420=>"111111111",
  9421=>"010101111",
  9422=>"010011111",
  9423=>"011010111",
  9424=>"111000000",
  9425=>"001101011",
  9426=>"100100000",
  9427=>"100111000",
  9428=>"001011010",
  9429=>"111110110",
  9430=>"101101111",
  9431=>"111110101",
  9432=>"110110100",
  9433=>"100000010",
  9434=>"000110010",
  9435=>"100010011",
  9436=>"011110110",
  9437=>"001101100",
  9438=>"011010001",
  9439=>"101110011",
  9440=>"001010000",
  9441=>"101001001",
  9442=>"011000111",
  9443=>"010001100",
  9444=>"111001100",
  9445=>"011011011",
  9446=>"000010011",
  9447=>"110101011",
  9448=>"010001100",
  9449=>"000010110",
  9450=>"001110010",
  9451=>"111100001",
  9452=>"000011110",
  9453=>"010000000",
  9454=>"101111111",
  9455=>"110111100",
  9456=>"010101011",
  9457=>"011010010",
  9458=>"101001111",
  9459=>"000000100",
  9460=>"101111101",
  9461=>"100101111",
  9462=>"001011000",
  9463=>"011111001",
  9464=>"011000101",
  9465=>"010001101",
  9466=>"111001100",
  9467=>"110011010",
  9468=>"100000110",
  9469=>"101001000",
  9470=>"000001110",
  9471=>"000011100",
  9472=>"110011101",
  9473=>"000110011",
  9474=>"100010001",
  9475=>"110010111",
  9476=>"011100111",
  9477=>"001110111",
  9478=>"101001010",
  9479=>"100010000",
  9480=>"100111110",
  9481=>"111010000",
  9482=>"010001110",
  9483=>"000111110",
  9484=>"001011010",
  9485=>"000100011",
  9486=>"010110100",
  9487=>"010100001",
  9488=>"101111000",
  9489=>"011011100",
  9490=>"000001010",
  9491=>"111010000",
  9492=>"001000010",
  9493=>"101101111",
  9494=>"101010000",
  9495=>"110011111",
  9496=>"001011110",
  9497=>"100000000",
  9498=>"100110100",
  9499=>"010000110",
  9500=>"101001010",
  9501=>"111101010",
  9502=>"110100111",
  9503=>"000001101",
  9504=>"111010001",
  9505=>"000000101",
  9506=>"000101001",
  9507=>"100100101",
  9508=>"110111010",
  9509=>"000010110",
  9510=>"011010111",
  9511=>"001001010",
  9512=>"001010001",
  9513=>"011100000",
  9514=>"011100000",
  9515=>"111010100",
  9516=>"101100001",
  9517=>"000111110",
  9518=>"110010100",
  9519=>"010110011",
  9520=>"010001001",
  9521=>"010010110",
  9522=>"110100011",
  9523=>"000010101",
  9524=>"101001010",
  9525=>"100101101",
  9526=>"000111101",
  9527=>"111100101",
  9528=>"000101101",
  9529=>"100101000",
  9530=>"110110011",
  9531=>"101011100",
  9532=>"001011001",
  9533=>"100001001",
  9534=>"110001010",
  9535=>"111001101",
  9536=>"010111110",
  9537=>"100001000",
  9538=>"100001101",
  9539=>"100011101",
  9540=>"010101101",
  9541=>"010110111",
  9542=>"111001011",
  9543=>"001001010",
  9544=>"111100110",
  9545=>"011001011",
  9546=>"100111110",
  9547=>"000111011",
  9548=>"001001010",
  9549=>"111111001",
  9550=>"010001010",
  9551=>"011000110",
  9552=>"100111110",
  9553=>"100000100",
  9554=>"010111110",
  9555=>"011101101",
  9556=>"010001101",
  9557=>"100101101",
  9558=>"110000111",
  9559=>"110001000",
  9560=>"100100101",
  9561=>"000001101",
  9562=>"001100110",
  9563=>"111100001",
  9564=>"100111101",
  9565=>"100101011",
  9566=>"110111111",
  9567=>"011010001",
  9568=>"110110100",
  9569=>"010110001",
  9570=>"000001001",
  9571=>"001000110",
  9572=>"100001101",
  9573=>"100000100",
  9574=>"100011111",
  9575=>"000101110",
  9576=>"101110001",
  9577=>"001010111",
  9578=>"011000010",
  9579=>"011011011",
  9580=>"111100001",
  9581=>"101101011",
  9582=>"101001011",
  9583=>"000110100",
  9584=>"100110011",
  9585=>"000001111",
  9586=>"110001111",
  9587=>"111011011",
  9588=>"101000100",
  9589=>"010001111",
  9590=>"001101011",
  9591=>"000010101",
  9592=>"011101101",
  9593=>"111001010",
  9594=>"101111111",
  9595=>"111011100",
  9596=>"000000110",
  9597=>"111110111",
  9598=>"101010010",
  9599=>"111100001",
  9600=>"001010011",
  9601=>"110000010",
  9602=>"101011101",
  9603=>"001110101",
  9604=>"111000111",
  9605=>"110101101",
  9606=>"110011101",
  9607=>"011111101",
  9608=>"010100010",
  9609=>"011010111",
  9610=>"011111111",
  9611=>"011010101",
  9612=>"010101001",
  9613=>"100010000",
  9614=>"010010101",
  9615=>"010110000",
  9616=>"100001101",
  9617=>"000111111",
  9618=>"101101000",
  9619=>"010111111",
  9620=>"110010111",
  9621=>"100000001",
  9622=>"101000001",
  9623=>"101010100",
  9624=>"111010111",
  9625=>"101001000",
  9626=>"111111101",
  9627=>"111011000",
  9628=>"010010100",
  9629=>"001000100",
  9630=>"000110100",
  9631=>"100110011",
  9632=>"010101100",
  9633=>"011001101",
  9634=>"100010000",
  9635=>"010001000",
  9636=>"111000111",
  9637=>"100000001",
  9638=>"110001000",
  9639=>"010010111",
  9640=>"010110111",
  9641=>"100001101",
  9642=>"000111000",
  9643=>"010110111",
  9644=>"000001011",
  9645=>"000101011",
  9646=>"010100010",
  9647=>"011000100",
  9648=>"101110110",
  9649=>"000001100",
  9650=>"011101001",
  9651=>"001110111",
  9652=>"001111100",
  9653=>"111101101",
  9654=>"001100011",
  9655=>"111011011",
  9656=>"101011001",
  9657=>"110000000",
  9658=>"010011111",
  9659=>"000110001",
  9660=>"000010010",
  9661=>"101000000",
  9662=>"010000010",
  9663=>"110110100",
  9664=>"110000001",
  9665=>"101111101",
  9666=>"001010000",
  9667=>"101001011",
  9668=>"011100100",
  9669=>"000001100",
  9670=>"111010010",
  9671=>"101001001",
  9672=>"010100110",
  9673=>"001101011",
  9674=>"011111000",
  9675=>"101110111",
  9676=>"100001011",
  9677=>"100010001",
  9678=>"010110000",
  9679=>"111110100",
  9680=>"101001111",
  9681=>"100100101",
  9682=>"010110101",
  9683=>"000110010",
  9684=>"011110001",
  9685=>"000010011",
  9686=>"110011110",
  9687=>"110011110",
  9688=>"001000111",
  9689=>"101110001",
  9690=>"111110001",
  9691=>"100011100",
  9692=>"101110011",
  9693=>"000011100",
  9694=>"101100000",
  9695=>"110110100",
  9696=>"000010101",
  9697=>"000101110",
  9698=>"111100001",
  9699=>"111100110",
  9700=>"000010001",
  9701=>"001011111",
  9702=>"010000001",
  9703=>"001001101",
  9704=>"010110001",
  9705=>"101101110",
  9706=>"000101110",
  9707=>"010000000",
  9708=>"000001011",
  9709=>"111010111",
  9710=>"000110010",
  9711=>"000011101",
  9712=>"101100000",
  9713=>"101100000",
  9714=>"100110111",
  9715=>"010010101",
  9716=>"101010011",
  9717=>"001111110",
  9718=>"100100101",
  9719=>"011110100",
  9720=>"100010100",
  9721=>"110110001",
  9722=>"001111001",
  9723=>"101100101",
  9724=>"000000010",
  9725=>"100001010",
  9726=>"001111111",
  9727=>"100101001",
  9728=>"011111001",
  9729=>"001101001",
  9730=>"110110111",
  9731=>"111011111",
  9732=>"011000110",
  9733=>"000010000",
  9734=>"101011011",
  9735=>"000110011",
  9736=>"000110000",
  9737=>"111111001",
  9738=>"100001100",
  9739=>"110001100",
  9740=>"001111010",
  9741=>"000011000",
  9742=>"110100000",
  9743=>"110001111",
  9744=>"100110010",
  9745=>"000000101",
  9746=>"111111100",
  9747=>"100111010",
  9748=>"000000000",
  9749=>"010000000",
  9750=>"100100101",
  9751=>"000110111",
  9752=>"001111001",
  9753=>"001101100",
  9754=>"101110101",
  9755=>"001100101",
  9756=>"010110101",
  9757=>"110011000",
  9758=>"001011000",
  9759=>"001000100",
  9760=>"011010010",
  9761=>"100001110",
  9762=>"001001100",
  9763=>"010010111",
  9764=>"001111010",
  9765=>"110001000",
  9766=>"000000001",
  9767=>"101100111",
  9768=>"011110001",
  9769=>"100010000",
  9770=>"011011001",
  9771=>"011000010",
  9772=>"110011010",
  9773=>"000100000",
  9774=>"111111000",
  9775=>"000101001",
  9776=>"110001110",
  9777=>"101110111",
  9778=>"010001000",
  9779=>"000101001",
  9780=>"101011101",
  9781=>"110100110",
  9782=>"000001011",
  9783=>"110111100",
  9784=>"111100101",
  9785=>"101011110",
  9786=>"110110010",
  9787=>"110100010",
  9788=>"001001110",
  9789=>"011001001",
  9790=>"111110001",
  9791=>"011101000",
  9792=>"100011011",
  9793=>"001110100",
  9794=>"010101011",
  9795=>"000100101",
  9796=>"001101001",
  9797=>"110100000",
  9798=>"100110100",
  9799=>"001001101",
  9800=>"111110111",
  9801=>"111110011",
  9802=>"101110111",
  9803=>"111101010",
  9804=>"110100000",
  9805=>"001110110",
  9806=>"100111011",
  9807=>"000000110",
  9808=>"101111000",
  9809=>"110111111",
  9810=>"100000111",
  9811=>"111101000",
  9812=>"011100101",
  9813=>"001010111",
  9814=>"001000101",
  9815=>"101111100",
  9816=>"011001110",
  9817=>"010111000",
  9818=>"010101100",
  9819=>"101000100",
  9820=>"000111000",
  9821=>"001011111",
  9822=>"000000101",
  9823=>"000111100",
  9824=>"101000010",
  9825=>"000011000",
  9826=>"111011100",
  9827=>"000111000",
  9828=>"001111101",
  9829=>"111011100",
  9830=>"100111001",
  9831=>"011000001",
  9832=>"000100101",
  9833=>"000011010",
  9834=>"001110111",
  9835=>"111010010",
  9836=>"111101100",
  9837=>"000010101",
  9838=>"011101111",
  9839=>"100011101",
  9840=>"010101100",
  9841=>"000010100",
  9842=>"000100000",
  9843=>"000000000",
  9844=>"001000010",
  9845=>"110111011",
  9846=>"001111000",
  9847=>"001101110",
  9848=>"001011111",
  9849=>"011101100",
  9850=>"101010101",
  9851=>"000111111",
  9852=>"000100000",
  9853=>"001111011",
  9854=>"010100011",
  9855=>"000111110",
  9856=>"011110100",
  9857=>"110011111",
  9858=>"000000001",
  9859=>"111000010",
  9860=>"011000000",
  9861=>"000100011",
  9862=>"011011101",
  9863=>"001010100",
  9864=>"111010010",
  9865=>"000000010",
  9866=>"110111101",
  9867=>"010111011",
  9868=>"010100001",
  9869=>"011001101",
  9870=>"111000010",
  9871=>"011101011",
  9872=>"100101010",
  9873=>"000100000",
  9874=>"111101111",
  9875=>"101001110",
  9876=>"000110100",
  9877=>"111111111",
  9878=>"001111100",
  9879=>"001110100",
  9880=>"011110001",
  9881=>"100101001",
  9882=>"110000111",
  9883=>"011111000",
  9884=>"111111100",
  9885=>"100000000",
  9886=>"000011000",
  9887=>"101000111",
  9888=>"101000000",
  9889=>"110000101",
  9890=>"010110111",
  9891=>"110111111",
  9892=>"100111101",
  9893=>"010101101",
  9894=>"010100001",
  9895=>"111001101",
  9896=>"111000110",
  9897=>"111000101",
  9898=>"001000110",
  9899=>"110000010",
  9900=>"110000110",
  9901=>"101000010",
  9902=>"010001011",
  9903=>"101111100",
  9904=>"111010101",
  9905=>"011011011",
  9906=>"001111000",
  9907=>"101110101",
  9908=>"100001000",
  9909=>"010010110",
  9910=>"111111011",
  9911=>"100110100",
  9912=>"011101000",
  9913=>"010001100",
  9914=>"110100010",
  9915=>"101010010",
  9916=>"111001110",
  9917=>"010101011",
  9918=>"001000010",
  9919=>"011111100",
  9920=>"110000110",
  9921=>"010010110",
  9922=>"110001001",
  9923=>"110001111",
  9924=>"001111010",
  9925=>"100100110",
  9926=>"111110111",
  9927=>"000001000",
  9928=>"100001110",
  9929=>"111010001",
  9930=>"101110100",
  9931=>"110111011",
  9932=>"001101000",
  9933=>"011011001",
  9934=>"101010111",
  9935=>"011100000",
  9936=>"000010001",
  9937=>"000100000",
  9938=>"101101000",
  9939=>"010100011",
  9940=>"011010100",
  9941=>"110111100",
  9942=>"101011001",
  9943=>"101010011",
  9944=>"100101000",
  9945=>"000001011",
  9946=>"011001000",
  9947=>"101010111",
  9948=>"001100111",
  9949=>"001000000",
  9950=>"011101010",
  9951=>"100010100",
  9952=>"010110001",
  9953=>"111111000",
  9954=>"010101000",
  9955=>"000101111",
  9956=>"000111111",
  9957=>"101111001",
  9958=>"100011001",
  9959=>"001000000",
  9960=>"011010011",
  9961=>"111010111",
  9962=>"110111110",
  9963=>"100100111",
  9964=>"110001010",
  9965=>"101111111",
  9966=>"001111110",
  9967=>"111101111",
  9968=>"111000110",
  9969=>"111101011",
  9970=>"101000110",
  9971=>"100000001",
  9972=>"000110100",
  9973=>"101100000",
  9974=>"000100100",
  9975=>"101011111",
  9976=>"001000010",
  9977=>"111100000",
  9978=>"000101100",
  9979=>"110001011",
  9980=>"001111111",
  9981=>"010101101",
  9982=>"111000011",
  9983=>"011010110",
  9984=>"001011000",
  9985=>"000010101",
  9986=>"000010010",
  9987=>"011000010",
  9988=>"000001101",
  9989=>"001010110",
  9990=>"100110110",
  9991=>"000000010",
  9992=>"011110101",
  9993=>"010110111",
  9994=>"101001010",
  9995=>"000000000",
  9996=>"000011101",
  9997=>"111010001",
  9998=>"000000000",
  9999=>"111011110",
  10000=>"011100110",
  10001=>"100100011",
  10002=>"100001010",
  10003=>"000101100",
  10004=>"111011000",
  10005=>"100100101",
  10006=>"000000011",
  10007=>"111001010",
  10008=>"011111001",
  10009=>"010010001",
  10010=>"111101111",
  10011=>"010010101",
  10012=>"110111011",
  10013=>"111111001",
  10014=>"010100001",
  10015=>"010000000",
  10016=>"111001010",
  10017=>"101001111",
  10018=>"101110001",
  10019=>"010101111",
  10020=>"011101011",
  10021=>"111101001",
  10022=>"010100011",
  10023=>"100110010",
  10024=>"101010101",
  10025=>"101000110",
  10026=>"011110001",
  10027=>"001101001",
  10028=>"000011110",
  10029=>"000000001",
  10030=>"000011110",
  10031=>"011000001",
  10032=>"101000101",
  10033=>"110101011",
  10034=>"110010000",
  10035=>"001100110",
  10036=>"111111010",
  10037=>"111100100",
  10038=>"100001100",
  10039=>"000000011",
  10040=>"000011000",
  10041=>"001001111",
  10042=>"101110010",
  10043=>"000110000",
  10044=>"001010110",
  10045=>"101010011",
  10046=>"011111011",
  10047=>"011111100",
  10048=>"100111101",
  10049=>"100101011",
  10050=>"101111011",
  10051=>"001011111",
  10052=>"010101111",
  10053=>"111111111",
  10054=>"110011010",
  10055=>"010011010",
  10056=>"100101011",
  10057=>"010111000",
  10058=>"100110010",
  10059=>"111010000",
  10060=>"011101100",
  10061=>"101110111",
  10062=>"001100100",
  10063=>"101111101",
  10064=>"000111010",
  10065=>"000010110",
  10066=>"001101111",
  10067=>"001111011",
  10068=>"111101011",
  10069=>"010101011",
  10070=>"000001010",
  10071=>"001111011",
  10072=>"001110000",
  10073=>"110110000",
  10074=>"000100101",
  10075=>"000000001",
  10076=>"110001000",
  10077=>"001101000",
  10078=>"010001010",
  10079=>"100011110",
  10080=>"000110111",
  10081=>"001101011",
  10082=>"100101011",
  10083=>"111000001",
  10084=>"111101000",
  10085=>"001001100",
  10086=>"001000000",
  10087=>"011011011",
  10088=>"111111001",
  10089=>"010000111",
  10090=>"011110001",
  10091=>"101000110",
  10092=>"110111110",
  10093=>"011110010",
  10094=>"110001011",
  10095=>"110101111",
  10096=>"110101000",
  10097=>"110101010",
  10098=>"111000110",
  10099=>"000011000",
  10100=>"010001000",
  10101=>"111001111",
  10102=>"000011010",
  10103=>"101000000",
  10104=>"111110010",
  10105=>"110110000",
  10106=>"101101000",
  10107=>"100011101",
  10108=>"010011001",
  10109=>"001000110",
  10110=>"101001001",
  10111=>"011010101",
  10112=>"100101001",
  10113=>"001100110",
  10114=>"010100110",
  10115=>"011010000",
  10116=>"011101110",
  10117=>"100010010",
  10118=>"100001111",
  10119=>"111001011",
  10120=>"010011111",
  10121=>"100001100",
  10122=>"011011001",
  10123=>"101000000",
  10124=>"010011001",
  10125=>"011011101",
  10126=>"100110000",
  10127=>"011001100",
  10128=>"011011010",
  10129=>"010011010",
  10130=>"000001000",
  10131=>"000011110",
  10132=>"001101100",
  10133=>"001111100",
  10134=>"111100101",
  10135=>"101111111",
  10136=>"000010100",
  10137=>"111101101",
  10138=>"100111000",
  10139=>"000000010",
  10140=>"100101010",
  10141=>"111111101",
  10142=>"010101100",
  10143=>"011010000",
  10144=>"011110011",
  10145=>"100010000",
  10146=>"011001000",
  10147=>"110001100",
  10148=>"001100010",
  10149=>"001111101",
  10150=>"010110011",
  10151=>"010110111",
  10152=>"001010011",
  10153=>"000010000",
  10154=>"101010110",
  10155=>"010010100",
  10156=>"101100110",
  10157=>"000111010",
  10158=>"000101101",
  10159=>"101110111",
  10160=>"110110001",
  10161=>"101111100",
  10162=>"110010010",
  10163=>"011101000",
  10164=>"011001000",
  10165=>"101011000",
  10166=>"000110111",
  10167=>"011000111",
  10168=>"001101001",
  10169=>"011110001",
  10170=>"010111110",
  10171=>"100111000",
  10172=>"010010000",
  10173=>"000100101",
  10174=>"111110110",
  10175=>"110100000",
  10176=>"101010101",
  10177=>"100111011",
  10178=>"100110010",
  10179=>"101100100",
  10180=>"111111110",
  10181=>"000011011",
  10182=>"001011010",
  10183=>"000110000",
  10184=>"111001101",
  10185=>"100011001",
  10186=>"011011101",
  10187=>"010010100",
  10188=>"110011101",
  10189=>"010010000",
  10190=>"001000110",
  10191=>"110100000",
  10192=>"000011011",
  10193=>"110100111",
  10194=>"010101101",
  10195=>"101111010",
  10196=>"000010010",
  10197=>"111011110",
  10198=>"100001100",
  10199=>"000010010",
  10200=>"101000101",
  10201=>"001010101",
  10202=>"000111000",
  10203=>"110101111",
  10204=>"100100011",
  10205=>"110011000",
  10206=>"111000101",
  10207=>"011101100",
  10208=>"000000010",
  10209=>"100001111",
  10210=>"001001100",
  10211=>"000101100",
  10212=>"000001000",
  10213=>"111111111",
  10214=>"011011111",
  10215=>"011000001",
  10216=>"010001001",
  10217=>"101010110",
  10218=>"001010001",
  10219=>"111010001",
  10220=>"000100001",
  10221=>"001101011",
  10222=>"000100101",
  10223=>"010110011",
  10224=>"011000010",
  10225=>"001001001",
  10226=>"000001001",
  10227=>"110010001",
  10228=>"001111101",
  10229=>"000111011",
  10230=>"111101001",
  10231=>"111010101",
  10232=>"101100101",
  10233=>"000001110",
  10234=>"100100111",
  10235=>"100100111",
  10236=>"111001110",
  10237=>"110100000",
  10238=>"010011000",
  10239=>"100010111",
  10240=>"100110111",
  10241=>"010100100",
  10242=>"111101001",
  10243=>"000111001",
  10244=>"010110011",
  10245=>"101000001",
  10246=>"100110001",
  10247=>"011110010",
  10248=>"101010110",
  10249=>"011010001",
  10250=>"000001101",
  10251=>"001011100",
  10252=>"000000000",
  10253=>"011001101",
  10254=>"001000110",
  10255=>"000100011",
  10256=>"001010110",
  10257=>"101101111",
  10258=>"100011100",
  10259=>"010010101",
  10260=>"001111000",
  10261=>"111111001",
  10262=>"110000111",
  10263=>"100100011",
  10264=>"110110100",
  10265=>"100110111",
  10266=>"101100101",
  10267=>"100100001",
  10268=>"010010111",
  10269=>"111001011",
  10270=>"111110001",
  10271=>"110100111",
  10272=>"000111000",
  10273=>"001110111",
  10274=>"000010000",
  10275=>"001001101",
  10276=>"111110111",
  10277=>"011101000",
  10278=>"001001000",
  10279=>"100000011",
  10280=>"010010010",
  10281=>"101011010",
  10282=>"010011101",
  10283=>"101010100",
  10284=>"000100101",
  10285=>"101001000",
  10286=>"100111000",
  10287=>"001100110",
  10288=>"111110010",
  10289=>"000001110",
  10290=>"000001110",
  10291=>"100000110",
  10292=>"101000010",
  10293=>"110000100",
  10294=>"111010010",
  10295=>"110101111",
  10296=>"011110101",
  10297=>"111111111",
  10298=>"111000001",
  10299=>"110100110",
  10300=>"010101101",
  10301=>"101010111",
  10302=>"100000100",
  10303=>"010001000",
  10304=>"111101000",
  10305=>"010011101",
  10306=>"000001000",
  10307=>"000101011",
  10308=>"010101001",
  10309=>"101101110",
  10310=>"000110101",
  10311=>"000010000",
  10312=>"011100110",
  10313=>"100111001",
  10314=>"100010111",
  10315=>"000111011",
  10316=>"111101100",
  10317=>"000001000",
  10318=>"000000110",
  10319=>"111001101",
  10320=>"110100101",
  10321=>"000010000",
  10322=>"010000010",
  10323=>"111100100",
  10324=>"010000000",
  10325=>"100000001",
  10326=>"010110001",
  10327=>"001000001",
  10328=>"111101001",
  10329=>"101011000",
  10330=>"010101100",
  10331=>"011101111",
  10332=>"000111110",
  10333=>"101110000",
  10334=>"011000010",
  10335=>"110100101",
  10336=>"001110110",
  10337=>"100100101",
  10338=>"001111111",
  10339=>"001000001",
  10340=>"111111001",
  10341=>"111010110",
  10342=>"001011000",
  10343=>"000010111",
  10344=>"011001111",
  10345=>"010101000",
  10346=>"100000010",
  10347=>"101011011",
  10348=>"110000110",
  10349=>"010111110",
  10350=>"010101100",
  10351=>"111010001",
  10352=>"010101011",
  10353=>"111000100",
  10354=>"001010100",
  10355=>"000010100",
  10356=>"101001011",
  10357=>"001111111",
  10358=>"101000011",
  10359=>"011100100",
  10360=>"110010011",
  10361=>"101000000",
  10362=>"100011101",
  10363=>"000101111",
  10364=>"100110000",
  10365=>"010111001",
  10366=>"110100011",
  10367=>"000000011",
  10368=>"100011101",
  10369=>"011101101",
  10370=>"000011100",
  10371=>"101100101",
  10372=>"010101010",
  10373=>"011100010",
  10374=>"001011011",
  10375=>"111111111",
  10376=>"100100011",
  10377=>"100100010",
  10378=>"111000010",
  10379=>"111001001",
  10380=>"111100100",
  10381=>"000010000",
  10382=>"100101010",
  10383=>"110111101",
  10384=>"111111101",
  10385=>"111001011",
  10386=>"011011110",
  10387=>"011110110",
  10388=>"111101011",
  10389=>"100100111",
  10390=>"001100001",
  10391=>"101110011",
  10392=>"000010111",
  10393=>"100110001",
  10394=>"010110001",
  10395=>"011011011",
  10396=>"000101010",
  10397=>"101111111",
  10398=>"000011111",
  10399=>"111101110",
  10400=>"101010001",
  10401=>"100000101",
  10402=>"001110000",
  10403=>"011111010",
  10404=>"111111110",
  10405=>"010101001",
  10406=>"100110000",
  10407=>"111100110",
  10408=>"001001101",
  10409=>"011010000",
  10410=>"000011010",
  10411=>"101000100",
  10412=>"111000000",
  10413=>"110101101",
  10414=>"110111111",
  10415=>"110000010",
  10416=>"011001111",
  10417=>"110111110",
  10418=>"001010011",
  10419=>"001111010",
  10420=>"110111111",
  10421=>"100111111",
  10422=>"110001010",
  10423=>"110111110",
  10424=>"110001011",
  10425=>"100100100",
  10426=>"110100000",
  10427=>"001101101",
  10428=>"011001000",
  10429=>"110011110",
  10430=>"110011100",
  10431=>"101100101",
  10432=>"111001100",
  10433=>"011101000",
  10434=>"001001100",
  10435=>"011010001",
  10436=>"010000100",
  10437=>"100010111",
  10438=>"000111010",
  10439=>"101101101",
  10440=>"100011010",
  10441=>"011101010",
  10442=>"001010100",
  10443=>"001011111",
  10444=>"001000000",
  10445=>"100000010",
  10446=>"011101111",
  10447=>"111011110",
  10448=>"110001011",
  10449=>"110000010",
  10450=>"100001100",
  10451=>"111111110",
  10452=>"101001100",
  10453=>"000101010",
  10454=>"000000001",
  10455=>"010001011",
  10456=>"010011000",
  10457=>"001000110",
  10458=>"101100011",
  10459=>"010100001",
  10460=>"111100101",
  10461=>"001101110",
  10462=>"001101001",
  10463=>"010001100",
  10464=>"101000110",
  10465=>"100000001",
  10466=>"101110111",
  10467=>"100000100",
  10468=>"100000001",
  10469=>"111010010",
  10470=>"111111101",
  10471=>"110110110",
  10472=>"000000000",
  10473=>"100100100",
  10474=>"111110111",
  10475=>"110010011",
  10476=>"001110000",
  10477=>"101000010",
  10478=>"111000010",
  10479=>"000110101",
  10480=>"111001100",
  10481=>"010111111",
  10482=>"111100111",
  10483=>"111101001",
  10484=>"000001010",
  10485=>"010000000",
  10486=>"010111110",
  10487=>"000000000",
  10488=>"000001100",
  10489=>"110011111",
  10490=>"001011110",
  10491=>"001101110",
  10492=>"010011011",
  10493=>"000011100",
  10494=>"011000010",
  10495=>"000000111",
  10496=>"001011011",
  10497=>"100110000",
  10498=>"100001011",
  10499=>"100010111",
  10500=>"111110101",
  10501=>"000101101",
  10502=>"010111111",
  10503=>"000010111",
  10504=>"101111111",
  10505=>"000010111",
  10506=>"110011010",
  10507=>"000100111",
  10508=>"000111101",
  10509=>"010101100",
  10510=>"110101001",
  10511=>"111010011",
  10512=>"011111000",
  10513=>"000010110",
  10514=>"110001100",
  10515=>"111101101",
  10516=>"001100011",
  10517=>"001100110",
  10518=>"110110000",
  10519=>"010110101",
  10520=>"100010000",
  10521=>"001000101",
  10522=>"100100110",
  10523=>"111101010",
  10524=>"110000001",
  10525=>"101010100",
  10526=>"000001110",
  10527=>"000001010",
  10528=>"110111000",
  10529=>"011101100",
  10530=>"011000000",
  10531=>"000001011",
  10532=>"101110110",
  10533=>"111100101",
  10534=>"110101110",
  10535=>"010100001",
  10536=>"101000100",
  10537=>"010010001",
  10538=>"011010011",
  10539=>"000011111",
  10540=>"011011100",
  10541=>"101001010",
  10542=>"100110000",
  10543=>"101100000",
  10544=>"001111100",
  10545=>"001110110",
  10546=>"010001111",
  10547=>"000101001",
  10548=>"011011001",
  10549=>"000001101",
  10550=>"101001110",
  10551=>"110011111",
  10552=>"010000101",
  10553=>"011011100",
  10554=>"101100010",
  10555=>"000100110",
  10556=>"001100110",
  10557=>"111101000",
  10558=>"110111100",
  10559=>"101010111",
  10560=>"000001110",
  10561=>"011110011",
  10562=>"000001011",
  10563=>"010111011",
  10564=>"111001000",
  10565=>"001000110",
  10566=>"000001100",
  10567=>"101101111",
  10568=>"111101000",
  10569=>"000111111",
  10570=>"010111001",
  10571=>"111111001",
  10572=>"000010101",
  10573=>"001110101",
  10574=>"011011101",
  10575=>"001100110",
  10576=>"010111100",
  10577=>"101000011",
  10578=>"111010011",
  10579=>"110110011",
  10580=>"000110001",
  10581=>"000001011",
  10582=>"000110000",
  10583=>"011000010",
  10584=>"101010111",
  10585=>"100100000",
  10586=>"011101001",
  10587=>"111001111",
  10588=>"111011100",
  10589=>"011110110",
  10590=>"101100000",
  10591=>"011011100",
  10592=>"010001110",
  10593=>"010010001",
  10594=>"011111110",
  10595=>"010101011",
  10596=>"111110010",
  10597=>"110011101",
  10598=>"011010101",
  10599=>"000001110",
  10600=>"000010011",
  10601=>"001111000",
  10602=>"001011010",
  10603=>"110010111",
  10604=>"101101001",
  10605=>"101000100",
  10606=>"100001010",
  10607=>"110010100",
  10608=>"110011111",
  10609=>"010000101",
  10610=>"010000011",
  10611=>"000011000",
  10612=>"010001000",
  10613=>"111101111",
  10614=>"011010111",
  10615=>"111001100",
  10616=>"011011101",
  10617=>"000101110",
  10618=>"111000011",
  10619=>"010011110",
  10620=>"111011010",
  10621=>"101111101",
  10622=>"101110110",
  10623=>"111001101",
  10624=>"010100010",
  10625=>"100101110",
  10626=>"011011010",
  10627=>"011101000",
  10628=>"111111101",
  10629=>"001000010",
  10630=>"011110001",
  10631=>"011000001",
  10632=>"101101010",
  10633=>"101110100",
  10634=>"011111000",
  10635=>"111111011",
  10636=>"011000001",
  10637=>"111100100",
  10638=>"000011100",
  10639=>"101100101",
  10640=>"110101101",
  10641=>"010101011",
  10642=>"001011111",
  10643=>"100001101",
  10644=>"011011011",
  10645=>"100000110",
  10646=>"100100101",
  10647=>"110111111",
  10648=>"100011010",
  10649=>"110000001",
  10650=>"101111111",
  10651=>"100010100",
  10652=>"010111011",
  10653=>"111001111",
  10654=>"110100010",
  10655=>"110100101",
  10656=>"101100001",
  10657=>"111000001",
  10658=>"100001111",
  10659=>"000001111",
  10660=>"111101111",
  10661=>"110000100",
  10662=>"000111010",
  10663=>"001000111",
  10664=>"101000011",
  10665=>"000111011",
  10666=>"010001001",
  10667=>"000010101",
  10668=>"101011100",
  10669=>"111001010",
  10670=>"111111111",
  10671=>"010010111",
  10672=>"011101111",
  10673=>"001111111",
  10674=>"101000100",
  10675=>"111001010",
  10676=>"001111111",
  10677=>"110100111",
  10678=>"100110100",
  10679=>"101101101",
  10680=>"010100000",
  10681=>"001010011",
  10682=>"001000111",
  10683=>"101000000",
  10684=>"100010100",
  10685=>"010101101",
  10686=>"101011000",
  10687=>"101100000",
  10688=>"101100101",
  10689=>"111001111",
  10690=>"111011001",
  10691=>"111110110",
  10692=>"110000011",
  10693=>"001111100",
  10694=>"111111111",
  10695=>"101010101",
  10696=>"110110110",
  10697=>"111111010",
  10698=>"000000110",
  10699=>"100010011",
  10700=>"100101001",
  10701=>"000010011",
  10702=>"110100000",
  10703=>"011000000",
  10704=>"010010001",
  10705=>"111011110",
  10706=>"111100111",
  10707=>"110000101",
  10708=>"010011010",
  10709=>"100010100",
  10710=>"111011100",
  10711=>"001001001",
  10712=>"000001000",
  10713=>"011111111",
  10714=>"111101010",
  10715=>"111111010",
  10716=>"100000111",
  10717=>"101001011",
  10718=>"000010110",
  10719=>"100110010",
  10720=>"011000111",
  10721=>"110110101",
  10722=>"001011011",
  10723=>"100010111",
  10724=>"110000110",
  10725=>"110110110",
  10726=>"101010100",
  10727=>"010111010",
  10728=>"000001110",
  10729=>"011101110",
  10730=>"000100100",
  10731=>"100001011",
  10732=>"111010101",
  10733=>"101011110",
  10734=>"110000111",
  10735=>"001000100",
  10736=>"000111101",
  10737=>"110101010",
  10738=>"111000000",
  10739=>"101011101",
  10740=>"010001000",
  10741=>"000010001",
  10742=>"011101100",
  10743=>"111000101",
  10744=>"111111000",
  10745=>"000101001",
  10746=>"010000100",
  10747=>"010110000",
  10748=>"000010111",
  10749=>"101100011",
  10750=>"011111000",
  10751=>"001000010",
  10752=>"111011101",
  10753=>"000001111",
  10754=>"110100111",
  10755=>"010110011",
  10756=>"111100001",
  10757=>"100111011",
  10758=>"110011010",
  10759=>"000110110",
  10760=>"011011001",
  10761=>"010000000",
  10762=>"011111010",
  10763=>"010110000",
  10764=>"010100100",
  10765=>"001100010",
  10766=>"000100001",
  10767=>"000001011",
  10768=>"111010000",
  10769=>"000010010",
  10770=>"111001100",
  10771=>"010011111",
  10772=>"110000000",
  10773=>"110000110",
  10774=>"111001101",
  10775=>"001100101",
  10776=>"001101111",
  10777=>"010011110",
  10778=>"000001001",
  10779=>"010101110",
  10780=>"011011000",
  10781=>"001001110",
  10782=>"110001100",
  10783=>"011100110",
  10784=>"010010001",
  10785=>"000010000",
  10786=>"010000010",
  10787=>"100101111",
  10788=>"110100101",
  10789=>"111001101",
  10790=>"100001110",
  10791=>"111110100",
  10792=>"011110100",
  10793=>"011011111",
  10794=>"101000001",
  10795=>"111111111",
  10796=>"110101101",
  10797=>"011100000",
  10798=>"010011111",
  10799=>"010001001",
  10800=>"011011110",
  10801=>"111001111",
  10802=>"000100011",
  10803=>"101101111",
  10804=>"100000001",
  10805=>"101111010",
  10806=>"010110110",
  10807=>"100011001",
  10808=>"110101001",
  10809=>"100110011",
  10810=>"010101101",
  10811=>"000000011",
  10812=>"011110101",
  10813=>"000110101",
  10814=>"010000000",
  10815=>"001101111",
  10816=>"011010111",
  10817=>"001111110",
  10818=>"101001001",
  10819=>"101101000",
  10820=>"100001010",
  10821=>"101000100",
  10822=>"001000010",
  10823=>"101001001",
  10824=>"001000000",
  10825=>"001110100",
  10826=>"100101101",
  10827=>"111111001",
  10828=>"010110001",
  10829=>"010100100",
  10830=>"111111100",
  10831=>"110010000",
  10832=>"110100111",
  10833=>"011001000",
  10834=>"110100110",
  10835=>"001101111",
  10836=>"001100111",
  10837=>"000110011",
  10838=>"101110000",
  10839=>"111000111",
  10840=>"010111001",
  10841=>"010001110",
  10842=>"100010100",
  10843=>"010101010",
  10844=>"000111110",
  10845=>"011010111",
  10846=>"110001010",
  10847=>"100010001",
  10848=>"111011000",
  10849=>"010010010",
  10850=>"010010011",
  10851=>"010010010",
  10852=>"110010110",
  10853=>"101001000",
  10854=>"010001111",
  10855=>"010110000",
  10856=>"010010000",
  10857=>"101010011",
  10858=>"010111001",
  10859=>"101111001",
  10860=>"001101110",
  10861=>"010001100",
  10862=>"011000001",
  10863=>"000110111",
  10864=>"010011000",
  10865=>"010101001",
  10866=>"110111101",
  10867=>"100110101",
  10868=>"100101101",
  10869=>"110101100",
  10870=>"111011101",
  10871=>"111100101",
  10872=>"100011010",
  10873=>"000001101",
  10874=>"111011000",
  10875=>"111011001",
  10876=>"011000000",
  10877=>"000110000",
  10878=>"001100000",
  10879=>"011101001",
  10880=>"110110010",
  10881=>"100101110",
  10882=>"101101101",
  10883=>"110101001",
  10884=>"100111010",
  10885=>"011000110",
  10886=>"110010000",
  10887=>"010101001",
  10888=>"000010010",
  10889=>"011011110",
  10890=>"100011100",
  10891=>"010010101",
  10892=>"101000111",
  10893=>"111100101",
  10894=>"010000000",
  10895=>"100111001",
  10896=>"101100010",
  10897=>"111111111",
  10898=>"000000010",
  10899=>"011001101",
  10900=>"011111011",
  10901=>"011111001",
  10902=>"111010110",
  10903=>"011010001",
  10904=>"100000100",
  10905=>"100100101",
  10906=>"101011110",
  10907=>"010110001",
  10908=>"001100100",
  10909=>"101101110",
  10910=>"111110010",
  10911=>"010011101",
  10912=>"100000111",
  10913=>"111110010",
  10914=>"101111010",
  10915=>"100101011",
  10916=>"111100000",
  10917=>"001101111",
  10918=>"110011111",
  10919=>"010000100",
  10920=>"011100110",
  10921=>"101011010",
  10922=>"100110101",
  10923=>"110000100",
  10924=>"001010001",
  10925=>"101000100",
  10926=>"110010110",
  10927=>"110110100",
  10928=>"001010000",
  10929=>"101110101",
  10930=>"110010001",
  10931=>"101011101",
  10932=>"010100010",
  10933=>"011001110",
  10934=>"100001010",
  10935=>"001010101",
  10936=>"000011010",
  10937=>"101101111",
  10938=>"000111010",
  10939=>"110011000",
  10940=>"101110001",
  10941=>"000101000",
  10942=>"110101011",
  10943=>"010011000",
  10944=>"111010111",
  10945=>"011110011",
  10946=>"110001010",
  10947=>"101011000",
  10948=>"000100001",
  10949=>"111000010",
  10950=>"001101101",
  10951=>"000110001",
  10952=>"010000101",
  10953=>"111110100",
  10954=>"110111110",
  10955=>"000010011",
  10956=>"111100101",
  10957=>"100100010",
  10958=>"111000011",
  10959=>"101001011",
  10960=>"110000000",
  10961=>"001100011",
  10962=>"010000001",
  10963=>"101110001",
  10964=>"001010100",
  10965=>"110001101",
  10966=>"110100101",
  10967=>"000111110",
  10968=>"010101111",
  10969=>"010011000",
  10970=>"000000101",
  10971=>"011100111",
  10972=>"010000101",
  10973=>"011001000",
  10974=>"010010000",
  10975=>"100011100",
  10976=>"100000000",
  10977=>"001001110",
  10978=>"011110001",
  10979=>"011010101",
  10980=>"000111100",
  10981=>"001100100",
  10982=>"100101110",
  10983=>"000111010",
  10984=>"011001110",
  10985=>"111110010",
  10986=>"111110110",
  10987=>"011110110",
  10988=>"111110011",
  10989=>"111000011",
  10990=>"010100000",
  10991=>"111001101",
  10992=>"100110010",
  10993=>"010100010",
  10994=>"001101100",
  10995=>"010100010",
  10996=>"010100110",
  10997=>"100011101",
  10998=>"011011111",
  10999=>"011101111",
  11000=>"101001001",
  11001=>"101001111",
  11002=>"001011101",
  11003=>"000001001",
  11004=>"110110101",
  11005=>"010111011",
  11006=>"111000100",
  11007=>"101101110",
  11008=>"001100101",
  11009=>"000101111",
  11010=>"110001001",
  11011=>"001100010",
  11012=>"111001001",
  11013=>"010011011",
  11014=>"100110111",
  11015=>"111010110",
  11016=>"000100010",
  11017=>"010110011",
  11018=>"101111011",
  11019=>"000001000",
  11020=>"001111111",
  11021=>"010011001",
  11022=>"110110101",
  11023=>"000011100",
  11024=>"111101101",
  11025=>"111111111",
  11026=>"010101010",
  11027=>"100010000",
  11028=>"000110001",
  11029=>"100011110",
  11030=>"010011101",
  11031=>"000000101",
  11032=>"001000001",
  11033=>"001100010",
  11034=>"101101100",
  11035=>"101010001",
  11036=>"000011000",
  11037=>"101100001",
  11038=>"111011101",
  11039=>"000010000",
  11040=>"000001100",
  11041=>"010100001",
  11042=>"000100011",
  11043=>"000000101",
  11044=>"101000101",
  11045=>"100111100",
  11046=>"011001000",
  11047=>"001101100",
  11048=>"000001010",
  11049=>"110001011",
  11050=>"010001110",
  11051=>"110001101",
  11052=>"001100111",
  11053=>"000001011",
  11054=>"011011110",
  11055=>"001010010",
  11056=>"010001010",
  11057=>"010101101",
  11058=>"001100100",
  11059=>"100001001",
  11060=>"111101111",
  11061=>"011110111",
  11062=>"101110101",
  11063=>"100110010",
  11064=>"110001001",
  11065=>"110100101",
  11066=>"000100011",
  11067=>"001111111",
  11068=>"011110101",
  11069=>"001001001",
  11070=>"001010011",
  11071=>"101111010",
  11072=>"010011011",
  11073=>"000011011",
  11074=>"010111101",
  11075=>"010010110",
  11076=>"000000010",
  11077=>"111111111",
  11078=>"001001110",
  11079=>"011011000",
  11080=>"111101101",
  11081=>"000111100",
  11082=>"011110100",
  11083=>"000001010",
  11084=>"111001101",
  11085=>"011000100",
  11086=>"110011001",
  11087=>"001010101",
  11088=>"101001101",
  11089=>"000011101",
  11090=>"001001111",
  11091=>"011001111",
  11092=>"100100110",
  11093=>"000010111",
  11094=>"111000001",
  11095=>"010100111",
  11096=>"100011110",
  11097=>"010000000",
  11098=>"111010010",
  11099=>"101010100",
  11100=>"110011001",
  11101=>"010101001",
  11102=>"111010000",
  11103=>"000110110",
  11104=>"000001000",
  11105=>"010010111",
  11106=>"011001110",
  11107=>"111011110",
  11108=>"011000101",
  11109=>"111110101",
  11110=>"111010110",
  11111=>"001001111",
  11112=>"101101000",
  11113=>"010100100",
  11114=>"001101100",
  11115=>"010110111",
  11116=>"011100001",
  11117=>"100100111",
  11118=>"101001001",
  11119=>"100010011",
  11120=>"111010110",
  11121=>"010100001",
  11122=>"011101111",
  11123=>"110000011",
  11124=>"001110100",
  11125=>"001000100",
  11126=>"110011100",
  11127=>"001011111",
  11128=>"101010111",
  11129=>"011111100",
  11130=>"011101001",
  11131=>"100101100",
  11132=>"101111111",
  11133=>"000011101",
  11134=>"110010101",
  11135=>"010010010",
  11136=>"110001000",
  11137=>"110111011",
  11138=>"001011010",
  11139=>"000110010",
  11140=>"101100111",
  11141=>"111010111",
  11142=>"000110000",
  11143=>"110010000",
  11144=>"110011010",
  11145=>"000100101",
  11146=>"111000000",
  11147=>"111101111",
  11148=>"101001001",
  11149=>"010011110",
  11150=>"001000111",
  11151=>"011011110",
  11152=>"000000001",
  11153=>"111010100",
  11154=>"000001100",
  11155=>"110101001",
  11156=>"010010111",
  11157=>"000010011",
  11158=>"011101001",
  11159=>"100110011",
  11160=>"011011011",
  11161=>"000100000",
  11162=>"001001110",
  11163=>"100101100",
  11164=>"110000011",
  11165=>"011010000",
  11166=>"110010000",
  11167=>"001110010",
  11168=>"110011001",
  11169=>"110000011",
  11170=>"101101111",
  11171=>"000101000",
  11172=>"010001000",
  11173=>"011111010",
  11174=>"011111111",
  11175=>"011011011",
  11176=>"100100000",
  11177=>"010011001",
  11178=>"011011111",
  11179=>"010011001",
  11180=>"100011110",
  11181=>"101110011",
  11182=>"101010000",
  11183=>"001001000",
  11184=>"011000111",
  11185=>"010001111",
  11186=>"100100001",
  11187=>"111111111",
  11188=>"111101011",
  11189=>"011011001",
  11190=>"110001000",
  11191=>"110001000",
  11192=>"111110110",
  11193=>"011100111",
  11194=>"001100111",
  11195=>"100101010",
  11196=>"000001000",
  11197=>"001111110",
  11198=>"100100110",
  11199=>"101111100",
  11200=>"100111000",
  11201=>"111110100",
  11202=>"100010111",
  11203=>"011000101",
  11204=>"010000001",
  11205=>"100100001",
  11206=>"011100101",
  11207=>"111111101",
  11208=>"100100100",
  11209=>"001000101",
  11210=>"101101011",
  11211=>"101100100",
  11212=>"000101001",
  11213=>"110110000",
  11214=>"101111010",
  11215=>"000100001",
  11216=>"001101100",
  11217=>"010110001",
  11218=>"100111010",
  11219=>"100101001",
  11220=>"100111010",
  11221=>"100001010",
  11222=>"000001101",
  11223=>"000110111",
  11224=>"110100011",
  11225=>"001101010",
  11226=>"100100100",
  11227=>"001111010",
  11228=>"100000001",
  11229=>"100011010",
  11230=>"100011101",
  11231=>"011001010",
  11232=>"100001101",
  11233=>"110001100",
  11234=>"111001111",
  11235=>"101011110",
  11236=>"000101011",
  11237=>"111101011",
  11238=>"101001000",
  11239=>"011001010",
  11240=>"101100100",
  11241=>"001010101",
  11242=>"001100101",
  11243=>"011111001",
  11244=>"010101010",
  11245=>"111001100",
  11246=>"011001110",
  11247=>"111101110",
  11248=>"101101011",
  11249=>"001111101",
  11250=>"101010001",
  11251=>"100110110",
  11252=>"001110110",
  11253=>"010000100",
  11254=>"001101001",
  11255=>"000100110",
  11256=>"000111111",
  11257=>"010101011",
  11258=>"000010000",
  11259=>"101010000",
  11260=>"110100000",
  11261=>"111110111",
  11262=>"100100111",
  11263=>"011001000",
  11264=>"111101111",
  11265=>"110011011",
  11266=>"110111101",
  11267=>"110101101",
  11268=>"011011010",
  11269=>"100101111",
  11270=>"111111111",
  11271=>"010010011",
  11272=>"100001111",
  11273=>"001100111",
  11274=>"000000010",
  11275=>"011001110",
  11276=>"001001101",
  11277=>"110100001",
  11278=>"010100000",
  11279=>"010010000",
  11280=>"111010001",
  11281=>"110011111",
  11282=>"110001001",
  11283=>"111001100",
  11284=>"001110100",
  11285=>"110100010",
  11286=>"001110101",
  11287=>"010100110",
  11288=>"111011000",
  11289=>"010011010",
  11290=>"001010010",
  11291=>"100010011",
  11292=>"101100111",
  11293=>"010101001",
  11294=>"100011101",
  11295=>"101110111",
  11296=>"110101001",
  11297=>"101000100",
  11298=>"000011011",
  11299=>"000100110",
  11300=>"111000000",
  11301=>"101111001",
  11302=>"111011111",
  11303=>"010100011",
  11304=>"010111000",
  11305=>"111000100",
  11306=>"111010101",
  11307=>"100000101",
  11308=>"001010100",
  11309=>"100010111",
  11310=>"011100111",
  11311=>"111000010",
  11312=>"101001000",
  11313=>"100001000",
  11314=>"011000010",
  11315=>"110111010",
  11316=>"000001100",
  11317=>"000000001",
  11318=>"000100101",
  11319=>"011000110",
  11320=>"111010101",
  11321=>"101010000",
  11322=>"000001110",
  11323=>"110000110",
  11324=>"110111010",
  11325=>"000111111",
  11326=>"111110110",
  11327=>"001101110",
  11328=>"011001110",
  11329=>"010000101",
  11330=>"100000111",
  11331=>"111111101",
  11332=>"100011110",
  11333=>"100100111",
  11334=>"111000000",
  11335=>"100000101",
  11336=>"111111001",
  11337=>"111010000",
  11338=>"001101101",
  11339=>"101011011",
  11340=>"111111110",
  11341=>"001011111",
  11342=>"100011000",
  11343=>"110000011",
  11344=>"101011110",
  11345=>"111000110",
  11346=>"010110100",
  11347=>"100000110",
  11348=>"111100010",
  11349=>"110111001",
  11350=>"001100110",
  11351=>"011000111",
  11352=>"010101100",
  11353=>"101111001",
  11354=>"110111101",
  11355=>"001100000",
  11356=>"101011100",
  11357=>"011111100",
  11358=>"000000111",
  11359=>"011101000",
  11360=>"010101010",
  11361=>"101111010",
  11362=>"010111101",
  11363=>"010100101",
  11364=>"100001101",
  11365=>"000000010",
  11366=>"101100001",
  11367=>"001100100",
  11368=>"001011001",
  11369=>"100101010",
  11370=>"011100111",
  11371=>"111001000",
  11372=>"110001101",
  11373=>"011111011",
  11374=>"000100010",
  11375=>"010110000",
  11376=>"010000010",
  11377=>"110001111",
  11378=>"110000111",
  11379=>"011101111",
  11380=>"010100011",
  11381=>"010100000",
  11382=>"011000101",
  11383=>"111000101",
  11384=>"001000001",
  11385=>"010100000",
  11386=>"101000001",
  11387=>"111110011",
  11388=>"100101010",
  11389=>"001110011",
  11390=>"111101000",
  11391=>"011011111",
  11392=>"000010010",
  11393=>"111011101",
  11394=>"110101000",
  11395=>"011001100",
  11396=>"101001101",
  11397=>"001001001",
  11398=>"111010101",
  11399=>"010110111",
  11400=>"011010100",
  11401=>"000000101",
  11402=>"010010011",
  11403=>"101011011",
  11404=>"011001100",
  11405=>"100000001",
  11406=>"111101010",
  11407=>"010111011",
  11408=>"001001110",
  11409=>"001110000",
  11410=>"011110101",
  11411=>"101010010",
  11412=>"000000000",
  11413=>"011010011",
  11414=>"110011010",
  11415=>"100001001",
  11416=>"100000110",
  11417=>"101111101",
  11418=>"001101101",
  11419=>"010010111",
  11420=>"110011100",
  11421=>"100011001",
  11422=>"100011011",
  11423=>"100000000",
  11424=>"111101011",
  11425=>"111101110",
  11426=>"111110001",
  11427=>"000000011",
  11428=>"100001011",
  11429=>"110010011",
  11430=>"001010000",
  11431=>"100110101",
  11432=>"000010111",
  11433=>"111001000",
  11434=>"110110000",
  11435=>"100010110",
  11436=>"110100011",
  11437=>"110111111",
  11438=>"010000111",
  11439=>"001100010",
  11440=>"000100100",
  11441=>"001000111",
  11442=>"110101011",
  11443=>"110001000",
  11444=>"110100010",
  11445=>"001100011",
  11446=>"111001110",
  11447=>"000011110",
  11448=>"000111101",
  11449=>"011001100",
  11450=>"101111101",
  11451=>"110011011",
  11452=>"110011000",
  11453=>"111011110",
  11454=>"000110000",
  11455=>"000101111",
  11456=>"111101000",
  11457=>"001110010",
  11458=>"110110110",
  11459=>"110011110",
  11460=>"101110101",
  11461=>"000101110",
  11462=>"010101111",
  11463=>"010100101",
  11464=>"110011101",
  11465=>"001111110",
  11466=>"111100101",
  11467=>"011001110",
  11468=>"011000010",
  11469=>"101100111",
  11470=>"011001000",
  11471=>"010001011",
  11472=>"111110111",
  11473=>"011110100",
  11474=>"101111010",
  11475=>"001011000",
  11476=>"000001001",
  11477=>"001110100",
  11478=>"010101010",
  11479=>"001111110",
  11480=>"000110111",
  11481=>"100011100",
  11482=>"010010001",
  11483=>"001011111",
  11484=>"101111001",
  11485=>"011101111",
  11486=>"001000001",
  11487=>"010110000",
  11488=>"110001011",
  11489=>"100011001",
  11490=>"010100011",
  11491=>"001110111",
  11492=>"010010111",
  11493=>"010111011",
  11494=>"011101000",
  11495=>"101001010",
  11496=>"001001000",
  11497=>"100100100",
  11498=>"111010100",
  11499=>"001010000",
  11500=>"101001100",
  11501=>"111001000",
  11502=>"010101101",
  11503=>"111000111",
  11504=>"111010101",
  11505=>"101000001",
  11506=>"010001100",
  11507=>"000100101",
  11508=>"011010101",
  11509=>"011001100",
  11510=>"001100001",
  11511=>"000011101",
  11512=>"101111101",
  11513=>"000001100",
  11514=>"010111100",
  11515=>"110111101",
  11516=>"011111011",
  11517=>"101000010",
  11518=>"110000101",
  11519=>"000111111",
  11520=>"110100001",
  11521=>"110010001",
  11522=>"110101111",
  11523=>"101100011",
  11524=>"100010100",
  11525=>"010011010",
  11526=>"110000101",
  11527=>"000110000",
  11528=>"001010110",
  11529=>"111010010",
  11530=>"110001111",
  11531=>"101000111",
  11532=>"010000100",
  11533=>"110000110",
  11534=>"000000000",
  11535=>"111010111",
  11536=>"001001011",
  11537=>"001000001",
  11538=>"101111111",
  11539=>"011110111",
  11540=>"001111111",
  11541=>"100110111",
  11542=>"001000100",
  11543=>"100101100",
  11544=>"100010100",
  11545=>"000101101",
  11546=>"100000111",
  11547=>"011001011",
  11548=>"010110011",
  11549=>"010100111",
  11550=>"000110100",
  11551=>"110101110",
  11552=>"111010010",
  11553=>"101110001",
  11554=>"000000110",
  11555=>"011111101",
  11556=>"110101110",
  11557=>"111100100",
  11558=>"111100100",
  11559=>"011101000",
  11560=>"100110110",
  11561=>"001001001",
  11562=>"110000010",
  11563=>"010110010",
  11564=>"011111010",
  11565=>"101011111",
  11566=>"001111110",
  11567=>"011000111",
  11568=>"111001011",
  11569=>"000010001",
  11570=>"111011011",
  11571=>"111110001",
  11572=>"011101000",
  11573=>"000000011",
  11574=>"111000111",
  11575=>"010101111",
  11576=>"000100101",
  11577=>"000110000",
  11578=>"100000000",
  11579=>"110111110",
  11580=>"000000100",
  11581=>"111001000",
  11582=>"000000100",
  11583=>"101011011",
  11584=>"111100000",
  11585=>"010001110",
  11586=>"100000001",
  11587=>"001010011",
  11588=>"101110010",
  11589=>"111001001",
  11590=>"101000001",
  11591=>"001111000",
  11592=>"000101000",
  11593=>"010101100",
  11594=>"110110010",
  11595=>"000110011",
  11596=>"010101110",
  11597=>"110100000",
  11598=>"000110110",
  11599=>"001000010",
  11600=>"011100001",
  11601=>"001110100",
  11602=>"100111110",
  11603=>"000111000",
  11604=>"000110101",
  11605=>"110010111",
  11606=>"111010001",
  11607=>"111010110",
  11608=>"111111010",
  11609=>"000001000",
  11610=>"000101111",
  11611=>"001011100",
  11612=>"010100101",
  11613=>"010111110",
  11614=>"111101101",
  11615=>"000011001",
  11616=>"100011001",
  11617=>"101000110",
  11618=>"001000111",
  11619=>"000000000",
  11620=>"001100000",
  11621=>"111000100",
  11622=>"110101100",
  11623=>"001101001",
  11624=>"011101000",
  11625=>"111011001",
  11626=>"101100101",
  11627=>"001000110",
  11628=>"100110011",
  11629=>"000100111",
  11630=>"111010000",
  11631=>"001111111",
  11632=>"011001010",
  11633=>"000000100",
  11634=>"100010101",
  11635=>"000000100",
  11636=>"000001000",
  11637=>"101111011",
  11638=>"010001000",
  11639=>"101000001",
  11640=>"001011111",
  11641=>"111000101",
  11642=>"010000101",
  11643=>"010011101",
  11644=>"111100010",
  11645=>"100001010",
  11646=>"111010111",
  11647=>"111011101",
  11648=>"111101111",
  11649=>"111100000",
  11650=>"000011011",
  11651=>"101001101",
  11652=>"000111111",
  11653=>"010000001",
  11654=>"001101101",
  11655=>"000100110",
  11656=>"110000110",
  11657=>"001110100",
  11658=>"001010111",
  11659=>"100110001",
  11660=>"111111011",
  11661=>"111010001",
  11662=>"001110010",
  11663=>"110000010",
  11664=>"010001111",
  11665=>"010001011",
  11666=>"000010010",
  11667=>"100000000",
  11668=>"110001001",
  11669=>"001010100",
  11670=>"111110111",
  11671=>"111010001",
  11672=>"000101101",
  11673=>"100110101",
  11674=>"000110100",
  11675=>"011111011",
  11676=>"101011111",
  11677=>"010110000",
  11678=>"100100101",
  11679=>"000101100",
  11680=>"000000001",
  11681=>"110000000",
  11682=>"100101111",
  11683=>"010000001",
  11684=>"101011001",
  11685=>"110111000",
  11686=>"101111111",
  11687=>"000010010",
  11688=>"000010111",
  11689=>"111111101",
  11690=>"000100000",
  11691=>"111100111",
  11692=>"100010001",
  11693=>"110110111",
  11694=>"010001011",
  11695=>"100010100",
  11696=>"000010001",
  11697=>"010001001",
  11698=>"101101001",
  11699=>"110111010",
  11700=>"011101001",
  11701=>"011110100",
  11702=>"111100011",
  11703=>"111001001",
  11704=>"000001100",
  11705=>"010101111",
  11706=>"111000011",
  11707=>"111010011",
  11708=>"111101011",
  11709=>"101110000",
  11710=>"101001001",
  11711=>"011110100",
  11712=>"010010100",
  11713=>"001011011",
  11714=>"010101001",
  11715=>"010001010",
  11716=>"100001110",
  11717=>"110101011",
  11718=>"011100100",
  11719=>"000101000",
  11720=>"100000100",
  11721=>"001001100",
  11722=>"011010100",
  11723=>"000101111",
  11724=>"100110111",
  11725=>"100110100",
  11726=>"111101011",
  11727=>"011011011",
  11728=>"100001111",
  11729=>"111110110",
  11730=>"010011100",
  11731=>"110101101",
  11732=>"100000000",
  11733=>"101101011",
  11734=>"101000110",
  11735=>"011101010",
  11736=>"001110001",
  11737=>"010101110",
  11738=>"101101010",
  11739=>"000100111",
  11740=>"100011001",
  11741=>"011011000",
  11742=>"110000010",
  11743=>"000010011",
  11744=>"000010111",
  11745=>"000110010",
  11746=>"000001110",
  11747=>"000000001",
  11748=>"110111111",
  11749=>"000010101",
  11750=>"010111101",
  11751=>"011001111",
  11752=>"000111000",
  11753=>"010000110",
  11754=>"011000000",
  11755=>"011111111",
  11756=>"011101010",
  11757=>"101011111",
  11758=>"110011011",
  11759=>"101110000",
  11760=>"000000001",
  11761=>"001000000",
  11762=>"011100011",
  11763=>"101110100",
  11764=>"100011000",
  11765=>"011110100",
  11766=>"110100010",
  11767=>"010101011",
  11768=>"010001000",
  11769=>"110010001",
  11770=>"101111010",
  11771=>"011111111",
  11772=>"010001000",
  11773=>"101111001",
  11774=>"110111011",
  11775=>"101110100",
  11776=>"010011111",
  11777=>"100011101",
  11778=>"110111001",
  11779=>"000110011",
  11780=>"011101010",
  11781=>"011100011",
  11782=>"111101101",
  11783=>"000000001",
  11784=>"011011010",
  11785=>"111011000",
  11786=>"010101100",
  11787=>"111110100",
  11788=>"101111010",
  11789=>"010011010",
  11790=>"000101100",
  11791=>"000110011",
  11792=>"001001010",
  11793=>"000100111",
  11794=>"110010011",
  11795=>"010011100",
  11796=>"011001110",
  11797=>"011001011",
  11798=>"000001111",
  11799=>"100101010",
  11800=>"001010000",
  11801=>"011111110",
  11802=>"111101010",
  11803=>"101110100",
  11804=>"010000001",
  11805=>"011010110",
  11806=>"100111100",
  11807=>"000000001",
  11808=>"001101111",
  11809=>"000100011",
  11810=>"100011100",
  11811=>"001001100",
  11812=>"000000000",
  11813=>"110001010",
  11814=>"100011111",
  11815=>"110100101",
  11816=>"011100100",
  11817=>"001110000",
  11818=>"101111011",
  11819=>"001101100",
  11820=>"010010000",
  11821=>"010000010",
  11822=>"101011010",
  11823=>"010000001",
  11824=>"110111100",
  11825=>"011110000",
  11826=>"011111001",
  11827=>"100011001",
  11828=>"011111000",
  11829=>"111100000",
  11830=>"100010100",
  11831=>"001100110",
  11832=>"101101010",
  11833=>"000100110",
  11834=>"000010011",
  11835=>"011101000",
  11836=>"111110100",
  11837=>"001000111",
  11838=>"111010110",
  11839=>"111110001",
  11840=>"100010110",
  11841=>"110101000",
  11842=>"001111011",
  11843=>"111110111",
  11844=>"101000010",
  11845=>"001011001",
  11846=>"010111010",
  11847=>"001000100",
  11848=>"000100101",
  11849=>"010010110",
  11850=>"101100111",
  11851=>"110110110",
  11852=>"001011110",
  11853=>"001011010",
  11854=>"101000110",
  11855=>"111000101",
  11856=>"000001100",
  11857=>"001100100",
  11858=>"010100101",
  11859=>"001001101",
  11860=>"100101010",
  11861=>"000110000",
  11862=>"011101110",
  11863=>"111100100",
  11864=>"111101001",
  11865=>"000011010",
  11866=>"000101010",
  11867=>"000001001",
  11868=>"001000111",
  11869=>"100010000",
  11870=>"110101010",
  11871=>"100000011",
  11872=>"011000011",
  11873=>"010011101",
  11874=>"010000111",
  11875=>"111000011",
  11876=>"010100111",
  11877=>"100101010",
  11878=>"001101010",
  11879=>"111011111",
  11880=>"111001100",
  11881=>"100110011",
  11882=>"001011001",
  11883=>"110110001",
  11884=>"001010011",
  11885=>"010110100",
  11886=>"100000110",
  11887=>"101000001",
  11888=>"111001101",
  11889=>"101011111",
  11890=>"101011100",
  11891=>"110100010",
  11892=>"101001000",
  11893=>"101111101",
  11894=>"010010100",
  11895=>"000001111",
  11896=>"010110000",
  11897=>"000000011",
  11898=>"010111001",
  11899=>"100011111",
  11900=>"000000111",
  11901=>"001000110",
  11902=>"011101001",
  11903=>"010110101",
  11904=>"100001101",
  11905=>"010101001",
  11906=>"000101011",
  11907=>"111001100",
  11908=>"100000111",
  11909=>"010010011",
  11910=>"001110000",
  11911=>"000010110",
  11912=>"010100000",
  11913=>"111100011",
  11914=>"100110101",
  11915=>"001010111",
  11916=>"111111100",
  11917=>"111100110",
  11918=>"000001111",
  11919=>"000001000",
  11920=>"110110111",
  11921=>"010010011",
  11922=>"011100100",
  11923=>"100100010",
  11924=>"010001011",
  11925=>"110110010",
  11926=>"110110011",
  11927=>"100000010",
  11928=>"100011101",
  11929=>"000011011",
  11930=>"101010110",
  11931=>"101001111",
  11932=>"010110010",
  11933=>"111101011",
  11934=>"110101111",
  11935=>"000011001",
  11936=>"010001010",
  11937=>"000001111",
  11938=>"011011110",
  11939=>"101010110",
  11940=>"100011111",
  11941=>"001010110",
  11942=>"000010010",
  11943=>"101001000",
  11944=>"010101101",
  11945=>"011000010",
  11946=>"001100001",
  11947=>"110001000",
  11948=>"110110001",
  11949=>"000111010",
  11950=>"111111111",
  11951=>"001101011",
  11952=>"001000100",
  11953=>"101001111",
  11954=>"000110101",
  11955=>"111111110",
  11956=>"101001100",
  11957=>"100000000",
  11958=>"111000101",
  11959=>"111110011",
  11960=>"010000101",
  11961=>"011001101",
  11962=>"101110110",
  11963=>"001000001",
  11964=>"110011011",
  11965=>"110010000",
  11966=>"110111111",
  11967=>"001011000",
  11968=>"000110001",
  11969=>"100011000",
  11970=>"000001100",
  11971=>"001101001",
  11972=>"001001101",
  11973=>"010010000",
  11974=>"100001000",
  11975=>"001010011",
  11976=>"110100101",
  11977=>"011010111",
  11978=>"100001110",
  11979=>"110111101",
  11980=>"100010000",
  11981=>"010011011",
  11982=>"100000001",
  11983=>"000011000",
  11984=>"011111010",
  11985=>"010011111",
  11986=>"011011111",
  11987=>"101010101",
  11988=>"000000101",
  11989=>"000110000",
  11990=>"100001001",
  11991=>"100011101",
  11992=>"011000000",
  11993=>"101001011",
  11994=>"100010101",
  11995=>"100101100",
  11996=>"010011111",
  11997=>"010110110",
  11998=>"110110111",
  11999=>"100100111",
  12000=>"010000101",
  12001=>"011010000",
  12002=>"101110111",
  12003=>"010101101",
  12004=>"010111001",
  12005=>"110110100",
  12006=>"101001111",
  12007=>"010010010",
  12008=>"010111111",
  12009=>"001000010",
  12010=>"110100100",
  12011=>"101111010",
  12012=>"001000000",
  12013=>"011111101",
  12014=>"100111110",
  12015=>"001100010",
  12016=>"111001000",
  12017=>"000100000",
  12018=>"010100111",
  12019=>"100000100",
  12020=>"010100001",
  12021=>"001111011",
  12022=>"101000100",
  12023=>"100110000",
  12024=>"000011010",
  12025=>"111110010",
  12026=>"011111110",
  12027=>"000111001",
  12028=>"100000011",
  12029=>"111100001",
  12030=>"001010100",
  12031=>"111011111",
  12032=>"100010010",
  12033=>"101100011",
  12034=>"010100111",
  12035=>"001001101",
  12036=>"010001110",
  12037=>"001000011",
  12038=>"010010101",
  12039=>"110011000",
  12040=>"101000000",
  12041=>"100010111",
  12042=>"011100110",
  12043=>"111111111",
  12044=>"101000110",
  12045=>"100011100",
  12046=>"111100101",
  12047=>"001110100",
  12048=>"111101010",
  12049=>"111101101",
  12050=>"110110111",
  12051=>"101001101",
  12052=>"101000110",
  12053=>"000011011",
  12054=>"001001000",
  12055=>"100111001",
  12056=>"001101101",
  12057=>"110111000",
  12058=>"000000100",
  12059=>"111111011",
  12060=>"000101011",
  12061=>"010011100",
  12062=>"001110000",
  12063=>"111110100",
  12064=>"111001101",
  12065=>"011111101",
  12066=>"001100011",
  12067=>"010100110",
  12068=>"000110000",
  12069=>"011100010",
  12070=>"110101000",
  12071=>"010100000",
  12072=>"111011101",
  12073=>"010000011",
  12074=>"101101001",
  12075=>"111011110",
  12076=>"011110100",
  12077=>"110000001",
  12078=>"100101000",
  12079=>"000001100",
  12080=>"110010100",
  12081=>"001010011",
  12082=>"001100101",
  12083=>"101111001",
  12084=>"000100000",
  12085=>"111001010",
  12086=>"011001001",
  12087=>"011111100",
  12088=>"011100011",
  12089=>"010011110",
  12090=>"010110111",
  12091=>"010110100",
  12092=>"011011100",
  12093=>"000110100",
  12094=>"011000010",
  12095=>"010110100",
  12096=>"010110101",
  12097=>"010001100",
  12098=>"010000001",
  12099=>"111100111",
  12100=>"010111010",
  12101=>"011000110",
  12102=>"110100110",
  12103=>"000111111",
  12104=>"110110010",
  12105=>"111101000",
  12106=>"011110011",
  12107=>"000100110",
  12108=>"010010000",
  12109=>"100110110",
  12110=>"010111000",
  12111=>"100011111",
  12112=>"111001101",
  12113=>"001101100",
  12114=>"010001000",
  12115=>"000011100",
  12116=>"001010110",
  12117=>"111000001",
  12118=>"110010000",
  12119=>"111001001",
  12120=>"000011110",
  12121=>"000100101",
  12122=>"000001111",
  12123=>"110010100",
  12124=>"100110000",
  12125=>"000001000",
  12126=>"011011010",
  12127=>"000100001",
  12128=>"001111010",
  12129=>"110000101",
  12130=>"001110110",
  12131=>"011101110",
  12132=>"011011111",
  12133=>"011100110",
  12134=>"111111011",
  12135=>"001011000",
  12136=>"100100100",
  12137=>"110111101",
  12138=>"001000111",
  12139=>"010110011",
  12140=>"001111110",
  12141=>"001010111",
  12142=>"111100000",
  12143=>"101101111",
  12144=>"010101100",
  12145=>"101001101",
  12146=>"101001000",
  12147=>"010000100",
  12148=>"000000000",
  12149=>"101100001",
  12150=>"111101110",
  12151=>"010011101",
  12152=>"000100011",
  12153=>"101001100",
  12154=>"100110010",
  12155=>"110111111",
  12156=>"000110111",
  12157=>"010111100",
  12158=>"100101011",
  12159=>"010110101",
  12160=>"111111110",
  12161=>"010011110",
  12162=>"011000011",
  12163=>"000100110",
  12164=>"011000001",
  12165=>"001010111",
  12166=>"010000000",
  12167=>"010011101",
  12168=>"100101010",
  12169=>"110110100",
  12170=>"110010010",
  12171=>"000001100",
  12172=>"001100100",
  12173=>"110010111",
  12174=>"101011111",
  12175=>"101001011",
  12176=>"010010111",
  12177=>"111111010",
  12178=>"001101100",
  12179=>"000111110",
  12180=>"110101000",
  12181=>"010110010",
  12182=>"000001000",
  12183=>"001110111",
  12184=>"011110100",
  12185=>"001010001",
  12186=>"010010101",
  12187=>"100110011",
  12188=>"101000010",
  12189=>"000011011",
  12190=>"000000111",
  12191=>"100001011",
  12192=>"110101001",
  12193=>"000011000",
  12194=>"110011001",
  12195=>"100100000",
  12196=>"000111111",
  12197=>"111101000",
  12198=>"100110111",
  12199=>"001000100",
  12200=>"101011110",
  12201=>"001111001",
  12202=>"111111000",
  12203=>"110100100",
  12204=>"110100100",
  12205=>"110111011",
  12206=>"001011111",
  12207=>"001001110",
  12208=>"011010000",
  12209=>"011001111",
  12210=>"101000010",
  12211=>"000011010",
  12212=>"001001001",
  12213=>"001010101",
  12214=>"100111100",
  12215=>"100010100",
  12216=>"010111100",
  12217=>"111010101",
  12218=>"100111100",
  12219=>"011000110",
  12220=>"110110101",
  12221=>"111101101",
  12222=>"011111001",
  12223=>"101010001",
  12224=>"101011111",
  12225=>"111011001",
  12226=>"110000001",
  12227=>"010000010",
  12228=>"111100110",
  12229=>"000010111",
  12230=>"011100000",
  12231=>"111010101",
  12232=>"101011001",
  12233=>"000100100",
  12234=>"011000001",
  12235=>"010001101",
  12236=>"110110011",
  12237=>"111111111",
  12238=>"010000001",
  12239=>"000101111",
  12240=>"001111100",
  12241=>"001001101",
  12242=>"001100001",
  12243=>"110101000",
  12244=>"001001101",
  12245=>"001000001",
  12246=>"000100010",
  12247=>"110010110",
  12248=>"111000000",
  12249=>"100111100",
  12250=>"111001000",
  12251=>"101110000",
  12252=>"110101100",
  12253=>"000111100",
  12254=>"000010000",
  12255=>"110101000",
  12256=>"010100000",
  12257=>"110101000",
  12258=>"111111110",
  12259=>"111100001",
  12260=>"001010010",
  12261=>"001011010",
  12262=>"001001101",
  12263=>"101001011",
  12264=>"101011001",
  12265=>"110011011",
  12266=>"100100111",
  12267=>"100011000",
  12268=>"001101001",
  12269=>"100111111",
  12270=>"101010101",
  12271=>"000110111",
  12272=>"001001011",
  12273=>"010001010",
  12274=>"010110011",
  12275=>"011100000",
  12276=>"010111000",
  12277=>"000101100",
  12278=>"000110100",
  12279=>"011111111",
  12280=>"011001101",
  12281=>"010100110",
  12282=>"011010001",
  12283=>"111011001",
  12284=>"011111101",
  12285=>"101101011",
  12286=>"010001011",
  12287=>"110011000",
  12288=>"000001001",
  12289=>"110100101",
  12290=>"100111100",
  12291=>"000111110",
  12292=>"001010011",
  12293=>"011100011",
  12294=>"101000010",
  12295=>"000000001",
  12296=>"111010011",
  12297=>"000000000",
  12298=>"111110111",
  12299=>"111111001",
  12300=>"111001111",
  12301=>"110101111",
  12302=>"110011001",
  12303=>"101001101",
  12304=>"110000000",
  12305=>"001000011",
  12306=>"111000010",
  12307=>"110101010",
  12308=>"101000100",
  12309=>"111000111",
  12310=>"110111011",
  12311=>"001011010",
  12312=>"111100000",
  12313=>"110011001",
  12314=>"100100110",
  12315=>"000111010",
  12316=>"001110110",
  12317=>"111010111",
  12318=>"001011100",
  12319=>"000010101",
  12320=>"000100000",
  12321=>"101100111",
  12322=>"101101110",
  12323=>"101101000",
  12324=>"011011001",
  12325=>"000110001",
  12326=>"000101111",
  12327=>"101111111",
  12328=>"010010010",
  12329=>"010011111",
  12330=>"011001100",
  12331=>"101101100",
  12332=>"011011100",
  12333=>"010011011",
  12334=>"011001010",
  12335=>"100100101",
  12336=>"000101100",
  12337=>"110111101",
  12338=>"101110010",
  12339=>"000010010",
  12340=>"000011000",
  12341=>"011001111",
  12342=>"111000111",
  12343=>"110001001",
  12344=>"000111011",
  12345=>"000100011",
  12346=>"001100000",
  12347=>"100011100",
  12348=>"010010001",
  12349=>"111111011",
  12350=>"010011110",
  12351=>"001111110",
  12352=>"001000011",
  12353=>"011001011",
  12354=>"110011010",
  12355=>"110111011",
  12356=>"101101011",
  12357=>"010110100",
  12358=>"101110111",
  12359=>"000011010",
  12360=>"001101111",
  12361=>"111100111",
  12362=>"110101000",
  12363=>"111011011",
  12364=>"001101111",
  12365=>"100100011",
  12366=>"111111111",
  12367=>"001000010",
  12368=>"110111001",
  12369=>"111111100",
  12370=>"010000110",
  12371=>"000010001",
  12372=>"110111001",
  12373=>"101111110",
  12374=>"011010101",
  12375=>"111010101",
  12376=>"000000011",
  12377=>"111001101",
  12378=>"001010001",
  12379=>"110101101",
  12380=>"001001000",
  12381=>"100000011",
  12382=>"100011001",
  12383=>"100010001",
  12384=>"000000010",
  12385=>"010000011",
  12386=>"100101110",
  12387=>"010100111",
  12388=>"010001000",
  12389=>"000000110",
  12390=>"110111010",
  12391=>"111101101",
  12392=>"101110100",
  12393=>"000010000",
  12394=>"110111100",
  12395=>"010001101",
  12396=>"000100111",
  12397=>"100010011",
  12398=>"100101001",
  12399=>"001100111",
  12400=>"100101111",
  12401=>"111111111",
  12402=>"111010000",
  12403=>"000101011",
  12404=>"100001110",
  12405=>"111001100",
  12406=>"101011011",
  12407=>"101110001",
  12408=>"100011100",
  12409=>"000110001",
  12410=>"001001111",
  12411=>"111011101",
  12412=>"101101001",
  12413=>"110111011",
  12414=>"011110000",
  12415=>"100010011",
  12416=>"000011000",
  12417=>"100000001",
  12418=>"000010110",
  12419=>"101110111",
  12420=>"010011110",
  12421=>"111101101",
  12422=>"111100101",
  12423=>"110100110",
  12424=>"011100010",
  12425=>"100101000",
  12426=>"011011111",
  12427=>"011111000",
  12428=>"001000111",
  12429=>"000100011",
  12430=>"000101001",
  12431=>"100001110",
  12432=>"101111010",
  12433=>"011001101",
  12434=>"100001001",
  12435=>"000011010",
  12436=>"100001011",
  12437=>"000110010",
  12438=>"000000111",
  12439=>"111011010",
  12440=>"101101011",
  12441=>"010101110",
  12442=>"111100000",
  12443=>"011010111",
  12444=>"111000111",
  12445=>"111100101",
  12446=>"010011111",
  12447=>"111010011",
  12448=>"110101010",
  12449=>"001110000",
  12450=>"000100001",
  12451=>"111110110",
  12452=>"100111111",
  12453=>"011110101",
  12454=>"101001010",
  12455=>"000100111",
  12456=>"001000011",
  12457=>"010101110",
  12458=>"001011011",
  12459=>"000111110",
  12460=>"011100010",
  12461=>"100100101",
  12462=>"000100000",
  12463=>"111111101",
  12464=>"110001001",
  12465=>"001010101",
  12466=>"011101100",
  12467=>"011010101",
  12468=>"010110000",
  12469=>"110001011",
  12470=>"000001011",
  12471=>"001001000",
  12472=>"110100010",
  12473=>"110101010",
  12474=>"010101101",
  12475=>"110111100",
  12476=>"011011100",
  12477=>"101101001",
  12478=>"100110101",
  12479=>"110111110",
  12480=>"101110010",
  12481=>"001011010",
  12482=>"110100010",
  12483=>"111000110",
  12484=>"100000001",
  12485=>"101000110",
  12486=>"011110111",
  12487=>"011001010",
  12488=>"011011110",
  12489=>"111101111",
  12490=>"001010111",
  12491=>"100000111",
  12492=>"101000101",
  12493=>"111000100",
  12494=>"011111110",
  12495=>"011110010",
  12496=>"010100010",
  12497=>"111111100",
  12498=>"100000001",
  12499=>"011110011",
  12500=>"001000100",
  12501=>"000001100",
  12502=>"110001011",
  12503=>"111000101",
  12504=>"000010001",
  12505=>"011010001",
  12506=>"000000111",
  12507=>"011110110",
  12508=>"001100111",
  12509=>"110010001",
  12510=>"011111111",
  12511=>"100011001",
  12512=>"110110110",
  12513=>"000111111",
  12514=>"000111100",
  12515=>"000100001",
  12516=>"111110111",
  12517=>"110000110",
  12518=>"000011100",
  12519=>"110100011",
  12520=>"001001011",
  12521=>"000101010",
  12522=>"111111001",
  12523=>"010001101",
  12524=>"111001010",
  12525=>"010011110",
  12526=>"011111001",
  12527=>"111101001",
  12528=>"010100100",
  12529=>"100111111",
  12530=>"110000000",
  12531=>"000110000",
  12532=>"101011000",
  12533=>"011010001",
  12534=>"101101100",
  12535=>"100110010",
  12536=>"001110011",
  12537=>"000000100",
  12538=>"000001101",
  12539=>"101011110",
  12540=>"111001111",
  12541=>"101111001",
  12542=>"110110011",
  12543=>"101001110",
  12544=>"101010101",
  12545=>"111110100",
  12546=>"001010000",
  12547=>"110010111",
  12548=>"111110010",
  12549=>"100110101",
  12550=>"100001001",
  12551=>"100110011",
  12552=>"010101001",
  12553=>"001000000",
  12554=>"100010000",
  12555=>"000000001",
  12556=>"001110001",
  12557=>"101111010",
  12558=>"100011111",
  12559=>"101101010",
  12560=>"101111011",
  12561=>"101010011",
  12562=>"010110000",
  12563=>"010101001",
  12564=>"011011111",
  12565=>"011100010",
  12566=>"100010111",
  12567=>"000011110",
  12568=>"111111011",
  12569=>"101110010",
  12570=>"000010000",
  12571=>"010000100",
  12572=>"101001101",
  12573=>"010000000",
  12574=>"110111101",
  12575=>"110101010",
  12576=>"000010111",
  12577=>"100111101",
  12578=>"101011110",
  12579=>"100011111",
  12580=>"000101100",
  12581=>"111111100",
  12582=>"000100000",
  12583=>"001100011",
  12584=>"110100010",
  12585=>"111001101",
  12586=>"100100100",
  12587=>"010101100",
  12588=>"000101001",
  12589=>"101110010",
  12590=>"111010010",
  12591=>"000111100",
  12592=>"111111101",
  12593=>"111000010",
  12594=>"001000011",
  12595=>"110010111",
  12596=>"101100100",
  12597=>"011011000",
  12598=>"010001001",
  12599=>"000001101",
  12600=>"010011110",
  12601=>"101100111",
  12602=>"100011111",
  12603=>"100001110",
  12604=>"010100111",
  12605=>"000110001",
  12606=>"100111110",
  12607=>"110111010",
  12608=>"110100100",
  12609=>"100100011",
  12610=>"011110100",
  12611=>"010110100",
  12612=>"010011111",
  12613=>"110100011",
  12614=>"100100011",
  12615=>"011011110",
  12616=>"111011101",
  12617=>"000100001",
  12618=>"000101110",
  12619=>"000000010",
  12620=>"110110110",
  12621=>"010101010",
  12622=>"101110101",
  12623=>"000000111",
  12624=>"111000101",
  12625=>"000001011",
  12626=>"001011100",
  12627=>"111111001",
  12628=>"001010110",
  12629=>"110001110",
  12630=>"110110100",
  12631=>"100001000",
  12632=>"010000011",
  12633=>"011001100",
  12634=>"101110010",
  12635=>"101100011",
  12636=>"000100100",
  12637=>"101011011",
  12638=>"011001100",
  12639=>"011111001",
  12640=>"110100110",
  12641=>"110011101",
  12642=>"101110100",
  12643=>"111000101",
  12644=>"000010000",
  12645=>"000111110",
  12646=>"001101111",
  12647=>"011111101",
  12648=>"111101001",
  12649=>"100011011",
  12650=>"111000001",
  12651=>"100001010",
  12652=>"110110111",
  12653=>"111100011",
  12654=>"111110100",
  12655=>"001010101",
  12656=>"000011100",
  12657=>"010100011",
  12658=>"101010000",
  12659=>"110100110",
  12660=>"111010111",
  12661=>"101101001",
  12662=>"111101000",
  12663=>"000101111",
  12664=>"100010000",
  12665=>"100111001",
  12666=>"000011110",
  12667=>"001110000",
  12668=>"100001000",
  12669=>"111111101",
  12670=>"111011011",
  12671=>"000001100",
  12672=>"000100111",
  12673=>"011001011",
  12674=>"011011100",
  12675=>"011101111",
  12676=>"111110111",
  12677=>"000000110",
  12678=>"110111111",
  12679=>"101000000",
  12680=>"010000101",
  12681=>"110101011",
  12682=>"100101110",
  12683=>"001110101",
  12684=>"011111010",
  12685=>"101110111",
  12686=>"001001110",
  12687=>"010110011",
  12688=>"011011000",
  12689=>"000001100",
  12690=>"001100101",
  12691=>"110100001",
  12692=>"110000111",
  12693=>"110000000",
  12694=>"100110010",
  12695=>"101100101",
  12696=>"001001011",
  12697=>"000000000",
  12698=>"011000000",
  12699=>"111000000",
  12700=>"111111110",
  12701=>"100101110",
  12702=>"110100110",
  12703=>"110100000",
  12704=>"010100101",
  12705=>"111000001",
  12706=>"111101001",
  12707=>"110001010",
  12708=>"100000110",
  12709=>"011000111",
  12710=>"001000000",
  12711=>"010101101",
  12712=>"100001111",
  12713=>"001101000",
  12714=>"011110100",
  12715=>"011010101",
  12716=>"100000110",
  12717=>"111000010",
  12718=>"110010110",
  12719=>"000010000",
  12720=>"100010001",
  12721=>"111100010",
  12722=>"110111000",
  12723=>"100010100",
  12724=>"000100101",
  12725=>"111100100",
  12726=>"001101101",
  12727=>"001110100",
  12728=>"111111010",
  12729=>"000011101",
  12730=>"000000111",
  12731=>"010010101",
  12732=>"110001000",
  12733=>"111101100",
  12734=>"000001110",
  12735=>"011000000",
  12736=>"011010000",
  12737=>"001101111",
  12738=>"001110111",
  12739=>"110001001",
  12740=>"110010001",
  12741=>"011001101",
  12742=>"110110111",
  12743=>"101010011",
  12744=>"110010010",
  12745=>"000100011",
  12746=>"000011111",
  12747=>"001000111",
  12748=>"111101010",
  12749=>"011001100",
  12750=>"111110110",
  12751=>"001011101",
  12752=>"110100101",
  12753=>"100111011",
  12754=>"001011110",
  12755=>"101000000",
  12756=>"001011111",
  12757=>"000000111",
  12758=>"111110111",
  12759=>"001110011",
  12760=>"000111101",
  12761=>"010100010",
  12762=>"110010001",
  12763=>"011011001",
  12764=>"001101111",
  12765=>"101010111",
  12766=>"110101001",
  12767=>"111100000",
  12768=>"110100010",
  12769=>"101011101",
  12770=>"110010000",
  12771=>"001100101",
  12772=>"010000010",
  12773=>"111100111",
  12774=>"100011100",
  12775=>"000111011",
  12776=>"010011000",
  12777=>"001010011",
  12778=>"101000001",
  12779=>"001111001",
  12780=>"000011000",
  12781=>"001100101",
  12782=>"011010111",
  12783=>"110011100",
  12784=>"010011010",
  12785=>"110001001",
  12786=>"011010010",
  12787=>"100001111",
  12788=>"010010100",
  12789=>"000101010",
  12790=>"111100110",
  12791=>"101110010",
  12792=>"000100001",
  12793=>"000000011",
  12794=>"010000011",
  12795=>"111111010",
  12796=>"100001001",
  12797=>"010110100",
  12798=>"010100011",
  12799=>"111100010",
  12800=>"011110001",
  12801=>"110111011",
  12802=>"101011111",
  12803=>"101100100",
  12804=>"111100000",
  12805=>"100011111",
  12806=>"111111011",
  12807=>"100001100",
  12808=>"100111001",
  12809=>"001101111",
  12810=>"111101100",
  12811=>"000101001",
  12812=>"001111001",
  12813=>"001110000",
  12814=>"010001000",
  12815=>"100101000",
  12816=>"001010010",
  12817=>"011111111",
  12818=>"000100011",
  12819=>"101000011",
  12820=>"100010011",
  12821=>"101111100",
  12822=>"110100010",
  12823=>"001100000",
  12824=>"001110111",
  12825=>"100101111",
  12826=>"011011001",
  12827=>"010011011",
  12828=>"011100100",
  12829=>"001000110",
  12830=>"011011101",
  12831=>"100101001",
  12832=>"001101001",
  12833=>"100010101",
  12834=>"010110100",
  12835=>"101011110",
  12836=>"111110111",
  12837=>"110100101",
  12838=>"011100000",
  12839=>"101111001",
  12840=>"101110111",
  12841=>"111110101",
  12842=>"110101100",
  12843=>"011101011",
  12844=>"001000111",
  12845=>"000101000",
  12846=>"110001110",
  12847=>"111110010",
  12848=>"100001111",
  12849=>"111111111",
  12850=>"111101110",
  12851=>"101101001",
  12852=>"111101100",
  12853=>"011000100",
  12854=>"010000101",
  12855=>"111001100",
  12856=>"110101101",
  12857=>"101000011",
  12858=>"010101110",
  12859=>"100100111",
  12860=>"001100111",
  12861=>"010100100",
  12862=>"111101110",
  12863=>"001111110",
  12864=>"101001001",
  12865=>"100110101",
  12866=>"000101111",
  12867=>"001011010",
  12868=>"110100001",
  12869=>"010100011",
  12870=>"001011111",
  12871=>"001100100",
  12872=>"000100010",
  12873=>"100100011",
  12874=>"000111001",
  12875=>"111101000",
  12876=>"000000001",
  12877=>"111111001",
  12878=>"111101111",
  12879=>"011110100",
  12880=>"100100110",
  12881=>"111011101",
  12882=>"111010000",
  12883=>"001000110",
  12884=>"010000001",
  12885=>"000011100",
  12886=>"001001110",
  12887=>"101011001",
  12888=>"110011000",
  12889=>"111011100",
  12890=>"110010110",
  12891=>"110010010",
  12892=>"110011101",
  12893=>"001001000",
  12894=>"101101110",
  12895=>"100010000",
  12896=>"110110010",
  12897=>"000001010",
  12898=>"011110111",
  12899=>"110111000",
  12900=>"011111010",
  12901=>"100011101",
  12902=>"011111000",
  12903=>"100010011",
  12904=>"011010110",
  12905=>"110010011",
  12906=>"111110001",
  12907=>"010010010",
  12908=>"000101001",
  12909=>"001001111",
  12910=>"101111001",
  12911=>"100111101",
  12912=>"101100010",
  12913=>"000000010",
  12914=>"001111010",
  12915=>"111001001",
  12916=>"011111010",
  12917=>"101011100",
  12918=>"101010101",
  12919=>"001111101",
  12920=>"001000011",
  12921=>"010111110",
  12922=>"100101100",
  12923=>"001001000",
  12924=>"111010001",
  12925=>"010110000",
  12926=>"000001111",
  12927=>"100110110",
  12928=>"101111100",
  12929=>"001000110",
  12930=>"000001101",
  12931=>"010010010",
  12932=>"001001100",
  12933=>"101010100",
  12934=>"001110001",
  12935=>"000110111",
  12936=>"010011001",
  12937=>"010110010",
  12938=>"100101110",
  12939=>"000000101",
  12940=>"111011111",
  12941=>"101010000",
  12942=>"000110100",
  12943=>"111101111",
  12944=>"010111100",
  12945=>"011101111",
  12946=>"011110011",
  12947=>"100000100",
  12948=>"000010100",
  12949=>"101011100",
  12950=>"011001001",
  12951=>"101100000",
  12952=>"001010001",
  12953=>"001000000",
  12954=>"101011011",
  12955=>"110100111",
  12956=>"111011000",
  12957=>"000000010",
  12958=>"101011111",
  12959=>"100110100",
  12960=>"100011001",
  12961=>"000000010",
  12962=>"101000111",
  12963=>"010101100",
  12964=>"011010000",
  12965=>"100111101",
  12966=>"111100111",
  12967=>"110000100",
  12968=>"110111000",
  12969=>"000010001",
  12970=>"000000101",
  12971=>"110111010",
  12972=>"110001100",
  12973=>"011100000",
  12974=>"101111110",
  12975=>"011111011",
  12976=>"111001000",
  12977=>"000010100",
  12978=>"010100000",
  12979=>"000001011",
  12980=>"011000110",
  12981=>"110110001",
  12982=>"001000110",
  12983=>"001011000",
  12984=>"100011011",
  12985=>"110000101",
  12986=>"111001001",
  12987=>"011110111",
  12988=>"111111100",
  12989=>"000001100",
  12990=>"010001100",
  12991=>"010111100",
  12992=>"000010010",
  12993=>"111000001",
  12994=>"001100000",
  12995=>"111110011",
  12996=>"001110000",
  12997=>"110100110",
  12998=>"010100101",
  12999=>"101110011",
  13000=>"000000000",
  13001=>"001011101",
  13002=>"011010101",
  13003=>"000111000",
  13004=>"000000001",
  13005=>"100110110",
  13006=>"110110011",
  13007=>"010000110",
  13008=>"011010001",
  13009=>"000110011",
  13010=>"011010000",
  13011=>"000100111",
  13012=>"111101000",
  13013=>"000111011",
  13014=>"110000000",
  13015=>"011111100",
  13016=>"000110111",
  13017=>"110100101",
  13018=>"010000011",
  13019=>"100111010",
  13020=>"101101011",
  13021=>"000010000",
  13022=>"101100100",
  13023=>"101010001",
  13024=>"100011000",
  13025=>"011001011",
  13026=>"011110010",
  13027=>"100010101",
  13028=>"110011000",
  13029=>"100110101",
  13030=>"101101001",
  13031=>"000111101",
  13032=>"001000001",
  13033=>"010011001",
  13034=>"010100110",
  13035=>"101010010",
  13036=>"000010001",
  13037=>"000100100",
  13038=>"000111100",
  13039=>"000100010",
  13040=>"001110101",
  13041=>"001111101",
  13042=>"011001001",
  13043=>"101001100",
  13044=>"101001011",
  13045=>"011110101",
  13046=>"010000001",
  13047=>"100111101",
  13048=>"101100100",
  13049=>"010001001",
  13050=>"100010110",
  13051=>"000110010",
  13052=>"001111111",
  13053=>"010000101",
  13054=>"000001000",
  13055=>"010101011",
  13056=>"010000011",
  13057=>"001011000",
  13058=>"001110000",
  13059=>"000010111",
  13060=>"100110000",
  13061=>"010001100",
  13062=>"000100110",
  13063=>"101100001",
  13064=>"011011101",
  13065=>"010101110",
  13066=>"111110111",
  13067=>"111000010",
  13068=>"100000000",
  13069=>"110010101",
  13070=>"110110001",
  13071=>"000000011",
  13072=>"110110011",
  13073=>"010110001",
  13074=>"101010010",
  13075=>"001011100",
  13076=>"001010001",
  13077=>"001000111",
  13078=>"100010101",
  13079=>"100111110",
  13080=>"000010011",
  13081=>"010101001",
  13082=>"100010111",
  13083=>"010010000",
  13084=>"000010000",
  13085=>"100001001",
  13086=>"111110100",
  13087=>"000011100",
  13088=>"100001110",
  13089=>"100000011",
  13090=>"100010001",
  13091=>"001001000",
  13092=>"001100000",
  13093=>"000001011",
  13094=>"111100000",
  13095=>"011000010",
  13096=>"101110011",
  13097=>"100010000",
  13098=>"010010010",
  13099=>"100000100",
  13100=>"010100110",
  13101=>"011010111",
  13102=>"010000110",
  13103=>"111010101",
  13104=>"100001111",
  13105=>"111010101",
  13106=>"011010101",
  13107=>"110110111",
  13108=>"100110011",
  13109=>"001001100",
  13110=>"100000000",
  13111=>"101101111",
  13112=>"011101100",
  13113=>"000101011",
  13114=>"001101010",
  13115=>"111111001",
  13116=>"000010110",
  13117=>"000011111",
  13118=>"111100100",
  13119=>"011010001",
  13120=>"100100110",
  13121=>"011110111",
  13122=>"111101101",
  13123=>"111101000",
  13124=>"000011110",
  13125=>"000011011",
  13126=>"111001101",
  13127=>"110111111",
  13128=>"000111000",
  13129=>"100001000",
  13130=>"100110101",
  13131=>"000001000",
  13132=>"001001001",
  13133=>"010001110",
  13134=>"000111010",
  13135=>"111011000",
  13136=>"011011000",
  13137=>"111011111",
  13138=>"000101000",
  13139=>"011000010",
  13140=>"000010000",
  13141=>"111000111",
  13142=>"110001100",
  13143=>"010000100",
  13144=>"010001101",
  13145=>"001110010",
  13146=>"011001001",
  13147=>"000111111",
  13148=>"010010100",
  13149=>"110011001",
  13150=>"110010001",
  13151=>"001000111",
  13152=>"011111100",
  13153=>"100011101",
  13154=>"000000111",
  13155=>"010011101",
  13156=>"111101011",
  13157=>"100010001",
  13158=>"011110000",
  13159=>"100100111",
  13160=>"010001000",
  13161=>"111111111",
  13162=>"111110001",
  13163=>"011100001",
  13164=>"011111001",
  13165=>"110100010",
  13166=>"000000100",
  13167=>"111010001",
  13168=>"110011101",
  13169=>"111101110",
  13170=>"000100001",
  13171=>"110100011",
  13172=>"011100100",
  13173=>"001101111",
  13174=>"100110101",
  13175=>"011111011",
  13176=>"001111011",
  13177=>"100100000",
  13178=>"000100001",
  13179=>"001110100",
  13180=>"001100001",
  13181=>"001111011",
  13182=>"010001010",
  13183=>"001001101",
  13184=>"101010001",
  13185=>"010001001",
  13186=>"101010011",
  13187=>"000011000",
  13188=>"111011011",
  13189=>"000010100",
  13190=>"101001010",
  13191=>"101011000",
  13192=>"010110100",
  13193=>"010111101",
  13194=>"001001010",
  13195=>"001000000",
  13196=>"111111000",
  13197=>"111100011",
  13198=>"111110101",
  13199=>"010111111",
  13200=>"110011001",
  13201=>"111111111",
  13202=>"100110101",
  13203=>"110010001",
  13204=>"000101111",
  13205=>"100111001",
  13206=>"000111111",
  13207=>"101000000",
  13208=>"011111011",
  13209=>"110010110",
  13210=>"000110110",
  13211=>"100110111",
  13212=>"010000011",
  13213=>"001111111",
  13214=>"001011101",
  13215=>"011000100",
  13216=>"100101001",
  13217=>"001101011",
  13218=>"011111111",
  13219=>"100011100",
  13220=>"111111111",
  13221=>"110101101",
  13222=>"000000010",
  13223=>"011000000",
  13224=>"100011100",
  13225=>"100001011",
  13226=>"111100111",
  13227=>"101011000",
  13228=>"111011010",
  13229=>"101111010",
  13230=>"000100111",
  13231=>"001111111",
  13232=>"101001011",
  13233=>"100111100",
  13234=>"000110101",
  13235=>"101010100",
  13236=>"000110011",
  13237=>"010110111",
  13238=>"000011100",
  13239=>"111001001",
  13240=>"101010110",
  13241=>"101110010",
  13242=>"110010010",
  13243=>"100111001",
  13244=>"010110110",
  13245=>"010010101",
  13246=>"101001111",
  13247=>"010111001",
  13248=>"100001000",
  13249=>"101001001",
  13250=>"111000001",
  13251=>"001111101",
  13252=>"100001111",
  13253=>"011011100",
  13254=>"100101111",
  13255=>"001000000",
  13256=>"101010010",
  13257=>"011011100",
  13258=>"101111011",
  13259=>"000001000",
  13260=>"110011101",
  13261=>"001100000",
  13262=>"101111000",
  13263=>"100010010",
  13264=>"000110101",
  13265=>"001000001",
  13266=>"000000000",
  13267=>"000111110",
  13268=>"000110100",
  13269=>"000001001",
  13270=>"101001010",
  13271=>"001011011",
  13272=>"010111101",
  13273=>"110000001",
  13274=>"110011100",
  13275=>"000101011",
  13276=>"111101100",
  13277=>"011001000",
  13278=>"001111000",
  13279=>"000101010",
  13280=>"010001000",
  13281=>"111100111",
  13282=>"000011101",
  13283=>"000000110",
  13284=>"011111111",
  13285=>"010001010",
  13286=>"001000110",
  13287=>"110001110",
  13288=>"011001111",
  13289=>"010100101",
  13290=>"101010000",
  13291=>"010011010",
  13292=>"111011111",
  13293=>"100000000",
  13294=>"100110101",
  13295=>"101001101",
  13296=>"011010000",
  13297=>"000110100",
  13298=>"100001100",
  13299=>"110100001",
  13300=>"111110101",
  13301=>"010110000",
  13302=>"100100010",
  13303=>"100011000",
  13304=>"101011111",
  13305=>"011011111",
  13306=>"001110101",
  13307=>"110001101",
  13308=>"011110000",
  13309=>"001001000",
  13310=>"000010100",
  13311=>"010001000",
  13312=>"011011000",
  13313=>"100001101",
  13314=>"011001010",
  13315=>"010101011",
  13316=>"010110111",
  13317=>"010010101",
  13318=>"001011111",
  13319=>"111001011",
  13320=>"110101101",
  13321=>"111000110",
  13322=>"011001111",
  13323=>"000111001",
  13324=>"111101111",
  13325=>"001010010",
  13326=>"111001001",
  13327=>"001001110",
  13328=>"110111001",
  13329=>"000100111",
  13330=>"000011000",
  13331=>"000001000",
  13332=>"010101011",
  13333=>"000110100",
  13334=>"001100110",
  13335=>"101101000",
  13336=>"101100100",
  13337=>"001001000",
  13338=>"001110100",
  13339=>"011011001",
  13340=>"111011101",
  13341=>"101110101",
  13342=>"101011000",
  13343=>"100100010",
  13344=>"010000100",
  13345=>"010000011",
  13346=>"100001110",
  13347=>"101111101",
  13348=>"010111001",
  13349=>"001001111",
  13350=>"011011001",
  13351=>"100110101",
  13352=>"101010111",
  13353=>"010100000",
  13354=>"001000011",
  13355=>"000101111",
  13356=>"000110110",
  13357=>"111110100",
  13358=>"000001101",
  13359=>"001001011",
  13360=>"010111001",
  13361=>"011100111",
  13362=>"000010011",
  13363=>"101101100",
  13364=>"111101111",
  13365=>"110101110",
  13366=>"010110001",
  13367=>"101000111",
  13368=>"000000100",
  13369=>"000101110",
  13370=>"001001101",
  13371=>"011000100",
  13372=>"111001011",
  13373=>"001011011",
  13374=>"011001100",
  13375=>"000100000",
  13376=>"110000110",
  13377=>"010111100",
  13378=>"101110000",
  13379=>"001110110",
  13380=>"000000000",
  13381=>"000010001",
  13382=>"011010111",
  13383=>"011011000",
  13384=>"001100111",
  13385=>"010111101",
  13386=>"111100000",
  13387=>"000000011",
  13388=>"000011001",
  13389=>"001001111",
  13390=>"001100110",
  13391=>"111001100",
  13392=>"000011101",
  13393=>"010000000",
  13394=>"110111101",
  13395=>"010000000",
  13396=>"101000110",
  13397=>"111111000",
  13398=>"010110101",
  13399=>"000000001",
  13400=>"100000111",
  13401=>"000000111",
  13402=>"001100111",
  13403=>"010101110",
  13404=>"101000100",
  13405=>"100100111",
  13406=>"011100011",
  13407=>"011001000",
  13408=>"111011011",
  13409=>"101111001",
  13410=>"111100011",
  13411=>"011001001",
  13412=>"000000000",
  13413=>"011011101",
  13414=>"111011000",
  13415=>"100011001",
  13416=>"000000011",
  13417=>"110101010",
  13418=>"011000111",
  13419=>"101010110",
  13420=>"111110111",
  13421=>"111010100",
  13422=>"010000000",
  13423=>"001101001",
  13424=>"101010100",
  13425=>"010011110",
  13426=>"000011000",
  13427=>"100110001",
  13428=>"010100110",
  13429=>"000100001",
  13430=>"111010001",
  13431=>"000011101",
  13432=>"110101011",
  13433=>"010111111",
  13434=>"111100101",
  13435=>"110110010",
  13436=>"110100111",
  13437=>"101001011",
  13438=>"000000010",
  13439=>"101111001",
  13440=>"001100000",
  13441=>"000010010",
  13442=>"000000000",
  13443=>"001010110",
  13444=>"011110011",
  13445=>"010100010",
  13446=>"101100101",
  13447=>"111001110",
  13448=>"101011100",
  13449=>"011001101",
  13450=>"010100010",
  13451=>"000000000",
  13452=>"001001000",
  13453=>"100100101",
  13454=>"011011001",
  13455=>"101111010",
  13456=>"111111010",
  13457=>"100001110",
  13458=>"000011110",
  13459=>"111001000",
  13460=>"001011011",
  13461=>"011111110",
  13462=>"010111111",
  13463=>"111010001",
  13464=>"000010100",
  13465=>"100010011",
  13466=>"011101010",
  13467=>"111101110",
  13468=>"100001001",
  13469=>"111001000",
  13470=>"101000100",
  13471=>"110110000",
  13472=>"100011000",
  13473=>"000110011",
  13474=>"110100100",
  13475=>"100111010",
  13476=>"110101011",
  13477=>"000010110",
  13478=>"101110111",
  13479=>"010111010",
  13480=>"110001100",
  13481=>"110010110",
  13482=>"100011100",
  13483=>"110111001",
  13484=>"100000111",
  13485=>"100001001",
  13486=>"110001101",
  13487=>"001111011",
  13488=>"000000000",
  13489=>"101000010",
  13490=>"001110111",
  13491=>"001110100",
  13492=>"001111001",
  13493=>"111001000",
  13494=>"011010010",
  13495=>"010011100",
  13496=>"011010001",
  13497=>"101010000",
  13498=>"011000110",
  13499=>"001111001",
  13500=>"101100011",
  13501=>"111101111",
  13502=>"000000011",
  13503=>"000111111",
  13504=>"011110100",
  13505=>"011101010",
  13506=>"011100111",
  13507=>"011111011",
  13508=>"001101001",
  13509=>"010000010",
  13510=>"000111100",
  13511=>"110000100",
  13512=>"111011101",
  13513=>"011000101",
  13514=>"011101011",
  13515=>"011110100",
  13516=>"001001101",
  13517=>"111001010",
  13518=>"010001001",
  13519=>"101100001",
  13520=>"110111011",
  13521=>"101011110",
  13522=>"110100110",
  13523=>"001000001",
  13524=>"001000111",
  13525=>"100111001",
  13526=>"101100111",
  13527=>"110100101",
  13528=>"110110101",
  13529=>"000101010",
  13530=>"101001111",
  13531=>"001111000",
  13532=>"111011111",
  13533=>"111101110",
  13534=>"010011101",
  13535=>"001111000",
  13536=>"110100110",
  13537=>"000011010",
  13538=>"100011111",
  13539=>"001101010",
  13540=>"011100101",
  13541=>"000101001",
  13542=>"000110001",
  13543=>"000100010",
  13544=>"111010011",
  13545=>"110111011",
  13546=>"010100011",
  13547=>"111010100",
  13548=>"001101011",
  13549=>"100000110",
  13550=>"001111110",
  13551=>"110001001",
  13552=>"001011101",
  13553=>"110110111",
  13554=>"011111011",
  13555=>"111001111",
  13556=>"100000001",
  13557=>"011000111",
  13558=>"111001011",
  13559=>"011001000",
  13560=>"000010010",
  13561=>"000000000",
  13562=>"110111010",
  13563=>"111000011",
  13564=>"011100110",
  13565=>"101010001",
  13566=>"001000011",
  13567=>"000011100",
  13568=>"000110001",
  13569=>"010010101",
  13570=>"001110010",
  13571=>"011011001",
  13572=>"101011010",
  13573=>"001000011",
  13574=>"001010101",
  13575=>"111001010",
  13576=>"110010100",
  13577=>"000100101",
  13578=>"111000010",
  13579=>"100110001",
  13580=>"011010010",
  13581=>"000100110",
  13582=>"101111111",
  13583=>"111101111",
  13584=>"010011011",
  13585=>"000101010",
  13586=>"000000000",
  13587=>"110110000",
  13588=>"001010110",
  13589=>"100001110",
  13590=>"010111001",
  13591=>"000000010",
  13592=>"011101111",
  13593=>"110110100",
  13594=>"111100110",
  13595=>"011001111",
  13596=>"011101010",
  13597=>"010010000",
  13598=>"011011101",
  13599=>"010001011",
  13600=>"011000110",
  13601=>"110010000",
  13602=>"110100100",
  13603=>"010101100",
  13604=>"111011101",
  13605=>"100000010",
  13606=>"111010000",
  13607=>"010010010",
  13608=>"000101101",
  13609=>"111010111",
  13610=>"001101110",
  13611=>"010011110",
  13612=>"110100010",
  13613=>"000000111",
  13614=>"110000110",
  13615=>"011100011",
  13616=>"010101100",
  13617=>"000100110",
  13618=>"001011101",
  13619=>"010111110",
  13620=>"111011011",
  13621=>"000101100",
  13622=>"001100000",
  13623=>"001001100",
  13624=>"110001010",
  13625=>"111010011",
  13626=>"101100100",
  13627=>"000111100",
  13628=>"000001001",
  13629=>"000001001",
  13630=>"100111110",
  13631=>"100111001",
  13632=>"110001010",
  13633=>"010001000",
  13634=>"101000010",
  13635=>"011111001",
  13636=>"101001001",
  13637=>"001111001",
  13638=>"011011011",
  13639=>"110001011",
  13640=>"100110010",
  13641=>"110101010",
  13642=>"111001010",
  13643=>"101010010",
  13644=>"011111111",
  13645=>"001111100",
  13646=>"000000010",
  13647=>"001010100",
  13648=>"111001001",
  13649=>"100101011",
  13650=>"011001100",
  13651=>"000010000",
  13652=>"000101000",
  13653=>"101101101",
  13654=>"110111000",
  13655=>"001100000",
  13656=>"000010000",
  13657=>"000010000",
  13658=>"010010111",
  13659=>"011000111",
  13660=>"100111010",
  13661=>"101011010",
  13662=>"011111100",
  13663=>"101111100",
  13664=>"010111110",
  13665=>"010111000",
  13666=>"111010100",
  13667=>"100010111",
  13668=>"011110001",
  13669=>"010111001",
  13670=>"100111100",
  13671=>"010101111",
  13672=>"010001001",
  13673=>"011101111",
  13674=>"010110010",
  13675=>"110011110",
  13676=>"100001001",
  13677=>"111000001",
  13678=>"000100101",
  13679=>"101111001",
  13680=>"111011000",
  13681=>"100000100",
  13682=>"101100001",
  13683=>"001110100",
  13684=>"110100010",
  13685=>"011000000",
  13686=>"010011111",
  13687=>"011011100",
  13688=>"001001100",
  13689=>"101010110",
  13690=>"000101111",
  13691=>"101100100",
  13692=>"010111010",
  13693=>"101101000",
  13694=>"100001011",
  13695=>"011001101",
  13696=>"100101001",
  13697=>"000001110",
  13698=>"001111000",
  13699=>"000111001",
  13700=>"001000110",
  13701=>"001110000",
  13702=>"011001100",
  13703=>"011111010",
  13704=>"111001011",
  13705=>"100010100",
  13706=>"001010111",
  13707=>"001100000",
  13708=>"001110001",
  13709=>"011001000",
  13710=>"111010101",
  13711=>"111010110",
  13712=>"010111110",
  13713=>"011011000",
  13714=>"101010000",
  13715=>"000000010",
  13716=>"001000010",
  13717=>"000111001",
  13718=>"101111011",
  13719=>"111000111",
  13720=>"110100010",
  13721=>"000101011",
  13722=>"011010100",
  13723=>"111011111",
  13724=>"001001110",
  13725=>"001001101",
  13726=>"000101111",
  13727=>"011110010",
  13728=>"000001000",
  13729=>"001101110",
  13730=>"001101000",
  13731=>"110111001",
  13732=>"010010101",
  13733=>"111101001",
  13734=>"010111111",
  13735=>"011110101",
  13736=>"001111110",
  13737=>"000001111",
  13738=>"001001100",
  13739=>"111000010",
  13740=>"001000110",
  13741=>"110100100",
  13742=>"001001010",
  13743=>"010011000",
  13744=>"010101100",
  13745=>"001111000",
  13746=>"110001110",
  13747=>"111101000",
  13748=>"111101010",
  13749=>"000010000",
  13750=>"101011000",
  13751=>"110110010",
  13752=>"110000010",
  13753=>"011101010",
  13754=>"000011010",
  13755=>"100000010",
  13756=>"010100011",
  13757=>"101001011",
  13758=>"001101001",
  13759=>"000001110",
  13760=>"001010100",
  13761=>"110011010",
  13762=>"111011100",
  13763=>"100110111",
  13764=>"000001000",
  13765=>"100001011",
  13766=>"100010011",
  13767=>"111011011",
  13768=>"110011010",
  13769=>"001100100",
  13770=>"000110001",
  13771=>"010000010",
  13772=>"011010000",
  13773=>"001001100",
  13774=>"011000101",
  13775=>"111010100",
  13776=>"101000000",
  13777=>"010101000",
  13778=>"010110011",
  13779=>"000000001",
  13780=>"001111110",
  13781=>"111110000",
  13782=>"010001010",
  13783=>"110001011",
  13784=>"011010110",
  13785=>"011110110",
  13786=>"011011101",
  13787=>"100111000",
  13788=>"111101000",
  13789=>"001111100",
  13790=>"000011111",
  13791=>"011001001",
  13792=>"100111000",
  13793=>"001100110",
  13794=>"101011001",
  13795=>"000100111",
  13796=>"011111101",
  13797=>"001011000",
  13798=>"111110110",
  13799=>"110101101",
  13800=>"100100110",
  13801=>"001000111",
  13802=>"100000001",
  13803=>"011101011",
  13804=>"100001101",
  13805=>"001011101",
  13806=>"010111101",
  13807=>"101110100",
  13808=>"111111111",
  13809=>"101000111",
  13810=>"010100001",
  13811=>"101010101",
  13812=>"100100111",
  13813=>"100100110",
  13814=>"001011001",
  13815=>"100011001",
  13816=>"111111111",
  13817=>"011011111",
  13818=>"001001111",
  13819=>"000011111",
  13820=>"100000001",
  13821=>"001011000",
  13822=>"111101111",
  13823=>"110110101",
  13824=>"100111011",
  13825=>"010011110",
  13826=>"101000111",
  13827=>"011100000",
  13828=>"001001011",
  13829=>"110111000",
  13830=>"111010011",
  13831=>"100110101",
  13832=>"110011001",
  13833=>"100011001",
  13834=>"011001011",
  13835=>"101010111",
  13836=>"100110110",
  13837=>"111000110",
  13838=>"111000001",
  13839=>"111100011",
  13840=>"111001110",
  13841=>"110000000",
  13842=>"011000011",
  13843=>"011111111",
  13844=>"101101110",
  13845=>"111000001",
  13846=>"100110111",
  13847=>"001010101",
  13848=>"010110100",
  13849=>"011111100",
  13850=>"001001111",
  13851=>"101001101",
  13852=>"011111000",
  13853=>"010011011",
  13854=>"000101111",
  13855=>"111010110",
  13856=>"011001111",
  13857=>"001100011",
  13858=>"100110010",
  13859=>"011000111",
  13860=>"111011011",
  13861=>"001000110",
  13862=>"000101010",
  13863=>"101001001",
  13864=>"100110100",
  13865=>"000101110",
  13866=>"111100110",
  13867=>"011110010",
  13868=>"010110000",
  13869=>"100110111",
  13870=>"000100001",
  13871=>"001010110",
  13872=>"111011011",
  13873=>"111101010",
  13874=>"000111000",
  13875=>"110010101",
  13876=>"111000110",
  13877=>"000001110",
  13878=>"000000101",
  13879=>"110011001",
  13880=>"011011101",
  13881=>"011100100",
  13882=>"000010001",
  13883=>"111111001",
  13884=>"001101011",
  13885=>"110110110",
  13886=>"001010000",
  13887=>"111111001",
  13888=>"011100011",
  13889=>"111001001",
  13890=>"101100110",
  13891=>"001100100",
  13892=>"101110000",
  13893=>"001110110",
  13894=>"001000100",
  13895=>"010001101",
  13896=>"001010010",
  13897=>"001100010",
  13898=>"111110001",
  13899=>"101000001",
  13900=>"010001011",
  13901=>"100010101",
  13902=>"010010110",
  13903=>"011001111",
  13904=>"000110010",
  13905=>"000100101",
  13906=>"001011011",
  13907=>"000001100",
  13908=>"101000101",
  13909=>"000011100",
  13910=>"010000101",
  13911=>"111110000",
  13912=>"000101010",
  13913=>"011111101",
  13914=>"001100101",
  13915=>"100000110",
  13916=>"011111011",
  13917=>"110010100",
  13918=>"100000100",
  13919=>"010001001",
  13920=>"110011111",
  13921=>"010011001",
  13922=>"111011111",
  13923=>"001011000",
  13924=>"011110000",
  13925=>"110011001",
  13926=>"110000000",
  13927=>"000011001",
  13928=>"011001010",
  13929=>"111111001",
  13930=>"000010111",
  13931=>"101101001",
  13932=>"000110001",
  13933=>"101110100",
  13934=>"101110100",
  13935=>"111110001",
  13936=>"010000110",
  13937=>"010000000",
  13938=>"010110001",
  13939=>"100010010",
  13940=>"111110001",
  13941=>"111111000",
  13942=>"111100011",
  13943=>"001100000",
  13944=>"100011001",
  13945=>"010110110",
  13946=>"110111001",
  13947=>"011000001",
  13948=>"011001011",
  13949=>"010101011",
  13950=>"110101100",
  13951=>"110000000",
  13952=>"001101111",
  13953=>"111111101",
  13954=>"010111001",
  13955=>"000000001",
  13956=>"011101010",
  13957=>"000100010",
  13958=>"101100100",
  13959=>"111100110",
  13960=>"011100101",
  13961=>"001110110",
  13962=>"000010000",
  13963=>"011001011",
  13964=>"011001001",
  13965=>"000001010",
  13966=>"111001101",
  13967=>"011101001",
  13968=>"010110001",
  13969=>"111011011",
  13970=>"011001101",
  13971=>"010101011",
  13972=>"010000001",
  13973=>"111011011",
  13974=>"110101011",
  13975=>"101111000",
  13976=>"000111111",
  13977=>"001000010",
  13978=>"001011110",
  13979=>"010100000",
  13980=>"111000110",
  13981=>"001100111",
  13982=>"000100010",
  13983=>"100101000",
  13984=>"100000111",
  13985=>"100001001",
  13986=>"000011100",
  13987=>"101011000",
  13988=>"011111000",
  13989=>"000000111",
  13990=>"000101010",
  13991=>"011010010",
  13992=>"111000000",
  13993=>"100001110",
  13994=>"001000011",
  13995=>"110010111",
  13996=>"110011001",
  13997=>"111001011",
  13998=>"111101000",
  13999=>"010010111",
  14000=>"011011101",
  14001=>"010100011",
  14002=>"110000001",
  14003=>"011011001",
  14004=>"011000101",
  14005=>"000101011",
  14006=>"000001111",
  14007=>"111001101",
  14008=>"001110100",
  14009=>"111101101",
  14010=>"100011011",
  14011=>"011111000",
  14012=>"110101100",
  14013=>"001100001",
  14014=>"111110000",
  14015=>"001111110",
  14016=>"111010010",
  14017=>"001000010",
  14018=>"001001101",
  14019=>"111101111",
  14020=>"011101011",
  14021=>"111001111",
  14022=>"111011101",
  14023=>"110110011",
  14024=>"001011111",
  14025=>"110000111",
  14026=>"011011101",
  14027=>"010000100",
  14028=>"100001110",
  14029=>"111000010",
  14030=>"011010111",
  14031=>"110011011",
  14032=>"100100110",
  14033=>"011010010",
  14034=>"100001000",
  14035=>"100111011",
  14036=>"001101011",
  14037=>"000010000",
  14038=>"011111001",
  14039=>"100011001",
  14040=>"001001101",
  14041=>"010111011",
  14042=>"010111111",
  14043=>"111011001",
  14044=>"011110100",
  14045=>"111010110",
  14046=>"001111100",
  14047=>"100000100",
  14048=>"111010100",
  14049=>"111110110",
  14050=>"000110111",
  14051=>"011000110",
  14052=>"011100100",
  14053=>"110000100",
  14054=>"000101100",
  14055=>"010101000",
  14056=>"000100101",
  14057=>"001001100",
  14058=>"100000000",
  14059=>"001111101",
  14060=>"000010001",
  14061=>"011001000",
  14062=>"010000000",
  14063=>"001010111",
  14064=>"111111101",
  14065=>"000110010",
  14066=>"101110101",
  14067=>"101001000",
  14068=>"001010110",
  14069=>"011101101",
  14070=>"001011000",
  14071=>"001111101",
  14072=>"110001110",
  14073=>"100011110",
  14074=>"101001101",
  14075=>"111000010",
  14076=>"000001100",
  14077=>"000001101",
  14078=>"111001111",
  14079=>"000010010",
  14080=>"110000100",
  14081=>"011100101",
  14082=>"100101000",
  14083=>"000001001",
  14084=>"100001101",
  14085=>"000100001",
  14086=>"000001100",
  14087=>"110111011",
  14088=>"101111010",
  14089=>"101110100",
  14090=>"110100001",
  14091=>"001100110",
  14092=>"100011010",
  14093=>"010100011",
  14094=>"001000000",
  14095=>"100010000",
  14096=>"111010010",
  14097=>"000001011",
  14098=>"000100100",
  14099=>"011010110",
  14100=>"111101011",
  14101=>"111011101",
  14102=>"010111001",
  14103=>"110110111",
  14104=>"010001111",
  14105=>"011011001",
  14106=>"001111010",
  14107=>"110010000",
  14108=>"011100001",
  14109=>"010100010",
  14110=>"001111010",
  14111=>"001100101",
  14112=>"100110000",
  14113=>"111110011",
  14114=>"001101010",
  14115=>"100111100",
  14116=>"100011001",
  14117=>"011101010",
  14118=>"000011010",
  14119=>"001000110",
  14120=>"111011001",
  14121=>"111111111",
  14122=>"001100111",
  14123=>"000011001",
  14124=>"101011110",
  14125=>"001001011",
  14126=>"000011000",
  14127=>"001110101",
  14128=>"111010101",
  14129=>"000110110",
  14130=>"110010110",
  14131=>"011001100",
  14132=>"011101011",
  14133=>"010001100",
  14134=>"000111110",
  14135=>"000000100",
  14136=>"111010001",
  14137=>"011000001",
  14138=>"000000110",
  14139=>"110101101",
  14140=>"000100101",
  14141=>"010000011",
  14142=>"111100001",
  14143=>"111001000",
  14144=>"100000000",
  14145=>"110100111",
  14146=>"110111100",
  14147=>"000110111",
  14148=>"000000111",
  14149=>"010110101",
  14150=>"100010000",
  14151=>"100101101",
  14152=>"011110111",
  14153=>"101111111",
  14154=>"000100110",
  14155=>"010011100",
  14156=>"001101110",
  14157=>"111111001",
  14158=>"111110000",
  14159=>"010011010",
  14160=>"000010110",
  14161=>"111100110",
  14162=>"100000110",
  14163=>"111100000",
  14164=>"110001100",
  14165=>"111010010",
  14166=>"010001000",
  14167=>"010010010",
  14168=>"011001100",
  14169=>"110000111",
  14170=>"111101100",
  14171=>"100111010",
  14172=>"011100011",
  14173=>"010000000",
  14174=>"111000001",
  14175=>"100110001",
  14176=>"100010111",
  14177=>"111110011",
  14178=>"000000101",
  14179=>"110100010",
  14180=>"001101001",
  14181=>"011101101",
  14182=>"101100111",
  14183=>"010011011",
  14184=>"011111011",
  14185=>"110010100",
  14186=>"101101100",
  14187=>"111111000",
  14188=>"110000001",
  14189=>"100100101",
  14190=>"100110101",
  14191=>"010101100",
  14192=>"100011110",
  14193=>"111110110",
  14194=>"101100010",
  14195=>"001010001",
  14196=>"011110000",
  14197=>"100011101",
  14198=>"011110110",
  14199=>"100100110",
  14200=>"100001000",
  14201=>"101100001",
  14202=>"101101100",
  14203=>"011010010",
  14204=>"011011001",
  14205=>"001011100",
  14206=>"000000111",
  14207=>"110011110",
  14208=>"010111110",
  14209=>"111100001",
  14210=>"010011110",
  14211=>"100001111",
  14212=>"101000111",
  14213=>"101010111",
  14214=>"100001000",
  14215=>"111010010",
  14216=>"110010111",
  14217=>"010000111",
  14218=>"111111011",
  14219=>"010100011",
  14220=>"111010011",
  14221=>"111001011",
  14222=>"100001000",
  14223=>"101010110",
  14224=>"000110010",
  14225=>"110010011",
  14226=>"110110000",
  14227=>"011111010",
  14228=>"001001010",
  14229=>"000011000",
  14230=>"111110110",
  14231=>"011010000",
  14232=>"001110101",
  14233=>"001001111",
  14234=>"000011000",
  14235=>"000011001",
  14236=>"001000110",
  14237=>"110011000",
  14238=>"001101000",
  14239=>"011101100",
  14240=>"111010001",
  14241=>"111111111",
  14242=>"011110111",
  14243=>"110001000",
  14244=>"000000011",
  14245=>"010001001",
  14246=>"011001010",
  14247=>"101111101",
  14248=>"111011000",
  14249=>"100000011",
  14250=>"011000001",
  14251=>"011000011",
  14252=>"001011100",
  14253=>"101000010",
  14254=>"000010001",
  14255=>"010110101",
  14256=>"001000011",
  14257=>"000010101",
  14258=>"000011001",
  14259=>"101110100",
  14260=>"110100110",
  14261=>"010001000",
  14262=>"001100011",
  14263=>"010101110",
  14264=>"011011111",
  14265=>"001000010",
  14266=>"000111000",
  14267=>"000011011",
  14268=>"111111011",
  14269=>"000111111",
  14270=>"111110101",
  14271=>"101001111",
  14272=>"011110111",
  14273=>"000100101",
  14274=>"000001101",
  14275=>"111010111",
  14276=>"010001110",
  14277=>"100101101",
  14278=>"100100001",
  14279=>"101011011",
  14280=>"100101000",
  14281=>"101110100",
  14282=>"000001000",
  14283=>"101000101",
  14284=>"100100100",
  14285=>"110001101",
  14286=>"000000111",
  14287=>"011000001",
  14288=>"110110010",
  14289=>"100101101",
  14290=>"101110111",
  14291=>"011101000",
  14292=>"000000000",
  14293=>"101111010",
  14294=>"101001000",
  14295=>"011110110",
  14296=>"111100001",
  14297=>"000100111",
  14298=>"110111100",
  14299=>"111000001",
  14300=>"010101010",
  14301=>"110101110",
  14302=>"010100001",
  14303=>"111011010",
  14304=>"010011111",
  14305=>"011000011",
  14306=>"111001010",
  14307=>"010011100",
  14308=>"111000110",
  14309=>"001110101",
  14310=>"000110111",
  14311=>"110011000",
  14312=>"101100000",
  14313=>"110001110",
  14314=>"010101101",
  14315=>"111110010",
  14316=>"101010011",
  14317=>"011010011",
  14318=>"010000001",
  14319=>"011111000",
  14320=>"010010100",
  14321=>"010011100",
  14322=>"000101110",
  14323=>"010001011",
  14324=>"111100100",
  14325=>"111011011",
  14326=>"001111110",
  14327=>"100001001",
  14328=>"100011111",
  14329=>"001001001",
  14330=>"110100100",
  14331=>"100100110",
  14332=>"101110000",
  14333=>"000110011",
  14334=>"110110001",
  14335=>"111101011",
  14336=>"101101011",
  14337=>"110100101",
  14338=>"001010111",
  14339=>"001011111",
  14340=>"101000111",
  14341=>"101010110",
  14342=>"001000101",
  14343=>"001010000",
  14344=>"111010110",
  14345=>"010001001",
  14346=>"001010101",
  14347=>"100111110",
  14348=>"000010011",
  14349=>"101110010",
  14350=>"000001000",
  14351=>"011100000",
  14352=>"110110001",
  14353=>"100111011",
  14354=>"101110100",
  14355=>"011110110",
  14356=>"110110011",
  14357=>"011001000",
  14358=>"001000000",
  14359=>"111100100",
  14360=>"011101000",
  14361=>"111111100",
  14362=>"010001011",
  14363=>"000000001",
  14364=>"000011111",
  14365=>"001001011",
  14366=>"011010001",
  14367=>"000000011",
  14368=>"000101111",
  14369=>"010101001",
  14370=>"101000101",
  14371=>"110111010",
  14372=>"101101001",
  14373=>"110101111",
  14374=>"011111111",
  14375=>"010111100",
  14376=>"000001000",
  14377=>"100010010",
  14378=>"001111001",
  14379=>"110100011",
  14380=>"110111001",
  14381=>"011011000",
  14382=>"001101101",
  14383=>"001001001",
  14384=>"111010100",
  14385=>"000110111",
  14386=>"001011100",
  14387=>"011100100",
  14388=>"010000101",
  14389=>"111000100",
  14390=>"100001000",
  14391=>"100100000",
  14392=>"000010111",
  14393=>"010000011",
  14394=>"000110110",
  14395=>"101001011",
  14396=>"111010011",
  14397=>"100111111",
  14398=>"110000111",
  14399=>"110010001",
  14400=>"111001000",
  14401=>"101010011",
  14402=>"100100000",
  14403=>"000010100",
  14404=>"011111101",
  14405=>"100101100",
  14406=>"100111001",
  14407=>"001000000",
  14408=>"010111000",
  14409=>"000001010",
  14410=>"111001010",
  14411=>"100101101",
  14412=>"101110010",
  14413=>"100111000",
  14414=>"011001000",
  14415=>"000010101",
  14416=>"001111111",
  14417=>"111111111",
  14418=>"000110110",
  14419=>"111100001",
  14420=>"011111010",
  14421=>"100011010",
  14422=>"100100110",
  14423=>"101100101",
  14424=>"101100000",
  14425=>"001000000",
  14426=>"100100000",
  14427=>"011001000",
  14428=>"001011000",
  14429=>"000101100",
  14430=>"100011000",
  14431=>"100010101",
  14432=>"000110011",
  14433=>"001000010",
  14434=>"011010011",
  14435=>"001010101",
  14436=>"111010010",
  14437=>"110110100",
  14438=>"000011000",
  14439=>"101011110",
  14440=>"110000100",
  14441=>"110110110",
  14442=>"001101111",
  14443=>"010101010",
  14444=>"101111110",
  14445=>"110000111",
  14446=>"010110001",
  14447=>"111001110",
  14448=>"000101101",
  14449=>"001100101",
  14450=>"001001101",
  14451=>"000110011",
  14452=>"100110011",
  14453=>"001010010",
  14454=>"101111011",
  14455=>"110111100",
  14456=>"010001000",
  14457=>"111110101",
  14458=>"111000001",
  14459=>"011110100",
  14460=>"011101000",
  14461=>"000010101",
  14462=>"111011000",
  14463=>"111001010",
  14464=>"010100000",
  14465=>"010010001",
  14466=>"100000100",
  14467=>"000101010",
  14468=>"100000111",
  14469=>"010101101",
  14470=>"011000111",
  14471=>"000010100",
  14472=>"111101110",
  14473=>"110011001",
  14474=>"110000110",
  14475=>"000000111",
  14476=>"000111111",
  14477=>"010101110",
  14478=>"101000110",
  14479=>"100001000",
  14480=>"011111110",
  14481=>"101001100",
  14482=>"001000001",
  14483=>"101010000",
  14484=>"001100010",
  14485=>"010011001",
  14486=>"000001110",
  14487=>"001011010",
  14488=>"011000100",
  14489=>"110001000",
  14490=>"101010000",
  14491=>"101111101",
  14492=>"000011101",
  14493=>"110100010",
  14494=>"100001110",
  14495=>"001010001",
  14496=>"011010001",
  14497=>"101111011",
  14498=>"111000010",
  14499=>"000001001",
  14500=>"110011110",
  14501=>"110110110",
  14502=>"100101011",
  14503=>"110101111",
  14504=>"111111000",
  14505=>"000110010",
  14506=>"111001101",
  14507=>"010101100",
  14508=>"010111100",
  14509=>"101010101",
  14510=>"110001100",
  14511=>"010101110",
  14512=>"001110001",
  14513=>"100011001",
  14514=>"011011110",
  14515=>"011100010",
  14516=>"010000010",
  14517=>"100101111",
  14518=>"101110101",
  14519=>"100001010",
  14520=>"010110111",
  14521=>"100011010",
  14522=>"011111111",
  14523=>"110100110",
  14524=>"011101011",
  14525=>"111000111",
  14526=>"000000010",
  14527=>"110100110",
  14528=>"010010110",
  14529=>"101010000",
  14530=>"111100000",
  14531=>"010011010",
  14532=>"111100110",
  14533=>"010100101",
  14534=>"001101110",
  14535=>"000110111",
  14536=>"010110110",
  14537=>"010110101",
  14538=>"010110000",
  14539=>"100101110",
  14540=>"111010010",
  14541=>"100010111",
  14542=>"110101010",
  14543=>"111011011",
  14544=>"000101110",
  14545=>"001010011",
  14546=>"110100101",
  14547=>"111000110",
  14548=>"010000100",
  14549=>"011101110",
  14550=>"011000101",
  14551=>"010000110",
  14552=>"100100100",
  14553=>"000001000",
  14554=>"001001011",
  14555=>"000101101",
  14556=>"011101010",
  14557=>"110000111",
  14558=>"010001011",
  14559=>"110011010",
  14560=>"000100011",
  14561=>"110101111",
  14562=>"010001001",
  14563=>"101101110",
  14564=>"000111100",
  14565=>"100010010",
  14566=>"101110000",
  14567=>"001001111",
  14568=>"110100001",
  14569=>"011111010",
  14570=>"010110111",
  14571=>"000010011",
  14572=>"010000110",
  14573=>"100111001",
  14574=>"100001101",
  14575=>"100110100",
  14576=>"000110111",
  14577=>"101101101",
  14578=>"001010000",
  14579=>"110110100",
  14580=>"110100000",
  14581=>"001111011",
  14582=>"000011000",
  14583=>"101001000",
  14584=>"100101111",
  14585=>"000100110",
  14586=>"101000100",
  14587=>"001110011",
  14588=>"000101000",
  14589=>"101011111",
  14590=>"110010010",
  14591=>"011111000",
  14592=>"010000110",
  14593=>"111101111",
  14594=>"010010011",
  14595=>"000000100",
  14596=>"010011000",
  14597=>"110101111",
  14598=>"010110100",
  14599=>"100100001",
  14600=>"101110001",
  14601=>"010110010",
  14602=>"010000111",
  14603=>"010000000",
  14604=>"111011100",
  14605=>"110111010",
  14606=>"101101010",
  14607=>"101000110",
  14608=>"111010110",
  14609=>"011111010",
  14610=>"010000111",
  14611=>"010000011",
  14612=>"000010011",
  14613=>"001000101",
  14614=>"010110001",
  14615=>"100011000",
  14616=>"100111000",
  14617=>"110100010",
  14618=>"001000001",
  14619=>"110011000",
  14620=>"010011011",
  14621=>"101110110",
  14622=>"101101110",
  14623=>"001001010",
  14624=>"010010111",
  14625=>"001001010",
  14626=>"101011010",
  14627=>"101011000",
  14628=>"001000110",
  14629=>"111110011",
  14630=>"011010010",
  14631=>"000010011",
  14632=>"000100111",
  14633=>"101111000",
  14634=>"100000011",
  14635=>"000011001",
  14636=>"111110001",
  14637=>"011000100",
  14638=>"010100111",
  14639=>"001010000",
  14640=>"000000011",
  14641=>"011101101",
  14642=>"100010100",
  14643=>"101111111",
  14644=>"001101011",
  14645=>"100101011",
  14646=>"001010100",
  14647=>"100010010",
  14648=>"000001000",
  14649=>"011110100",
  14650=>"001010001",
  14651=>"010110010",
  14652=>"000000111",
  14653=>"001010111",
  14654=>"100101101",
  14655=>"001101011",
  14656=>"001001010",
  14657=>"000000011",
  14658=>"001010100",
  14659=>"111100110",
  14660=>"011101111",
  14661=>"000111110",
  14662=>"111000001",
  14663=>"111110111",
  14664=>"101011001",
  14665=>"000110001",
  14666=>"101000110",
  14667=>"100000001",
  14668=>"010100110",
  14669=>"010001011",
  14670=>"111010011",
  14671=>"101101111",
  14672=>"111010101",
  14673=>"011001100",
  14674=>"111111000",
  14675=>"011011110",
  14676=>"101100001",
  14677=>"000100110",
  14678=>"101110101",
  14679=>"110110101",
  14680=>"001000001",
  14681=>"001100001",
  14682=>"011001100",
  14683=>"101110111",
  14684=>"100010000",
  14685=>"111010110",
  14686=>"001101000",
  14687=>"001100011",
  14688=>"000000100",
  14689=>"000110011",
  14690=>"011101000",
  14691=>"100000110",
  14692=>"111100110",
  14693=>"101011000",
  14694=>"111111100",
  14695=>"000110110",
  14696=>"111000011",
  14697=>"110001001",
  14698=>"010110100",
  14699=>"100101110",
  14700=>"011011010",
  14701=>"010101010",
  14702=>"000000101",
  14703=>"010100001",
  14704=>"101000000",
  14705=>"100011101",
  14706=>"011001011",
  14707=>"110011000",
  14708=>"101000011",
  14709=>"100111011",
  14710=>"000000100",
  14711=>"010001000",
  14712=>"010010000",
  14713=>"110111101",
  14714=>"010001011",
  14715=>"110011000",
  14716=>"100101111",
  14717=>"110010010",
  14718=>"111110100",
  14719=>"010100001",
  14720=>"010001101",
  14721=>"000100010",
  14722=>"101110100",
  14723=>"011111011",
  14724=>"000110000",
  14725=>"110111011",
  14726=>"000111101",
  14727=>"111011011",
  14728=>"101001111",
  14729=>"111101101",
  14730=>"011001100",
  14731=>"001101111",
  14732=>"100000000",
  14733=>"111110001",
  14734=>"001100100",
  14735=>"001110100",
  14736=>"101010100",
  14737=>"000000000",
  14738=>"101101111",
  14739=>"001100001",
  14740=>"100001101",
  14741=>"110001101",
  14742=>"001100001",
  14743=>"010010111",
  14744=>"101100111",
  14745=>"001011100",
  14746=>"011101010",
  14747=>"111111010",
  14748=>"101101111",
  14749=>"001100001",
  14750=>"111111010",
  14751=>"011011000",
  14752=>"001101101",
  14753=>"001000011",
  14754=>"100100110",
  14755=>"100101010",
  14756=>"010110000",
  14757=>"100010111",
  14758=>"011001000",
  14759=>"010110100",
  14760=>"011111101",
  14761=>"010111000",
  14762=>"000001111",
  14763=>"111011000",
  14764=>"000101011",
  14765=>"101010001",
  14766=>"001000101",
  14767=>"010010000",
  14768=>"011001101",
  14769=>"110111101",
  14770=>"000101111",
  14771=>"011100101",
  14772=>"100001101",
  14773=>"011101110",
  14774=>"101010101",
  14775=>"001110100",
  14776=>"111010011",
  14777=>"000001101",
  14778=>"101001011",
  14779=>"011000000",
  14780=>"000011110",
  14781=>"010001100",
  14782=>"001000010",
  14783=>"001111110",
  14784=>"110101010",
  14785=>"100011010",
  14786=>"010110111",
  14787=>"010100101",
  14788=>"000000110",
  14789=>"110110010",
  14790=>"011100011",
  14791=>"010100011",
  14792=>"100001101",
  14793=>"101101001",
  14794=>"101010111",
  14795=>"010010010",
  14796=>"001010100",
  14797=>"010111101",
  14798=>"110010111",
  14799=>"100010010",
  14800=>"001111110",
  14801=>"100101001",
  14802=>"001101001",
  14803=>"100001100",
  14804=>"011000100",
  14805=>"001011111",
  14806=>"100011011",
  14807=>"111111101",
  14808=>"110111111",
  14809=>"110000100",
  14810=>"010011101",
  14811=>"001000100",
  14812=>"011101011",
  14813=>"000110011",
  14814=>"110000011",
  14815=>"000110111",
  14816=>"010000101",
  14817=>"100110000",
  14818=>"110111000",
  14819=>"110001000",
  14820=>"000110010",
  14821=>"011110101",
  14822=>"101011000",
  14823=>"001001001",
  14824=>"011100010",
  14825=>"110000110",
  14826=>"110011100",
  14827=>"101010001",
  14828=>"000000110",
  14829=>"111101111",
  14830=>"011101011",
  14831=>"111000001",
  14832=>"010110111",
  14833=>"110001010",
  14834=>"101111111",
  14835=>"000010001",
  14836=>"100010010",
  14837=>"010010110",
  14838=>"000110011",
  14839=>"110000101",
  14840=>"011101011",
  14841=>"100100000",
  14842=>"111000000",
  14843=>"111111101",
  14844=>"000010011",
  14845=>"110101100",
  14846=>"011111110",
  14847=>"010101101",
  14848=>"110110100",
  14849=>"101001101",
  14850=>"111111111",
  14851=>"101010101",
  14852=>"110010000",
  14853=>"101010000",
  14854=>"001011011",
  14855=>"111100100",
  14856=>"011001110",
  14857=>"101111111",
  14858=>"101010000",
  14859=>"011000001",
  14860=>"101010011",
  14861=>"001101010",
  14862=>"111001010",
  14863=>"001001111",
  14864=>"100111000",
  14865=>"101011010",
  14866=>"111100000",
  14867=>"011110010",
  14868=>"101101110",
  14869=>"110100001",
  14870=>"011111101",
  14871=>"000100001",
  14872=>"001101010",
  14873=>"000001011",
  14874=>"010101011",
  14875=>"100100010",
  14876=>"110100001",
  14877=>"011100101",
  14878=>"000010000",
  14879=>"010001100",
  14880=>"001101011",
  14881=>"110000000",
  14882=>"001000001",
  14883=>"011101111",
  14884=>"001010010",
  14885=>"101001000",
  14886=>"001011001",
  14887=>"111111010",
  14888=>"100101001",
  14889=>"001110111",
  14890=>"000011110",
  14891=>"000111111",
  14892=>"111100011",
  14893=>"111111101",
  14894=>"010000101",
  14895=>"001110101",
  14896=>"110000010",
  14897=>"100010100",
  14898=>"111100011",
  14899=>"110101010",
  14900=>"001001100",
  14901=>"000010010",
  14902=>"000011100",
  14903=>"101000010",
  14904=>"011111001",
  14905=>"011101101",
  14906=>"101110001",
  14907=>"111110100",
  14908=>"000010000",
  14909=>"000001111",
  14910=>"010101111",
  14911=>"111000111",
  14912=>"110011111",
  14913=>"101010000",
  14914=>"110011010",
  14915=>"111101100",
  14916=>"101010010",
  14917=>"010010001",
  14918=>"001000010",
  14919=>"111000101",
  14920=>"100011110",
  14921=>"000110110",
  14922=>"100101001",
  14923=>"111011010",
  14924=>"111011110",
  14925=>"101000000",
  14926=>"111111101",
  14927=>"000101001",
  14928=>"001000000",
  14929=>"110010100",
  14930=>"010000011",
  14931=>"010101011",
  14932=>"110101110",
  14933=>"000001101",
  14934=>"111000010",
  14935=>"100111111",
  14936=>"010100100",
  14937=>"110100111",
  14938=>"110000110",
  14939=>"101011011",
  14940=>"001100001",
  14941=>"000101100",
  14942=>"010110010",
  14943=>"010000011",
  14944=>"101000110",
  14945=>"010110001",
  14946=>"111100011",
  14947=>"010100111",
  14948=>"011100100",
  14949=>"101000010",
  14950=>"001100001",
  14951=>"110011100",
  14952=>"000101010",
  14953=>"010100010",
  14954=>"100110100",
  14955=>"000100000",
  14956=>"100010000",
  14957=>"111101011",
  14958=>"001011110",
  14959=>"001111110",
  14960=>"101110101",
  14961=>"110100010",
  14962=>"000000001",
  14963=>"011111010",
  14964=>"110101101",
  14965=>"000001010",
  14966=>"111111000",
  14967=>"011111100",
  14968=>"010001100",
  14969=>"110101110",
  14970=>"110100110",
  14971=>"011000100",
  14972=>"001111111",
  14973=>"000001111",
  14974=>"110010100",
  14975=>"101001001",
  14976=>"111010010",
  14977=>"001001111",
  14978=>"110110101",
  14979=>"001010001",
  14980=>"001000001",
  14981=>"110110101",
  14982=>"100010100",
  14983=>"100110010",
  14984=>"101000010",
  14985=>"001001110",
  14986=>"110010001",
  14987=>"011001110",
  14988=>"001000111",
  14989=>"011111101",
  14990=>"000011110",
  14991=>"110110110",
  14992=>"011101011",
  14993=>"111010011",
  14994=>"111010111",
  14995=>"001100101",
  14996=>"110100001",
  14997=>"111001110",
  14998=>"110101000",
  14999=>"101010111",
  15000=>"111101010",
  15001=>"001101011",
  15002=>"000010000",
  15003=>"011100001",
  15004=>"101111010",
  15005=>"111101011",
  15006=>"011100001",
  15007=>"000010100",
  15008=>"111111111",
  15009=>"111001000",
  15010=>"000010000",
  15011=>"110010101",
  15012=>"101110101",
  15013=>"001010000",
  15014=>"110000101",
  15015=>"000000100",
  15016=>"110011110",
  15017=>"000100101",
  15018=>"011100100",
  15019=>"011001010",
  15020=>"100000001",
  15021=>"000010101",
  15022=>"000111111",
  15023=>"010010110",
  15024=>"010011010",
  15025=>"110011000",
  15026=>"000100011",
  15027=>"101001000",
  15028=>"110111011",
  15029=>"000100101",
  15030=>"110011011",
  15031=>"110011110",
  15032=>"110000011",
  15033=>"100000111",
  15034=>"001001000",
  15035=>"000000110",
  15036=>"000101111",
  15037=>"111101011",
  15038=>"000000001",
  15039=>"001100110",
  15040=>"010011111",
  15041=>"000011001",
  15042=>"010010011",
  15043=>"000010110",
  15044=>"001000100",
  15045=>"010000101",
  15046=>"011111000",
  15047=>"010000011",
  15048=>"010110111",
  15049=>"110111001",
  15050=>"001111100",
  15051=>"010101000",
  15052=>"000100101",
  15053=>"110101011",
  15054=>"010010110",
  15055=>"111001001",
  15056=>"000011111",
  15057=>"011000000",
  15058=>"000010111",
  15059=>"101011101",
  15060=>"111101001",
  15061=>"010101110",
  15062=>"010100100",
  15063=>"010110100",
  15064=>"100010101",
  15065=>"000010011",
  15066=>"101101001",
  15067=>"010100111",
  15068=>"000101110",
  15069=>"110000000",
  15070=>"100010111",
  15071=>"100101111",
  15072=>"010000110",
  15073=>"011100111",
  15074=>"001110001",
  15075=>"101100110",
  15076=>"001001010",
  15077=>"010110110",
  15078=>"101101000",
  15079=>"001101101",
  15080=>"110111001",
  15081=>"101001011",
  15082=>"001011000",
  15083=>"110101111",
  15084=>"101001001",
  15085=>"001100011",
  15086=>"001110011",
  15087=>"001001011",
  15088=>"000000100",
  15089=>"111100100",
  15090=>"101001000",
  15091=>"011110010",
  15092=>"110100100",
  15093=>"101100010",
  15094=>"000000001",
  15095=>"001100001",
  15096=>"100111011",
  15097=>"001001110",
  15098=>"110101011",
  15099=>"100100110",
  15100=>"011001111",
  15101=>"110101000",
  15102=>"110001011",
  15103=>"111110111",
  15104=>"010111110",
  15105=>"100000000",
  15106=>"100101000",
  15107=>"010100000",
  15108=>"011010100",
  15109=>"100000001",
  15110=>"100001001",
  15111=>"011111001",
  15112=>"101100101",
  15113=>"111001000",
  15114=>"001010101",
  15115=>"100000001",
  15116=>"101000010",
  15117=>"101111010",
  15118=>"111101110",
  15119=>"001100100",
  15120=>"011001100",
  15121=>"111001101",
  15122=>"001100000",
  15123=>"011100000",
  15124=>"000100101",
  15125=>"001111100",
  15126=>"110100111",
  15127=>"001110111",
  15128=>"101001101",
  15129=>"011010110",
  15130=>"101110001",
  15131=>"110100011",
  15132=>"100001001",
  15133=>"000000001",
  15134=>"110011000",
  15135=>"101001100",
  15136=>"111011100",
  15137=>"101010110",
  15138=>"010010000",
  15139=>"011000110",
  15140=>"100111001",
  15141=>"111101011",
  15142=>"011111111",
  15143=>"001001011",
  15144=>"011011101",
  15145=>"000011000",
  15146=>"001000001",
  15147=>"111111010",
  15148=>"011110101",
  15149=>"000110011",
  15150=>"111001001",
  15151=>"111010000",
  15152=>"000011111",
  15153=>"110011010",
  15154=>"001100101",
  15155=>"000010010",
  15156=>"011101111",
  15157=>"000101001",
  15158=>"111010110",
  15159=>"000111000",
  15160=>"101010110",
  15161=>"000111101",
  15162=>"101110101",
  15163=>"000000010",
  15164=>"011111110",
  15165=>"110010000",
  15166=>"000001010",
  15167=>"101010000",
  15168=>"100110100",
  15169=>"100010011",
  15170=>"101011000",
  15171=>"101001110",
  15172=>"111110111",
  15173=>"000011101",
  15174=>"101111101",
  15175=>"011110101",
  15176=>"101101011",
  15177=>"010100110",
  15178=>"000001001",
  15179=>"100011010",
  15180=>"001100110",
  15181=>"001111011",
  15182=>"101101001",
  15183=>"000100100",
  15184=>"101101100",
  15185=>"001101000",
  15186=>"001011100",
  15187=>"101000101",
  15188=>"110111110",
  15189=>"010100000",
  15190=>"111011100",
  15191=>"001010000",
  15192=>"000000001",
  15193=>"001001100",
  15194=>"100001110",
  15195=>"000001110",
  15196=>"010111110",
  15197=>"011000111",
  15198=>"100101100",
  15199=>"100111000",
  15200=>"010011100",
  15201=>"101111100",
  15202=>"001111110",
  15203=>"010111101",
  15204=>"110110001",
  15205=>"010100010",
  15206=>"001011001",
  15207=>"000111111",
  15208=>"111101110",
  15209=>"001100100",
  15210=>"000001000",
  15211=>"010110110",
  15212=>"000000010",
  15213=>"001000111",
  15214=>"111001000",
  15215=>"010000111",
  15216=>"010101100",
  15217=>"111011010",
  15218=>"010101110",
  15219=>"011111010",
  15220=>"100100111",
  15221=>"010110111",
  15222=>"000111001",
  15223=>"100101101",
  15224=>"011100000",
  15225=>"111001011",
  15226=>"011010111",
  15227=>"111011100",
  15228=>"111100101",
  15229=>"100110111",
  15230=>"100010000",
  15231=>"111010110",
  15232=>"101000001",
  15233=>"101110100",
  15234=>"100000011",
  15235=>"000101010",
  15236=>"000100110",
  15237=>"110100001",
  15238=>"010011000",
  15239=>"010011101",
  15240=>"000010011",
  15241=>"010010100",
  15242=>"100010111",
  15243=>"000101010",
  15244=>"111110100",
  15245=>"110101011",
  15246=>"110000011",
  15247=>"101100110",
  15248=>"101100101",
  15249=>"110000100",
  15250=>"100101011",
  15251=>"110011011",
  15252=>"010101000",
  15253=>"000101110",
  15254=>"010100101",
  15255=>"110010111",
  15256=>"110100011",
  15257=>"001111101",
  15258=>"101110000",
  15259=>"101011111",
  15260=>"001100011",
  15261=>"001000011",
  15262=>"000010000",
  15263=>"111110000",
  15264=>"000001111",
  15265=>"111101101",
  15266=>"011001000",
  15267=>"011100001",
  15268=>"000100111",
  15269=>"110011000",
  15270=>"100010111",
  15271=>"101100000",
  15272=>"010010011",
  15273=>"000001000",
  15274=>"100000010",
  15275=>"000010111",
  15276=>"101111100",
  15277=>"111111000",
  15278=>"000100011",
  15279=>"001000111",
  15280=>"101010110",
  15281=>"110100111",
  15282=>"010001101",
  15283=>"000100110",
  15284=>"001011110",
  15285=>"111011111",
  15286=>"010011110",
  15287=>"111001111",
  15288=>"100100101",
  15289=>"001010110",
  15290=>"110111111",
  15291=>"111111111",
  15292=>"100100011",
  15293=>"101001101",
  15294=>"010010111",
  15295=>"011001001",
  15296=>"011010100",
  15297=>"101010011",
  15298=>"111111000",
  15299=>"100110100",
  15300=>"100010110",
  15301=>"000001111",
  15302=>"101000010",
  15303=>"000000100",
  15304=>"010000000",
  15305=>"011101001",
  15306=>"111110000",
  15307=>"110110100",
  15308=>"010100011",
  15309=>"000100110",
  15310=>"100110110",
  15311=>"000010100",
  15312=>"110111011",
  15313=>"000011111",
  15314=>"101000000",
  15315=>"110010101",
  15316=>"111011111",
  15317=>"010011010",
  15318=>"000010111",
  15319=>"100110010",
  15320=>"001011011",
  15321=>"001001100",
  15322=>"101100100",
  15323=>"011010000",
  15324=>"001101110",
  15325=>"111111100",
  15326=>"000000010",
  15327=>"110011100",
  15328=>"100111011",
  15329=>"011110110",
  15330=>"010110011",
  15331=>"010101101",
  15332=>"101011011",
  15333=>"000000000",
  15334=>"100110010",
  15335=>"101110001",
  15336=>"000101111",
  15337=>"010111011",
  15338=>"011110000",
  15339=>"000010111",
  15340=>"001000000",
  15341=>"101010010",
  15342=>"000011101",
  15343=>"000110111",
  15344=>"011000010",
  15345=>"100101100",
  15346=>"100001000",
  15347=>"111001011",
  15348=>"111111001",
  15349=>"000101111",
  15350=>"010011000",
  15351=>"101000010",
  15352=>"110110011",
  15353=>"110110100",
  15354=>"100100110",
  15355=>"101011111",
  15356=>"111111001",
  15357=>"011010110",
  15358=>"000010000",
  15359=>"011001000",
  15360=>"000110000",
  15361=>"111010101",
  15362=>"101001011",
  15363=>"101100001",
  15364=>"111100010",
  15365=>"010010111",
  15366=>"101011010",
  15367=>"001110001",
  15368=>"000010010",
  15369=>"110100011",
  15370=>"011101011",
  15371=>"111010101",
  15372=>"011000100",
  15373=>"110100011",
  15374=>"001111000",
  15375=>"001010111",
  15376=>"010101111",
  15377=>"101001111",
  15378=>"101001000",
  15379=>"110001110",
  15380=>"101000100",
  15381=>"100010001",
  15382=>"101011001",
  15383=>"000011001",
  15384=>"000110100",
  15385=>"100001011",
  15386=>"001000110",
  15387=>"011111011",
  15388=>"000101010",
  15389=>"001001001",
  15390=>"111000100",
  15391=>"101010100",
  15392=>"110000101",
  15393=>"110000100",
  15394=>"011001110",
  15395=>"110011010",
  15396=>"000011001",
  15397=>"001101101",
  15398=>"000100010",
  15399=>"111010010",
  15400=>"011101111",
  15401=>"010001111",
  15402=>"010010011",
  15403=>"101000101",
  15404=>"000011001",
  15405=>"111110001",
  15406=>"001001100",
  15407=>"001110111",
  15408=>"011011101",
  15409=>"001010101",
  15410=>"101111100",
  15411=>"010000100",
  15412=>"101000000",
  15413=>"110000001",
  15414=>"100001101",
  15415=>"000110101",
  15416=>"100000101",
  15417=>"001100110",
  15418=>"111111111",
  15419=>"000101001",
  15420=>"001001110",
  15421=>"011010000",
  15422=>"101000101",
  15423=>"000010111",
  15424=>"010110100",
  15425=>"100110111",
  15426=>"100011111",
  15427=>"011110011",
  15428=>"111011101",
  15429=>"101001110",
  15430=>"110011101",
  15431=>"100000011",
  15432=>"011100011",
  15433=>"011101100",
  15434=>"001111010",
  15435=>"010111110",
  15436=>"101100010",
  15437=>"011101001",
  15438=>"000001101",
  15439=>"010010000",
  15440=>"000001011",
  15441=>"100100010",
  15442=>"001110101",
  15443=>"001001100",
  15444=>"111111100",
  15445=>"001110001",
  15446=>"101001100",
  15447=>"101010000",
  15448=>"011010101",
  15449=>"110100111",
  15450=>"100100100",
  15451=>"101000100",
  15452=>"000000100",
  15453=>"000000010",
  15454=>"001000000",
  15455=>"110100001",
  15456=>"011101111",
  15457=>"110101110",
  15458=>"100010011",
  15459=>"111101001",
  15460=>"010100001",
  15461=>"010011101",
  15462=>"111111101",
  15463=>"011001111",
  15464=>"101001101",
  15465=>"111111010",
  15466=>"101010010",
  15467=>"111000010",
  15468=>"011000110",
  15469=>"000001110",
  15470=>"111000011",
  15471=>"001000001",
  15472=>"111111000",
  15473=>"100100101",
  15474=>"011011011",
  15475=>"001000000",
  15476=>"011000100",
  15477=>"101110001",
  15478=>"101111100",
  15479=>"000011000",
  15480=>"011110111",
  15481=>"011001111",
  15482=>"101110011",
  15483=>"000101011",
  15484=>"000010100",
  15485=>"110011110",
  15486=>"000010000",
  15487=>"011001000",
  15488=>"111000011",
  15489=>"000010100",
  15490=>"011101000",
  15491=>"010110011",
  15492=>"100101011",
  15493=>"110111110",
  15494=>"011001110",
  15495=>"000100010",
  15496=>"000111000",
  15497=>"011000101",
  15498=>"101001011",
  15499=>"111101100",
  15500=>"000101010",
  15501=>"110101000",
  15502=>"100111101",
  15503=>"100011000",
  15504=>"001010101",
  15505=>"100001000",
  15506=>"110101100",
  15507=>"011010001",
  15508=>"101000000",
  15509=>"100101000",
  15510=>"011101010",
  15511=>"011000110",
  15512=>"010010110",
  15513=>"101100001",
  15514=>"100010011",
  15515=>"010110011",
  15516=>"011101111",
  15517=>"101001111",
  15518=>"110000011",
  15519=>"011010110",
  15520=>"101011100",
  15521=>"111011001",
  15522=>"111110000",
  15523=>"011111011",
  15524=>"101010100",
  15525=>"111101111",
  15526=>"011011110",
  15527=>"110011110",
  15528=>"100100000",
  15529=>"010011110",
  15530=>"110100011",
  15531=>"000100000",
  15532=>"111110111",
  15533=>"111000000",
  15534=>"100010100",
  15535=>"111000101",
  15536=>"001010110",
  15537=>"011100111",
  15538=>"000100010",
  15539=>"111010100",
  15540=>"010101111",
  15541=>"111100001",
  15542=>"111000100",
  15543=>"000000100",
  15544=>"010010110",
  15545=>"001110111",
  15546=>"111111000",
  15547=>"100000111",
  15548=>"110010010",
  15549=>"101111110",
  15550=>"001001100",
  15551=>"110011101",
  15552=>"001011010",
  15553=>"110000010",
  15554=>"001011100",
  15555=>"111010001",
  15556=>"000100001",
  15557=>"100111110",
  15558=>"111011101",
  15559=>"100111011",
  15560=>"110010011",
  15561=>"101001100",
  15562=>"010101010",
  15563=>"110001000",
  15564=>"010100110",
  15565=>"010110101",
  15566=>"010100111",
  15567=>"110110101",
  15568=>"001000010",
  15569=>"111000101",
  15570=>"000000011",
  15571=>"100000001",
  15572=>"111110111",
  15573=>"011101100",
  15574=>"111000111",
  15575=>"111000101",
  15576=>"011101101",
  15577=>"110101010",
  15578=>"001111111",
  15579=>"101101000",
  15580=>"110001100",
  15581=>"000010010",
  15582=>"101001110",
  15583=>"011011100",
  15584=>"111110011",
  15585=>"010111010",
  15586=>"001101010",
  15587=>"011001111",
  15588=>"101111000",
  15589=>"010000011",
  15590=>"101001011",
  15591=>"010111100",
  15592=>"010101110",
  15593=>"010011011",
  15594=>"101110101",
  15595=>"001010000",
  15596=>"001001000",
  15597=>"100000011",
  15598=>"001100100",
  15599=>"000111100",
  15600=>"111001101",
  15601=>"011110111",
  15602=>"001100010",
  15603=>"110110000",
  15604=>"011010110",
  15605=>"111001111",
  15606=>"011010110",
  15607=>"111001001",
  15608=>"101110110",
  15609=>"010101101",
  15610=>"110011100",
  15611=>"000001100",
  15612=>"110111111",
  15613=>"100000001",
  15614=>"001010010",
  15615=>"111000010",
  15616=>"010000101",
  15617=>"110011000",
  15618=>"101000011",
  15619=>"111100000",
  15620=>"011000010",
  15621=>"100001100",
  15622=>"010000101",
  15623=>"101010010",
  15624=>"100111010",
  15625=>"011100100",
  15626=>"011011000",
  15627=>"101111111",
  15628=>"101011001",
  15629=>"000100000",
  15630=>"000000010",
  15631=>"000000111",
  15632=>"110100100",
  15633=>"011000000",
  15634=>"011010000",
  15635=>"110111100",
  15636=>"011011001",
  15637=>"000111011",
  15638=>"101111110",
  15639=>"111000110",
  15640=>"111001010",
  15641=>"000100000",
  15642=>"010010100",
  15643=>"011010111",
  15644=>"001100000",
  15645=>"100000010",
  15646=>"010010001",
  15647=>"010001000",
  15648=>"110111010",
  15649=>"100111101",
  15650=>"101111000",
  15651=>"000010000",
  15652=>"101010001",
  15653=>"011111011",
  15654=>"001001001",
  15655=>"111101100",
  15656=>"111111001",
  15657=>"010110000",
  15658=>"001111011",
  15659=>"000100011",
  15660=>"110000110",
  15661=>"000000000",
  15662=>"101110000",
  15663=>"001001001",
  15664=>"100101100",
  15665=>"010001000",
  15666=>"110111101",
  15667=>"010011101",
  15668=>"110101110",
  15669=>"010100001",
  15670=>"110100110",
  15671=>"001001111",
  15672=>"000000111",
  15673=>"110110101",
  15674=>"101110000",
  15675=>"111110001",
  15676=>"110101101",
  15677=>"001100011",
  15678=>"011110000",
  15679=>"100100111",
  15680=>"111111111",
  15681=>"110001010",
  15682=>"101010001",
  15683=>"111000101",
  15684=>"011001111",
  15685=>"001101101",
  15686=>"010100011",
  15687=>"110000000",
  15688=>"111011011",
  15689=>"110010010",
  15690=>"111100100",
  15691=>"011000010",
  15692=>"011011100",
  15693=>"111100101",
  15694=>"101110000",
  15695=>"111101101",
  15696=>"011110111",
  15697=>"000110000",
  15698=>"001011011",
  15699=>"010100011",
  15700=>"101000001",
  15701=>"100011000",
  15702=>"010011011",
  15703=>"000011011",
  15704=>"010001110",
  15705=>"011101111",
  15706=>"100110000",
  15707=>"100101110",
  15708=>"101010010",
  15709=>"111110111",
  15710=>"000011011",
  15711=>"101101101",
  15712=>"010001010",
  15713=>"010000011",
  15714=>"010110010",
  15715=>"011110011",
  15716=>"001000111",
  15717=>"100101011",
  15718=>"101111011",
  15719=>"111011111",
  15720=>"010101101",
  15721=>"000011110",
  15722=>"110001100",
  15723=>"001111000",
  15724=>"110011101",
  15725=>"110110110",
  15726=>"110011001",
  15727=>"010100011",
  15728=>"111111101",
  15729=>"000010111",
  15730=>"100111100",
  15731=>"101101110",
  15732=>"011111001",
  15733=>"010011000",
  15734=>"101001111",
  15735=>"100010110",
  15736=>"001110111",
  15737=>"100110111",
  15738=>"111010110",
  15739=>"100000000",
  15740=>"111001101",
  15741=>"001111010",
  15742=>"100100101",
  15743=>"111001110",
  15744=>"110111110",
  15745=>"001111100",
  15746=>"000001100",
  15747=>"100010111",
  15748=>"001000001",
  15749=>"010000111",
  15750=>"011101111",
  15751=>"100100111",
  15752=>"101101101",
  15753=>"010001111",
  15754=>"111101100",
  15755=>"001111010",
  15756=>"010010100",
  15757=>"001010100",
  15758=>"001001000",
  15759=>"010011111",
  15760=>"101110100",
  15761=>"011101100",
  15762=>"111110111",
  15763=>"111100001",
  15764=>"110101011",
  15765=>"010101011",
  15766=>"010000010",
  15767=>"000010010",
  15768=>"010111010",
  15769=>"010101100",
  15770=>"110011101",
  15771=>"111011011",
  15772=>"010010010",
  15773=>"001000000",
  15774=>"110001010",
  15775=>"100001101",
  15776=>"011100000",
  15777=>"110111110",
  15778=>"010110100",
  15779=>"100110110",
  15780=>"011100001",
  15781=>"010010110",
  15782=>"000011010",
  15783=>"010000010",
  15784=>"111100000",
  15785=>"011001111",
  15786=>"110010001",
  15787=>"010110100",
  15788=>"111111000",
  15789=>"100101101",
  15790=>"000110010",
  15791=>"111110101",
  15792=>"111001001",
  15793=>"101100010",
  15794=>"111100110",
  15795=>"101100001",
  15796=>"101001010",
  15797=>"001111010",
  15798=>"101000110",
  15799=>"000011101",
  15800=>"101111100",
  15801=>"000101111",
  15802=>"101010011",
  15803=>"011001101",
  15804=>"011000001",
  15805=>"000011011",
  15806=>"001101001",
  15807=>"100010011",
  15808=>"110100000",
  15809=>"000100111",
  15810=>"000010001",
  15811=>"100010110",
  15812=>"110110010",
  15813=>"001001111",
  15814=>"011010110",
  15815=>"001000110",
  15816=>"001010101",
  15817=>"110000011",
  15818=>"001000011",
  15819=>"110100100",
  15820=>"010101001",
  15821=>"000011100",
  15822=>"100111111",
  15823=>"011110010",
  15824=>"001010011",
  15825=>"010000110",
  15826=>"010100110",
  15827=>"000100001",
  15828=>"111101101",
  15829=>"011101001",
  15830=>"011001001",
  15831=>"000011111",
  15832=>"010110110",
  15833=>"010110001",
  15834=>"000010001",
  15835=>"011100000",
  15836=>"110111011",
  15837=>"101100000",
  15838=>"110110010",
  15839=>"101011000",
  15840=>"010100111",
  15841=>"000011100",
  15842=>"110000101",
  15843=>"110110111",
  15844=>"011111101",
  15845=>"101000101",
  15846=>"100111000",
  15847=>"000011111",
  15848=>"010001100",
  15849=>"001010010",
  15850=>"101011110",
  15851=>"110001101",
  15852=>"000110110",
  15853=>"110111110",
  15854=>"100011011",
  15855=>"100100001",
  15856=>"111000000",
  15857=>"111000011",
  15858=>"101100101",
  15859=>"000001100",
  15860=>"110100111",
  15861=>"011010110",
  15862=>"001010010",
  15863=>"101000101",
  15864=>"100101101",
  15865=>"100000000",
  15866=>"011010110",
  15867=>"101011001",
  15868=>"000100011",
  15869=>"101011010",
  15870=>"001101001",
  15871=>"110111111",
  15872=>"100011000",
  15873=>"100101011",
  15874=>"000111011",
  15875=>"101101111",
  15876=>"011101010",
  15877=>"101111111",
  15878=>"110001011",
  15879=>"111001110",
  15880=>"110110001",
  15881=>"101011101",
  15882=>"000010100",
  15883=>"111111101",
  15884=>"001011000",
  15885=>"011001100",
  15886=>"101111110",
  15887=>"100010010",
  15888=>"111101011",
  15889=>"000100001",
  15890=>"011011011",
  15891=>"111111001",
  15892=>"111001100",
  15893=>"110100001",
  15894=>"011011101",
  15895=>"001000101",
  15896=>"100000010",
  15897=>"101100110",
  15898=>"001110010",
  15899=>"111110010",
  15900=>"001110101",
  15901=>"010110011",
  15902=>"011110111",
  15903=>"111101010",
  15904=>"111110100",
  15905=>"001010100",
  15906=>"111101111",
  15907=>"001010111",
  15908=>"011010011",
  15909=>"111101001",
  15910=>"111111001",
  15911=>"000001010",
  15912=>"010001100",
  15913=>"101100010",
  15914=>"010100101",
  15915=>"101011010",
  15916=>"010001111",
  15917=>"001001111",
  15918=>"010001000",
  15919=>"110011000",
  15920=>"010010100",
  15921=>"010011100",
  15922=>"001111110",
  15923=>"100000010",
  15924=>"000011111",
  15925=>"000110010",
  15926=>"010101001",
  15927=>"010011100",
  15928=>"110101111",
  15929=>"101100111",
  15930=>"011000111",
  15931=>"000011101",
  15932=>"011111000",
  15933=>"000110110",
  15934=>"101100111",
  15935=>"101011101",
  15936=>"100100001",
  15937=>"010001000",
  15938=>"000011011",
  15939=>"111100100",
  15940=>"001000111",
  15941=>"100010010",
  15942=>"010000001",
  15943=>"101001100",
  15944=>"101001000",
  15945=>"110001000",
  15946=>"110001001",
  15947=>"001001011",
  15948=>"100011011",
  15949=>"001111100",
  15950=>"111111111",
  15951=>"110111110",
  15952=>"001101110",
  15953=>"011100011",
  15954=>"010001111",
  15955=>"001110001",
  15956=>"110000110",
  15957=>"101100101",
  15958=>"111111101",
  15959=>"001101100",
  15960=>"101000010",
  15961=>"001001011",
  15962=>"011100011",
  15963=>"001000011",
  15964=>"010101001",
  15965=>"011011011",
  15966=>"111011010",
  15967=>"100001011",
  15968=>"100101111",
  15969=>"000100110",
  15970=>"010100100",
  15971=>"011011111",
  15972=>"110001101",
  15973=>"000010101",
  15974=>"100011010",
  15975=>"101001110",
  15976=>"100111111",
  15977=>"000100001",
  15978=>"101010000",
  15979=>"101110000",
  15980=>"010110010",
  15981=>"111111001",
  15982=>"101001000",
  15983=>"001100100",
  15984=>"010101010",
  15985=>"000101111",
  15986=>"111000110",
  15987=>"011100101",
  15988=>"100011011",
  15989=>"111101011",
  15990=>"111001001",
  15991=>"001110000",
  15992=>"011100111",
  15993=>"011100100",
  15994=>"011110110",
  15995=>"101101100",
  15996=>"010101011",
  15997=>"010111111",
  15998=>"001100000",
  15999=>"111010010",
  16000=>"110100011",
  16001=>"110100011",
  16002=>"001111111",
  16003=>"101011111",
  16004=>"111111101",
  16005=>"000110111",
  16006=>"011111000",
  16007=>"110001000",
  16008=>"100000101",
  16009=>"111100001",
  16010=>"110000011",
  16011=>"010001011",
  16012=>"100100000",
  16013=>"001000001",
  16014=>"010000100",
  16015=>"000001111",
  16016=>"110001101",
  16017=>"110001111",
  16018=>"101010010",
  16019=>"101001101",
  16020=>"011110100",
  16021=>"010011110",
  16022=>"010001011",
  16023=>"010111111",
  16024=>"111011111",
  16025=>"010011100",
  16026=>"000010011",
  16027=>"010011010",
  16028=>"100000010",
  16029=>"000111000",
  16030=>"010001111",
  16031=>"000101111",
  16032=>"011001111",
  16033=>"101001001",
  16034=>"110111001",
  16035=>"100100010",
  16036=>"000000001",
  16037=>"111110110",
  16038=>"000100011",
  16039=>"000111100",
  16040=>"111100001",
  16041=>"101100000",
  16042=>"100000010",
  16043=>"011100010",
  16044=>"101001010",
  16045=>"000010011",
  16046=>"001110010",
  16047=>"010000010",
  16048=>"000000110",
  16049=>"000011010",
  16050=>"101111100",
  16051=>"101011110",
  16052=>"110010001",
  16053=>"101011100",
  16054=>"100100100",
  16055=>"100101101",
  16056=>"011101010",
  16057=>"110000000",
  16058=>"111111100",
  16059=>"100011000",
  16060=>"110111110",
  16061=>"100000011",
  16062=>"010010110",
  16063=>"011110100",
  16064=>"010110100",
  16065=>"010110101",
  16066=>"011001110",
  16067=>"011001000",
  16068=>"101101110",
  16069=>"001100110",
  16070=>"010110100",
  16071=>"111111101",
  16072=>"001100011",
  16073=>"000010110",
  16074=>"110010000",
  16075=>"000100110",
  16076=>"010001111",
  16077=>"011000111",
  16078=>"010100010",
  16079=>"100000110",
  16080=>"111010101",
  16081=>"110100010",
  16082=>"110011110",
  16083=>"101010100",
  16084=>"010110010",
  16085=>"000110001",
  16086=>"011010010",
  16087=>"000100101",
  16088=>"101011111",
  16089=>"011010100",
  16090=>"101010001",
  16091=>"001010000",
  16092=>"100110010",
  16093=>"110110111",
  16094=>"100010010",
  16095=>"110111000",
  16096=>"110111111",
  16097=>"000110001",
  16098=>"111100110",
  16099=>"001110111",
  16100=>"100000001",
  16101=>"100000011",
  16102=>"111110001",
  16103=>"101011111",
  16104=>"100101111",
  16105=>"110001001",
  16106=>"000010100",
  16107=>"000000001",
  16108=>"000110001",
  16109=>"001110011",
  16110=>"111101001",
  16111=>"010100010",
  16112=>"010100011",
  16113=>"101010010",
  16114=>"011101001",
  16115=>"110110111",
  16116=>"001011101",
  16117=>"011111111",
  16118=>"011001111",
  16119=>"110010110",
  16120=>"010011001",
  16121=>"000010110",
  16122=>"000010011",
  16123=>"100010111",
  16124=>"000110011",
  16125=>"000111001",
  16126=>"011001111",
  16127=>"101100100",
  16128=>"010011011",
  16129=>"111100011",
  16130=>"010000101",
  16131=>"110011011",
  16132=>"010010000",
  16133=>"111100101",
  16134=>"001111000",
  16135=>"100000110",
  16136=>"001101010",
  16137=>"110110110",
  16138=>"010110001",
  16139=>"001101111",
  16140=>"000111101",
  16141=>"010101100",
  16142=>"011011111",
  16143=>"001111011",
  16144=>"001111101",
  16145=>"100001111",
  16146=>"111101011",
  16147=>"011110101",
  16148=>"001011000",
  16149=>"101010110",
  16150=>"011100001",
  16151=>"110110010",
  16152=>"001001111",
  16153=>"001001101",
  16154=>"011000010",
  16155=>"101011111",
  16156=>"101100010",
  16157=>"101110000",
  16158=>"000000011",
  16159=>"001000111",
  16160=>"100001111",
  16161=>"010101110",
  16162=>"101010100",
  16163=>"010110101",
  16164=>"000101010",
  16165=>"011100001",
  16166=>"111101001",
  16167=>"111111101",
  16168=>"011001011",
  16169=>"000010100",
  16170=>"111011010",
  16171=>"100110100",
  16172=>"001001000",
  16173=>"001100110",
  16174=>"111110011",
  16175=>"001110111",
  16176=>"001100110",
  16177=>"110101111",
  16178=>"100101100",
  16179=>"110001011",
  16180=>"011100101",
  16181=>"110010111",
  16182=>"001000000",
  16183=>"000010101",
  16184=>"001011010",
  16185=>"111110010",
  16186=>"000101010",
  16187=>"001001011",
  16188=>"101000000",
  16189=>"001110111",
  16190=>"101111101",
  16191=>"000001111",
  16192=>"110001111",
  16193=>"110100000",
  16194=>"010100101",
  16195=>"010000010",
  16196=>"010111000",
  16197=>"110011000",
  16198=>"110000000",
  16199=>"101100111",
  16200=>"100111110",
  16201=>"100110001",
  16202=>"000001111",
  16203=>"111101110",
  16204=>"010100100",
  16205=>"011000100",
  16206=>"110111110",
  16207=>"001101111",
  16208=>"010101011",
  16209=>"001111101",
  16210=>"101110100",
  16211=>"000000011",
  16212=>"110100000",
  16213=>"010111111",
  16214=>"000010111",
  16215=>"100110011",
  16216=>"101000000",
  16217=>"001100111",
  16218=>"001101011",
  16219=>"000010011",
  16220=>"101000001",
  16221=>"000000100",
  16222=>"101011001",
  16223=>"111100111",
  16224=>"011110011",
  16225=>"011111111",
  16226=>"000011011",
  16227=>"111111101",
  16228=>"010111111",
  16229=>"000001110",
  16230=>"000011111",
  16231=>"111000111",
  16232=>"000001111",
  16233=>"101101001",
  16234=>"101011000",
  16235=>"110101111",
  16236=>"100010110",
  16237=>"000010000",
  16238=>"011011101",
  16239=>"110101111",
  16240=>"110000010",
  16241=>"101010111",
  16242=>"001101110",
  16243=>"100001100",
  16244=>"011100011",
  16245=>"101111100",
  16246=>"001110110",
  16247=>"111101111",
  16248=>"101101011",
  16249=>"001011000",
  16250=>"000110000",
  16251=>"101110010",
  16252=>"011100001",
  16253=>"101111011",
  16254=>"011010000",
  16255=>"001001001",
  16256=>"001110111",
  16257=>"110101000",
  16258=>"111111000",
  16259=>"100001001",
  16260=>"100000110",
  16261=>"101110000",
  16262=>"001001000",
  16263=>"111001110",
  16264=>"101011100",
  16265=>"011101011",
  16266=>"111111111",
  16267=>"100101101",
  16268=>"000110000",
  16269=>"101100001",
  16270=>"111001111",
  16271=>"111010011",
  16272=>"111100000",
  16273=>"101111001",
  16274=>"111111000",
  16275=>"011101111",
  16276=>"111110110",
  16277=>"010010001",
  16278=>"000110100",
  16279=>"001010010",
  16280=>"001111111",
  16281=>"111100101",
  16282=>"101111011",
  16283=>"101110111",
  16284=>"111011100",
  16285=>"000000110",
  16286=>"110100000",
  16287=>"010000011",
  16288=>"010010101",
  16289=>"011100100",
  16290=>"000110001",
  16291=>"011010100",
  16292=>"100011010",
  16293=>"011101101",
  16294=>"000011111",
  16295=>"101111011",
  16296=>"110001110",
  16297=>"000010011",
  16298=>"001001101",
  16299=>"100000100",
  16300=>"001010100",
  16301=>"111100001",
  16302=>"101111101",
  16303=>"101100111",
  16304=>"000001010",
  16305=>"000100010",
  16306=>"101101010",
  16307=>"111110110",
  16308=>"110100111",
  16309=>"000001111",
  16310=>"000010000",
  16311=>"001111101",
  16312=>"011111101",
  16313=>"110001110",
  16314=>"011001010",
  16315=>"110110110",
  16316=>"010000000",
  16317=>"001000101",
  16318=>"101101000",
  16319=>"110001111",
  16320=>"110000000",
  16321=>"100111111",
  16322=>"111011010",
  16323=>"011001010",
  16324=>"111001000",
  16325=>"000111111",
  16326=>"000001000",
  16327=>"100001101",
  16328=>"010111010",
  16329=>"001111000",
  16330=>"010010011",
  16331=>"000010001",
  16332=>"111011001",
  16333=>"101110011",
  16334=>"100110111",
  16335=>"100111001",
  16336=>"101000110",
  16337=>"100111111",
  16338=>"000110010",
  16339=>"010111011",
  16340=>"000011000",
  16341=>"101101001",
  16342=>"101011100",
  16343=>"111110001",
  16344=>"010111101",
  16345=>"101100010",
  16346=>"101001101",
  16347=>"100111000",
  16348=>"110011000",
  16349=>"000101011",
  16350=>"000000000",
  16351=>"011001110",
  16352=>"110111011",
  16353=>"000000101",
  16354=>"110111001",
  16355=>"011010001",
  16356=>"110010010",
  16357=>"000111101",
  16358=>"111011100",
  16359=>"001110101",
  16360=>"001110111",
  16361=>"100011001",
  16362=>"101000100",
  16363=>"000001101",
  16364=>"010111110",
  16365=>"111111010",
  16366=>"110010010",
  16367=>"011110110",
  16368=>"011111000",
  16369=>"010111111",
  16370=>"101000100",
  16371=>"000011001",
  16372=>"111001100",
  16373=>"100111101",
  16374=>"010001100",
  16375=>"101011111",
  16376=>"100110000",
  16377=>"000000110",
  16378=>"111100101",
  16379=>"000010111",
  16380=>"011101001",
  16381=>"001010110",
  16382=>"000011101",
  16383=>"011100011",
  16384=>"111110111",
  16385=>"100001111",
  16386=>"111010111",
  16387=>"011110100",
  16388=>"101101100",
  16389=>"111001111",
  16390=>"011010010",
  16391=>"111110010",
  16392=>"011001001",
  16393=>"100000000",
  16394=>"011111111",
  16395=>"110101111",
  16396=>"010010001",
  16397=>"100110101",
  16398=>"111010001",
  16399=>"010110011",
  16400=>"110000100",
  16401=>"110110011",
  16402=>"100001000",
  16403=>"000011000",
  16404=>"111111011",
  16405=>"110001101",
  16406=>"001110010",
  16407=>"001010101",
  16408=>"010111001",
  16409=>"111100101",
  16410=>"001001100",
  16411=>"100101100",
  16412=>"011100101",
  16413=>"011111001",
  16414=>"110100001",
  16415=>"001000001",
  16416=>"111011111",
  16417=>"101111110",
  16418=>"100000010",
  16419=>"010000101",
  16420=>"111101001",
  16421=>"011001100",
  16422=>"010010010",
  16423=>"110011001",
  16424=>"000111001",
  16425=>"000101111",
  16426=>"100000111",
  16427=>"011110010",
  16428=>"001011001",
  16429=>"000000100",
  16430=>"101010010",
  16431=>"110100001",
  16432=>"010110100",
  16433=>"111010101",
  16434=>"011100110",
  16435=>"100110001",
  16436=>"101101111",
  16437=>"001011101",
  16438=>"111011101",
  16439=>"110000000",
  16440=>"001100101",
  16441=>"111111010",
  16442=>"001101110",
  16443=>"000000010",
  16444=>"101001110",
  16445=>"001100101",
  16446=>"011011111",
  16447=>"111111100",
  16448=>"000010100",
  16449=>"111001110",
  16450=>"001010110",
  16451=>"100100101",
  16452=>"000000010",
  16453=>"001101101",
  16454=>"100010110",
  16455=>"010011000",
  16456=>"101111010",
  16457=>"111001111",
  16458=>"100101111",
  16459=>"011001010",
  16460=>"110010111",
  16461=>"000110010",
  16462=>"100000011",
  16463=>"111010010",
  16464=>"101110110",
  16465=>"010111001",
  16466=>"110110010",
  16467=>"100110100",
  16468=>"000011001",
  16469=>"101100000",
  16470=>"110100100",
  16471=>"001101110",
  16472=>"101010101",
  16473=>"111100101",
  16474=>"001000101",
  16475=>"101111011",
  16476=>"011101010",
  16477=>"110010001",
  16478=>"111001111",
  16479=>"000110011",
  16480=>"001001111",
  16481=>"110000000",
  16482=>"011011001",
  16483=>"110001001",
  16484=>"100001101",
  16485=>"110011001",
  16486=>"110000110",
  16487=>"000011100",
  16488=>"011000001",
  16489=>"110001010",
  16490=>"001110110",
  16491=>"100111110",
  16492=>"101110001",
  16493=>"101101111",
  16494=>"110101000",
  16495=>"111110111",
  16496=>"111011110",
  16497=>"110101101",
  16498=>"000000100",
  16499=>"011010111",
  16500=>"010111100",
  16501=>"010011010",
  16502=>"110111011",
  16503=>"110101011",
  16504=>"111010110",
  16505=>"001001011",
  16506=>"111101011",
  16507=>"001100001",
  16508=>"111110100",
  16509=>"010000100",
  16510=>"101000101",
  16511=>"111100010",
  16512=>"100000010",
  16513=>"100111010",
  16514=>"000100010",
  16515=>"101100001",
  16516=>"000101101",
  16517=>"101011100",
  16518=>"100111111",
  16519=>"100011000",
  16520=>"110110011",
  16521=>"001101111",
  16522=>"011011101",
  16523=>"110111101",
  16524=>"110101111",
  16525=>"001111000",
  16526=>"010001010",
  16527=>"011101101",
  16528=>"011010011",
  16529=>"101111010",
  16530=>"000101000",
  16531=>"011110101",
  16532=>"111101001",
  16533=>"000000011",
  16534=>"101000010",
  16535=>"101010100",
  16536=>"100001110",
  16537=>"110111110",
  16538=>"100011110",
  16539=>"110011100",
  16540=>"111110101",
  16541=>"000000110",
  16542=>"010110110",
  16543=>"000010010",
  16544=>"111111011",
  16545=>"111110000",
  16546=>"100111111",
  16547=>"001010101",
  16548=>"001010010",
  16549=>"111011001",
  16550=>"101001010",
  16551=>"000000101",
  16552=>"001111010",
  16553=>"000101011",
  16554=>"000000111",
  16555=>"111100010",
  16556=>"000000001",
  16557=>"101111110",
  16558=>"001101100",
  16559=>"010110111",
  16560=>"011100100",
  16561=>"001111111",
  16562=>"000111001",
  16563=>"010001111",
  16564=>"000011111",
  16565=>"100101011",
  16566=>"011101111",
  16567=>"100101101",
  16568=>"011010110",
  16569=>"010101110",
  16570=>"101101111",
  16571=>"110001010",
  16572=>"001011011",
  16573=>"000001111",
  16574=>"011000011",
  16575=>"010111101",
  16576=>"001111000",
  16577=>"000111110",
  16578=>"001100000",
  16579=>"100101001",
  16580=>"011011001",
  16581=>"101101111",
  16582=>"110110001",
  16583=>"001111101",
  16584=>"110000100",
  16585=>"110000000",
  16586=>"100011001",
  16587=>"000000110",
  16588=>"010110111",
  16589=>"001000100",
  16590=>"111011101",
  16591=>"011000111",
  16592=>"110001001",
  16593=>"100110101",
  16594=>"011001110",
  16595=>"101001111",
  16596=>"001010111",
  16597=>"001011011",
  16598=>"011001111",
  16599=>"101011010",
  16600=>"010000100",
  16601=>"111110010",
  16602=>"111110011",
  16603=>"011101101",
  16604=>"010011011",
  16605=>"000100001",
  16606=>"110010100",
  16607=>"000000011",
  16608=>"100011011",
  16609=>"000011011",
  16610=>"011001100",
  16611=>"111100110",
  16612=>"111101101",
  16613=>"001111111",
  16614=>"000101011",
  16615=>"111111101",
  16616=>"110001001",
  16617=>"000010010",
  16618=>"010010001",
  16619=>"101101100",
  16620=>"000011000",
  16621=>"111111010",
  16622=>"001000110",
  16623=>"111000000",
  16624=>"100110011",
  16625=>"001010011",
  16626=>"110011111",
  16627=>"110010010",
  16628=>"101100010",
  16629=>"100010111",
  16630=>"111110110",
  16631=>"001011011",
  16632=>"101011001",
  16633=>"000111000",
  16634=>"000110000",
  16635=>"010001000",
  16636=>"011011100",
  16637=>"011110001",
  16638=>"110001000",
  16639=>"100001110",
  16640=>"000110011",
  16641=>"100110000",
  16642=>"111101000",
  16643=>"011110100",
  16644=>"100000001",
  16645=>"001010110",
  16646=>"101101111",
  16647=>"100100110",
  16648=>"100100100",
  16649=>"010110000",
  16650=>"110100101",
  16651=>"110011111",
  16652=>"101011100",
  16653=>"000101110",
  16654=>"000100001",
  16655=>"111111011",
  16656=>"000011100",
  16657=>"110111111",
  16658=>"110110001",
  16659=>"010010011",
  16660=>"011001010",
  16661=>"110110000",
  16662=>"010111010",
  16663=>"101001010",
  16664=>"111010100",
  16665=>"011000010",
  16666=>"001110111",
  16667=>"000010001",
  16668=>"111000101",
  16669=>"000110011",
  16670=>"101001111",
  16671=>"111011111",
  16672=>"011100110",
  16673=>"001110010",
  16674=>"001111100",
  16675=>"010001010",
  16676=>"111111110",
  16677=>"100011110",
  16678=>"000110101",
  16679=>"100111000",
  16680=>"001010111",
  16681=>"010100000",
  16682=>"101101101",
  16683=>"110010100",
  16684=>"010000001",
  16685=>"001110000",
  16686=>"110111011",
  16687=>"111011011",
  16688=>"001111011",
  16689=>"101111101",
  16690=>"110011010",
  16691=>"100101101",
  16692=>"011001001",
  16693=>"100010000",
  16694=>"101000001",
  16695=>"111111000",
  16696=>"000101100",
  16697=>"111010011",
  16698=>"001110111",
  16699=>"010000010",
  16700=>"111011110",
  16701=>"011111001",
  16702=>"010100001",
  16703=>"110011010",
  16704=>"111110101",
  16705=>"000010000",
  16706=>"011100011",
  16707=>"111010111",
  16708=>"101101111",
  16709=>"111010111",
  16710=>"011011110",
  16711=>"101000011",
  16712=>"010111011",
  16713=>"110011010",
  16714=>"101000110",
  16715=>"110011001",
  16716=>"011100111",
  16717=>"101110110",
  16718=>"110011001",
  16719=>"111111111",
  16720=>"101111111",
  16721=>"111001000",
  16722=>"100011000",
  16723=>"111010010",
  16724=>"000111000",
  16725=>"100101011",
  16726=>"110010000",
  16727=>"101100010",
  16728=>"100001101",
  16729=>"101111000",
  16730=>"110000101",
  16731=>"000111111",
  16732=>"011001101",
  16733=>"011000001",
  16734=>"101100011",
  16735=>"011101100",
  16736=>"000100110",
  16737=>"001110101",
  16738=>"001110110",
  16739=>"101101000",
  16740=>"011100111",
  16741=>"110110111",
  16742=>"101010001",
  16743=>"111011011",
  16744=>"001000100",
  16745=>"111111111",
  16746=>"100101101",
  16747=>"111011110",
  16748=>"000001000",
  16749=>"000001011",
  16750=>"001011110",
  16751=>"001110110",
  16752=>"101100110",
  16753=>"111011000",
  16754=>"111100000",
  16755=>"110110111",
  16756=>"110011101",
  16757=>"001101111",
  16758=>"101011010",
  16759=>"011111110",
  16760=>"111001011",
  16761=>"100101001",
  16762=>"011010010",
  16763=>"101001011",
  16764=>"011101010",
  16765=>"100100011",
  16766=>"111110110",
  16767=>"001100011",
  16768=>"000001011",
  16769=>"011000100",
  16770=>"111001110",
  16771=>"100110100",
  16772=>"111110011",
  16773=>"111101101",
  16774=>"100000011",
  16775=>"110011000",
  16776=>"101001011",
  16777=>"000010111",
  16778=>"101111101",
  16779=>"010100001",
  16780=>"101001001",
  16781=>"100101011",
  16782=>"111100111",
  16783=>"001110000",
  16784=>"111010100",
  16785=>"110010101",
  16786=>"010011010",
  16787=>"001100010",
  16788=>"111100100",
  16789=>"100000010",
  16790=>"011010011",
  16791=>"100110001",
  16792=>"101000110",
  16793=>"001101111",
  16794=>"100000011",
  16795=>"000010011",
  16796=>"110110100",
  16797=>"010100100",
  16798=>"010101110",
  16799=>"010110000",
  16800=>"110111011",
  16801=>"001100111",
  16802=>"100100110",
  16803=>"010000001",
  16804=>"000000101",
  16805=>"001110100",
  16806=>"000001111",
  16807=>"101111111",
  16808=>"100011010",
  16809=>"001000111",
  16810=>"011011110",
  16811=>"111110111",
  16812=>"111101111",
  16813=>"100010010",
  16814=>"101000101",
  16815=>"011110011",
  16816=>"000101110",
  16817=>"001000001",
  16818=>"001000100",
  16819=>"011111111",
  16820=>"001010010",
  16821=>"101001000",
  16822=>"100100001",
  16823=>"100110101",
  16824=>"111111000",
  16825=>"101111010",
  16826=>"111101111",
  16827=>"101111000",
  16828=>"000000000",
  16829=>"100011010",
  16830=>"111100101",
  16831=>"010011100",
  16832=>"000101110",
  16833=>"111110001",
  16834=>"011000110",
  16835=>"000011110",
  16836=>"001010110",
  16837=>"011110100",
  16838=>"110001111",
  16839=>"000111111",
  16840=>"000011011",
  16841=>"001100101",
  16842=>"010101110",
  16843=>"000111100",
  16844=>"100110000",
  16845=>"010100011",
  16846=>"011001101",
  16847=>"110011000",
  16848=>"101101001",
  16849=>"111011101",
  16850=>"011001010",
  16851=>"111011010",
  16852=>"101011001",
  16853=>"110010111",
  16854=>"000101001",
  16855=>"111101111",
  16856=>"111001101",
  16857=>"100011110",
  16858=>"111010100",
  16859=>"111110010",
  16860=>"011110111",
  16861=>"011010110",
  16862=>"110000010",
  16863=>"000101110",
  16864=>"110110001",
  16865=>"100100001",
  16866=>"101110011",
  16867=>"011100100",
  16868=>"010101011",
  16869=>"001010010",
  16870=>"111010111",
  16871=>"111111001",
  16872=>"111101110",
  16873=>"100111111",
  16874=>"110111111",
  16875=>"011010101",
  16876=>"101011010",
  16877=>"010011101",
  16878=>"111001001",
  16879=>"010000110",
  16880=>"101001010",
  16881=>"000100000",
  16882=>"111000010",
  16883=>"111101110",
  16884=>"011011010",
  16885=>"110010000",
  16886=>"010001011",
  16887=>"000000000",
  16888=>"011110110",
  16889=>"100001010",
  16890=>"111101000",
  16891=>"011001000",
  16892=>"011010001",
  16893=>"111111001",
  16894=>"001010101",
  16895=>"000101111",
  16896=>"011100011",
  16897=>"101101110",
  16898=>"000010010",
  16899=>"001101100",
  16900=>"010110101",
  16901=>"010011111",
  16902=>"110010010",
  16903=>"110010001",
  16904=>"111001001",
  16905=>"100110000",
  16906=>"001100101",
  16907=>"110110110",
  16908=>"001111011",
  16909=>"011101011",
  16910=>"011010110",
  16911=>"110110011",
  16912=>"011110001",
  16913=>"000000000",
  16914=>"010000100",
  16915=>"111111001",
  16916=>"001110001",
  16917=>"101101110",
  16918=>"010001010",
  16919=>"111000000",
  16920=>"010100111",
  16921=>"110101000",
  16922=>"011101010",
  16923=>"110110110",
  16924=>"110110000",
  16925=>"111011100",
  16926=>"101110000",
  16927=>"011111100",
  16928=>"101100001",
  16929=>"001010010",
  16930=>"011111110",
  16931=>"110011111",
  16932=>"111101011",
  16933=>"010100100",
  16934=>"011011010",
  16935=>"000001110",
  16936=>"000010010",
  16937=>"101000000",
  16938=>"011001011",
  16939=>"101010011",
  16940=>"011101010",
  16941=>"101011111",
  16942=>"111111010",
  16943=>"101111010",
  16944=>"100100101",
  16945=>"011000010",
  16946=>"001110011",
  16947=>"011111111",
  16948=>"101111101",
  16949=>"111110110",
  16950=>"011100010",
  16951=>"001101000",
  16952=>"100110110",
  16953=>"111011111",
  16954=>"000100011",
  16955=>"101011111",
  16956=>"111001100",
  16957=>"110000110",
  16958=>"110000010",
  16959=>"001001100",
  16960=>"000110010",
  16961=>"011111010",
  16962=>"001100011",
  16963=>"101011011",
  16964=>"001100101",
  16965=>"001111011",
  16966=>"111011111",
  16967=>"001111000",
  16968=>"110100011",
  16969=>"101111010",
  16970=>"100100001",
  16971=>"010000010",
  16972=>"110000000",
  16973=>"100100100",
  16974=>"000001010",
  16975=>"001111100",
  16976=>"011011010",
  16977=>"010011000",
  16978=>"001111111",
  16979=>"010101111",
  16980=>"110111111",
  16981=>"111100010",
  16982=>"011111111",
  16983=>"100100001",
  16984=>"101000010",
  16985=>"000101001",
  16986=>"100111111",
  16987=>"110100011",
  16988=>"001111000",
  16989=>"000100110",
  16990=>"111000011",
  16991=>"011100010",
  16992=>"001100101",
  16993=>"010101000",
  16994=>"011111110",
  16995=>"100010001",
  16996=>"000111101",
  16997=>"110111110",
  16998=>"110100111",
  16999=>"011010011",
  17000=>"011001001",
  17001=>"100010010",
  17002=>"100100100",
  17003=>"111010011",
  17004=>"101101001",
  17005=>"001110110",
  17006=>"111100010",
  17007=>"010010001",
  17008=>"011111101",
  17009=>"000101001",
  17010=>"011101011",
  17011=>"110111110",
  17012=>"001111001",
  17013=>"001000101",
  17014=>"101011000",
  17015=>"100011100",
  17016=>"001010011",
  17017=>"111110011",
  17018=>"111111111",
  17019=>"101111001",
  17020=>"001111101",
  17021=>"110110001",
  17022=>"100001010",
  17023=>"010100000",
  17024=>"011010110",
  17025=>"110001011",
  17026=>"111000010",
  17027=>"110100011",
  17028=>"110100001",
  17029=>"110110010",
  17030=>"000101000",
  17031=>"011000000",
  17032=>"001001000",
  17033=>"100111111",
  17034=>"110011111",
  17035=>"000011010",
  17036=>"011101001",
  17037=>"000010010",
  17038=>"011000110",
  17039=>"010111011",
  17040=>"111011011",
  17041=>"011000001",
  17042=>"111100111",
  17043=>"000000111",
  17044=>"111001000",
  17045=>"011100001",
  17046=>"001001101",
  17047=>"100110111",
  17048=>"110111000",
  17049=>"110100011",
  17050=>"100101100",
  17051=>"010101101",
  17052=>"010000000",
  17053=>"100011110",
  17054=>"000110010",
  17055=>"001000000",
  17056=>"010100010",
  17057=>"011000101",
  17058=>"100011111",
  17059=>"000001001",
  17060=>"111010100",
  17061=>"110101111",
  17062=>"000011110",
  17063=>"000000100",
  17064=>"000111100",
  17065=>"101111111",
  17066=>"100111010",
  17067=>"111111101",
  17068=>"100001100",
  17069=>"111000100",
  17070=>"001101101",
  17071=>"100110101",
  17072=>"000101010",
  17073=>"100110111",
  17074=>"101001111",
  17075=>"111110110",
  17076=>"011011100",
  17077=>"001100000",
  17078=>"000111101",
  17079=>"110011100",
  17080=>"011110110",
  17081=>"001101111",
  17082=>"011010010",
  17083=>"000000000",
  17084=>"100100111",
  17085=>"010110101",
  17086=>"000101011",
  17087=>"100011000",
  17088=>"111000010",
  17089=>"001011000",
  17090=>"010110001",
  17091=>"100110000",
  17092=>"011111011",
  17093=>"100000001",
  17094=>"000010110",
  17095=>"000101010",
  17096=>"010100011",
  17097=>"010100010",
  17098=>"011111110",
  17099=>"101011001",
  17100=>"100110111",
  17101=>"011000010",
  17102=>"010010001",
  17103=>"111011101",
  17104=>"111000111",
  17105=>"010010011",
  17106=>"110011011",
  17107=>"001111101",
  17108=>"000101110",
  17109=>"010111101",
  17110=>"100010100",
  17111=>"101000111",
  17112=>"010111111",
  17113=>"111000111",
  17114=>"110001011",
  17115=>"011101111",
  17116=>"100001110",
  17117=>"101010100",
  17118=>"111011000",
  17119=>"100010010",
  17120=>"110000000",
  17121=>"011101110",
  17122=>"111111101",
  17123=>"110110111",
  17124=>"111111011",
  17125=>"010010000",
  17126=>"001100011",
  17127=>"110011111",
  17128=>"111101011",
  17129=>"000100001",
  17130=>"101010110",
  17131=>"011100011",
  17132=>"111001100",
  17133=>"110100000",
  17134=>"011010000",
  17135=>"110010000",
  17136=>"001000000",
  17137=>"101110110",
  17138=>"010100010",
  17139=>"000101110",
  17140=>"110011110",
  17141=>"000001000",
  17142=>"101110101",
  17143=>"101110001",
  17144=>"100100111",
  17145=>"101010001",
  17146=>"010000100",
  17147=>"100100111",
  17148=>"010011110",
  17149=>"010101000",
  17150=>"010011111",
  17151=>"101001110",
  17152=>"001011111",
  17153=>"111101011",
  17154=>"000000111",
  17155=>"010111000",
  17156=>"111100101",
  17157=>"010011011",
  17158=>"110100110",
  17159=>"101111101",
  17160=>"001111010",
  17161=>"100000011",
  17162=>"110000110",
  17163=>"001111110",
  17164=>"110110101",
  17165=>"011110010",
  17166=>"111010110",
  17167=>"101111100",
  17168=>"011010001",
  17169=>"011011011",
  17170=>"100111010",
  17171=>"011111000",
  17172=>"101010111",
  17173=>"010001001",
  17174=>"110000111",
  17175=>"101010111",
  17176=>"001110110",
  17177=>"001110000",
  17178=>"110101000",
  17179=>"100001110",
  17180=>"000011010",
  17181=>"000110011",
  17182=>"001111010",
  17183=>"011100001",
  17184=>"101011000",
  17185=>"100110010",
  17186=>"000000001",
  17187=>"001010011",
  17188=>"101110110",
  17189=>"000010011",
  17190=>"000011011",
  17191=>"001000110",
  17192=>"011100011",
  17193=>"011000100",
  17194=>"110101001",
  17195=>"101111101",
  17196=>"111000011",
  17197=>"000011110",
  17198=>"101101110",
  17199=>"001011100",
  17200=>"111011101",
  17201=>"010111001",
  17202=>"000010100",
  17203=>"101100010",
  17204=>"000110001",
  17205=>"001100010",
  17206=>"011000010",
  17207=>"100010111",
  17208=>"111111011",
  17209=>"011100111",
  17210=>"001111111",
  17211=>"000101101",
  17212=>"010010010",
  17213=>"001011101",
  17214=>"110001001",
  17215=>"010101011",
  17216=>"111101000",
  17217=>"100110000",
  17218=>"010110011",
  17219=>"000111010",
  17220=>"011011001",
  17221=>"101000001",
  17222=>"101000000",
  17223=>"011101100",
  17224=>"010011111",
  17225=>"011010110",
  17226=>"011011111",
  17227=>"011001000",
  17228=>"101011010",
  17229=>"110111100",
  17230=>"011111101",
  17231=>"110100011",
  17232=>"001101101",
  17233=>"011110010",
  17234=>"100101110",
  17235=>"000010100",
  17236=>"010100001",
  17237=>"011110100",
  17238=>"100001010",
  17239=>"110011011",
  17240=>"110101011",
  17241=>"111010011",
  17242=>"100011111",
  17243=>"000100110",
  17244=>"111011010",
  17245=>"100010101",
  17246=>"111000110",
  17247=>"011111111",
  17248=>"010000011",
  17249=>"111101011",
  17250=>"100110100",
  17251=>"100001110",
  17252=>"001110000",
  17253=>"101000100",
  17254=>"000011001",
  17255=>"010001010",
  17256=>"010110101",
  17257=>"011111110",
  17258=>"101011111",
  17259=>"000000101",
  17260=>"101111001",
  17261=>"101001101",
  17262=>"010100101",
  17263=>"100101110",
  17264=>"111001101",
  17265=>"100000000",
  17266=>"011001101",
  17267=>"000111010",
  17268=>"111111010",
  17269=>"010110011",
  17270=>"011000011",
  17271=>"000001010",
  17272=>"111011100",
  17273=>"110001000",
  17274=>"000110000",
  17275=>"100010011",
  17276=>"001111101",
  17277=>"101110100",
  17278=>"000000011",
  17279=>"010100000",
  17280=>"001111010",
  17281=>"111110001",
  17282=>"100110011",
  17283=>"101011101",
  17284=>"010011000",
  17285=>"011100001",
  17286=>"000111010",
  17287=>"100000010",
  17288=>"001000010",
  17289=>"001101011",
  17290=>"101010101",
  17291=>"000000111",
  17292=>"001101001",
  17293=>"001111101",
  17294=>"101000111",
  17295=>"011111011",
  17296=>"001000100",
  17297=>"111111011",
  17298=>"000010110",
  17299=>"101111110",
  17300=>"111001010",
  17301=>"110000100",
  17302=>"101000111",
  17303=>"101100101",
  17304=>"001101100",
  17305=>"001000101",
  17306=>"100111011",
  17307=>"101011001",
  17308=>"110010111",
  17309=>"011111100",
  17310=>"000010001",
  17311=>"101010011",
  17312=>"000010001",
  17313=>"001010001",
  17314=>"111100001",
  17315=>"101111101",
  17316=>"001100110",
  17317=>"000001011",
  17318=>"001011111",
  17319=>"111001101",
  17320=>"011001111",
  17321=>"001010111",
  17322=>"001101001",
  17323=>"101101101",
  17324=>"010011011",
  17325=>"001010100",
  17326=>"100000001",
  17327=>"101100101",
  17328=>"011011111",
  17329=>"111000111",
  17330=>"110110001",
  17331=>"100110011",
  17332=>"011101110",
  17333=>"100101011",
  17334=>"001011100",
  17335=>"010111100",
  17336=>"110110110",
  17337=>"111001011",
  17338=>"000001100",
  17339=>"111111100",
  17340=>"111111111",
  17341=>"111000000",
  17342=>"011001011",
  17343=>"101101111",
  17344=>"010000000",
  17345=>"001101011",
  17346=>"111111111",
  17347=>"001101110",
  17348=>"110011010",
  17349=>"010010101",
  17350=>"011001000",
  17351=>"100000000",
  17352=>"010000101",
  17353=>"001011001",
  17354=>"001010001",
  17355=>"000111111",
  17356=>"100110010",
  17357=>"000001101",
  17358=>"100001010",
  17359=>"010110010",
  17360=>"110110010",
  17361=>"111001101",
  17362=>"011110011",
  17363=>"001111111",
  17364=>"000101101",
  17365=>"011011111",
  17366=>"101111000",
  17367=>"111100101",
  17368=>"011111110",
  17369=>"111011101",
  17370=>"100101100",
  17371=>"001101000",
  17372=>"100111110",
  17373=>"111001001",
  17374=>"000101111",
  17375=>"110010011",
  17376=>"001111011",
  17377=>"100110011",
  17378=>"100010111",
  17379=>"100101000",
  17380=>"100111011",
  17381=>"000010000",
  17382=>"100010101",
  17383=>"011110100",
  17384=>"110111000",
  17385=>"001001011",
  17386=>"100011000",
  17387=>"000101001",
  17388=>"111110010",
  17389=>"001111000",
  17390=>"111001100",
  17391=>"101000111",
  17392=>"001010010",
  17393=>"001000011",
  17394=>"001110000",
  17395=>"001000010",
  17396=>"011100010",
  17397=>"100001100",
  17398=>"101111110",
  17399=>"011001110",
  17400=>"111101101",
  17401=>"000111010",
  17402=>"000001000",
  17403=>"001001111",
  17404=>"100010110",
  17405=>"011101100",
  17406=>"110111101",
  17407=>"000011101",
  17408=>"010000110",
  17409=>"111101000",
  17410=>"111000110",
  17411=>"100110110",
  17412=>"100011110",
  17413=>"111110001",
  17414=>"110111000",
  17415=>"011110100",
  17416=>"100100001",
  17417=>"101001111",
  17418=>"000000001",
  17419=>"100101000",
  17420=>"000001111",
  17421=>"001011110",
  17422=>"111100110",
  17423=>"110101000",
  17424=>"101010110",
  17425=>"110100101",
  17426=>"101010001",
  17427=>"110101100",
  17428=>"100110011",
  17429=>"111100001",
  17430=>"110001011",
  17431=>"010101000",
  17432=>"010111000",
  17433=>"001011101",
  17434=>"011110100",
  17435=>"001100001",
  17436=>"011001010",
  17437=>"001000000",
  17438=>"101010111",
  17439=>"101111000",
  17440=>"101010111",
  17441=>"001111010",
  17442=>"001100101",
  17443=>"001000000",
  17444=>"100010101",
  17445=>"111000101",
  17446=>"010100110",
  17447=>"000001110",
  17448=>"111100000",
  17449=>"100000100",
  17450=>"101001111",
  17451=>"000110011",
  17452=>"000110000",
  17453=>"011000000",
  17454=>"000110010",
  17455=>"111111101",
  17456=>"100011111",
  17457=>"111011011",
  17458=>"110111110",
  17459=>"111000100",
  17460=>"110011001",
  17461=>"001100111",
  17462=>"101010001",
  17463=>"110100010",
  17464=>"110001011",
  17465=>"011011011",
  17466=>"000011111",
  17467=>"111101011",
  17468=>"111100101",
  17469=>"101001101",
  17470=>"110111001",
  17471=>"011101010",
  17472=>"100100101",
  17473=>"000010001",
  17474=>"000011010",
  17475=>"111010111",
  17476=>"000010001",
  17477=>"010001101",
  17478=>"011001111",
  17479=>"000001011",
  17480=>"100100100",
  17481=>"111010001",
  17482=>"010100000",
  17483=>"110100110",
  17484=>"111110110",
  17485=>"100000000",
  17486=>"100000011",
  17487=>"000100001",
  17488=>"111011001",
  17489=>"000100111",
  17490=>"110001010",
  17491=>"101000000",
  17492=>"100110100",
  17493=>"000110010",
  17494=>"000111000",
  17495=>"001101000",
  17496=>"010100101",
  17497=>"000111100",
  17498=>"101111110",
  17499=>"000010001",
  17500=>"101011101",
  17501=>"010101010",
  17502=>"011000100",
  17503=>"011111000",
  17504=>"000001100",
  17505=>"110101111",
  17506=>"011010000",
  17507=>"111111100",
  17508=>"100110010",
  17509=>"100101110",
  17510=>"011000100",
  17511=>"110110010",
  17512=>"111110000",
  17513=>"110011000",
  17514=>"100110111",
  17515=>"010000001",
  17516=>"000101111",
  17517=>"111110001",
  17518=>"000110001",
  17519=>"001000111",
  17520=>"001101110",
  17521=>"110101010",
  17522=>"101011101",
  17523=>"001010100",
  17524=>"000000110",
  17525=>"000110010",
  17526=>"010111100",
  17527=>"011010010",
  17528=>"000100001",
  17529=>"011010110",
  17530=>"100101111",
  17531=>"100000000",
  17532=>"101000100",
  17533=>"011000000",
  17534=>"010110101",
  17535=>"001001100",
  17536=>"000110011",
  17537=>"011110110",
  17538=>"000110010",
  17539=>"110011011",
  17540=>"000100010",
  17541=>"101000111",
  17542=>"111010010",
  17543=>"000000000",
  17544=>"111100010",
  17545=>"110010011",
  17546=>"100100101",
  17547=>"000011010",
  17548=>"000011001",
  17549=>"010001100",
  17550=>"001001011",
  17551=>"000110100",
  17552=>"101010001",
  17553=>"101011110",
  17554=>"100000100",
  17555=>"100001101",
  17556=>"111111110",
  17557=>"111100111",
  17558=>"111101011",
  17559=>"111110010",
  17560=>"111001001",
  17561=>"001100000",
  17562=>"000001011",
  17563=>"001100101",
  17564=>"000010111",
  17565=>"001010100",
  17566=>"101010001",
  17567=>"010101100",
  17568=>"000100110",
  17569=>"111011011",
  17570=>"110011001",
  17571=>"100000010",
  17572=>"010010011",
  17573=>"011101101",
  17574=>"100100100",
  17575=>"010000111",
  17576=>"100000000",
  17577=>"000000110",
  17578=>"111011000",
  17579=>"001001000",
  17580=>"011010100",
  17581=>"010100101",
  17582=>"110100110",
  17583=>"111001111",
  17584=>"110000011",
  17585=>"010010111",
  17586=>"110010010",
  17587=>"000110110",
  17588=>"011000111",
  17589=>"100000101",
  17590=>"110111001",
  17591=>"000100000",
  17592=>"010011111",
  17593=>"011001000",
  17594=>"011011110",
  17595=>"101011110",
  17596=>"000111100",
  17597=>"011010110",
  17598=>"101001111",
  17599=>"000011001",
  17600=>"001111100",
  17601=>"100111110",
  17602=>"111000111",
  17603=>"010010011",
  17604=>"101101011",
  17605=>"011000101",
  17606=>"010100000",
  17607=>"001010010",
  17608=>"000101001",
  17609=>"000001100",
  17610=>"100110000",
  17611=>"100000010",
  17612=>"101111100",
  17613=>"110111100",
  17614=>"011111110",
  17615=>"000110010",
  17616=>"100011100",
  17617=>"100000100",
  17618=>"000100000",
  17619=>"111001101",
  17620=>"110110011",
  17621=>"111111111",
  17622=>"011000110",
  17623=>"101111100",
  17624=>"100001011",
  17625=>"010111010",
  17626=>"111010101",
  17627=>"110111001",
  17628=>"010110111",
  17629=>"111111000",
  17630=>"101001001",
  17631=>"101000001",
  17632=>"101010001",
  17633=>"110000001",
  17634=>"111010001",
  17635=>"000000110",
  17636=>"101100101",
  17637=>"001000000",
  17638=>"110000101",
  17639=>"111111000",
  17640=>"001010101",
  17641=>"010101110",
  17642=>"000100001",
  17643=>"010010100",
  17644=>"011110000",
  17645=>"000000000",
  17646=>"001001011",
  17647=>"111111110",
  17648=>"111010111",
  17649=>"101000001",
  17650=>"100000001",
  17651=>"100011100",
  17652=>"010100111",
  17653=>"010010101",
  17654=>"010000100",
  17655=>"000010001",
  17656=>"000100000",
  17657=>"000111011",
  17658=>"101111010",
  17659=>"000101000",
  17660=>"100111000",
  17661=>"111000000",
  17662=>"101101001",
  17663=>"000011111",
  17664=>"010111010",
  17665=>"100111110",
  17666=>"100100000",
  17667=>"111000010",
  17668=>"100000010",
  17669=>"000000000",
  17670=>"111001001",
  17671=>"101100100",
  17672=>"011001000",
  17673=>"111011111",
  17674=>"100111011",
  17675=>"000010100",
  17676=>"100110011",
  17677=>"111001111",
  17678=>"010100110",
  17679=>"001001110",
  17680=>"100110000",
  17681=>"010111010",
  17682=>"111111110",
  17683=>"110100000",
  17684=>"011111110",
  17685=>"100010111",
  17686=>"011110111",
  17687=>"101110000",
  17688=>"101000100",
  17689=>"100010000",
  17690=>"000000010",
  17691=>"001010000",
  17692=>"001011100",
  17693=>"110000011",
  17694=>"000110110",
  17695=>"110101111",
  17696=>"001001101",
  17697=>"111100111",
  17698=>"010010000",
  17699=>"100100111",
  17700=>"010011101",
  17701=>"011110000",
  17702=>"100001001",
  17703=>"011010011",
  17704=>"111111001",
  17705=>"011000101",
  17706=>"001000100",
  17707=>"101001000",
  17708=>"111110001",
  17709=>"111110000",
  17710=>"110101110",
  17711=>"000111000",
  17712=>"101001111",
  17713=>"010000101",
  17714=>"001100100",
  17715=>"110000010",
  17716=>"011111000",
  17717=>"010101010",
  17718=>"001000011",
  17719=>"111100101",
  17720=>"000001001",
  17721=>"011111101",
  17722=>"111101001",
  17723=>"001000011",
  17724=>"001000110",
  17725=>"001000011",
  17726=>"011000000",
  17727=>"111011011",
  17728=>"111101111",
  17729=>"011111111",
  17730=>"111111010",
  17731=>"010010100",
  17732=>"101001011",
  17733=>"111110000",
  17734=>"110100101",
  17735=>"010100111",
  17736=>"011110101",
  17737=>"000010110",
  17738=>"100110001",
  17739=>"111110111",
  17740=>"110110000",
  17741=>"000111100",
  17742=>"110000111",
  17743=>"011110110",
  17744=>"011010100",
  17745=>"000000111",
  17746=>"000000001",
  17747=>"111000010",
  17748=>"001111010",
  17749=>"001100010",
  17750=>"000000101",
  17751=>"000001010",
  17752=>"010000011",
  17753=>"010111101",
  17754=>"011111100",
  17755=>"000000010",
  17756=>"000101011",
  17757=>"010001111",
  17758=>"111000001",
  17759=>"111001000",
  17760=>"000011010",
  17761=>"111101101",
  17762=>"000000010",
  17763=>"001001001",
  17764=>"011010000",
  17765=>"111001110",
  17766=>"010110011",
  17767=>"000111010",
  17768=>"000010011",
  17769=>"000011101",
  17770=>"100000001",
  17771=>"001011101",
  17772=>"010011100",
  17773=>"100001001",
  17774=>"110111010",
  17775=>"011100000",
  17776=>"000110011",
  17777=>"101110101",
  17778=>"101110111",
  17779=>"000000100",
  17780=>"000100101",
  17781=>"010000100",
  17782=>"001101000",
  17783=>"000101100",
  17784=>"100100101",
  17785=>"000000000",
  17786=>"001001100",
  17787=>"110100001",
  17788=>"010111001",
  17789=>"000111100",
  17790=>"111100101",
  17791=>"001001000",
  17792=>"101110001",
  17793=>"110100010",
  17794=>"111101001",
  17795=>"001101000",
  17796=>"001111111",
  17797=>"001111111",
  17798=>"011010101",
  17799=>"111001011",
  17800=>"101100110",
  17801=>"010100100",
  17802=>"101010101",
  17803=>"100101110",
  17804=>"101100000",
  17805=>"111001001",
  17806=>"010111011",
  17807=>"000011110",
  17808=>"010110011",
  17809=>"011101101",
  17810=>"101111100",
  17811=>"100100101",
  17812=>"100101100",
  17813=>"101011100",
  17814=>"000111101",
  17815=>"111010100",
  17816=>"101110100",
  17817=>"000110011",
  17818=>"001001111",
  17819=>"110000000",
  17820=>"010101111",
  17821=>"011001000",
  17822=>"101001111",
  17823=>"100000001",
  17824=>"000110111",
  17825=>"010010101",
  17826=>"110110110",
  17827=>"010101000",
  17828=>"100010011",
  17829=>"000001111",
  17830=>"000000100",
  17831=>"100001000",
  17832=>"010000000",
  17833=>"111000101",
  17834=>"101001000",
  17835=>"010100011",
  17836=>"001110001",
  17837=>"111010111",
  17838=>"110110001",
  17839=>"001011111",
  17840=>"001101110",
  17841=>"101100011",
  17842=>"110001101",
  17843=>"100101100",
  17844=>"001000011",
  17845=>"000010010",
  17846=>"011111011",
  17847=>"100011111",
  17848=>"001001100",
  17849=>"011001100",
  17850=>"110000000",
  17851=>"101111010",
  17852=>"101100110",
  17853=>"111010001",
  17854=>"010011101",
  17855=>"111100001",
  17856=>"011010110",
  17857=>"110100111",
  17858=>"000100111",
  17859=>"011011110",
  17860=>"001001110",
  17861=>"101011111",
  17862=>"011100100",
  17863=>"101100000",
  17864=>"111101111",
  17865=>"101100111",
  17866=>"001011011",
  17867=>"000111000",
  17868=>"011110111",
  17869=>"000110100",
  17870=>"001101100",
  17871=>"000100100",
  17872=>"100001110",
  17873=>"100101001",
  17874=>"000000111",
  17875=>"010000110",
  17876=>"000001100",
  17877=>"011010000",
  17878=>"100001110",
  17879=>"111110101",
  17880=>"011000000",
  17881=>"111111110",
  17882=>"111110111",
  17883=>"000110110",
  17884=>"101111111",
  17885=>"001000010",
  17886=>"011010100",
  17887=>"110110111",
  17888=>"010011001",
  17889=>"001100100",
  17890=>"011100101",
  17891=>"110000100",
  17892=>"100100110",
  17893=>"000011100",
  17894=>"010110000",
  17895=>"001000110",
  17896=>"001100110",
  17897=>"000110011",
  17898=>"000110100",
  17899=>"100111100",
  17900=>"011011100",
  17901=>"100110101",
  17902=>"010000100",
  17903=>"000000011",
  17904=>"101000011",
  17905=>"010011000",
  17906=>"011010101",
  17907=>"101100111",
  17908=>"001011001",
  17909=>"011000000",
  17910=>"110111010",
  17911=>"001110011",
  17912=>"010110010",
  17913=>"111110011",
  17914=>"011101010",
  17915=>"001001001",
  17916=>"010111011",
  17917=>"110010100",
  17918=>"100100001",
  17919=>"010000011",
  17920=>"000111101",
  17921=>"011011110",
  17922=>"001011011",
  17923=>"011011011",
  17924=>"001111111",
  17925=>"001001001",
  17926=>"110000001",
  17927=>"000001000",
  17928=>"011010001",
  17929=>"000111101",
  17930=>"100101010",
  17931=>"101010110",
  17932=>"000100011",
  17933=>"101100010",
  17934=>"000001100",
  17935=>"000010000",
  17936=>"011000000",
  17937=>"011111010",
  17938=>"111010011",
  17939=>"111010011",
  17940=>"110111110",
  17941=>"011110001",
  17942=>"011001111",
  17943=>"001010110",
  17944=>"000101100",
  17945=>"001000111",
  17946=>"101101001",
  17947=>"100011000",
  17948=>"001001010",
  17949=>"001000100",
  17950=>"110110111",
  17951=>"000100011",
  17952=>"111100101",
  17953=>"101010001",
  17954=>"111101011",
  17955=>"000000101",
  17956=>"101001001",
  17957=>"101110010",
  17958=>"111101001",
  17959=>"001000010",
  17960=>"001110000",
  17961=>"001000001",
  17962=>"011100100",
  17963=>"011111111",
  17964=>"001001110",
  17965=>"000001011",
  17966=>"011010011",
  17967=>"000101111",
  17968=>"111101101",
  17969=>"101110000",
  17970=>"011000101",
  17971=>"111111111",
  17972=>"111010100",
  17973=>"110111011",
  17974=>"101011110",
  17975=>"011100101",
  17976=>"101100100",
  17977=>"110100110",
  17978=>"111011111",
  17979=>"101011010",
  17980=>"011111111",
  17981=>"000010000",
  17982=>"000000010",
  17983=>"111000010",
  17984=>"010010100",
  17985=>"000001000",
  17986=>"111100000",
  17987=>"100000011",
  17988=>"000101111",
  17989=>"110101011",
  17990=>"100010111",
  17991=>"101010100",
  17992=>"111010000",
  17993=>"100100101",
  17994=>"011101110",
  17995=>"110001001",
  17996=>"010111111",
  17997=>"111000011",
  17998=>"111011011",
  17999=>"000101010",
  18000=>"000100000",
  18001=>"110001011",
  18002=>"101101101",
  18003=>"000100000",
  18004=>"001000011",
  18005=>"011110001",
  18006=>"111100001",
  18007=>"001100110",
  18008=>"111111000",
  18009=>"011100110",
  18010=>"110101010",
  18011=>"101101100",
  18012=>"000101101",
  18013=>"001101010",
  18014=>"000010010",
  18015=>"011100111",
  18016=>"011011110",
  18017=>"101100010",
  18018=>"101010111",
  18019=>"101000010",
  18020=>"000010010",
  18021=>"111100111",
  18022=>"000101011",
  18023=>"100000011",
  18024=>"101010111",
  18025=>"100001000",
  18026=>"010110010",
  18027=>"001111111",
  18028=>"101110100",
  18029=>"110000001",
  18030=>"101001100",
  18031=>"000101101",
  18032=>"101011100",
  18033=>"000100101",
  18034=>"001011101",
  18035=>"001001101",
  18036=>"111010011",
  18037=>"100110000",
  18038=>"110100100",
  18039=>"100100001",
  18040=>"111110000",
  18041=>"100100001",
  18042=>"100111101",
  18043=>"010011100",
  18044=>"111010001",
  18045=>"101110111",
  18046=>"110110110",
  18047=>"110010111",
  18048=>"101011001",
  18049=>"001110001",
  18050=>"001101100",
  18051=>"001001001",
  18052=>"110001101",
  18053=>"010001111",
  18054=>"010011011",
  18055=>"100111000",
  18056=>"001101001",
  18057=>"001010011",
  18058=>"111110010",
  18059=>"110101100",
  18060=>"001100000",
  18061=>"110111000",
  18062=>"100100100",
  18063=>"010111010",
  18064=>"100001011",
  18065=>"000111111",
  18066=>"101010000",
  18067=>"001110010",
  18068=>"000000101",
  18069=>"010101010",
  18070=>"100110111",
  18071=>"101001110",
  18072=>"011110011",
  18073=>"011110100",
  18074=>"101110000",
  18075=>"111101010",
  18076=>"001101010",
  18077=>"111101101",
  18078=>"100111110",
  18079=>"010010011",
  18080=>"100000110",
  18081=>"000001001",
  18082=>"010100110",
  18083=>"011100010",
  18084=>"010101101",
  18085=>"011010100",
  18086=>"100101110",
  18087=>"100011011",
  18088=>"110000000",
  18089=>"111101101",
  18090=>"010110101",
  18091=>"000000101",
  18092=>"100101111",
  18093=>"100010001",
  18094=>"110111100",
  18095=>"010111011",
  18096=>"101111101",
  18097=>"111111100",
  18098=>"010100101",
  18099=>"001111111",
  18100=>"001101110",
  18101=>"000110100",
  18102=>"110101101",
  18103=>"110100101",
  18104=>"010001011",
  18105=>"101101011",
  18106=>"100001111",
  18107=>"000101111",
  18108=>"100011000",
  18109=>"010000010",
  18110=>"000110101",
  18111=>"100110111",
  18112=>"110010010",
  18113=>"001110111",
  18114=>"001111000",
  18115=>"100100001",
  18116=>"001101001",
  18117=>"010111111",
  18118=>"111000000",
  18119=>"000001010",
  18120=>"000110101",
  18121=>"001110111",
  18122=>"101000111",
  18123=>"011010111",
  18124=>"100100001",
  18125=>"000011100",
  18126=>"011010000",
  18127=>"000100001",
  18128=>"111010101",
  18129=>"010001001",
  18130=>"110110111",
  18131=>"001100100",
  18132=>"110110100",
  18133=>"100010011",
  18134=>"101110101",
  18135=>"101111010",
  18136=>"111101100",
  18137=>"011110001",
  18138=>"010110000",
  18139=>"110010001",
  18140=>"000000000",
  18141=>"011001011",
  18142=>"110111110",
  18143=>"001010001",
  18144=>"001001011",
  18145=>"110000100",
  18146=>"100010101",
  18147=>"011110001",
  18148=>"010010001",
  18149=>"001110100",
  18150=>"010110101",
  18151=>"011100000",
  18152=>"011101111",
  18153=>"111001110",
  18154=>"111110010",
  18155=>"011101111",
  18156=>"001000100",
  18157=>"010110001",
  18158=>"011101101",
  18159=>"100011111",
  18160=>"000110001",
  18161=>"010000001",
  18162=>"101111000",
  18163=>"101010001",
  18164=>"101110111",
  18165=>"101000111",
  18166=>"101111100",
  18167=>"100100010",
  18168=>"000100101",
  18169=>"101111010",
  18170=>"000010110",
  18171=>"010000100",
  18172=>"011111000",
  18173=>"001111011",
  18174=>"011111101",
  18175=>"000000011",
  18176=>"111000011",
  18177=>"100101101",
  18178=>"011111000",
  18179=>"001100101",
  18180=>"001101000",
  18181=>"010111110",
  18182=>"011111011",
  18183=>"100011111",
  18184=>"010011001",
  18185=>"110110000",
  18186=>"001011100",
  18187=>"111100111",
  18188=>"100000101",
  18189=>"101010110",
  18190=>"100101000",
  18191=>"111101010",
  18192=>"000101101",
  18193=>"100111110",
  18194=>"100001100",
  18195=>"110000101",
  18196=>"110010100",
  18197=>"101100000",
  18198=>"000001001",
  18199=>"101111100",
  18200=>"111111111",
  18201=>"000000001",
  18202=>"000000001",
  18203=>"110110011",
  18204=>"100101010",
  18205=>"000001010",
  18206=>"011000000",
  18207=>"111010100",
  18208=>"011100001",
  18209=>"001000011",
  18210=>"100011000",
  18211=>"011110110",
  18212=>"110101010",
  18213=>"010001001",
  18214=>"111000111",
  18215=>"000100011",
  18216=>"000110011",
  18217=>"110101001",
  18218=>"111010101",
  18219=>"010110001",
  18220=>"111010101",
  18221=>"000110000",
  18222=>"111110011",
  18223=>"111101110",
  18224=>"001000111",
  18225=>"001011101",
  18226=>"101100110",
  18227=>"101000100",
  18228=>"010110101",
  18229=>"010001110",
  18230=>"111110101",
  18231=>"001100110",
  18232=>"000001001",
  18233=>"010110111",
  18234=>"001111001",
  18235=>"111010010",
  18236=>"101111111",
  18237=>"110101110",
  18238=>"000100000",
  18239=>"110000100",
  18240=>"001001110",
  18241=>"101000100",
  18242=>"111110001",
  18243=>"010000010",
  18244=>"000000000",
  18245=>"011110011",
  18246=>"111101110",
  18247=>"001010001",
  18248=>"001111001",
  18249=>"111110001",
  18250=>"000001110",
  18251=>"010001000",
  18252=>"101001100",
  18253=>"000000111",
  18254=>"110110001",
  18255=>"001110100",
  18256=>"111010111",
  18257=>"101010111",
  18258=>"100010000",
  18259=>"100010110",
  18260=>"011001101",
  18261=>"001000111",
  18262=>"000001001",
  18263=>"000111111",
  18264=>"110101101",
  18265=>"100101011",
  18266=>"011100011",
  18267=>"101110110",
  18268=>"101001110",
  18269=>"110011010",
  18270=>"011110010",
  18271=>"100010000",
  18272=>"000010010",
  18273=>"110111011",
  18274=>"101100000",
  18275=>"111011000",
  18276=>"111010000",
  18277=>"010111001",
  18278=>"111000110",
  18279=>"000001101",
  18280=>"000101000",
  18281=>"101101100",
  18282=>"011010100",
  18283=>"110001100",
  18284=>"000111111",
  18285=>"101111010",
  18286=>"111101011",
  18287=>"011000101",
  18288=>"000111100",
  18289=>"010101001",
  18290=>"110100111",
  18291=>"001001100",
  18292=>"111000010",
  18293=>"000001100",
  18294=>"110111111",
  18295=>"011110111",
  18296=>"101010100",
  18297=>"011000001",
  18298=>"111111010",
  18299=>"101101001",
  18300=>"001110011",
  18301=>"101110000",
  18302=>"111001101",
  18303=>"000010100",
  18304=>"100110010",
  18305=>"001000011",
  18306=>"010011010",
  18307=>"111101110",
  18308=>"011000011",
  18309=>"011000000",
  18310=>"110001111",
  18311=>"000000101",
  18312=>"001010100",
  18313=>"011010010",
  18314=>"110111110",
  18315=>"011101101",
  18316=>"101100011",
  18317=>"010011111",
  18318=>"111111000",
  18319=>"011111000",
  18320=>"111110010",
  18321=>"011100000",
  18322=>"101011010",
  18323=>"101100001",
  18324=>"101111101",
  18325=>"010011011",
  18326=>"110011110",
  18327=>"101111011",
  18328=>"001000010",
  18329=>"011111001",
  18330=>"111010110",
  18331=>"001101111",
  18332=>"101000010",
  18333=>"010110110",
  18334=>"100111110",
  18335=>"101001101",
  18336=>"000000001",
  18337=>"101100000",
  18338=>"111100110",
  18339=>"110111000",
  18340=>"111101111",
  18341=>"011010010",
  18342=>"110001011",
  18343=>"110111001",
  18344=>"101111110",
  18345=>"101000000",
  18346=>"010110111",
  18347=>"111011111",
  18348=>"010010001",
  18349=>"101000000",
  18350=>"001011100",
  18351=>"101001111",
  18352=>"001011111",
  18353=>"000110010",
  18354=>"100000011",
  18355=>"001001001",
  18356=>"011001010",
  18357=>"111010001",
  18358=>"110010101",
  18359=>"101011101",
  18360=>"111111111",
  18361=>"111011010",
  18362=>"111111111",
  18363=>"001000111",
  18364=>"011101000",
  18365=>"111001101",
  18366=>"111111110",
  18367=>"011011111",
  18368=>"001001100",
  18369=>"111000100",
  18370=>"010011011",
  18371=>"000001000",
  18372=>"001000110",
  18373=>"001011000",
  18374=>"111110100",
  18375=>"111110101",
  18376=>"011111101",
  18377=>"100000110",
  18378=>"010101110",
  18379=>"001100000",
  18380=>"011111010",
  18381=>"110001111",
  18382=>"111111000",
  18383=>"110000110",
  18384=>"110111110",
  18385=>"000100111",
  18386=>"000100000",
  18387=>"000111101",
  18388=>"000001001",
  18389=>"101110010",
  18390=>"011001110",
  18391=>"011001010",
  18392=>"011011101",
  18393=>"011111011",
  18394=>"000110111",
  18395=>"000100001",
  18396=>"101001111",
  18397=>"010101100",
  18398=>"011001110",
  18399=>"010000001",
  18400=>"000000100",
  18401=>"110100110",
  18402=>"001100101",
  18403=>"110100011",
  18404=>"101111011",
  18405=>"000011010",
  18406=>"111111110",
  18407=>"101101000",
  18408=>"100010101",
  18409=>"000111001",
  18410=>"111011100",
  18411=>"111001111",
  18412=>"001100011",
  18413=>"110110010",
  18414=>"111000100",
  18415=>"000010010",
  18416=>"011011001",
  18417=>"111010111",
  18418=>"100000101",
  18419=>"010000001",
  18420=>"100001100",
  18421=>"011111111",
  18422=>"111111001",
  18423=>"001011011",
  18424=>"111110101",
  18425=>"011011011",
  18426=>"011101001",
  18427=>"000001000",
  18428=>"111111100",
  18429=>"000000100",
  18430=>"111101000",
  18431=>"010011001",
  18432=>"100011010",
  18433=>"111110010",
  18434=>"011010001",
  18435=>"000001010",
  18436=>"100000111",
  18437=>"100011011",
  18438=>"001000100",
  18439=>"100000000",
  18440=>"010011010",
  18441=>"000110110",
  18442=>"101000001",
  18443=>"111001100",
  18444=>"010101101",
  18445=>"111011000",
  18446=>"111000101",
  18447=>"010000110",
  18448=>"000011100",
  18449=>"000101010",
  18450=>"110100100",
  18451=>"111100001",
  18452=>"110000101",
  18453=>"111010100",
  18454=>"110010101",
  18455=>"001101110",
  18456=>"011000001",
  18457=>"101110110",
  18458=>"111011010",
  18459=>"011010111",
  18460=>"111101100",
  18461=>"110111011",
  18462=>"000000000",
  18463=>"001000111",
  18464=>"000101110",
  18465=>"100111111",
  18466=>"110101110",
  18467=>"010000000",
  18468=>"110001010",
  18469=>"001101010",
  18470=>"010010000",
  18471=>"101101001",
  18472=>"011010010",
  18473=>"100001001",
  18474=>"011000100",
  18475=>"011011110",
  18476=>"000100101",
  18477=>"110101100",
  18478=>"110011111",
  18479=>"010111001",
  18480=>"011100001",
  18481=>"100101001",
  18482=>"011101000",
  18483=>"101000011",
  18484=>"001000001",
  18485=>"010010110",
  18486=>"010000011",
  18487=>"010001010",
  18488=>"100101101",
  18489=>"100011100",
  18490=>"101111101",
  18491=>"111101000",
  18492=>"011111010",
  18493=>"001010010",
  18494=>"100100011",
  18495=>"001111011",
  18496=>"010111111",
  18497=>"000010111",
  18498=>"001111110",
  18499=>"001001000",
  18500=>"110110000",
  18501=>"110110011",
  18502=>"101011010",
  18503=>"100100011",
  18504=>"101101111",
  18505=>"010011100",
  18506=>"100011011",
  18507=>"000011111",
  18508=>"101000000",
  18509=>"000000100",
  18510=>"010000111",
  18511=>"101110011",
  18512=>"100111101",
  18513=>"010000100",
  18514=>"100001010",
  18515=>"100010111",
  18516=>"111101100",
  18517=>"101000010",
  18518=>"000111001",
  18519=>"000111100",
  18520=>"101100100",
  18521=>"011001111",
  18522=>"001101100",
  18523=>"111101101",
  18524=>"010100000",
  18525=>"001100010",
  18526=>"000110001",
  18527=>"010101000",
  18528=>"001000001",
  18529=>"000101010",
  18530=>"101000001",
  18531=>"001010010",
  18532=>"000101001",
  18533=>"001010001",
  18534=>"100001000",
  18535=>"000100000",
  18536=>"110101111",
  18537=>"011110101",
  18538=>"000100011",
  18539=>"100101011",
  18540=>"010110000",
  18541=>"110001001",
  18542=>"101101100",
  18543=>"001011110",
  18544=>"000111100",
  18545=>"010010011",
  18546=>"110100111",
  18547=>"110011100",
  18548=>"001000011",
  18549=>"111111111",
  18550=>"010101001",
  18551=>"100000011",
  18552=>"000100111",
  18553=>"111110110",
  18554=>"111011000",
  18555=>"101000101",
  18556=>"010011101",
  18557=>"100001111",
  18558=>"101111100",
  18559=>"101000100",
  18560=>"101011010",
  18561=>"010101111",
  18562=>"111110100",
  18563=>"011111010",
  18564=>"100001110",
  18565=>"000001110",
  18566=>"000110001",
  18567=>"101001110",
  18568=>"101101110",
  18569=>"000110011",
  18570=>"000001011",
  18571=>"000011001",
  18572=>"101010011",
  18573=>"101101110",
  18574=>"000001100",
  18575=>"111001111",
  18576=>"100100000",
  18577=>"000000100",
  18578=>"111100000",
  18579=>"001010110",
  18580=>"101111110",
  18581=>"110100010",
  18582=>"000111011",
  18583=>"001101010",
  18584=>"100111010",
  18585=>"001100000",
  18586=>"100010100",
  18587=>"111001101",
  18588=>"000010111",
  18589=>"111000001",
  18590=>"001100000",
  18591=>"111000101",
  18592=>"111000000",
  18593=>"001011010",
  18594=>"000100001",
  18595=>"011000101",
  18596=>"110101100",
  18597=>"101111000",
  18598=>"101110011",
  18599=>"100100100",
  18600=>"111100100",
  18601=>"011100011",
  18602=>"101000010",
  18603=>"110111010",
  18604=>"001110100",
  18605=>"111100000",
  18606=>"011000100",
  18607=>"111100001",
  18608=>"110100000",
  18609=>"011100110",
  18610=>"100011110",
  18611=>"100111000",
  18612=>"101111001",
  18613=>"101101001",
  18614=>"010010010",
  18615=>"011111100",
  18616=>"011000100",
  18617=>"010010000",
  18618=>"101001101",
  18619=>"111111110",
  18620=>"110001001",
  18621=>"111100111",
  18622=>"001110100",
  18623=>"100101111",
  18624=>"100111110",
  18625=>"111010011",
  18626=>"000001010",
  18627=>"010011000",
  18628=>"010011001",
  18629=>"000010100",
  18630=>"001011110",
  18631=>"110010001",
  18632=>"011100001",
  18633=>"010000001",
  18634=>"001011101",
  18635=>"101101101",
  18636=>"100111010",
  18637=>"000011111",
  18638=>"001000101",
  18639=>"111001000",
  18640=>"000011110",
  18641=>"111000000",
  18642=>"000010101",
  18643=>"101110110",
  18644=>"010000010",
  18645=>"011100110",
  18646=>"100111000",
  18647=>"100001111",
  18648=>"100000001",
  18649=>"010010100",
  18650=>"010000001",
  18651=>"111101110",
  18652=>"011110100",
  18653=>"001000000",
  18654=>"100101010",
  18655=>"000110000",
  18656=>"100011110",
  18657=>"111111001",
  18658=>"001000011",
  18659=>"000000100",
  18660=>"110001100",
  18661=>"100111001",
  18662=>"101000100",
  18663=>"001100101",
  18664=>"010111011",
  18665=>"111101011",
  18666=>"100011101",
  18667=>"011111000",
  18668=>"101010101",
  18669=>"000011111",
  18670=>"001111010",
  18671=>"110110110",
  18672=>"111101101",
  18673=>"110000111",
  18674=>"100110110",
  18675=>"100111001",
  18676=>"000100100",
  18677=>"100110001",
  18678=>"100110110",
  18679=>"001000100",
  18680=>"100000010",
  18681=>"101011101",
  18682=>"001001010",
  18683=>"000000110",
  18684=>"010000110",
  18685=>"100000100",
  18686=>"110111011",
  18687=>"110110011",
  18688=>"110100010",
  18689=>"111100100",
  18690=>"111000001",
  18691=>"101110010",
  18692=>"010111000",
  18693=>"101110100",
  18694=>"000010110",
  18695=>"111011100",
  18696=>"000111011",
  18697=>"110101100",
  18698=>"011011101",
  18699=>"001001001",
  18700=>"110110100",
  18701=>"010110001",
  18702=>"001110101",
  18703=>"000000011",
  18704=>"011001111",
  18705=>"101001010",
  18706=>"100011110",
  18707=>"100111100",
  18708=>"111000110",
  18709=>"110000110",
  18710=>"100000001",
  18711=>"011101010",
  18712=>"110101110",
  18713=>"011100100",
  18714=>"110110101",
  18715=>"110111001",
  18716=>"001010000",
  18717=>"001111111",
  18718=>"110001101",
  18719=>"000001100",
  18720=>"111101001",
  18721=>"111100110",
  18722=>"000011011",
  18723=>"010101010",
  18724=>"110010100",
  18725=>"000111010",
  18726=>"100101111",
  18727=>"110100011",
  18728=>"010111010",
  18729=>"000100111",
  18730=>"010001000",
  18731=>"011001011",
  18732=>"101101110",
  18733=>"101000010",
  18734=>"011011000",
  18735=>"010111101",
  18736=>"100111101",
  18737=>"000000001",
  18738=>"111011111",
  18739=>"010000000",
  18740=>"001001101",
  18741=>"000010000",
  18742=>"011101100",
  18743=>"011011110",
  18744=>"000010100",
  18745=>"001000101",
  18746=>"010011100",
  18747=>"010101110",
  18748=>"000011000",
  18749=>"110100100",
  18750=>"100110001",
  18751=>"110011111",
  18752=>"111111001",
  18753=>"001110111",
  18754=>"111010100",
  18755=>"010101101",
  18756=>"100110101",
  18757=>"010110000",
  18758=>"000010001",
  18759=>"001000001",
  18760=>"101101001",
  18761=>"100100001",
  18762=>"010101100",
  18763=>"011111100",
  18764=>"000001000",
  18765=>"001000100",
  18766=>"110010111",
  18767=>"011100111",
  18768=>"111001100",
  18769=>"110000010",
  18770=>"100011001",
  18771=>"000010001",
  18772=>"001000001",
  18773=>"010100110",
  18774=>"000010100",
  18775=>"000011011",
  18776=>"000011010",
  18777=>"100110011",
  18778=>"110011101",
  18779=>"001011011",
  18780=>"001001000",
  18781=>"100100101",
  18782=>"110001011",
  18783=>"000111000",
  18784=>"010001110",
  18785=>"010000000",
  18786=>"001001100",
  18787=>"100011000",
  18788=>"001000101",
  18789=>"111010100",
  18790=>"101110110",
  18791=>"100111101",
  18792=>"011100101",
  18793=>"001111001",
  18794=>"101111111",
  18795=>"001101100",
  18796=>"101100011",
  18797=>"000011100",
  18798=>"001110111",
  18799=>"111011000",
  18800=>"000010000",
  18801=>"110001010",
  18802=>"011111010",
  18803=>"100100110",
  18804=>"000011110",
  18805=>"111001100",
  18806=>"010100011",
  18807=>"010000000",
  18808=>"110000100",
  18809=>"000110101",
  18810=>"000000010",
  18811=>"101100100",
  18812=>"111001110",
  18813=>"110001100",
  18814=>"000100111",
  18815=>"111011110",
  18816=>"111011101",
  18817=>"001000000",
  18818=>"010111101",
  18819=>"010100011",
  18820=>"001000110",
  18821=>"011110110",
  18822=>"100010101",
  18823=>"010000001",
  18824=>"001000111",
  18825=>"010110110",
  18826=>"010110100",
  18827=>"001101100",
  18828=>"000110100",
  18829=>"000000110",
  18830=>"100000100",
  18831=>"111000111",
  18832=>"110010110",
  18833=>"100100001",
  18834=>"011111010",
  18835=>"011000110",
  18836=>"101010010",
  18837=>"110000011",
  18838=>"011000101",
  18839=>"011001011",
  18840=>"011001111",
  18841=>"010110111",
  18842=>"110001010",
  18843=>"010001100",
  18844=>"101010110",
  18845=>"000000010",
  18846=>"011000000",
  18847=>"100110000",
  18848=>"001010110",
  18849=>"010100110",
  18850=>"001111111",
  18851=>"101010101",
  18852=>"011100100",
  18853=>"110010000",
  18854=>"100000000",
  18855=>"000010100",
  18856=>"001110110",
  18857=>"011000101",
  18858=>"001010111",
  18859=>"110010100",
  18860=>"000101010",
  18861=>"101000011",
  18862=>"001000100",
  18863=>"110100101",
  18864=>"111001110",
  18865=>"011110100",
  18866=>"110010111",
  18867=>"000010111",
  18868=>"110011011",
  18869=>"000001101",
  18870=>"111100100",
  18871=>"110101011",
  18872=>"010111000",
  18873=>"010110000",
  18874=>"110010110",
  18875=>"011010110",
  18876=>"101101010",
  18877=>"101000100",
  18878=>"111001100",
  18879=>"001110111",
  18880=>"010011111",
  18881=>"000100101",
  18882=>"000001100",
  18883=>"010100011",
  18884=>"110101110",
  18885=>"100011101",
  18886=>"010110111",
  18887=>"100011000",
  18888=>"001000110",
  18889=>"000010000",
  18890=>"001110100",
  18891=>"111111100",
  18892=>"001000101",
  18893=>"000010001",
  18894=>"001000100",
  18895=>"111101111",
  18896=>"111010011",
  18897=>"010010000",
  18898=>"110000101",
  18899=>"000100101",
  18900=>"011111011",
  18901=>"001101011",
  18902=>"100000101",
  18903=>"000001101",
  18904=>"100001000",
  18905=>"111111010",
  18906=>"111001101",
  18907=>"100000111",
  18908=>"111110101",
  18909=>"101000111",
  18910=>"110111100",
  18911=>"110010010",
  18912=>"001000000",
  18913=>"000111000",
  18914=>"100010101",
  18915=>"101111001",
  18916=>"101000001",
  18917=>"111101000",
  18918=>"001011101",
  18919=>"001010011",
  18920=>"000011110",
  18921=>"110001111",
  18922=>"000010000",
  18923=>"000010001",
  18924=>"001011110",
  18925=>"101011101",
  18926=>"101011001",
  18927=>"100010010",
  18928=>"111100100",
  18929=>"101001101",
  18930=>"111010001",
  18931=>"101100101",
  18932=>"010100000",
  18933=>"011111111",
  18934=>"110111000",
  18935=>"000011100",
  18936=>"101100011",
  18937=>"000000010",
  18938=>"001011000",
  18939=>"010100001",
  18940=>"000011111",
  18941=>"001011111",
  18942=>"001101100",
  18943=>"000011011",
  18944=>"011001100",
  18945=>"110000011",
  18946=>"001001010",
  18947=>"000100010",
  18948=>"000100110",
  18949=>"110000101",
  18950=>"110110011",
  18951=>"000011101",
  18952=>"110010000",
  18953=>"111111111",
  18954=>"010010100",
  18955=>"000110001",
  18956=>"111001110",
  18957=>"001110110",
  18958=>"111101000",
  18959=>"011000001",
  18960=>"000101110",
  18961=>"000100001",
  18962=>"000111000",
  18963=>"111100110",
  18964=>"000010010",
  18965=>"100101111",
  18966=>"110101110",
  18967=>"101010011",
  18968=>"001111000",
  18969=>"110000000",
  18970=>"000000101",
  18971=>"111011111",
  18972=>"111001000",
  18973=>"111001110",
  18974=>"001101011",
  18975=>"111010011",
  18976=>"111110010",
  18977=>"000000101",
  18978=>"000100011",
  18979=>"100010111",
  18980=>"011101100",
  18981=>"101101110",
  18982=>"110000110",
  18983=>"110011011",
  18984=>"010110000",
  18985=>"010010101",
  18986=>"100011111",
  18987=>"010011101",
  18988=>"001101010",
  18989=>"001101101",
  18990=>"100110001",
  18991=>"011010010",
  18992=>"110000011",
  18993=>"111101001",
  18994=>"001011101",
  18995=>"000110100",
  18996=>"000000110",
  18997=>"100011010",
  18998=>"110011101",
  18999=>"101101011",
  19000=>"001100011",
  19001=>"110000111",
  19002=>"000110011",
  19003=>"010001011",
  19004=>"000011100",
  19005=>"111001110",
  19006=>"000001100",
  19007=>"010110110",
  19008=>"100000110",
  19009=>"001101110",
  19010=>"110000011",
  19011=>"011010110",
  19012=>"101110111",
  19013=>"100110010",
  19014=>"000011000",
  19015=>"010001100",
  19016=>"011111001",
  19017=>"010101110",
  19018=>"110010000",
  19019=>"111010000",
  19020=>"111100111",
  19021=>"000101011",
  19022=>"101111000",
  19023=>"000010100",
  19024=>"011101111",
  19025=>"101011011",
  19026=>"111001101",
  19027=>"101100110",
  19028=>"111011110",
  19029=>"001111001",
  19030=>"000100010",
  19031=>"110001110",
  19032=>"111001001",
  19033=>"011010000",
  19034=>"110100011",
  19035=>"000111110",
  19036=>"000000011",
  19037=>"000001100",
  19038=>"100111011",
  19039=>"011000100",
  19040=>"111111101",
  19041=>"100000100",
  19042=>"000101010",
  19043=>"001000010",
  19044=>"110111101",
  19045=>"111110011",
  19046=>"101111100",
  19047=>"001001011",
  19048=>"000000010",
  19049=>"001110011",
  19050=>"001001100",
  19051=>"111000000",
  19052=>"000000001",
  19053=>"000010111",
  19054=>"110100110",
  19055=>"010001000",
  19056=>"010001110",
  19057=>"001110011",
  19058=>"001000110",
  19059=>"101101110",
  19060=>"111011110",
  19061=>"111010100",
  19062=>"000001001",
  19063=>"010011011",
  19064=>"110000100",
  19065=>"100001100",
  19066=>"110010101",
  19067=>"100001100",
  19068=>"100100010",
  19069=>"101110000",
  19070=>"111011110",
  19071=>"110101001",
  19072=>"101101101",
  19073=>"000011101",
  19074=>"100011110",
  19075=>"000001111",
  19076=>"111110101",
  19077=>"110000010",
  19078=>"011101111",
  19079=>"001100101",
  19080=>"111101110",
  19081=>"001001010",
  19082=>"011000011",
  19083=>"010000011",
  19084=>"110110111",
  19085=>"111110010",
  19086=>"111100000",
  19087=>"000101000",
  19088=>"000010101",
  19089=>"010100001",
  19090=>"001010101",
  19091=>"001111110",
  19092=>"010100011",
  19093=>"111010000",
  19094=>"011001101",
  19095=>"101001111",
  19096=>"101010000",
  19097=>"111111100",
  19098=>"000010110",
  19099=>"010100111",
  19100=>"110010010",
  19101=>"100101100",
  19102=>"000011000",
  19103=>"011011110",
  19104=>"010010110",
  19105=>"001001110",
  19106=>"110100111",
  19107=>"001001111",
  19108=>"100011100",
  19109=>"010001100",
  19110=>"001101100",
  19111=>"011000001",
  19112=>"000110001",
  19113=>"101000101",
  19114=>"101111100",
  19115=>"010010000",
  19116=>"011011010",
  19117=>"001001001",
  19118=>"101101000",
  19119=>"000111000",
  19120=>"001110001",
  19121=>"100000000",
  19122=>"010111101",
  19123=>"110110100",
  19124=>"010110101",
  19125=>"011010110",
  19126=>"110110101",
  19127=>"001000001",
  19128=>"110000011",
  19129=>"001001101",
  19130=>"110101001",
  19131=>"111101111",
  19132=>"110111001",
  19133=>"001001001",
  19134=>"000001010",
  19135=>"111110100",
  19136=>"101010010",
  19137=>"001000011",
  19138=>"010011100",
  19139=>"011000111",
  19140=>"100011111",
  19141=>"000101100",
  19142=>"101001111",
  19143=>"101101000",
  19144=>"000100000",
  19145=>"001001011",
  19146=>"000000101",
  19147=>"100011100",
  19148=>"000000011",
  19149=>"010101001",
  19150=>"100010001",
  19151=>"011000110",
  19152=>"111110110",
  19153=>"011000010",
  19154=>"100000000",
  19155=>"011000000",
  19156=>"010100101",
  19157=>"110101011",
  19158=>"111100001",
  19159=>"000000010",
  19160=>"000100101",
  19161=>"001111001",
  19162=>"000000000",
  19163=>"110101011",
  19164=>"000110111",
  19165=>"100010101",
  19166=>"110000011",
  19167=>"111100000",
  19168=>"010011101",
  19169=>"111110010",
  19170=>"001011111",
  19171=>"010000101",
  19172=>"011111010",
  19173=>"111101111",
  19174=>"101111110",
  19175=>"000110100",
  19176=>"110100100",
  19177=>"101110001",
  19178=>"011011111",
  19179=>"111000011",
  19180=>"001101101",
  19181=>"011111010",
  19182=>"111100110",
  19183=>"000001000",
  19184=>"001101000",
  19185=>"000111010",
  19186=>"011111100",
  19187=>"101100110",
  19188=>"000011111",
  19189=>"110101010",
  19190=>"011111110",
  19191=>"101100011",
  19192=>"000010100",
  19193=>"111101000",
  19194=>"111101100",
  19195=>"001010101",
  19196=>"101110101",
  19197=>"001100001",
  19198=>"001100011",
  19199=>"000000111",
  19200=>"110111001",
  19201=>"010000111",
  19202=>"000001011",
  19203=>"101000111",
  19204=>"000011010",
  19205=>"011000110",
  19206=>"000011111",
  19207=>"111110101",
  19208=>"101111101",
  19209=>"100001101",
  19210=>"011010100",
  19211=>"000010110",
  19212=>"100101001",
  19213=>"110011011",
  19214=>"110100001",
  19215=>"101111000",
  19216=>"000100010",
  19217=>"110111100",
  19218=>"110101010",
  19219=>"101100011",
  19220=>"011010110",
  19221=>"101100100",
  19222=>"010100000",
  19223=>"100110010",
  19224=>"011100110",
  19225=>"011100111",
  19226=>"001010001",
  19227=>"000010010",
  19228=>"011101010",
  19229=>"110110011",
  19230=>"100111000",
  19231=>"001101011",
  19232=>"110000110",
  19233=>"100000100",
  19234=>"010000010",
  19235=>"100101110",
  19236=>"100011101",
  19237=>"011001011",
  19238=>"001100001",
  19239=>"100010011",
  19240=>"100100010",
  19241=>"110000101",
  19242=>"101100111",
  19243=>"110101100",
  19244=>"111100011",
  19245=>"000001000",
  19246=>"011111000",
  19247=>"111111000",
  19248=>"000001100",
  19249=>"000110011",
  19250=>"101000010",
  19251=>"011100110",
  19252=>"111000000",
  19253=>"111011110",
  19254=>"101001001",
  19255=>"101010011",
  19256=>"100111110",
  19257=>"101101110",
  19258=>"001011100",
  19259=>"010000001",
  19260=>"000011000",
  19261=>"001101000",
  19262=>"011010001",
  19263=>"010010101",
  19264=>"100110001",
  19265=>"111110001",
  19266=>"100011000",
  19267=>"110001110",
  19268=>"000110101",
  19269=>"111100110",
  19270=>"100111010",
  19271=>"100100100",
  19272=>"111011011",
  19273=>"011000111",
  19274=>"000111010",
  19275=>"000110100",
  19276=>"101101111",
  19277=>"101101000",
  19278=>"100010100",
  19279=>"110101100",
  19280=>"101011110",
  19281=>"010101110",
  19282=>"010010111",
  19283=>"000010010",
  19284=>"110011010",
  19285=>"000011100",
  19286=>"101000110",
  19287=>"010011011",
  19288=>"100100000",
  19289=>"100010101",
  19290=>"001011010",
  19291=>"110010010",
  19292=>"001000110",
  19293=>"100101011",
  19294=>"111110100",
  19295=>"001011010",
  19296=>"100100011",
  19297=>"101010110",
  19298=>"010010001",
  19299=>"101010011",
  19300=>"101111011",
  19301=>"001000010",
  19302=>"000001011",
  19303=>"111010001",
  19304=>"100111011",
  19305=>"110110001",
  19306=>"000000001",
  19307=>"010101000",
  19308=>"101110000",
  19309=>"011110010",
  19310=>"011100111",
  19311=>"000101110",
  19312=>"001011100",
  19313=>"110010110",
  19314=>"110000110",
  19315=>"000100010",
  19316=>"011110110",
  19317=>"101000001",
  19318=>"110011100",
  19319=>"011000110",
  19320=>"001000001",
  19321=>"111011101",
  19322=>"111011111",
  19323=>"110111101",
  19324=>"000000000",
  19325=>"001010000",
  19326=>"110000111",
  19327=>"100100011",
  19328=>"001000100",
  19329=>"000101011",
  19330=>"010011011",
  19331=>"111010011",
  19332=>"110110101",
  19333=>"110010010",
  19334=>"011110110",
  19335=>"100100101",
  19336=>"010001000",
  19337=>"010011011",
  19338=>"100011101",
  19339=>"101111111",
  19340=>"110100011",
  19341=>"101110111",
  19342=>"001110101",
  19343=>"111011110",
  19344=>"111111101",
  19345=>"111010011",
  19346=>"001010000",
  19347=>"111100100",
  19348=>"110001101",
  19349=>"010101011",
  19350=>"011000000",
  19351=>"100111110",
  19352=>"111010111",
  19353=>"110011110",
  19354=>"001011100",
  19355=>"100101000",
  19356=>"001000001",
  19357=>"101011001",
  19358=>"000011001",
  19359=>"000100001",
  19360=>"101100110",
  19361=>"111011010",
  19362=>"111100101",
  19363=>"111010000",
  19364=>"010100001",
  19365=>"100100101",
  19366=>"011111000",
  19367=>"110111010",
  19368=>"010001001",
  19369=>"110111111",
  19370=>"011000000",
  19371=>"101100100",
  19372=>"010010011",
  19373=>"000101010",
  19374=>"010010111",
  19375=>"001100011",
  19376=>"011000010",
  19377=>"011001100",
  19378=>"110011000",
  19379=>"001011010",
  19380=>"001000011",
  19381=>"010001011",
  19382=>"110001010",
  19383=>"110011111",
  19384=>"011000001",
  19385=>"010010010",
  19386=>"110010110",
  19387=>"001011011",
  19388=>"100011000",
  19389=>"100000011",
  19390=>"101110010",
  19391=>"111110110",
  19392=>"110100011",
  19393=>"000011011",
  19394=>"010110000",
  19395=>"111101100",
  19396=>"010101000",
  19397=>"011101011",
  19398=>"000110100",
  19399=>"101000000",
  19400=>"101011111",
  19401=>"110100100",
  19402=>"001111001",
  19403=>"110001100",
  19404=>"000001010",
  19405=>"110111010",
  19406=>"110111010",
  19407=>"110011001",
  19408=>"000000010",
  19409=>"101001101",
  19410=>"100111001",
  19411=>"101010100",
  19412=>"010000111",
  19413=>"111101101",
  19414=>"101000000",
  19415=>"000011010",
  19416=>"000001110",
  19417=>"110011011",
  19418=>"010010111",
  19419=>"000111111",
  19420=>"111101000",
  19421=>"111111100",
  19422=>"110011101",
  19423=>"110110100",
  19424=>"001100110",
  19425=>"011101111",
  19426=>"000000001",
  19427=>"111100110",
  19428=>"000001110",
  19429=>"011000001",
  19430=>"111101101",
  19431=>"111011000",
  19432=>"001000010",
  19433=>"110001000",
  19434=>"100101111",
  19435=>"000111001",
  19436=>"000100000",
  19437=>"110111100",
  19438=>"011010000",
  19439=>"110111011",
  19440=>"000101111",
  19441=>"110101101",
  19442=>"011111101",
  19443=>"010010001",
  19444=>"100110111",
  19445=>"000001010",
  19446=>"111010111",
  19447=>"000100010",
  19448=>"111010011",
  19449=>"111110001",
  19450=>"011010000",
  19451=>"110101100",
  19452=>"100110001",
  19453=>"001001010",
  19454=>"001110011",
  19455=>"000001110",
  19456=>"100100111",
  19457=>"000100011",
  19458=>"110001111",
  19459=>"001101111",
  19460=>"101010010",
  19461=>"100110010",
  19462=>"111110100",
  19463=>"011011010",
  19464=>"100110000",
  19465=>"000000000",
  19466=>"001011000",
  19467=>"001100111",
  19468=>"001001011",
  19469=>"100011110",
  19470=>"011000111",
  19471=>"011001111",
  19472=>"111110110",
  19473=>"011111111",
  19474=>"110000001",
  19475=>"101111001",
  19476=>"010010000",
  19477=>"110010111",
  19478=>"001011001",
  19479=>"110000111",
  19480=>"110100000",
  19481=>"001011111",
  19482=>"110110100",
  19483=>"111010111",
  19484=>"010001001",
  19485=>"111111010",
  19486=>"010000011",
  19487=>"110010000",
  19488=>"101000100",
  19489=>"001110101",
  19490=>"011110001",
  19491=>"010110000",
  19492=>"000001000",
  19493=>"100001101",
  19494=>"001110000",
  19495=>"010100001",
  19496=>"111011100",
  19497=>"000001100",
  19498=>"001010101",
  19499=>"101101011",
  19500=>"001000000",
  19501=>"011101010",
  19502=>"001100110",
  19503=>"100111110",
  19504=>"101011000",
  19505=>"100110111",
  19506=>"110000101",
  19507=>"010001000",
  19508=>"100001000",
  19509=>"100011000",
  19510=>"110000100",
  19511=>"011111110",
  19512=>"101010000",
  19513=>"100000000",
  19514=>"001100101",
  19515=>"101111111",
  19516=>"111110011",
  19517=>"001111000",
  19518=>"101011101",
  19519=>"001111010",
  19520=>"010110110",
  19521=>"011101111",
  19522=>"110000010",
  19523=>"110000000",
  19524=>"111110011",
  19525=>"000101100",
  19526=>"011001100",
  19527=>"100100011",
  19528=>"101000010",
  19529=>"011010011",
  19530=>"000001111",
  19531=>"111101111",
  19532=>"010100111",
  19533=>"101110000",
  19534=>"000101111",
  19535=>"011111001",
  19536=>"010011000",
  19537=>"011101001",
  19538=>"111111000",
  19539=>"011001010",
  19540=>"101011011",
  19541=>"111111100",
  19542=>"001110010",
  19543=>"011011011",
  19544=>"100100100",
  19545=>"001110101",
  19546=>"011111101",
  19547=>"001100010",
  19548=>"011101110",
  19549=>"000111101",
  19550=>"010100111",
  19551=>"100001100",
  19552=>"010111100",
  19553=>"111001111",
  19554=>"101101000",
  19555=>"110000011",
  19556=>"110011001",
  19557=>"111010000",
  19558=>"100000011",
  19559=>"000000011",
  19560=>"100101111",
  19561=>"110011111",
  19562=>"100011101",
  19563=>"010101001",
  19564=>"101101100",
  19565=>"000000111",
  19566=>"000000001",
  19567=>"100100000",
  19568=>"010101000",
  19569=>"001011110",
  19570=>"100101110",
  19571=>"110001001",
  19572=>"000000111",
  19573=>"010101101",
  19574=>"110110100",
  19575=>"111111100",
  19576=>"100110001",
  19577=>"101011111",
  19578=>"000100010",
  19579=>"000100001",
  19580=>"000110001",
  19581=>"111011111",
  19582=>"101100101",
  19583=>"001001001",
  19584=>"011010110",
  19585=>"111100011",
  19586=>"011011001",
  19587=>"101100001",
  19588=>"101100101",
  19589=>"100001101",
  19590=>"001000110",
  19591=>"011000111",
  19592=>"001100011",
  19593=>"001011100",
  19594=>"110010001",
  19595=>"000001100",
  19596=>"011110000",
  19597=>"110100110",
  19598=>"000000111",
  19599=>"110111110",
  19600=>"100110001",
  19601=>"010001010",
  19602=>"101010010",
  19603=>"001100001",
  19604=>"000000110",
  19605=>"111001101",
  19606=>"011001110",
  19607=>"100111101",
  19608=>"010011110",
  19609=>"110111011",
  19610=>"011011111",
  19611=>"111111010",
  19612=>"000001011",
  19613=>"000000100",
  19614=>"111110011",
  19615=>"110011010",
  19616=>"000100010",
  19617=>"111101010",
  19618=>"010001111",
  19619=>"010111110",
  19620=>"010101010",
  19621=>"010001000",
  19622=>"000111001",
  19623=>"110010010",
  19624=>"101011000",
  19625=>"001111100",
  19626=>"001001101",
  19627=>"110111110",
  19628=>"110111000",
  19629=>"000011001",
  19630=>"011001101",
  19631=>"000011101",
  19632=>"110101010",
  19633=>"000011000",
  19634=>"000100000",
  19635=>"001111001",
  19636=>"110110010",
  19637=>"100010010",
  19638=>"110000111",
  19639=>"101000010",
  19640=>"010111111",
  19641=>"010000110",
  19642=>"110101111",
  19643=>"111010110",
  19644=>"000111000",
  19645=>"001100000",
  19646=>"110001101",
  19647=>"000001101",
  19648=>"100110111",
  19649=>"110001011",
  19650=>"101000111",
  19651=>"011110110",
  19652=>"011110111",
  19653=>"000110011",
  19654=>"100000010",
  19655=>"101111111",
  19656=>"010101010",
  19657=>"011011000",
  19658=>"000101101",
  19659=>"100101100",
  19660=>"101011010",
  19661=>"000011000",
  19662=>"000110111",
  19663=>"111111110",
  19664=>"110110101",
  19665=>"010111100",
  19666=>"001001100",
  19667=>"011001010",
  19668=>"110001100",
  19669=>"001110010",
  19670=>"011011001",
  19671=>"111001010",
  19672=>"011000111",
  19673=>"000101000",
  19674=>"101000001",
  19675=>"101000000",
  19676=>"001100010",
  19677=>"101010000",
  19678=>"110110010",
  19679=>"010100010",
  19680=>"010010101",
  19681=>"011111001",
  19682=>"011001000",
  19683=>"101011010",
  19684=>"111001110",
  19685=>"011111001",
  19686=>"000001100",
  19687=>"010111001",
  19688=>"000110110",
  19689=>"000111001",
  19690=>"110001011",
  19691=>"001001011",
  19692=>"100101000",
  19693=>"110100100",
  19694=>"110110010",
  19695=>"111101111",
  19696=>"000111101",
  19697=>"100001011",
  19698=>"000101011",
  19699=>"111001111",
  19700=>"010011111",
  19701=>"100010101",
  19702=>"111100001",
  19703=>"001100011",
  19704=>"101011100",
  19705=>"000111001",
  19706=>"010100101",
  19707=>"100111111",
  19708=>"001000001",
  19709=>"000010010",
  19710=>"100001011",
  19711=>"111001010",
  19712=>"010100011",
  19713=>"000111001",
  19714=>"111010010",
  19715=>"111010111",
  19716=>"111101011",
  19717=>"111011110",
  19718=>"101111110",
  19719=>"111111001",
  19720=>"000110000",
  19721=>"110000101",
  19722=>"010010011",
  19723=>"100101110",
  19724=>"100100101",
  19725=>"101100010",
  19726=>"000000011",
  19727=>"111011100",
  19728=>"110010101",
  19729=>"001110110",
  19730=>"000110010",
  19731=>"000010110",
  19732=>"011010111",
  19733=>"011011101",
  19734=>"000001111",
  19735=>"100000100",
  19736=>"001000001",
  19737=>"111110111",
  19738=>"000100000",
  19739=>"010011101",
  19740=>"000001110",
  19741=>"011110111",
  19742=>"011001000",
  19743=>"110011110",
  19744=>"111110110",
  19745=>"101011001",
  19746=>"100001110",
  19747=>"001111010",
  19748=>"101101110",
  19749=>"111110010",
  19750=>"101011010",
  19751=>"101111110",
  19752=>"101100110",
  19753=>"111011010",
  19754=>"010110010",
  19755=>"001010110",
  19756=>"000000000",
  19757=>"000101100",
  19758=>"001000010",
  19759=>"011100010",
  19760=>"010000111",
  19761=>"111110101",
  19762=>"001100010",
  19763=>"110100010",
  19764=>"001000001",
  19765=>"010100010",
  19766=>"100010001",
  19767=>"011000000",
  19768=>"000010110",
  19769=>"110110011",
  19770=>"100001111",
  19771=>"000011000",
  19772=>"110000011",
  19773=>"000111010",
  19774=>"111100101",
  19775=>"111011011",
  19776=>"011111010",
  19777=>"110110100",
  19778=>"100110111",
  19779=>"011110010",
  19780=>"010000101",
  19781=>"010010100",
  19782=>"000000100",
  19783=>"011111110",
  19784=>"110110011",
  19785=>"010100000",
  19786=>"001110000",
  19787=>"111010001",
  19788=>"101011011",
  19789=>"110001111",
  19790=>"111010101",
  19791=>"101111000",
  19792=>"010011010",
  19793=>"010101111",
  19794=>"110110000",
  19795=>"011111011",
  19796=>"000011111",
  19797=>"001010101",
  19798=>"110001011",
  19799=>"101000011",
  19800=>"000110111",
  19801=>"101110100",
  19802=>"101101001",
  19803=>"010110011",
  19804=>"000001100",
  19805=>"011101010",
  19806=>"100010101",
  19807=>"011001100",
  19808=>"000100001",
  19809=>"011001110",
  19810=>"110101011",
  19811=>"000001101",
  19812=>"100101000",
  19813=>"100011010",
  19814=>"111111100",
  19815=>"010011000",
  19816=>"000001011",
  19817=>"000000001",
  19818=>"100001011",
  19819=>"011110111",
  19820=>"000100011",
  19821=>"010110011",
  19822=>"000111101",
  19823=>"111001110",
  19824=>"100100110",
  19825=>"001100111",
  19826=>"001001111",
  19827=>"111111101",
  19828=>"101101111",
  19829=>"011110111",
  19830=>"011010110",
  19831=>"111000001",
  19832=>"100111101",
  19833=>"111100000",
  19834=>"101110011",
  19835=>"110110011",
  19836=>"001101111",
  19837=>"100010101",
  19838=>"001000000",
  19839=>"111011010",
  19840=>"101101101",
  19841=>"010010111",
  19842=>"000011000",
  19843=>"100101110",
  19844=>"010011011",
  19845=>"001011011",
  19846=>"100011111",
  19847=>"011000100",
  19848=>"110010010",
  19849=>"110010100",
  19850=>"110011100",
  19851=>"010001111",
  19852=>"010110010",
  19853=>"010101011",
  19854=>"001010001",
  19855=>"001101000",
  19856=>"001110111",
  19857=>"010011010",
  19858=>"100100111",
  19859=>"000001110",
  19860=>"110111111",
  19861=>"101010111",
  19862=>"000000001",
  19863=>"011111100",
  19864=>"100010000",
  19865=>"001000010",
  19866=>"000000110",
  19867=>"001110100",
  19868=>"100000101",
  19869=>"011011110",
  19870=>"111100011",
  19871=>"010111111",
  19872=>"001011110",
  19873=>"011000000",
  19874=>"110000111",
  19875=>"011100101",
  19876=>"101011110",
  19877=>"001111001",
  19878=>"010010110",
  19879=>"110100111",
  19880=>"000000100",
  19881=>"000011111",
  19882=>"001001000",
  19883=>"111111000",
  19884=>"100101110",
  19885=>"110101010",
  19886=>"111010100",
  19887=>"000111000",
  19888=>"100001010",
  19889=>"101001000",
  19890=>"101111000",
  19891=>"111100101",
  19892=>"101101101",
  19893=>"111110111",
  19894=>"010101001",
  19895=>"101011111",
  19896=>"001100110",
  19897=>"110111100",
  19898=>"010100000",
  19899=>"011100100",
  19900=>"000111110",
  19901=>"100101001",
  19902=>"000000000",
  19903=>"001001010",
  19904=>"110000001",
  19905=>"011000111",
  19906=>"111111000",
  19907=>"100001010",
  19908=>"101001011",
  19909=>"101010110",
  19910=>"100010011",
  19911=>"010001011",
  19912=>"101110011",
  19913=>"001001111",
  19914=>"010100001",
  19915=>"101101110",
  19916=>"011100011",
  19917=>"000100100",
  19918=>"011110110",
  19919=>"101011110",
  19920=>"001100010",
  19921=>"000100011",
  19922=>"110110010",
  19923=>"001001010",
  19924=>"001011101",
  19925=>"111100111",
  19926=>"101010010",
  19927=>"110010001",
  19928=>"110111100",
  19929=>"110011001",
  19930=>"001000100",
  19931=>"100100111",
  19932=>"100010000",
  19933=>"000001001",
  19934=>"100100111",
  19935=>"011111111",
  19936=>"110110101",
  19937=>"000110000",
  19938=>"100000011",
  19939=>"000010011",
  19940=>"000100100",
  19941=>"011101111",
  19942=>"100101101",
  19943=>"000011010",
  19944=>"011110000",
  19945=>"011111110",
  19946=>"010000001",
  19947=>"100100011",
  19948=>"011110011",
  19949=>"001001100",
  19950=>"100110010",
  19951=>"000100101",
  19952=>"011010000",
  19953=>"110110000",
  19954=>"001000001",
  19955=>"101000000",
  19956=>"000000111",
  19957=>"000000010",
  19958=>"111001011",
  19959=>"100010010",
  19960=>"110111101",
  19961=>"011000100",
  19962=>"111001110",
  19963=>"000101111",
  19964=>"001000010",
  19965=>"001011100",
  19966=>"000001101",
  19967=>"111111010",
  19968=>"101001001",
  19969=>"110010000",
  19970=>"100111011",
  19971=>"111111111",
  19972=>"011110110",
  19973=>"100000111",
  19974=>"011111011",
  19975=>"010000011",
  19976=>"011001011",
  19977=>"101010000",
  19978=>"101111111",
  19979=>"010000110",
  19980=>"110111010",
  19981=>"110111001",
  19982=>"111010111",
  19983=>"110000101",
  19984=>"110100101",
  19985=>"011001111",
  19986=>"000010101",
  19987=>"011001111",
  19988=>"111100100",
  19989=>"000111010",
  19990=>"110010011",
  19991=>"101000010",
  19992=>"001010011",
  19993=>"001111101",
  19994=>"011001011",
  19995=>"111110100",
  19996=>"010000010",
  19997=>"101000011",
  19998=>"010000100",
  19999=>"001100100",
  20000=>"010000011",
  20001=>"011101000",
  20002=>"000011000",
  20003=>"111010001",
  20004=>"100110010",
  20005=>"110100011",
  20006=>"100110100",
  20007=>"000101110",
  20008=>"111010011",
  20009=>"111111111",
  20010=>"101100000",
  20011=>"100000100",
  20012=>"001001111",
  20013=>"110001000",
  20014=>"001110011",
  20015=>"011000010",
  20016=>"110101000",
  20017=>"111110000",
  20018=>"101111000",
  20019=>"101101111",
  20020=>"111110001",
  20021=>"110101101",
  20022=>"100111110",
  20023=>"010001111",
  20024=>"100100011",
  20025=>"010100000",
  20026=>"011010011",
  20027=>"000001101",
  20028=>"111110100",
  20029=>"011011000",
  20030=>"101010100",
  20031=>"110011000",
  20032=>"001000111",
  20033=>"001110110",
  20034=>"110000111",
  20035=>"010110011",
  20036=>"001011110",
  20037=>"000001110",
  20038=>"101001000",
  20039=>"101010010",
  20040=>"110001111",
  20041=>"010111010",
  20042=>"010001011",
  20043=>"011101011",
  20044=>"101101010",
  20045=>"000101011",
  20046=>"111000001",
  20047=>"101011110",
  20048=>"111110001",
  20049=>"110110001",
  20050=>"001011101",
  20051=>"010010001",
  20052=>"110100010",
  20053=>"000111111",
  20054=>"111001110",
  20055=>"000111110",
  20056=>"110110011",
  20057=>"001110101",
  20058=>"000101101",
  20059=>"100101111",
  20060=>"100000000",
  20061=>"000000101",
  20062=>"011010000",
  20063=>"010110001",
  20064=>"111111001",
  20065=>"101011010",
  20066=>"000100000",
  20067=>"001011110",
  20068=>"000100111",
  20069=>"101111111",
  20070=>"110000100",
  20071=>"000000101",
  20072=>"000011110",
  20073=>"010001011",
  20074=>"100110101",
  20075=>"000000101",
  20076=>"101000111",
  20077=>"010101100",
  20078=>"001011011",
  20079=>"110110110",
  20080=>"100100001",
  20081=>"100010110",
  20082=>"010011000",
  20083=>"100001110",
  20084=>"001100001",
  20085=>"100110111",
  20086=>"000001011",
  20087=>"001111000",
  20088=>"111001000",
  20089=>"011000101",
  20090=>"010000110",
  20091=>"101011010",
  20092=>"100001110",
  20093=>"011111101",
  20094=>"101110111",
  20095=>"101101110",
  20096=>"000111011",
  20097=>"111001001",
  20098=>"011000110",
  20099=>"101010000",
  20100=>"100100010",
  20101=>"110010011",
  20102=>"010101011",
  20103=>"010110001",
  20104=>"001110101",
  20105=>"001000111",
  20106=>"000011000",
  20107=>"111111001",
  20108=>"011100000",
  20109=>"110000110",
  20110=>"110001110",
  20111=>"010100110",
  20112=>"011001001",
  20113=>"110111110",
  20114=>"110110100",
  20115=>"000101011",
  20116=>"110001110",
  20117=>"110001100",
  20118=>"111011110",
  20119=>"011101110",
  20120=>"110111000",
  20121=>"110110110",
  20122=>"001100001",
  20123=>"000010011",
  20124=>"111001111",
  20125=>"100010111",
  20126=>"011110011",
  20127=>"011010001",
  20128=>"111100111",
  20129=>"010111101",
  20130=>"011111011",
  20131=>"111010001",
  20132=>"001110100",
  20133=>"111100001",
  20134=>"011001000",
  20135=>"011010011",
  20136=>"010100011",
  20137=>"011011001",
  20138=>"000111011",
  20139=>"110001010",
  20140=>"100110101",
  20141=>"001100010",
  20142=>"100010101",
  20143=>"111111000",
  20144=>"000001110",
  20145=>"001000001",
  20146=>"010001100",
  20147=>"100010111",
  20148=>"001010001",
  20149=>"011011100",
  20150=>"111110111",
  20151=>"000100111",
  20152=>"010101110",
  20153=>"101101000",
  20154=>"100101110",
  20155=>"001101100",
  20156=>"101010110",
  20157=>"011001110",
  20158=>"111111001",
  20159=>"011001001",
  20160=>"010101101",
  20161=>"000110101",
  20162=>"110011101",
  20163=>"111111001",
  20164=>"110110011",
  20165=>"100011111",
  20166=>"010011000",
  20167=>"000101100",
  20168=>"100110111",
  20169=>"111111100",
  20170=>"011010001",
  20171=>"101000111",
  20172=>"011000000",
  20173=>"011100001",
  20174=>"001001010",
  20175=>"010011111",
  20176=>"001101010",
  20177=>"001110111",
  20178=>"110100100",
  20179=>"100100101",
  20180=>"011011010",
  20181=>"001111001",
  20182=>"001100111",
  20183=>"011110101",
  20184=>"000000000",
  20185=>"000101111",
  20186=>"110110000",
  20187=>"000011110",
  20188=>"101001100",
  20189=>"000001011",
  20190=>"111101101",
  20191=>"111111110",
  20192=>"101101111",
  20193=>"101010100",
  20194=>"100010100",
  20195=>"100110001",
  20196=>"111101100",
  20197=>"111011101",
  20198=>"111111101",
  20199=>"010111101",
  20200=>"101001101",
  20201=>"111000100",
  20202=>"101000101",
  20203=>"001000100",
  20204=>"110000110",
  20205=>"000100010",
  20206=>"100011011",
  20207=>"011100011",
  20208=>"010001001",
  20209=>"100001001",
  20210=>"010010111",
  20211=>"000110001",
  20212=>"011010100",
  20213=>"001000100",
  20214=>"001000110",
  20215=>"011001010",
  20216=>"001111100",
  20217=>"101001100",
  20218=>"100011001",
  20219=>"100001100",
  20220=>"111111100",
  20221=>"111010001",
  20222=>"101111010",
  20223=>"111011101",
  20224=>"111110010",
  20225=>"010010110",
  20226=>"110011010",
  20227=>"011001010",
  20228=>"011011010",
  20229=>"110111000",
  20230=>"000111001",
  20231=>"100000000",
  20232=>"100001101",
  20233=>"001100011",
  20234=>"111111010",
  20235=>"001100110",
  20236=>"111011001",
  20237=>"000010011",
  20238=>"011001111",
  20239=>"010100110",
  20240=>"011001111",
  20241=>"000010111",
  20242=>"110010100",
  20243=>"101011000",
  20244=>"111100000",
  20245=>"110101011",
  20246=>"000100010",
  20247=>"010011001",
  20248=>"010011111",
  20249=>"111001111",
  20250=>"101100010",
  20251=>"110110101",
  20252=>"100000110",
  20253=>"011011010",
  20254=>"001111011",
  20255=>"001000000",
  20256=>"001101010",
  20257=>"100100000",
  20258=>"011101101",
  20259=>"110000001",
  20260=>"111111001",
  20261=>"011111111",
  20262=>"011000011",
  20263=>"010011011",
  20264=>"110011011",
  20265=>"000010000",
  20266=>"001011001",
  20267=>"001100100",
  20268=>"100011111",
  20269=>"011000011",
  20270=>"100000000",
  20271=>"001111001",
  20272=>"110101111",
  20273=>"001101111",
  20274=>"101001101",
  20275=>"101100110",
  20276=>"001000111",
  20277=>"000100100",
  20278=>"000011101",
  20279=>"011100000",
  20280=>"101100110",
  20281=>"111001111",
  20282=>"000110000",
  20283=>"001001010",
  20284=>"111111011",
  20285=>"011111100",
  20286=>"101101110",
  20287=>"010101110",
  20288=>"000011001",
  20289=>"011011100",
  20290=>"111110101",
  20291=>"001011010",
  20292=>"001100001",
  20293=>"001011110",
  20294=>"000001101",
  20295=>"011111101",
  20296=>"011111111",
  20297=>"110111000",
  20298=>"010101000",
  20299=>"000100011",
  20300=>"110001111",
  20301=>"101101101",
  20302=>"000110011",
  20303=>"010111011",
  20304=>"011000111",
  20305=>"101011110",
  20306=>"111011110",
  20307=>"000011111",
  20308=>"010001010",
  20309=>"000100110",
  20310=>"010110001",
  20311=>"011111010",
  20312=>"111010000",
  20313=>"100101111",
  20314=>"101101101",
  20315=>"110001001",
  20316=>"111011011",
  20317=>"100111111",
  20318=>"000010000",
  20319=>"001011110",
  20320=>"100001111",
  20321=>"110001100",
  20322=>"111001011",
  20323=>"101111001",
  20324=>"001110101",
  20325=>"111011100",
  20326=>"101101001",
  20327=>"110110001",
  20328=>"101011100",
  20329=>"110111011",
  20330=>"001000010",
  20331=>"000111111",
  20332=>"011010011",
  20333=>"111001001",
  20334=>"000110110",
  20335=>"000010111",
  20336=>"010010010",
  20337=>"010001110",
  20338=>"000011110",
  20339=>"111110100",
  20340=>"101111110",
  20341=>"001100111",
  20342=>"111100000",
  20343=>"000011010",
  20344=>"001001110",
  20345=>"010111110",
  20346=>"100000000",
  20347=>"100001111",
  20348=>"010010010",
  20349=>"001001111",
  20350=>"010011110",
  20351=>"111010100",
  20352=>"011000111",
  20353=>"001011000",
  20354=>"111110011",
  20355=>"110001110",
  20356=>"001110100",
  20357=>"000000010",
  20358=>"110000110",
  20359=>"001000100",
  20360=>"000001111",
  20361=>"100000110",
  20362=>"110111010",
  20363=>"111101110",
  20364=>"011011010",
  20365=>"110011010",
  20366=>"100111110",
  20367=>"000111011",
  20368=>"001010101",
  20369=>"001100001",
  20370=>"110100011",
  20371=>"010101000",
  20372=>"011000011",
  20373=>"011111010",
  20374=>"011011111",
  20375=>"110010000",
  20376=>"000000101",
  20377=>"100110101",
  20378=>"000011101",
  20379=>"000110111",
  20380=>"100000100",
  20381=>"011101001",
  20382=>"011101010",
  20383=>"011010001",
  20384=>"101001101",
  20385=>"000001100",
  20386=>"100111110",
  20387=>"100011011",
  20388=>"111100101",
  20389=>"100111100",
  20390=>"101101110",
  20391=>"000111111",
  20392=>"101111111",
  20393=>"000010111",
  20394=>"000100100",
  20395=>"011110111",
  20396=>"101010010",
  20397=>"001100010",
  20398=>"001111000",
  20399=>"001110011",
  20400=>"001010010",
  20401=>"110001111",
  20402=>"000110000",
  20403=>"100010010",
  20404=>"000011110",
  20405=>"100110110",
  20406=>"010001010",
  20407=>"110110110",
  20408=>"101000010",
  20409=>"001011010",
  20410=>"111011001",
  20411=>"100100101",
  20412=>"011110001",
  20413=>"001001000",
  20414=>"110111111",
  20415=>"101110010",
  20416=>"110001101",
  20417=>"000000111",
  20418=>"011100011",
  20419=>"100110000",
  20420=>"111000011",
  20421=>"100111000",
  20422=>"110011000",
  20423=>"100100000",
  20424=>"010111001",
  20425=>"100001011",
  20426=>"111110100",
  20427=>"011111001",
  20428=>"101000101",
  20429=>"110010001",
  20430=>"001100011",
  20431=>"110111001",
  20432=>"010111110",
  20433=>"110000011",
  20434=>"000001111",
  20435=>"011011000",
  20436=>"010001110",
  20437=>"011000110",
  20438=>"111000000",
  20439=>"100011000",
  20440=>"000100010",
  20441=>"001111111",
  20442=>"001010000",
  20443=>"110110100",
  20444=>"111000111",
  20445=>"101011001",
  20446=>"001010100",
  20447=>"101010011",
  20448=>"011010111",
  20449=>"111000010",
  20450=>"101101011",
  20451=>"101000101",
  20452=>"000111100",
  20453=>"011000111",
  20454=>"111011111",
  20455=>"110111111",
  20456=>"001000010",
  20457=>"110111010",
  20458=>"100100010",
  20459=>"101010101",
  20460=>"010011100",
  20461=>"111000001",
  20462=>"101101011",
  20463=>"100000011",
  20464=>"110101110",
  20465=>"000011101",
  20466=>"111011011",
  20467=>"001010011",
  20468=>"011001000",
  20469=>"010111000",
  20470=>"110110100",
  20471=>"011100111",
  20472=>"111100000",
  20473=>"100001101",
  20474=>"111010011",
  20475=>"100011000",
  20476=>"000001111",
  20477=>"101100001",
  20478=>"000010100",
  20479=>"010111100",
  20480=>"000100001",
  20481=>"111100100",
  20482=>"011011100",
  20483=>"111110000",
  20484=>"111100110",
  20485=>"100010100",
  20486=>"101010000",
  20487=>"011010001",
  20488=>"100101001",
  20489=>"101100011",
  20490=>"110100010",
  20491=>"111110011",
  20492=>"101110110",
  20493=>"001001111",
  20494=>"000101111",
  20495=>"111111101",
  20496=>"011000000",
  20497=>"001110000",
  20498=>"010101101",
  20499=>"101000011",
  20500=>"000010000",
  20501=>"010100000",
  20502=>"111101010",
  20503=>"110010000",
  20504=>"101100001",
  20505=>"001000001",
  20506=>"110100111",
  20507=>"000100011",
  20508=>"110001000",
  20509=>"000001101",
  20510=>"101111101",
  20511=>"001101001",
  20512=>"111100110",
  20513=>"101001010",
  20514=>"110111111",
  20515=>"000000101",
  20516=>"100010100",
  20517=>"110000101",
  20518=>"111001100",
  20519=>"110011111",
  20520=>"010111011",
  20521=>"001011111",
  20522=>"000010101",
  20523=>"101000011",
  20524=>"100000001",
  20525=>"101101101",
  20526=>"101101010",
  20527=>"010110100",
  20528=>"001001110",
  20529=>"110000001",
  20530=>"001001000",
  20531=>"101001001",
  20532=>"101111001",
  20533=>"100100011",
  20534=>"001011100",
  20535=>"100000000",
  20536=>"000001001",
  20537=>"111010000",
  20538=>"001011101",
  20539=>"011111101",
  20540=>"001110100",
  20541=>"011110000",
  20542=>"000111111",
  20543=>"110100101",
  20544=>"110001001",
  20545=>"110101111",
  20546=>"111001000",
  20547=>"000000001",
  20548=>"110100110",
  20549=>"010001100",
  20550=>"000011111",
  20551=>"100110100",
  20552=>"101100100",
  20553=>"100110000",
  20554=>"010010000",
  20555=>"001011111",
  20556=>"011000111",
  20557=>"000001111",
  20558=>"100001110",
  20559=>"100111011",
  20560=>"111010010",
  20561=>"100000100",
  20562=>"101000010",
  20563=>"001010111",
  20564=>"101010000",
  20565=>"011110011",
  20566=>"100100101",
  20567=>"001000110",
  20568=>"011010000",
  20569=>"110100101",
  20570=>"010010111",
  20571=>"010011101",
  20572=>"010011000",
  20573=>"100000110",
  20574=>"000111011",
  20575=>"010100010",
  20576=>"000011000",
  20577=>"001000001",
  20578=>"001001001",
  20579=>"111111110",
  20580=>"101001111",
  20581=>"011110010",
  20582=>"101010101",
  20583=>"000000001",
  20584=>"001100100",
  20585=>"001111001",
  20586=>"111110000",
  20587=>"000001000",
  20588=>"000001011",
  20589=>"001101010",
  20590=>"111111000",
  20591=>"001101010",
  20592=>"100001011",
  20593=>"000111011",
  20594=>"111111101",
  20595=>"000010000",
  20596=>"001111111",
  20597=>"100100110",
  20598=>"000100111",
  20599=>"000000100",
  20600=>"001000001",
  20601=>"101111001",
  20602=>"001110111",
  20603=>"000010011",
  20604=>"000100001",
  20605=>"101110101",
  20606=>"100010000",
  20607=>"101000111",
  20608=>"001000001",
  20609=>"010001010",
  20610=>"101000000",
  20611=>"010000001",
  20612=>"001001100",
  20613=>"011010110",
  20614=>"011101110",
  20615=>"010001011",
  20616=>"101101100",
  20617=>"000000010",
  20618=>"101111100",
  20619=>"101010010",
  20620=>"111000111",
  20621=>"110101101",
  20622=>"101111101",
  20623=>"001111101",
  20624=>"110100101",
  20625=>"000010010",
  20626=>"000001100",
  20627=>"111010101",
  20628=>"101011101",
  20629=>"000001100",
  20630=>"010101011",
  20631=>"001001111",
  20632=>"101001000",
  20633=>"001000001",
  20634=>"000011011",
  20635=>"110101010",
  20636=>"001101110",
  20637=>"000101000",
  20638=>"000001000",
  20639=>"001010011",
  20640=>"100100101",
  20641=>"000111100",
  20642=>"111100001",
  20643=>"100011111",
  20644=>"110111100",
  20645=>"101010111",
  20646=>"101110010",
  20647=>"101100010",
  20648=>"110011110",
  20649=>"010110111",
  20650=>"001010011",
  20651=>"010000011",
  20652=>"101000000",
  20653=>"100000000",
  20654=>"011111100",
  20655=>"111101110",
  20656=>"010100011",
  20657=>"011010000",
  20658=>"100111001",
  20659=>"000000001",
  20660=>"110010010",
  20661=>"010111000",
  20662=>"101101010",
  20663=>"101100110",
  20664=>"010001001",
  20665=>"101101010",
  20666=>"101011100",
  20667=>"001001000",
  20668=>"010100110",
  20669=>"010010010",
  20670=>"010011001",
  20671=>"111111111",
  20672=>"011101100",
  20673=>"010011101",
  20674=>"100011000",
  20675=>"101110000",
  20676=>"001101101",
  20677=>"111110100",
  20678=>"000000111",
  20679=>"001100100",
  20680=>"011011011",
  20681=>"001001110",
  20682=>"110001010",
  20683=>"110100000",
  20684=>"001100111",
  20685=>"001101011",
  20686=>"001110110",
  20687=>"111111111",
  20688=>"010001110",
  20689=>"100100010",
  20690=>"101001100",
  20691=>"001000001",
  20692=>"101100110",
  20693=>"000011110",
  20694=>"111011010",
  20695=>"101110010",
  20696=>"001100001",
  20697=>"011000111",
  20698=>"110101011",
  20699=>"000011000",
  20700=>"111110001",
  20701=>"000011100",
  20702=>"110001111",
  20703=>"010001011",
  20704=>"011101001",
  20705=>"100011110",
  20706=>"010001111",
  20707=>"110010011",
  20708=>"010111111",
  20709=>"101011000",
  20710=>"001011110",
  20711=>"000001100",
  20712=>"000100101",
  20713=>"110100101",
  20714=>"001111110",
  20715=>"000011111",
  20716=>"100000000",
  20717=>"101010001",
  20718=>"101010000",
  20719=>"011110011",
  20720=>"011100011",
  20721=>"011011111",
  20722=>"001001000",
  20723=>"100011001",
  20724=>"000110111",
  20725=>"110100110",
  20726=>"111011100",
  20727=>"100111010",
  20728=>"001101111",
  20729=>"001110000",
  20730=>"000001101",
  20731=>"100111001",
  20732=>"000101000",
  20733=>"111010101",
  20734=>"000111011",
  20735=>"110111010",
  20736=>"000001101",
  20737=>"111101111",
  20738=>"000000010",
  20739=>"101110010",
  20740=>"011100000",
  20741=>"010101001",
  20742=>"000001001",
  20743=>"001010110",
  20744=>"000010000",
  20745=>"010111000",
  20746=>"001101111",
  20747=>"000000111",
  20748=>"100100001",
  20749=>"101000000",
  20750=>"010110000",
  20751=>"000001100",
  20752=>"000100111",
  20753=>"011000010",
  20754=>"101000100",
  20755=>"110010110",
  20756=>"010110000",
  20757=>"110100011",
  20758=>"111101111",
  20759=>"001000100",
  20760=>"010011110",
  20761=>"100001010",
  20762=>"001010101",
  20763=>"001000101",
  20764=>"010110011",
  20765=>"101001100",
  20766=>"100101001",
  20767=>"111001101",
  20768=>"000100000",
  20769=>"011110000",
  20770=>"110100101",
  20771=>"111011111",
  20772=>"100111101",
  20773=>"110111010",
  20774=>"100010010",
  20775=>"100100100",
  20776=>"111001101",
  20777=>"110110011",
  20778=>"011110000",
  20779=>"100110000",
  20780=>"001110111",
  20781=>"110111111",
  20782=>"011110011",
  20783=>"100101110",
  20784=>"111011001",
  20785=>"110010010",
  20786=>"011001001",
  20787=>"111001000",
  20788=>"101100011",
  20789=>"010000001",
  20790=>"011110111",
  20791=>"000101010",
  20792=>"001001001",
  20793=>"110111001",
  20794=>"100110101",
  20795=>"000001000",
  20796=>"100011100",
  20797=>"001100011",
  20798=>"001110101",
  20799=>"110000100",
  20800=>"111101110",
  20801=>"101101101",
  20802=>"101101111",
  20803=>"101011111",
  20804=>"101111000",
  20805=>"011011101",
  20806=>"010000011",
  20807=>"101110101",
  20808=>"101011111",
  20809=>"111000101",
  20810=>"110111011",
  20811=>"000001010",
  20812=>"101010111",
  20813=>"110101010",
  20814=>"110001101",
  20815=>"001001010",
  20816=>"000010011",
  20817=>"010110101",
  20818=>"011000001",
  20819=>"000000101",
  20820=>"111011111",
  20821=>"000110111",
  20822=>"101000000",
  20823=>"111111111",
  20824=>"100000101",
  20825=>"110011010",
  20826=>"100001000",
  20827=>"111000000",
  20828=>"101000111",
  20829=>"011010010",
  20830=>"111000101",
  20831=>"011001000",
  20832=>"000001100",
  20833=>"111111111",
  20834=>"000011000",
  20835=>"001011110",
  20836=>"111100101",
  20837=>"111010100",
  20838=>"001110001",
  20839=>"111110100",
  20840=>"010100001",
  20841=>"100011111",
  20842=>"000101000",
  20843=>"111110001",
  20844=>"110111100",
  20845=>"111011010",
  20846=>"001000101",
  20847=>"001011001",
  20848=>"100000010",
  20849=>"000000011",
  20850=>"010101100",
  20851=>"111001111",
  20852=>"011111000",
  20853=>"100000100",
  20854=>"000101000",
  20855=>"001111011",
  20856=>"011010101",
  20857=>"100011001",
  20858=>"011111010",
  20859=>"001101010",
  20860=>"001000001",
  20861=>"011000110",
  20862=>"000100011",
  20863=>"010111000",
  20864=>"001011101",
  20865=>"010001001",
  20866=>"111010100",
  20867=>"110101101",
  20868=>"101011111",
  20869=>"110000011",
  20870=>"000111110",
  20871=>"000000101",
  20872=>"001000001",
  20873=>"100111100",
  20874=>"100111011",
  20875=>"110101100",
  20876=>"110111100",
  20877=>"111111100",
  20878=>"101101110",
  20879=>"101100111",
  20880=>"011101010",
  20881=>"111100110",
  20882=>"110100000",
  20883=>"110101011",
  20884=>"001100111",
  20885=>"100000011",
  20886=>"101111010",
  20887=>"110100010",
  20888=>"111000100",
  20889=>"010110111",
  20890=>"000100100",
  20891=>"010000000",
  20892=>"101101100",
  20893=>"111111010",
  20894=>"100000110",
  20895=>"001011001",
  20896=>"001111011",
  20897=>"011000101",
  20898=>"111010011",
  20899=>"110110110",
  20900=>"111010101",
  20901=>"010111101",
  20902=>"100000100",
  20903=>"111111111",
  20904=>"101111111",
  20905=>"101001110",
  20906=>"000100001",
  20907=>"010111101",
  20908=>"110011111",
  20909=>"010011101",
  20910=>"110000101",
  20911=>"110000101",
  20912=>"001010000",
  20913=>"000010001",
  20914=>"001011000",
  20915=>"101110111",
  20916=>"100110010",
  20917=>"100011000",
  20918=>"011001001",
  20919=>"010111010",
  20920=>"000001101",
  20921=>"011110101",
  20922=>"101011111",
  20923=>"010110000",
  20924=>"101001101",
  20925=>"011100101",
  20926=>"011100110",
  20927=>"110010100",
  20928=>"000000000",
  20929=>"111111000",
  20930=>"011011011",
  20931=>"110000011",
  20932=>"001110110",
  20933=>"110100100",
  20934=>"110110101",
  20935=>"000011000",
  20936=>"110101001",
  20937=>"110101011",
  20938=>"001110001",
  20939=>"000101100",
  20940=>"000000001",
  20941=>"001100101",
  20942=>"111111011",
  20943=>"100001001",
  20944=>"011011100",
  20945=>"001100110",
  20946=>"111111110",
  20947=>"001010100",
  20948=>"101001001",
  20949=>"101110101",
  20950=>"101110111",
  20951=>"110110111",
  20952=>"010010100",
  20953=>"101111101",
  20954=>"111111100",
  20955=>"010000001",
  20956=>"111011110",
  20957=>"101100111",
  20958=>"011101101",
  20959=>"111011011",
  20960=>"111101100",
  20961=>"111101011",
  20962=>"010101110",
  20963=>"100010100",
  20964=>"100010000",
  20965=>"111010010",
  20966=>"000101011",
  20967=>"010000010",
  20968=>"111011110",
  20969=>"100010100",
  20970=>"100000110",
  20971=>"101001111",
  20972=>"010110111",
  20973=>"100001110",
  20974=>"001000100",
  20975=>"101100011",
  20976=>"011010101",
  20977=>"110111011",
  20978=>"110010111",
  20979=>"110001111",
  20980=>"011101011",
  20981=>"101111111",
  20982=>"011110101",
  20983=>"110000100",
  20984=>"000000110",
  20985=>"010101011",
  20986=>"111111001",
  20987=>"011000110",
  20988=>"101000001",
  20989=>"000001101",
  20990=>"101110101",
  20991=>"000000000",
  20992=>"110001001",
  20993=>"010110001",
  20994=>"110011110",
  20995=>"101001001",
  20996=>"010010001",
  20997=>"000101001",
  20998=>"000101101",
  20999=>"010001001",
  21000=>"000101101",
  21001=>"101011101",
  21002=>"010011011",
  21003=>"000001001",
  21004=>"110001010",
  21005=>"110101101",
  21006=>"011001001",
  21007=>"011001101",
  21008=>"110100000",
  21009=>"110100010",
  21010=>"001100100",
  21011=>"110011110",
  21012=>"110111100",
  21013=>"111011010",
  21014=>"011110110",
  21015=>"111000000",
  21016=>"111110010",
  21017=>"011111000",
  21018=>"100110101",
  21019=>"100111110",
  21020=>"110111110",
  21021=>"011111100",
  21022=>"010101111",
  21023=>"000110110",
  21024=>"110000111",
  21025=>"001000101",
  21026=>"100110110",
  21027=>"010111111",
  21028=>"111011011",
  21029=>"000000110",
  21030=>"001110000",
  21031=>"100010010",
  21032=>"101101101",
  21033=>"101011101",
  21034=>"000100111",
  21035=>"001111010",
  21036=>"001101000",
  21037=>"001100010",
  21038=>"010000010",
  21039=>"100001100",
  21040=>"001110010",
  21041=>"010110000",
  21042=>"010000001",
  21043=>"111100111",
  21044=>"100100000",
  21045=>"000010111",
  21046=>"111011011",
  21047=>"001111110",
  21048=>"110011100",
  21049=>"010110110",
  21050=>"101000001",
  21051=>"111000110",
  21052=>"011100111",
  21053=>"001011100",
  21054=>"100001010",
  21055=>"101010100",
  21056=>"001000001",
  21057=>"110011000",
  21058=>"001000001",
  21059=>"100010110",
  21060=>"110111011",
  21061=>"101000001",
  21062=>"000001001",
  21063=>"001000010",
  21064=>"010111110",
  21065=>"010101101",
  21066=>"001000110",
  21067=>"100010011",
  21068=>"001001000",
  21069=>"010111100",
  21070=>"100000010",
  21071=>"101000011",
  21072=>"001011000",
  21073=>"010010000",
  21074=>"101011100",
  21075=>"111010111",
  21076=>"001101011",
  21077=>"101100000",
  21078=>"001000100",
  21079=>"001110001",
  21080=>"001010001",
  21081=>"101110010",
  21082=>"111110111",
  21083=>"000110110",
  21084=>"000011010",
  21085=>"000111000",
  21086=>"000010010",
  21087=>"000100100",
  21088=>"111001010",
  21089=>"000101101",
  21090=>"000001111",
  21091=>"110100110",
  21092=>"011111010",
  21093=>"111010000",
  21094=>"110111101",
  21095=>"110001111",
  21096=>"110010100",
  21097=>"111101000",
  21098=>"110010110",
  21099=>"110011011",
  21100=>"011100100",
  21101=>"101010000",
  21102=>"010101111",
  21103=>"100000100",
  21104=>"110111110",
  21105=>"010100110",
  21106=>"100000110",
  21107=>"110010101",
  21108=>"100000011",
  21109=>"010100000",
  21110=>"000101100",
  21111=>"010110011",
  21112=>"001000101",
  21113=>"111010011",
  21114=>"101001001",
  21115=>"111101011",
  21116=>"100101001",
  21117=>"000101111",
  21118=>"010000101",
  21119=>"110011101",
  21120=>"010001011",
  21121=>"111000100",
  21122=>"000111010",
  21123=>"001010001",
  21124=>"001110100",
  21125=>"001001000",
  21126=>"010101001",
  21127=>"110011011",
  21128=>"010111000",
  21129=>"001111001",
  21130=>"100000011",
  21131=>"111110100",
  21132=>"000001011",
  21133=>"101000010",
  21134=>"110111001",
  21135=>"011100010",
  21136=>"110001010",
  21137=>"000011000",
  21138=>"010100111",
  21139=>"000010101",
  21140=>"000100101",
  21141=>"001100001",
  21142=>"010101001",
  21143=>"001100000",
  21144=>"101011101",
  21145=>"000111001",
  21146=>"010101100",
  21147=>"001010101",
  21148=>"000011000",
  21149=>"011001010",
  21150=>"111100111",
  21151=>"111011100",
  21152=>"001011111",
  21153=>"000001110",
  21154=>"010001011",
  21155=>"101000101",
  21156=>"011110000",
  21157=>"110011000",
  21158=>"001100101",
  21159=>"011100110",
  21160=>"101001001",
  21161=>"011010110",
  21162=>"101111011",
  21163=>"101101001",
  21164=>"100001001",
  21165=>"101000011",
  21166=>"100111101",
  21167=>"011011101",
  21168=>"001000110",
  21169=>"110010101",
  21170=>"010101001",
  21171=>"001111010",
  21172=>"001010011",
  21173=>"101101101",
  21174=>"110010100",
  21175=>"001011000",
  21176=>"000111100",
  21177=>"010001000",
  21178=>"101111100",
  21179=>"001001101",
  21180=>"011001100",
  21181=>"111001100",
  21182=>"000111001",
  21183=>"111010010",
  21184=>"101101000",
  21185=>"100001010",
  21186=>"010000100",
  21187=>"001000100",
  21188=>"100011010",
  21189=>"011100010",
  21190=>"100101111",
  21191=>"110111010",
  21192=>"000000111",
  21193=>"000010101",
  21194=>"111110100",
  21195=>"111011100",
  21196=>"110000010",
  21197=>"000001110",
  21198=>"010000010",
  21199=>"001010011",
  21200=>"111111001",
  21201=>"110010101",
  21202=>"001101001",
  21203=>"010111011",
  21204=>"101101101",
  21205=>"010001011",
  21206=>"000100011",
  21207=>"101001001",
  21208=>"101011111",
  21209=>"011001110",
  21210=>"000000111",
  21211=>"011100001",
  21212=>"001100010",
  21213=>"000111100",
  21214=>"011100111",
  21215=>"000101001",
  21216=>"111101011",
  21217=>"001001011",
  21218=>"000101010",
  21219=>"110101101",
  21220=>"101111011",
  21221=>"111100000",
  21222=>"110010000",
  21223=>"000011101",
  21224=>"000001001",
  21225=>"110001100",
  21226=>"111000100",
  21227=>"101010101",
  21228=>"000000001",
  21229=>"000000110",
  21230=>"101101010",
  21231=>"100101110",
  21232=>"000011011",
  21233=>"101101000",
  21234=>"011001101",
  21235=>"110000000",
  21236=>"111100100",
  21237=>"010110110",
  21238=>"000100000",
  21239=>"111011111",
  21240=>"100011101",
  21241=>"111011110",
  21242=>"001101000",
  21243=>"110110101",
  21244=>"110101001",
  21245=>"001101111",
  21246=>"000100011",
  21247=>"010010010",
  21248=>"101111001",
  21249=>"010101000",
  21250=>"000101001",
  21251=>"101111100",
  21252=>"000010110",
  21253=>"000110101",
  21254=>"110111000",
  21255=>"111011011",
  21256=>"110101000",
  21257=>"100011010",
  21258=>"010010110",
  21259=>"000001000",
  21260=>"000110100",
  21261=>"101101010",
  21262=>"111100000",
  21263=>"110000101",
  21264=>"000010110",
  21265=>"000011000",
  21266=>"111100001",
  21267=>"001010000",
  21268=>"101001001",
  21269=>"000011000",
  21270=>"011010001",
  21271=>"000000001",
  21272=>"010101111",
  21273=>"000100110",
  21274=>"010100010",
  21275=>"101011101",
  21276=>"100111110",
  21277=>"101101000",
  21278=>"111100111",
  21279=>"111111100",
  21280=>"100110011",
  21281=>"101111100",
  21282=>"010010010",
  21283=>"101010010",
  21284=>"111111010",
  21285=>"010010110",
  21286=>"001101111",
  21287=>"010110010",
  21288=>"110111010",
  21289=>"011000010",
  21290=>"011111011",
  21291=>"111101110",
  21292=>"100000110",
  21293=>"000101100",
  21294=>"001111111",
  21295=>"001100111",
  21296=>"001001011",
  21297=>"001010010",
  21298=>"101111111",
  21299=>"100001110",
  21300=>"000001110",
  21301=>"001000011",
  21302=>"111001110",
  21303=>"000111111",
  21304=>"011111111",
  21305=>"100000101",
  21306=>"110100100",
  21307=>"111001110",
  21308=>"000000111",
  21309=>"010101100",
  21310=>"001110001",
  21311=>"010001011",
  21312=>"111111101",
  21313=>"100111000",
  21314=>"111010100",
  21315=>"111101010",
  21316=>"000001100",
  21317=>"001100010",
  21318=>"101110100",
  21319=>"000011101",
  21320=>"011100010",
  21321=>"100110010",
  21322=>"000100010",
  21323=>"110100101",
  21324=>"011101101",
  21325=>"010011000",
  21326=>"010010010",
  21327=>"111010001",
  21328=>"100101011",
  21329=>"000100111",
  21330=>"010011010",
  21331=>"011011010",
  21332=>"101100101",
  21333=>"001101010",
  21334=>"011101011",
  21335=>"110000101",
  21336=>"011110010",
  21337=>"101101110",
  21338=>"010100101",
  21339=>"001101100",
  21340=>"110101101",
  21341=>"110110011",
  21342=>"000111110",
  21343=>"000111010",
  21344=>"110001100",
  21345=>"100111001",
  21346=>"101001011",
  21347=>"010000110",
  21348=>"011111110",
  21349=>"111001001",
  21350=>"011100011",
  21351=>"000110101",
  21352=>"010101100",
  21353=>"001001011",
  21354=>"110001101",
  21355=>"110100010",
  21356=>"001111110",
  21357=>"000100110",
  21358=>"101100111",
  21359=>"100001111",
  21360=>"100100100",
  21361=>"111110101",
  21362=>"111011111",
  21363=>"000100101",
  21364=>"001110111",
  21365=>"110001000",
  21366=>"100110100",
  21367=>"100000100",
  21368=>"110111000",
  21369=>"101100011",
  21370=>"001110010",
  21371=>"111010110",
  21372=>"010101010",
  21373=>"100001001",
  21374=>"000100001",
  21375=>"110111011",
  21376=>"001011010",
  21377=>"111001111",
  21378=>"000011111",
  21379=>"011000111",
  21380=>"100100000",
  21381=>"010000010",
  21382=>"101111011",
  21383=>"000001101",
  21384=>"000111010",
  21385=>"011110101",
  21386=>"000111111",
  21387=>"101010101",
  21388=>"011100011",
  21389=>"001110000",
  21390=>"100111000",
  21391=>"010001011",
  21392=>"001000001",
  21393=>"000101110",
  21394=>"001110110",
  21395=>"101101111",
  21396=>"111000111",
  21397=>"111000110",
  21398=>"100000110",
  21399=>"101001001",
  21400=>"101111101",
  21401=>"110110110",
  21402=>"010101111",
  21403=>"010010100",
  21404=>"110000000",
  21405=>"101101001",
  21406=>"110000110",
  21407=>"111100001",
  21408=>"011101100",
  21409=>"000101101",
  21410=>"100011111",
  21411=>"001110111",
  21412=>"011100000",
  21413=>"111001011",
  21414=>"011111110",
  21415=>"001110100",
  21416=>"111000101",
  21417=>"000000010",
  21418=>"111110010",
  21419=>"001000001",
  21420=>"100110000",
  21421=>"101000110",
  21422=>"010001100",
  21423=>"010100000",
  21424=>"110000101",
  21425=>"011010111",
  21426=>"110111010",
  21427=>"011010111",
  21428=>"010011111",
  21429=>"000000100",
  21430=>"101001110",
  21431=>"011111000",
  21432=>"110010101",
  21433=>"001001000",
  21434=>"000101101",
  21435=>"101001010",
  21436=>"010100100",
  21437=>"110011010",
  21438=>"111001010",
  21439=>"000000000",
  21440=>"001110010",
  21441=>"001010111",
  21442=>"111111100",
  21443=>"011001111",
  21444=>"100101111",
  21445=>"101110011",
  21446=>"110011111",
  21447=>"000101011",
  21448=>"101001101",
  21449=>"000000000",
  21450=>"111000010",
  21451=>"110101000",
  21452=>"011101101",
  21453=>"000110110",
  21454=>"110011001",
  21455=>"111100011",
  21456=>"101101011",
  21457=>"000101000",
  21458=>"011100000",
  21459=>"001100000",
  21460=>"001010101",
  21461=>"011001001",
  21462=>"110010001",
  21463=>"001000011",
  21464=>"100001011",
  21465=>"101110110",
  21466=>"011111101",
  21467=>"000000001",
  21468=>"100100010",
  21469=>"111110110",
  21470=>"010011001",
  21471=>"001000010",
  21472=>"100110011",
  21473=>"101110010",
  21474=>"101010010",
  21475=>"000101011",
  21476=>"011001001",
  21477=>"001011101",
  21478=>"100011110",
  21479=>"111101000",
  21480=>"000000100",
  21481=>"100010100",
  21482=>"000100110",
  21483=>"100101101",
  21484=>"000010110",
  21485=>"011001100",
  21486=>"010110101",
  21487=>"001001011",
  21488=>"010011110",
  21489=>"110100101",
  21490=>"011001010",
  21491=>"011101010",
  21492=>"000000010",
  21493=>"110010100",
  21494=>"110110111",
  21495=>"110110100",
  21496=>"111000000",
  21497=>"000010011",
  21498=>"111000010",
  21499=>"110110011",
  21500=>"011001111",
  21501=>"111110011",
  21502=>"101000011",
  21503=>"110100011",
  21504=>"011111110",
  21505=>"010110010",
  21506=>"001010101",
  21507=>"111110111",
  21508=>"010110101",
  21509=>"111101110",
  21510=>"011001111",
  21511=>"110010000",
  21512=>"110101010",
  21513=>"101010111",
  21514=>"101011101",
  21515=>"111100111",
  21516=>"000011010",
  21517=>"110000100",
  21518=>"101000011",
  21519=>"101111101",
  21520=>"100110001",
  21521=>"100111111",
  21522=>"111110101",
  21523=>"101011111",
  21524=>"110000101",
  21525=>"011001101",
  21526=>"111101001",
  21527=>"000010000",
  21528=>"010000000",
  21529=>"001001000",
  21530=>"111111111",
  21531=>"100000111",
  21532=>"111010101",
  21533=>"101000110",
  21534=>"110000101",
  21535=>"110001000",
  21536=>"001000000",
  21537=>"011110100",
  21538=>"111101111",
  21539=>"010100101",
  21540=>"111001110",
  21541=>"010111000",
  21542=>"111010011",
  21543=>"100001001",
  21544=>"101000001",
  21545=>"000101111",
  21546=>"101101110",
  21547=>"110110011",
  21548=>"011100111",
  21549=>"000100010",
  21550=>"000000011",
  21551=>"111111111",
  21552=>"110000100",
  21553=>"100001111",
  21554=>"111011100",
  21555=>"100000000",
  21556=>"101011011",
  21557=>"010010110",
  21558=>"000101000",
  21559=>"001011001",
  21560=>"110001100",
  21561=>"000011010",
  21562=>"101111110",
  21563=>"010001011",
  21564=>"000000100",
  21565=>"100100001",
  21566=>"111011110",
  21567=>"011011000",
  21568=>"100011001",
  21569=>"010000111",
  21570=>"100101101",
  21571=>"101111111",
  21572=>"101100111",
  21573=>"000101101",
  21574=>"110000110",
  21575=>"110110000",
  21576=>"001100011",
  21577=>"011101111",
  21578=>"010111101",
  21579=>"000100100",
  21580=>"000101100",
  21581=>"101000111",
  21582=>"101111010",
  21583=>"010110111",
  21584=>"000110011",
  21585=>"000100000",
  21586=>"100011001",
  21587=>"110100100",
  21588=>"111110001",
  21589=>"111111010",
  21590=>"010110100",
  21591=>"010010011",
  21592=>"110101110",
  21593=>"010111001",
  21594=>"011011011",
  21595=>"000011101",
  21596=>"100110010",
  21597=>"111100011",
  21598=>"010110100",
  21599=>"111001100",
  21600=>"000000110",
  21601=>"100101011",
  21602=>"111101001",
  21603=>"100000110",
  21604=>"100111101",
  21605=>"100010011",
  21606=>"110010100",
  21607=>"011100000",
  21608=>"111001101",
  21609=>"010110000",
  21610=>"101111000",
  21611=>"001010100",
  21612=>"011000101",
  21613=>"100010101",
  21614=>"011110000",
  21615=>"000010010",
  21616=>"111001001",
  21617=>"110000011",
  21618=>"110101100",
  21619=>"011110001",
  21620=>"101000111",
  21621=>"000110100",
  21622=>"001010000",
  21623=>"110101010",
  21624=>"110010100",
  21625=>"101000011",
  21626=>"011110101",
  21627=>"111000011",
  21628=>"100100001",
  21629=>"101011010",
  21630=>"101010001",
  21631=>"000000000",
  21632=>"010101000",
  21633=>"111001111",
  21634=>"010000001",
  21635=>"101000110",
  21636=>"000100000",
  21637=>"101111101",
  21638=>"110100000",
  21639=>"110000111",
  21640=>"010000010",
  21641=>"000101010",
  21642=>"001001001",
  21643=>"000100100",
  21644=>"011011110",
  21645=>"011000100",
  21646=>"001101010",
  21647=>"111111101",
  21648=>"110000000",
  21649=>"011001101",
  21650=>"001101011",
  21651=>"001110000",
  21652=>"000110001",
  21653=>"011000100",
  21654=>"110011110",
  21655=>"011100101",
  21656=>"001111011",
  21657=>"110001110",
  21658=>"000110001",
  21659=>"000001100",
  21660=>"010011000",
  21661=>"011110001",
  21662=>"111101100",
  21663=>"001110100",
  21664=>"110101101",
  21665=>"100101010",
  21666=>"010101011",
  21667=>"010100101",
  21668=>"001011010",
  21669=>"010001111",
  21670=>"111101110",
  21671=>"100110110",
  21672=>"001001011",
  21673=>"100101101",
  21674=>"111101100",
  21675=>"010110111",
  21676=>"100000100",
  21677=>"110101010",
  21678=>"111000100",
  21679=>"010110010",
  21680=>"001100111",
  21681=>"001001110",
  21682=>"001001001",
  21683=>"110010100",
  21684=>"101101101",
  21685=>"010011101",
  21686=>"111000100",
  21687=>"111111001",
  21688=>"110111111",
  21689=>"001000010",
  21690=>"000001011",
  21691=>"111111110",
  21692=>"111110001",
  21693=>"101101011",
  21694=>"011110111",
  21695=>"111110101",
  21696=>"010000100",
  21697=>"100100011",
  21698=>"000001100",
  21699=>"010101000",
  21700=>"101011000",
  21701=>"000101001",
  21702=>"010001001",
  21703=>"001100101",
  21704=>"110111011",
  21705=>"001000101",
  21706=>"010001011",
  21707=>"010111101",
  21708=>"001011111",
  21709=>"111110010",
  21710=>"010011010",
  21711=>"011101001",
  21712=>"101000000",
  21713=>"110111011",
  21714=>"101000110",
  21715=>"101011100",
  21716=>"000011011",
  21717=>"010010110",
  21718=>"010101011",
  21719=>"000100010",
  21720=>"111101100",
  21721=>"000100010",
  21722=>"111100101",
  21723=>"000000110",
  21724=>"000111100",
  21725=>"110111100",
  21726=>"010110100",
  21727=>"010111010",
  21728=>"111000001",
  21729=>"011111001",
  21730=>"001101110",
  21731=>"010010111",
  21732=>"100001010",
  21733=>"100010000",
  21734=>"111101001",
  21735=>"101101010",
  21736=>"111110111",
  21737=>"101011011",
  21738=>"110110111",
  21739=>"010001000",
  21740=>"100100101",
  21741=>"100100111",
  21742=>"000001110",
  21743=>"010101100",
  21744=>"000001111",
  21745=>"111111110",
  21746=>"000111000",
  21747=>"000001111",
  21748=>"101111101",
  21749=>"100010010",
  21750=>"100011110",
  21751=>"001001001",
  21752=>"000101100",
  21753=>"000000100",
  21754=>"000010010",
  21755=>"100001101",
  21756=>"011000000",
  21757=>"101101000",
  21758=>"011111100",
  21759=>"010010000",
  21760=>"001001010",
  21761=>"011100010",
  21762=>"010001110",
  21763=>"110101010",
  21764=>"001001000",
  21765=>"100110100",
  21766=>"110010001",
  21767=>"000000011",
  21768=>"000001000",
  21769=>"100010010",
  21770=>"111011000",
  21771=>"111011111",
  21772=>"100010100",
  21773=>"010000100",
  21774=>"111100100",
  21775=>"011001001",
  21776=>"111110101",
  21777=>"000011010",
  21778=>"000010011",
  21779=>"010101001",
  21780=>"110100110",
  21781=>"011000111",
  21782=>"111001110",
  21783=>"010010000",
  21784=>"111101011",
  21785=>"100100010",
  21786=>"000010110",
  21787=>"111001111",
  21788=>"000111000",
  21789=>"111100011",
  21790=>"001000100",
  21791=>"010000100",
  21792=>"101101101",
  21793=>"000011010",
  21794=>"110000001",
  21795=>"001110000",
  21796=>"000011111",
  21797=>"101100100",
  21798=>"001001011",
  21799=>"100010011",
  21800=>"010001101",
  21801=>"000101001",
  21802=>"001100101",
  21803=>"111011110",
  21804=>"010011100",
  21805=>"010010000",
  21806=>"001111100",
  21807=>"010001111",
  21808=>"000010100",
  21809=>"001101101",
  21810=>"111101110",
  21811=>"100001111",
  21812=>"101100001",
  21813=>"001111000",
  21814=>"111100100",
  21815=>"011110001",
  21816=>"001010011",
  21817=>"011010100",
  21818=>"001011010",
  21819=>"001110100",
  21820=>"001101110",
  21821=>"100001110",
  21822=>"011101001",
  21823=>"010011010",
  21824=>"001000101",
  21825=>"011100111",
  21826=>"111101101",
  21827=>"010111110",
  21828=>"010100101",
  21829=>"010100010",
  21830=>"001111010",
  21831=>"000000100",
  21832=>"101101001",
  21833=>"111011001",
  21834=>"110011010",
  21835=>"000100001",
  21836=>"001110000",
  21837=>"000111010",
  21838=>"101100001",
  21839=>"101000000",
  21840=>"100110110",
  21841=>"111000101",
  21842=>"100110101",
  21843=>"110100011",
  21844=>"010101110",
  21845=>"100000011",
  21846=>"001100010",
  21847=>"100011100",
  21848=>"011001000",
  21849=>"111110110",
  21850=>"100000001",
  21851=>"010011100",
  21852=>"101100100",
  21853=>"110011001",
  21854=>"111111101",
  21855=>"101110110",
  21856=>"110010011",
  21857=>"101111001",
  21858=>"011101001",
  21859=>"010010000",
  21860=>"001001010",
  21861=>"100001001",
  21862=>"110001001",
  21863=>"011100000",
  21864=>"111100110",
  21865=>"111010101",
  21866=>"100001000",
  21867=>"011011101",
  21868=>"101000001",
  21869=>"100000001",
  21870=>"011100001",
  21871=>"110010010",
  21872=>"010001111",
  21873=>"001010111",
  21874=>"110010001",
  21875=>"101011000",
  21876=>"010000101",
  21877=>"111001101",
  21878=>"001010101",
  21879=>"010110100",
  21880=>"010111110",
  21881=>"110010110",
  21882=>"011000110",
  21883=>"111100011",
  21884=>"011000000",
  21885=>"110011111",
  21886=>"011110001",
  21887=>"000001000",
  21888=>"111100011",
  21889=>"110110011",
  21890=>"110100111",
  21891=>"110001100",
  21892=>"111100100",
  21893=>"011111001",
  21894=>"001010001",
  21895=>"111010101",
  21896=>"001001000",
  21897=>"000010110",
  21898=>"011010111",
  21899=>"110010101",
  21900=>"111111111",
  21901=>"111010001",
  21902=>"111010011",
  21903=>"000101011",
  21904=>"011000010",
  21905=>"001010111",
  21906=>"100110101",
  21907=>"111100111",
  21908=>"111011101",
  21909=>"100000000",
  21910=>"101101110",
  21911=>"001100110",
  21912=>"100001110",
  21913=>"110001101",
  21914=>"110111011",
  21915=>"100101000",
  21916=>"101000101",
  21917=>"010100001",
  21918=>"000111011",
  21919=>"010011010",
  21920=>"001100001",
  21921=>"011010011",
  21922=>"101001000",
  21923=>"111110010",
  21924=>"011010100",
  21925=>"110100000",
  21926=>"101111110",
  21927=>"001011110",
  21928=>"011110101",
  21929=>"010110010",
  21930=>"000000000",
  21931=>"010101010",
  21932=>"000111111",
  21933=>"110010100",
  21934=>"010010110",
  21935=>"010110111",
  21936=>"000000000",
  21937=>"111111001",
  21938=>"010110111",
  21939=>"000100000",
  21940=>"100011001",
  21941=>"100010110",
  21942=>"111110011",
  21943=>"000000011",
  21944=>"111010100",
  21945=>"011010000",
  21946=>"111010110",
  21947=>"111000001",
  21948=>"100111111",
  21949=>"100000111",
  21950=>"110001110",
  21951=>"001010001",
  21952=>"110111000",
  21953=>"110011011",
  21954=>"000000000",
  21955=>"000100010",
  21956=>"101110111",
  21957=>"000001111",
  21958=>"011111111",
  21959=>"011111000",
  21960=>"011001101",
  21961=>"010111111",
  21962=>"000111000",
  21963=>"101111101",
  21964=>"111111111",
  21965=>"000101110",
  21966=>"101001000",
  21967=>"011000000",
  21968=>"101100100",
  21969=>"000101111",
  21970=>"110001100",
  21971=>"011101100",
  21972=>"010011101",
  21973=>"001110010",
  21974=>"001011010",
  21975=>"010101001",
  21976=>"000000100",
  21977=>"111010001",
  21978=>"100111101",
  21979=>"100100001",
  21980=>"011110010",
  21981=>"010011100",
  21982=>"000001101",
  21983=>"000110111",
  21984=>"011011101",
  21985=>"011100100",
  21986=>"101101101",
  21987=>"110001011",
  21988=>"110011111",
  21989=>"110010001",
  21990=>"011011000",
  21991=>"011010000",
  21992=>"101111001",
  21993=>"010000111",
  21994=>"010001000",
  21995=>"101101000",
  21996=>"101010011",
  21997=>"010011001",
  21998=>"000001101",
  21999=>"011100001",
  22000=>"111101100",
  22001=>"010000101",
  22002=>"011000110",
  22003=>"000001100",
  22004=>"110000100",
  22005=>"011100000",
  22006=>"001100101",
  22007=>"101111000",
  22008=>"110000110",
  22009=>"000110000",
  22010=>"010001110",
  22011=>"110000001",
  22012=>"101101101",
  22013=>"111011111",
  22014=>"010010110",
  22015=>"011101110",
  22016=>"010111010",
  22017=>"100010111",
  22018=>"110000001",
  22019=>"011010010",
  22020=>"001110101",
  22021=>"111111011",
  22022=>"000010010",
  22023=>"100100110",
  22024=>"011000111",
  22025=>"100111110",
  22026=>"000001010",
  22027=>"110111001",
  22028=>"011001100",
  22029=>"110011101",
  22030=>"111110100",
  22031=>"110110011",
  22032=>"011100110",
  22033=>"110000110",
  22034=>"011100010",
  22035=>"010011000",
  22036=>"001110000",
  22037=>"010000010",
  22038=>"010101101",
  22039=>"010101111",
  22040=>"111100111",
  22041=>"010000011",
  22042=>"011010000",
  22043=>"110010000",
  22044=>"010011100",
  22045=>"011100000",
  22046=>"100100111",
  22047=>"111011011",
  22048=>"000011010",
  22049=>"000111111",
  22050=>"001101101",
  22051=>"011000010",
  22052=>"110100001",
  22053=>"100100010",
  22054=>"111010010",
  22055=>"111100111",
  22056=>"010110100",
  22057=>"000001111",
  22058=>"010010110",
  22059=>"110110111",
  22060=>"110111101",
  22061=>"110010100",
  22062=>"000010101",
  22063=>"110000001",
  22064=>"001011011",
  22065=>"110110100",
  22066=>"010001100",
  22067=>"110100101",
  22068=>"011001001",
  22069=>"000111100",
  22070=>"100100010",
  22071=>"001110101",
  22072=>"101010101",
  22073=>"000110111",
  22074=>"110001011",
  22075=>"001000000",
  22076=>"000011101",
  22077=>"111110101",
  22078=>"111001001",
  22079=>"110110001",
  22080=>"111101111",
  22081=>"011010110",
  22082=>"001010000",
  22083=>"110010001",
  22084=>"001110011",
  22085=>"101011011",
  22086=>"100111100",
  22087=>"111000001",
  22088=>"110101001",
  22089=>"001011011",
  22090=>"010101111",
  22091=>"110111000",
  22092=>"011101101",
  22093=>"001101101",
  22094=>"110010100",
  22095=>"000100100",
  22096=>"110111110",
  22097=>"110111010",
  22098=>"100111010",
  22099=>"001110100",
  22100=>"010010101",
  22101=>"111101000",
  22102=>"001110010",
  22103=>"111100011",
  22104=>"001101000",
  22105=>"000010001",
  22106=>"000000001",
  22107=>"000100100",
  22108=>"110011100",
  22109=>"110000010",
  22110=>"011000100",
  22111=>"011001010",
  22112=>"011111101",
  22113=>"100110000",
  22114=>"101001001",
  22115=>"101000001",
  22116=>"100101000",
  22117=>"001000111",
  22118=>"010110101",
  22119=>"111111010",
  22120=>"110100001",
  22121=>"011100110",
  22122=>"011110111",
  22123=>"110101100",
  22124=>"000000100",
  22125=>"000001100",
  22126=>"011101001",
  22127=>"111110011",
  22128=>"010011001",
  22129=>"010111110",
  22130=>"111111110",
  22131=>"011110101",
  22132=>"010010001",
  22133=>"011001010",
  22134=>"011110010",
  22135=>"000010101",
  22136=>"100101010",
  22137=>"010001001",
  22138=>"000100010",
  22139=>"000000010",
  22140=>"110111110",
  22141=>"110001011",
  22142=>"011100110",
  22143=>"100000001",
  22144=>"010111001",
  22145=>"011001100",
  22146=>"110011001",
  22147=>"111001100",
  22148=>"100101001",
  22149=>"010000001",
  22150=>"011001001",
  22151=>"111110101",
  22152=>"000000000",
  22153=>"011000101",
  22154=>"001001010",
  22155=>"000011110",
  22156=>"101001001",
  22157=>"000110101",
  22158=>"000110001",
  22159=>"111010101",
  22160=>"100001001",
  22161=>"111000111",
  22162=>"110111111",
  22163=>"110001000",
  22164=>"111000000",
  22165=>"001001010",
  22166=>"000000110",
  22167=>"111111000",
  22168=>"111101101",
  22169=>"011000010",
  22170=>"101001101",
  22171=>"110101011",
  22172=>"010100101",
  22173=>"111011110",
  22174=>"100111111",
  22175=>"111011110",
  22176=>"000100000",
  22177=>"100111001",
  22178=>"110101111",
  22179=>"100001001",
  22180=>"101011011",
  22181=>"110011001",
  22182=>"000000000",
  22183=>"000110010",
  22184=>"010011111",
  22185=>"101001111",
  22186=>"011010000",
  22187=>"101001001",
  22188=>"000101000",
  22189=>"100111011",
  22190=>"110100011",
  22191=>"011110010",
  22192=>"010100101",
  22193=>"101110101",
  22194=>"000011001",
  22195=>"110111101",
  22196=>"000101111",
  22197=>"011100011",
  22198=>"000110011",
  22199=>"100011111",
  22200=>"101000100",
  22201=>"010010010",
  22202=>"111010111",
  22203=>"010011110",
  22204=>"011111100",
  22205=>"111010101",
  22206=>"000001100",
  22207=>"000101111",
  22208=>"001110010",
  22209=>"111111000",
  22210=>"001111111",
  22211=>"100110000",
  22212=>"100000110",
  22213=>"010111100",
  22214=>"100011101",
  22215=>"000001000",
  22216=>"110101111",
  22217=>"110111100",
  22218=>"111011000",
  22219=>"100010010",
  22220=>"000011000",
  22221=>"101110101",
  22222=>"000000100",
  22223=>"001110010",
  22224=>"111010100",
  22225=>"010101101",
  22226=>"001100000",
  22227=>"101101011",
  22228=>"110111100",
  22229=>"001011000",
  22230=>"100110110",
  22231=>"111000011",
  22232=>"110000101",
  22233=>"100110000",
  22234=>"001111111",
  22235=>"011010011",
  22236=>"011000100",
  22237=>"001010010",
  22238=>"001011101",
  22239=>"001100101",
  22240=>"000000000",
  22241=>"010010010",
  22242=>"111010111",
  22243=>"111010101",
  22244=>"100000110",
  22245=>"111100000",
  22246=>"100010000",
  22247=>"010110000",
  22248=>"011001101",
  22249=>"000011100",
  22250=>"110110011",
  22251=>"001000110",
  22252=>"000000011",
  22253=>"111101000",
  22254=>"001110111",
  22255=>"111001100",
  22256=>"000111110",
  22257=>"010101000",
  22258=>"010111011",
  22259=>"001010110",
  22260=>"101111010",
  22261=>"100110010",
  22262=>"101101110",
  22263=>"101100110",
  22264=>"011000100",
  22265=>"100000100",
  22266=>"010111101",
  22267=>"000000011",
  22268=>"110011010",
  22269=>"010001110",
  22270=>"000101000",
  22271=>"110011111",
  22272=>"000111100",
  22273=>"001100001",
  22274=>"111100111",
  22275=>"101010001",
  22276=>"011001010",
  22277=>"000000010",
  22278=>"010011010",
  22279=>"010100101",
  22280=>"001110000",
  22281=>"000110111",
  22282=>"000110000",
  22283=>"101110001",
  22284=>"111100101",
  22285=>"101001000",
  22286=>"001001011",
  22287=>"000010000",
  22288=>"001101000",
  22289=>"000001011",
  22290=>"101111111",
  22291=>"100010111",
  22292=>"010100001",
  22293=>"011101110",
  22294=>"001100100",
  22295=>"000110000",
  22296=>"010011010",
  22297=>"001010011",
  22298=>"000100100",
  22299=>"001011111",
  22300=>"111110101",
  22301=>"001100100",
  22302=>"000000100",
  22303=>"101011101",
  22304=>"111111111",
  22305=>"100011011",
  22306=>"110101011",
  22307=>"100001011",
  22308=>"000001100",
  22309=>"110011000",
  22310=>"101101011",
  22311=>"001100100",
  22312=>"100110111",
  22313=>"111100001",
  22314=>"000100100",
  22315=>"101011111",
  22316=>"100000000",
  22317=>"000100000",
  22318=>"000101000",
  22319=>"011101010",
  22320=>"000111010",
  22321=>"111000010",
  22322=>"100101100",
  22323=>"111100100",
  22324=>"101001111",
  22325=>"010000001",
  22326=>"000001011",
  22327=>"111110001",
  22328=>"100101010",
  22329=>"101100100",
  22330=>"011001000",
  22331=>"011010001",
  22332=>"001111100",
  22333=>"011100000",
  22334=>"101011111",
  22335=>"101110101",
  22336=>"010000010",
  22337=>"000111100",
  22338=>"010011110",
  22339=>"111100110",
  22340=>"000010100",
  22341=>"010111101",
  22342=>"011111000",
  22343=>"100000011",
  22344=>"000001001",
  22345=>"011110110",
  22346=>"110111000",
  22347=>"010100011",
  22348=>"101011001",
  22349=>"000100001",
  22350=>"000000000",
  22351=>"100110111",
  22352=>"110001101",
  22353=>"100100011",
  22354=>"001000011",
  22355=>"011000101",
  22356=>"101100110",
  22357=>"110000001",
  22358=>"110000001",
  22359=>"100100111",
  22360=>"000001100",
  22361=>"100001111",
  22362=>"110001110",
  22363=>"011001110",
  22364=>"000001101",
  22365=>"100100111",
  22366=>"100100111",
  22367=>"000111101",
  22368=>"011010100",
  22369=>"111110111",
  22370=>"000111010",
  22371=>"011111110",
  22372=>"110000111",
  22373=>"000111100",
  22374=>"000101011",
  22375=>"001100100",
  22376=>"000000011",
  22377=>"010000100",
  22378=>"010011110",
  22379=>"100101100",
  22380=>"000001011",
  22381=>"101111111",
  22382=>"110110001",
  22383=>"110001011",
  22384=>"101110011",
  22385=>"010000001",
  22386=>"001101000",
  22387=>"000001111",
  22388=>"100000001",
  22389=>"011111111",
  22390=>"000101101",
  22391=>"011011101",
  22392=>"000100101",
  22393=>"011001001",
  22394=>"011101110",
  22395=>"000100001",
  22396=>"001000111",
  22397=>"110111010",
  22398=>"000110011",
  22399=>"100110101",
  22400=>"001110100",
  22401=>"001010000",
  22402=>"110000100",
  22403=>"001001001",
  22404=>"101010011",
  22405=>"000001001",
  22406=>"010000101",
  22407=>"010011111",
  22408=>"110100111",
  22409=>"011111110",
  22410=>"110110110",
  22411=>"000001100",
  22412=>"000101110",
  22413=>"111100001",
  22414=>"111111100",
  22415=>"101001000",
  22416=>"000111000",
  22417=>"000100011",
  22418=>"111101010",
  22419=>"000001100",
  22420=>"111010000",
  22421=>"110110111",
  22422=>"110101010",
  22423=>"110000000",
  22424=>"111100110",
  22425=>"111101001",
  22426=>"000100101",
  22427=>"110000000",
  22428=>"100000011",
  22429=>"111110000",
  22430=>"101101110",
  22431=>"000001101",
  22432=>"000000100",
  22433=>"011101011",
  22434=>"100100001",
  22435=>"011100001",
  22436=>"001001101",
  22437=>"010101101",
  22438=>"001111101",
  22439=>"110101111",
  22440=>"000100011",
  22441=>"111000010",
  22442=>"101101111",
  22443=>"000001000",
  22444=>"101111111",
  22445=>"010101110",
  22446=>"011000101",
  22447=>"111100100",
  22448=>"000000100",
  22449=>"110100010",
  22450=>"110100100",
  22451=>"110101011",
  22452=>"011101110",
  22453=>"101001000",
  22454=>"011100101",
  22455=>"000011111",
  22456=>"001000011",
  22457=>"101011110",
  22458=>"101010110",
  22459=>"001101100",
  22460=>"111001000",
  22461=>"011010110",
  22462=>"101101000",
  22463=>"001110000",
  22464=>"010010000",
  22465=>"110111110",
  22466=>"001101001",
  22467=>"110101011",
  22468=>"101001000",
  22469=>"111101110",
  22470=>"000010011",
  22471=>"111111010",
  22472=>"111011011",
  22473=>"001011101",
  22474=>"010010100",
  22475=>"001001111",
  22476=>"010010100",
  22477=>"010100001",
  22478=>"011010010",
  22479=>"011111110",
  22480=>"010000110",
  22481=>"000000001",
  22482=>"000110111",
  22483=>"101101011",
  22484=>"010011100",
  22485=>"101111001",
  22486=>"000011000",
  22487=>"010011101",
  22488=>"001101010",
  22489=>"001100011",
  22490=>"110101100",
  22491=>"110000110",
  22492=>"110010111",
  22493=>"100101100",
  22494=>"101010111",
  22495=>"111000000",
  22496=>"001001100",
  22497=>"010011010",
  22498=>"110110001",
  22499=>"100001010",
  22500=>"100110001",
  22501=>"111101101",
  22502=>"101101100",
  22503=>"001110111",
  22504=>"100101000",
  22505=>"100111111",
  22506=>"000110100",
  22507=>"100100110",
  22508=>"101101001",
  22509=>"100010000",
  22510=>"101011001",
  22511=>"000001011",
  22512=>"100010101",
  22513=>"100010100",
  22514=>"101000110",
  22515=>"010011001",
  22516=>"011010110",
  22517=>"010100111",
  22518=>"100011101",
  22519=>"001111100",
  22520=>"010011001",
  22521=>"000100110",
  22522=>"100001001",
  22523=>"101001000",
  22524=>"100101001",
  22525=>"101000110",
  22526=>"010011001",
  22527=>"011010011",
  22528=>"110111011",
  22529=>"111001100",
  22530=>"010111101",
  22531=>"111111110",
  22532=>"101110000",
  22533=>"110000000",
  22534=>"010000101",
  22535=>"100101100",
  22536=>"011100011",
  22537=>"101000001",
  22538=>"011111111",
  22539=>"011110011",
  22540=>"101011001",
  22541=>"111011000",
  22542=>"101111010",
  22543=>"100111000",
  22544=>"011010101",
  22545=>"100111110",
  22546=>"010110110",
  22547=>"111100001",
  22548=>"111101111",
  22549=>"000100110",
  22550=>"011001101",
  22551=>"110000110",
  22552=>"010000111",
  22553=>"011011011",
  22554=>"010000011",
  22555=>"101010010",
  22556=>"110011101",
  22557=>"001010101",
  22558=>"101010111",
  22559=>"101111000",
  22560=>"010101011",
  22561=>"001110001",
  22562=>"011000001",
  22563=>"000111010",
  22564=>"001100010",
  22565=>"110111100",
  22566=>"101111100",
  22567=>"111111111",
  22568=>"001000110",
  22569=>"100001110",
  22570=>"011000101",
  22571=>"101111010",
  22572=>"101110011",
  22573=>"110101100",
  22574=>"100101011",
  22575=>"010011100",
  22576=>"000111111",
  22577=>"100111001",
  22578=>"010010111",
  22579=>"010010110",
  22580=>"000000010",
  22581=>"111100111",
  22582=>"001100110",
  22583=>"000011010",
  22584=>"101101110",
  22585=>"110110010",
  22586=>"010100011",
  22587=>"001011011",
  22588=>"101000110",
  22589=>"000010000",
  22590=>"000010100",
  22591=>"000001001",
  22592=>"111011000",
  22593=>"000101001",
  22594=>"001111101",
  22595=>"100010010",
  22596=>"100010111",
  22597=>"010000111",
  22598=>"110000110",
  22599=>"101100001",
  22600=>"111010010",
  22601=>"101011001",
  22602=>"110111110",
  22603=>"111100011",
  22604=>"110100110",
  22605=>"011111000",
  22606=>"000100011",
  22607=>"010001100",
  22608=>"011111010",
  22609=>"100101011",
  22610=>"011100111",
  22611=>"101111100",
  22612=>"000011111",
  22613=>"011010111",
  22614=>"010101100",
  22615=>"100101110",
  22616=>"010101001",
  22617=>"111111110",
  22618=>"000111000",
  22619=>"100011001",
  22620=>"101101110",
  22621=>"110101000",
  22622=>"101000011",
  22623=>"111100101",
  22624=>"101110011",
  22625=>"111011010",
  22626=>"000001010",
  22627=>"000100000",
  22628=>"010100010",
  22629=>"001010000",
  22630=>"010111010",
  22631=>"111111010",
  22632=>"110100100",
  22633=>"110101010",
  22634=>"011000000",
  22635=>"111111100",
  22636=>"011000101",
  22637=>"110111110",
  22638=>"110110000",
  22639=>"001100111",
  22640=>"100001000",
  22641=>"011101011",
  22642=>"000000101",
  22643=>"101110111",
  22644=>"000111100",
  22645=>"100001000",
  22646=>"110011110",
  22647=>"001100001",
  22648=>"010010010",
  22649=>"111100100",
  22650=>"100111100",
  22651=>"000100101",
  22652=>"011110000",
  22653=>"101000111",
  22654=>"011010111",
  22655=>"000111011",
  22656=>"011110110",
  22657=>"111011000",
  22658=>"100001001",
  22659=>"010100011",
  22660=>"001100000",
  22661=>"000010001",
  22662=>"011100111",
  22663=>"000111100",
  22664=>"011001111",
  22665=>"000001000",
  22666=>"001001000",
  22667=>"001101011",
  22668=>"010001000",
  22669=>"001010101",
  22670=>"110010100",
  22671=>"010011001",
  22672=>"001000010",
  22673=>"000001001",
  22674=>"010100100",
  22675=>"010010000",
  22676=>"100111001",
  22677=>"011101010",
  22678=>"010000101",
  22679=>"010110001",
  22680=>"110110110",
  22681=>"000111000",
  22682=>"001001000",
  22683=>"101101011",
  22684=>"000111110",
  22685=>"111001011",
  22686=>"010110100",
  22687=>"010001010",
  22688=>"000111101",
  22689=>"011000110",
  22690=>"101010110",
  22691=>"000111000",
  22692=>"001001011",
  22693=>"101100001",
  22694=>"111100000",
  22695=>"101001001",
  22696=>"110101001",
  22697=>"000001010",
  22698=>"000111011",
  22699=>"110010101",
  22700=>"001110101",
  22701=>"100110010",
  22702=>"101111010",
  22703=>"001000001",
  22704=>"101000001",
  22705=>"110001010",
  22706=>"100001100",
  22707=>"111000000",
  22708=>"110011100",
  22709=>"000000010",
  22710=>"111101111",
  22711=>"101110001",
  22712=>"000011010",
  22713=>"001100100",
  22714=>"001110010",
  22715=>"110001100",
  22716=>"111110111",
  22717=>"000001101",
  22718=>"110000010",
  22719=>"101010011",
  22720=>"110010101",
  22721=>"011010111",
  22722=>"001101001",
  22723=>"010110000",
  22724=>"111000000",
  22725=>"000101011",
  22726=>"111111010",
  22727=>"010000000",
  22728=>"101101111",
  22729=>"011110100",
  22730=>"000101011",
  22731=>"000111011",
  22732=>"011001100",
  22733=>"011000011",
  22734=>"010001111",
  22735=>"010100000",
  22736=>"111110000",
  22737=>"010110001",
  22738=>"110010010",
  22739=>"001110000",
  22740=>"111000000",
  22741=>"100011001",
  22742=>"110101011",
  22743=>"101011111",
  22744=>"100111001",
  22745=>"001100001",
  22746=>"111001011",
  22747=>"011010010",
  22748=>"010101111",
  22749=>"001100000",
  22750=>"011101110",
  22751=>"110111110",
  22752=>"000010011",
  22753=>"001011000",
  22754=>"101001011",
  22755=>"110110110",
  22756=>"110000001",
  22757=>"000000010",
  22758=>"100011000",
  22759=>"010110110",
  22760=>"100000101",
  22761=>"100011010",
  22762=>"000101111",
  22763=>"100001111",
  22764=>"100101100",
  22765=>"000010100",
  22766=>"110011111",
  22767=>"001000110",
  22768=>"110101100",
  22769=>"100000001",
  22770=>"000010100",
  22771=>"111100010",
  22772=>"101000000",
  22773=>"100101010",
  22774=>"000100010",
  22775=>"100000100",
  22776=>"111111010",
  22777=>"100100011",
  22778=>"010111111",
  22779=>"100001100",
  22780=>"100000001",
  22781=>"100010001",
  22782=>"000001110",
  22783=>"000101100",
  22784=>"000111110",
  22785=>"100111010",
  22786=>"001000110",
  22787=>"110111111",
  22788=>"001100111",
  22789=>"110110101",
  22790=>"011110001",
  22791=>"100111011",
  22792=>"001110010",
  22793=>"110100001",
  22794=>"110100110",
  22795=>"000101000",
  22796=>"100100010",
  22797=>"111101111",
  22798=>"001011111",
  22799=>"111010111",
  22800=>"100010011",
  22801=>"100011101",
  22802=>"101101011",
  22803=>"100001100",
  22804=>"101110110",
  22805=>"110000011",
  22806=>"000100010",
  22807=>"101000011",
  22808=>"111010111",
  22809=>"111111010",
  22810=>"101011000",
  22811=>"000111010",
  22812=>"111100000",
  22813=>"001001011",
  22814=>"111000011",
  22815=>"001100000",
  22816=>"000011000",
  22817=>"000000000",
  22818=>"010111010",
  22819=>"010000110",
  22820=>"100101011",
  22821=>"000011101",
  22822=>"010110111",
  22823=>"000100001",
  22824=>"100000000",
  22825=>"011100011",
  22826=>"111011000",
  22827=>"100000001",
  22828=>"101101101",
  22829=>"101000000",
  22830=>"010000000",
  22831=>"011010110",
  22832=>"101100010",
  22833=>"011010011",
  22834=>"110000010",
  22835=>"011100010",
  22836=>"001011111",
  22837=>"001011111",
  22838=>"000001011",
  22839=>"011011100",
  22840=>"000100011",
  22841=>"101001110",
  22842=>"011000100",
  22843=>"111000011",
  22844=>"000011000",
  22845=>"010001111",
  22846=>"011011011",
  22847=>"111111000",
  22848=>"001100101",
  22849=>"100100000",
  22850=>"011010000",
  22851=>"010011110",
  22852=>"001011111",
  22853=>"110001101",
  22854=>"011010000",
  22855=>"101011111",
  22856=>"110011111",
  22857=>"101011100",
  22858=>"011101000",
  22859=>"101010001",
  22860=>"111000001",
  22861=>"000111110",
  22862=>"011000100",
  22863=>"100100111",
  22864=>"101111101",
  22865=>"110101000",
  22866=>"000111011",
  22867=>"011011010",
  22868=>"011100100",
  22869=>"101001011",
  22870=>"010001110",
  22871=>"110000110",
  22872=>"010110110",
  22873=>"100110010",
  22874=>"011011110",
  22875=>"110110011",
  22876=>"011100111",
  22877=>"001000000",
  22878=>"101111110",
  22879=>"000001000",
  22880=>"111000010",
  22881=>"001111000",
  22882=>"010010100",
  22883=>"001001111",
  22884=>"010001010",
  22885=>"101001010",
  22886=>"001110000",
  22887=>"100001101",
  22888=>"101011110",
  22889=>"011100011",
  22890=>"101010100",
  22891=>"100010010",
  22892=>"110000000",
  22893=>"000010000",
  22894=>"110101111",
  22895=>"011111111",
  22896=>"111000000",
  22897=>"010000110",
  22898=>"111010111",
  22899=>"000000011",
  22900=>"111100010",
  22901=>"000111001",
  22902=>"001000110",
  22903=>"001001001",
  22904=>"110110011",
  22905=>"111001000",
  22906=>"001111111",
  22907=>"010110111",
  22908=>"000100000",
  22909=>"111010011",
  22910=>"101001100",
  22911=>"111110110",
  22912=>"111000000",
  22913=>"001101010",
  22914=>"010110000",
  22915=>"111111010",
  22916=>"111100010",
  22917=>"001000100",
  22918=>"101111010",
  22919=>"000010000",
  22920=>"000010001",
  22921=>"111110011",
  22922=>"110001010",
  22923=>"010101111",
  22924=>"110111001",
  22925=>"100000100",
  22926=>"001011111",
  22927=>"100000011",
  22928=>"000011101",
  22929=>"110101101",
  22930=>"111011110",
  22931=>"001100100",
  22932=>"100010110",
  22933=>"101100001",
  22934=>"000001010",
  22935=>"111011101",
  22936=>"100111011",
  22937=>"010010100",
  22938=>"100010101",
  22939=>"100000110",
  22940=>"111001111",
  22941=>"000000001",
  22942=>"101100110",
  22943=>"000010001",
  22944=>"110001011",
  22945=>"010000101",
  22946=>"000101000",
  22947=>"101000111",
  22948=>"000001000",
  22949=>"101011010",
  22950=>"111001100",
  22951=>"011111101",
  22952=>"101000001",
  22953=>"010010110",
  22954=>"001001000",
  22955=>"001110000",
  22956=>"001011000",
  22957=>"111100111",
  22958=>"111011100",
  22959=>"111010010",
  22960=>"101110111",
  22961=>"111000101",
  22962=>"000011001",
  22963=>"111110101",
  22964=>"111110011",
  22965=>"001011101",
  22966=>"000011110",
  22967=>"100110101",
  22968=>"000101011",
  22969=>"001101110",
  22970=>"111011101",
  22971=>"100000111",
  22972=>"001101000",
  22973=>"010001000",
  22974=>"111011000",
  22975=>"111110111",
  22976=>"011101110",
  22977=>"100111100",
  22978=>"000100101",
  22979=>"110100010",
  22980=>"110000101",
  22981=>"000110001",
  22982=>"000101000",
  22983=>"000110111",
  22984=>"000001000",
  22985=>"001101101",
  22986=>"110101111",
  22987=>"111111111",
  22988=>"111100101",
  22989=>"010010100",
  22990=>"000001001",
  22991=>"001111100",
  22992=>"010001000",
  22993=>"011000111",
  22994=>"100110011",
  22995=>"101010110",
  22996=>"011001011",
  22997=>"010000011",
  22998=>"010111100",
  22999=>"011111010",
  23000=>"010001101",
  23001=>"111101000",
  23002=>"010000011",
  23003=>"101011000",
  23004=>"111110010",
  23005=>"000100010",
  23006=>"010011110",
  23007=>"000010011",
  23008=>"000100000",
  23009=>"000101100",
  23010=>"000010100",
  23011=>"101000101",
  23012=>"000011000",
  23013=>"110011100",
  23014=>"110111110",
  23015=>"111000101",
  23016=>"001101011",
  23017=>"100101000",
  23018=>"010110101",
  23019=>"001010001",
  23020=>"101100100",
  23021=>"000110001",
  23022=>"010100111",
  23023=>"010011111",
  23024=>"101010110",
  23025=>"111100101",
  23026=>"100100101",
  23027=>"000000000",
  23028=>"101001110",
  23029=>"010010101",
  23030=>"111001001",
  23031=>"110011110",
  23032=>"010100000",
  23033=>"001010000",
  23034=>"011110010",
  23035=>"101111010",
  23036=>"111011000",
  23037=>"010111110",
  23038=>"001000010",
  23039=>"101100110",
  23040=>"111001011",
  23041=>"000011011",
  23042=>"010011011",
  23043=>"010010110",
  23044=>"100001110",
  23045=>"000001111",
  23046=>"000010111",
  23047=>"111000011",
  23048=>"110100101",
  23049=>"111001100",
  23050=>"000011000",
  23051=>"010001011",
  23052=>"011001001",
  23053=>"010101111",
  23054=>"110010010",
  23055=>"001110111",
  23056=>"001010101",
  23057=>"000100011",
  23058=>"010011110",
  23059=>"100110100",
  23060=>"010100010",
  23061=>"011001001",
  23062=>"000011011",
  23063=>"000010100",
  23064=>"111111110",
  23065=>"001011101",
  23066=>"000011000",
  23067=>"001010000",
  23068=>"111101100",
  23069=>"111111001",
  23070=>"001101010",
  23071=>"111111111",
  23072=>"110001101",
  23073=>"001010100",
  23074=>"001100111",
  23075=>"110010101",
  23076=>"110001000",
  23077=>"100110100",
  23078=>"011001010",
  23079=>"100000110",
  23080=>"001011110",
  23081=>"100000101",
  23082=>"110101001",
  23083=>"110101110",
  23084=>"111101000",
  23085=>"100001011",
  23086=>"110000100",
  23087=>"001110000",
  23088=>"011000101",
  23089=>"011011010",
  23090=>"011001011",
  23091=>"000111010",
  23092=>"110011110",
  23093=>"101000100",
  23094=>"110111100",
  23095=>"110101110",
  23096=>"110010101",
  23097=>"100000110",
  23098=>"000100110",
  23099=>"001100011",
  23100=>"001010101",
  23101=>"110111011",
  23102=>"000111000",
  23103=>"011100000",
  23104=>"110011011",
  23105=>"010101010",
  23106=>"001100010",
  23107=>"001010100",
  23108=>"111111011",
  23109=>"111001110",
  23110=>"000010100",
  23111=>"000100011",
  23112=>"010000100",
  23113=>"101001011",
  23114=>"010100000",
  23115=>"000010110",
  23116=>"111000010",
  23117=>"010100100",
  23118=>"101011111",
  23119=>"110010011",
  23120=>"010111000",
  23121=>"000010010",
  23122=>"000011110",
  23123=>"010001010",
  23124=>"011010100",
  23125=>"010100000",
  23126=>"111000000",
  23127=>"000100111",
  23128=>"111110110",
  23129=>"010011010",
  23130=>"100001001",
  23131=>"101000101",
  23132=>"110100001",
  23133=>"100011000",
  23134=>"100111110",
  23135=>"000010110",
  23136=>"010111011",
  23137=>"001110001",
  23138=>"000010000",
  23139=>"010001111",
  23140=>"001001100",
  23141=>"000100001",
  23142=>"111001011",
  23143=>"001111010",
  23144=>"000100101",
  23145=>"000010000",
  23146=>"101110011",
  23147=>"101100010",
  23148=>"111101111",
  23149=>"001000110",
  23150=>"101111110",
  23151=>"110111100",
  23152=>"000000111",
  23153=>"000001111",
  23154=>"110100101",
  23155=>"110100101",
  23156=>"101100101",
  23157=>"001101110",
  23158=>"111000011",
  23159=>"111110101",
  23160=>"111000010",
  23161=>"110111000",
  23162=>"100011010",
  23163=>"001101111",
  23164=>"100110010",
  23165=>"110001010",
  23166=>"110011000",
  23167=>"101010110",
  23168=>"111111111",
  23169=>"110111001",
  23170=>"110100110",
  23171=>"000001101",
  23172=>"100110100",
  23173=>"111010100",
  23174=>"100001000",
  23175=>"001101010",
  23176=>"101110101",
  23177=>"000110110",
  23178=>"111000101",
  23179=>"100000010",
  23180=>"011100111",
  23181=>"110011101",
  23182=>"001110110",
  23183=>"100111101",
  23184=>"010110010",
  23185=>"010111111",
  23186=>"111111100",
  23187=>"000101101",
  23188=>"100001000",
  23189=>"011111001",
  23190=>"111101100",
  23191=>"100001000",
  23192=>"001101010",
  23193=>"010101100",
  23194=>"110111100",
  23195=>"001101011",
  23196=>"001010010",
  23197=>"000011001",
  23198=>"011000001",
  23199=>"100111110",
  23200=>"001010011",
  23201=>"001011011",
  23202=>"010111011",
  23203=>"100010000",
  23204=>"011110111",
  23205=>"011001011",
  23206=>"010101011",
  23207=>"110001101",
  23208=>"110100010",
  23209=>"110000111",
  23210=>"111011101",
  23211=>"010011100",
  23212=>"111111011",
  23213=>"011001000",
  23214=>"110110111",
  23215=>"110000111",
  23216=>"011000111",
  23217=>"011011100",
  23218=>"100000000",
  23219=>"010000101",
  23220=>"000101100",
  23221=>"001110000",
  23222=>"111001101",
  23223=>"110100111",
  23224=>"100011110",
  23225=>"101011111",
  23226=>"001001011",
  23227=>"111000000",
  23228=>"111010001",
  23229=>"010101101",
  23230=>"001000000",
  23231=>"011010010",
  23232=>"010000010",
  23233=>"011001011",
  23234=>"110101000",
  23235=>"110011111",
  23236=>"101011000",
  23237=>"110110100",
  23238=>"110011011",
  23239=>"011001101",
  23240=>"101110011",
  23241=>"000000101",
  23242=>"001000100",
  23243=>"100011111",
  23244=>"101000100",
  23245=>"101011010",
  23246=>"010001100",
  23247=>"010111101",
  23248=>"010000111",
  23249=>"101100011",
  23250=>"011010110",
  23251=>"000001010",
  23252=>"110000001",
  23253=>"101010110",
  23254=>"011010010",
  23255=>"010000011",
  23256=>"001011101",
  23257=>"100101110",
  23258=>"110100111",
  23259=>"100111000",
  23260=>"010101111",
  23261=>"000001010",
  23262=>"010100010",
  23263=>"100000110",
  23264=>"011000000",
  23265=>"000001010",
  23266=>"100111101",
  23267=>"011000111",
  23268=>"010111001",
  23269=>"011101111",
  23270=>"110010110",
  23271=>"011101010",
  23272=>"100101110",
  23273=>"111101101",
  23274=>"101000001",
  23275=>"000101000",
  23276=>"001011010",
  23277=>"101001010",
  23278=>"111000001",
  23279=>"010010110",
  23280=>"010110000",
  23281=>"000100011",
  23282=>"100001000",
  23283=>"100101010",
  23284=>"100001011",
  23285=>"101111111",
  23286=>"000110100",
  23287=>"010100001",
  23288=>"101011000",
  23289=>"110100100",
  23290=>"111000001",
  23291=>"100110000",
  23292=>"100001011",
  23293=>"101001110",
  23294=>"100100010",
  23295=>"110111101",
  23296=>"100101010",
  23297=>"001001011",
  23298=>"011001101",
  23299=>"100000111",
  23300=>"100000100",
  23301=>"110010001",
  23302=>"101010100",
  23303=>"110011110",
  23304=>"011110000",
  23305=>"000100000",
  23306=>"000110100",
  23307=>"010111000",
  23308=>"110110000",
  23309=>"111001001",
  23310=>"110101101",
  23311=>"111100110",
  23312=>"101011011",
  23313=>"101111110",
  23314=>"101110010",
  23315=>"000000100",
  23316=>"000001011",
  23317=>"000001011",
  23318=>"010101011",
  23319=>"110110101",
  23320=>"110111101",
  23321=>"111001001",
  23322=>"000101011",
  23323=>"010101111",
  23324=>"100111011",
  23325=>"101100001",
  23326=>"000001000",
  23327=>"011100110",
  23328=>"000010111",
  23329=>"111000001",
  23330=>"001101000",
  23331=>"001000111",
  23332=>"001101001",
  23333=>"011110111",
  23334=>"001001010",
  23335=>"010010100",
  23336=>"011100101",
  23337=>"110011011",
  23338=>"011000100",
  23339=>"111001111",
  23340=>"011011001",
  23341=>"100110101",
  23342=>"000000100",
  23343=>"010011010",
  23344=>"100001110",
  23345=>"100010111",
  23346=>"111101001",
  23347=>"011111001",
  23348=>"111010110",
  23349=>"111101100",
  23350=>"011010100",
  23351=>"000001011",
  23352=>"100000010",
  23353=>"001010010",
  23354=>"000111110",
  23355=>"111100010",
  23356=>"110111000",
  23357=>"111011111",
  23358=>"011000111",
  23359=>"101111101",
  23360=>"010111110",
  23361=>"101100101",
  23362=>"101001100",
  23363=>"010101010",
  23364=>"110000010",
  23365=>"001001101",
  23366=>"100111001",
  23367=>"100000111",
  23368=>"111101001",
  23369=>"011101100",
  23370=>"100001101",
  23371=>"010100100",
  23372=>"001010101",
  23373=>"001010100",
  23374=>"001001001",
  23375=>"110101111",
  23376=>"001101011",
  23377=>"101000000",
  23378=>"111101111",
  23379=>"100011110",
  23380=>"101100101",
  23381=>"110010111",
  23382=>"100001100",
  23383=>"101001110",
  23384=>"000111011",
  23385=>"010101001",
  23386=>"011111010",
  23387=>"011000101",
  23388=>"001011000",
  23389=>"101010010",
  23390=>"010100011",
  23391=>"010001010",
  23392=>"011010100",
  23393=>"011001101",
  23394=>"010100101",
  23395=>"010110111",
  23396=>"000011000",
  23397=>"000000100",
  23398=>"100011100",
  23399=>"000111001",
  23400=>"001010100",
  23401=>"110111101",
  23402=>"100001001",
  23403=>"001110111",
  23404=>"110000101",
  23405=>"000011011",
  23406=>"000000001",
  23407=>"011001111",
  23408=>"101101010",
  23409=>"100110111",
  23410=>"001001111",
  23411=>"000001000",
  23412=>"100000110",
  23413=>"111111011",
  23414=>"110101001",
  23415=>"000100010",
  23416=>"000010101",
  23417=>"001100010",
  23418=>"100101101",
  23419=>"000011001",
  23420=>"100110011",
  23421=>"010000101",
  23422=>"010010111",
  23423=>"110111101",
  23424=>"011110001",
  23425=>"101001011",
  23426=>"111100110",
  23427=>"000010000",
  23428=>"000110101",
  23429=>"010100000",
  23430=>"010111010",
  23431=>"010001101",
  23432=>"011101001",
  23433=>"110000110",
  23434=>"010100011",
  23435=>"101001001",
  23436=>"101111111",
  23437=>"101000000",
  23438=>"001110100",
  23439=>"011001001",
  23440=>"110110000",
  23441=>"010101100",
  23442=>"010110011",
  23443=>"000100010",
  23444=>"100010000",
  23445=>"100011111",
  23446=>"100100011",
  23447=>"101111100",
  23448=>"111001001",
  23449=>"011011000",
  23450=>"111001011",
  23451=>"111010010",
  23452=>"001000011",
  23453=>"111100110",
  23454=>"000001011",
  23455=>"110101111",
  23456=>"000101100",
  23457=>"011010100",
  23458=>"000011011",
  23459=>"110111001",
  23460=>"011001110",
  23461=>"101101111",
  23462=>"101100110",
  23463=>"001101101",
  23464=>"111100101",
  23465=>"001010000",
  23466=>"100000000",
  23467=>"011100111",
  23468=>"111100010",
  23469=>"101101010",
  23470=>"000100011",
  23471=>"000010011",
  23472=>"001001000",
  23473=>"111111011",
  23474=>"101011001",
  23475=>"000000010",
  23476=>"011010000",
  23477=>"110100101",
  23478=>"010010111",
  23479=>"110110101",
  23480=>"100000010",
  23481=>"110101101",
  23482=>"101110110",
  23483=>"110111101",
  23484=>"001101011",
  23485=>"001010001",
  23486=>"111011101",
  23487=>"001000001",
  23488=>"000000010",
  23489=>"000000001",
  23490=>"110101010",
  23491=>"101000011",
  23492=>"111110110",
  23493=>"111110011",
  23494=>"001110001",
  23495=>"000101011",
  23496=>"010010100",
  23497=>"011011101",
  23498=>"011110000",
  23499=>"111010111",
  23500=>"010110010",
  23501=>"111011101",
  23502=>"000100111",
  23503=>"011010000",
  23504=>"110001101",
  23505=>"110001101",
  23506=>"111100000",
  23507=>"110010000",
  23508=>"010110001",
  23509=>"000001001",
  23510=>"011111010",
  23511=>"000101001",
  23512=>"101010001",
  23513=>"100110001",
  23514=>"111001100",
  23515=>"011000001",
  23516=>"100101111",
  23517=>"100001011",
  23518=>"111010001",
  23519=>"001010000",
  23520=>"001110001",
  23521=>"000001111",
  23522=>"011000000",
  23523=>"001111001",
  23524=>"000010111",
  23525=>"010000000",
  23526=>"100110111",
  23527=>"111000001",
  23528=>"101100100",
  23529=>"101001000",
  23530=>"111100100",
  23531=>"111101010",
  23532=>"111111010",
  23533=>"100001111",
  23534=>"010001000",
  23535=>"010101101",
  23536=>"000011100",
  23537=>"010001111",
  23538=>"100110110",
  23539=>"100011101",
  23540=>"111101111",
  23541=>"100101111",
  23542=>"111000111",
  23543=>"011001001",
  23544=>"101010111",
  23545=>"100001000",
  23546=>"011110000",
  23547=>"111100010",
  23548=>"010110110",
  23549=>"101110000",
  23550=>"010110110",
  23551=>"110011000",
  23552=>"111000001",
  23553=>"000110010",
  23554=>"101100111",
  23555=>"101111000",
  23556=>"000011111",
  23557=>"110100101",
  23558=>"000110110",
  23559=>"011101101",
  23560=>"100000001",
  23561=>"000100010",
  23562=>"111101101",
  23563=>"011011101",
  23564=>"110010011",
  23565=>"110001101",
  23566=>"110000000",
  23567=>"100110100",
  23568=>"011101110",
  23569=>"100100000",
  23570=>"111111111",
  23571=>"010011000",
  23572=>"001000010",
  23573=>"100101101",
  23574=>"010001001",
  23575=>"111010110",
  23576=>"100010101",
  23577=>"011001111",
  23578=>"010111110",
  23579=>"110010010",
  23580=>"111011001",
  23581=>"000010111",
  23582=>"011100110",
  23583=>"011110000",
  23584=>"110111011",
  23585=>"000011100",
  23586=>"001001000",
  23587=>"101111000",
  23588=>"011100001",
  23589=>"100110011",
  23590=>"111001001",
  23591=>"001010010",
  23592=>"010001010",
  23593=>"011001010",
  23594=>"010111100",
  23595=>"001111111",
  23596=>"000100011",
  23597=>"011011111",
  23598=>"101110111",
  23599=>"001011101",
  23600=>"100100111",
  23601=>"011001011",
  23602=>"011011011",
  23603=>"110000101",
  23604=>"110010000",
  23605=>"000111001",
  23606=>"001000111",
  23607=>"000110000",
  23608=>"010111111",
  23609=>"101010100",
  23610=>"011011111",
  23611=>"110101011",
  23612=>"001101101",
  23613=>"100111111",
  23614=>"100010010",
  23615=>"000010010",
  23616=>"010101100",
  23617=>"100000100",
  23618=>"110001111",
  23619=>"111100011",
  23620=>"010110101",
  23621=>"001100100",
  23622=>"111011111",
  23623=>"011110100",
  23624=>"000101111",
  23625=>"101111000",
  23626=>"101001111",
  23627=>"001011110",
  23628=>"111110110",
  23629=>"011101111",
  23630=>"000000011",
  23631=>"111010001",
  23632=>"100111000",
  23633=>"010011000",
  23634=>"000010111",
  23635=>"111100010",
  23636=>"011000100",
  23637=>"101001011",
  23638=>"101111101",
  23639=>"101100001",
  23640=>"101001100",
  23641=>"011101111",
  23642=>"011100011",
  23643=>"101010110",
  23644=>"110111011",
  23645=>"000100001",
  23646=>"000000000",
  23647=>"010101011",
  23648=>"100101001",
  23649=>"110001100",
  23650=>"000010111",
  23651=>"011111000",
  23652=>"111100111",
  23653=>"001100111",
  23654=>"001110001",
  23655=>"100011110",
  23656=>"001111010",
  23657=>"110110011",
  23658=>"010110100",
  23659=>"111100010",
  23660=>"001100110",
  23661=>"011101010",
  23662=>"010100100",
  23663=>"000000000",
  23664=>"111100000",
  23665=>"000010100",
  23666=>"000111110",
  23667=>"110000110",
  23668=>"000111100",
  23669=>"100001010",
  23670=>"001100100",
  23671=>"000111001",
  23672=>"101100000",
  23673=>"011001111",
  23674=>"111010011",
  23675=>"011100100",
  23676=>"111110101",
  23677=>"110110011",
  23678=>"001000111",
  23679=>"001001101",
  23680=>"010110000",
  23681=>"011000100",
  23682=>"001000001",
  23683=>"001101000",
  23684=>"111110011",
  23685=>"011101101",
  23686=>"000110011",
  23687=>"101010111",
  23688=>"001011100",
  23689=>"100001001",
  23690=>"001011011",
  23691=>"011001001",
  23692=>"010011001",
  23693=>"001110100",
  23694=>"101111001",
  23695=>"000111110",
  23696=>"001010110",
  23697=>"100111100",
  23698=>"110111101",
  23699=>"101001101",
  23700=>"010001001",
  23701=>"001111110",
  23702=>"111001100",
  23703=>"101011100",
  23704=>"110010001",
  23705=>"100010100",
  23706=>"100111000",
  23707=>"000000101",
  23708=>"010100011",
  23709=>"010100100",
  23710=>"111100010",
  23711=>"001001010",
  23712=>"010000101",
  23713=>"100111111",
  23714=>"111100001",
  23715=>"010110100",
  23716=>"010010011",
  23717=>"100110110",
  23718=>"110111111",
  23719=>"000001101",
  23720=>"110100010",
  23721=>"001001010",
  23722=>"111110101",
  23723=>"100011010",
  23724=>"111100100",
  23725=>"001110110",
  23726=>"100001000",
  23727=>"000111011",
  23728=>"010011011",
  23729=>"100111001",
  23730=>"010111100",
  23731=>"001000000",
  23732=>"000101101",
  23733=>"011010101",
  23734=>"010001010",
  23735=>"101100110",
  23736=>"001110110",
  23737=>"110101110",
  23738=>"001111010",
  23739=>"001110101",
  23740=>"011010000",
  23741=>"000110010",
  23742=>"001010011",
  23743=>"110110011",
  23744=>"100011001",
  23745=>"000111101",
  23746=>"111001100",
  23747=>"111100101",
  23748=>"101110100",
  23749=>"010010000",
  23750=>"000111001",
  23751=>"001000010",
  23752=>"100110110",
  23753=>"000010010",
  23754=>"001111110",
  23755=>"101110100",
  23756=>"111100101",
  23757=>"011011010",
  23758=>"010001000",
  23759=>"010000000",
  23760=>"101101011",
  23761=>"110011101",
  23762=>"001000001",
  23763=>"000100011",
  23764=>"011110000",
  23765=>"101011001",
  23766=>"100001101",
  23767=>"111111111",
  23768=>"011111000",
  23769=>"001111000",
  23770=>"010001110",
  23771=>"010100100",
  23772=>"110000100",
  23773=>"111010011",
  23774=>"001001101",
  23775=>"100110000",
  23776=>"000111100",
  23777=>"110101011",
  23778=>"010011001",
  23779=>"001111000",
  23780=>"101011010",
  23781=>"000101000",
  23782=>"100011010",
  23783=>"110110100",
  23784=>"011011011",
  23785=>"111110000",
  23786=>"101001001",
  23787=>"011010010",
  23788=>"101111110",
  23789=>"001010001",
  23790=>"001101110",
  23791=>"100010010",
  23792=>"110011000",
  23793=>"010011010",
  23794=>"101000000",
  23795=>"101000100",
  23796=>"101010100",
  23797=>"001000000",
  23798=>"100111111",
  23799=>"110000110",
  23800=>"001010000",
  23801=>"000110000",
  23802=>"110010111",
  23803=>"010010010",
  23804=>"011101010",
  23805=>"010010001",
  23806=>"111111000",
  23807=>"001111000",
  23808=>"110011111",
  23809=>"001010100",
  23810=>"110101110",
  23811=>"101100101",
  23812=>"110100000",
  23813=>"100111000",
  23814=>"111010100",
  23815=>"100100111",
  23816=>"100011010",
  23817=>"110110111",
  23818=>"111000110",
  23819=>"110100000",
  23820=>"001001101",
  23821=>"101000001",
  23822=>"111101000",
  23823=>"000011100",
  23824=>"111011001",
  23825=>"011101001",
  23826=>"001111100",
  23827=>"110010110",
  23828=>"010101000",
  23829=>"000101110",
  23830=>"010100011",
  23831=>"100101011",
  23832=>"011110110",
  23833=>"010001101",
  23834=>"110100000",
  23835=>"011111101",
  23836=>"111110100",
  23837=>"010011000",
  23838=>"000100001",
  23839=>"011111001",
  23840=>"000010110",
  23841=>"110010100",
  23842=>"100100100",
  23843=>"111001110",
  23844=>"010111110",
  23845=>"100001100",
  23846=>"111100001",
  23847=>"001111100",
  23848=>"100001101",
  23849=>"000001000",
  23850=>"001001111",
  23851=>"111111100",
  23852=>"010001010",
  23853=>"001000011",
  23854=>"000110111",
  23855=>"111101100",
  23856=>"110010000",
  23857=>"011100010",
  23858=>"011100111",
  23859=>"101100111",
  23860=>"101101100",
  23861=>"111111011",
  23862=>"000011110",
  23863=>"010100100",
  23864=>"001011100",
  23865=>"011000100",
  23866=>"000101110",
  23867=>"000100110",
  23868=>"101000001",
  23869=>"111111110",
  23870=>"101100011",
  23871=>"110011100",
  23872=>"000110001",
  23873=>"001110111",
  23874=>"111001100",
  23875=>"101111111",
  23876=>"110001110",
  23877=>"100111000",
  23878=>"111001110",
  23879=>"111111000",
  23880=>"101000011",
  23881=>"001110000",
  23882=>"000111000",
  23883=>"001000000",
  23884=>"111100011",
  23885=>"110000010",
  23886=>"101111001",
  23887=>"010000010",
  23888=>"110110100",
  23889=>"001101110",
  23890=>"001111110",
  23891=>"111101010",
  23892=>"011011100",
  23893=>"110010010",
  23894=>"001010111",
  23895=>"101010010",
  23896=>"001000000",
  23897=>"100010101",
  23898=>"000111110",
  23899=>"111010100",
  23900=>"111010011",
  23901=>"000010110",
  23902=>"001000101",
  23903=>"110011100",
  23904=>"100101111",
  23905=>"000001011",
  23906=>"110000100",
  23907=>"110001001",
  23908=>"001101100",
  23909=>"000010100",
  23910=>"100101101",
  23911=>"111110000",
  23912=>"001110000",
  23913=>"110111101",
  23914=>"101000010",
  23915=>"010101111",
  23916=>"001011111",
  23917=>"011111011",
  23918=>"100000100",
  23919=>"100000010",
  23920=>"110101101",
  23921=>"010101010",
  23922=>"001110100",
  23923=>"000101110",
  23924=>"101010111",
  23925=>"000101111",
  23926=>"110011111",
  23927=>"000001010",
  23928=>"000110001",
  23929=>"011100110",
  23930=>"001100111",
  23931=>"010111010",
  23932=>"000000111",
  23933=>"011011011",
  23934=>"000011001",
  23935=>"101011100",
  23936=>"110101111",
  23937=>"100010110",
  23938=>"100001001",
  23939=>"111111110",
  23940=>"110000011",
  23941=>"111100010",
  23942=>"010010101",
  23943=>"100101001",
  23944=>"000000001",
  23945=>"000111110",
  23946=>"011100100",
  23947=>"111010001",
  23948=>"010111101",
  23949=>"101101100",
  23950=>"101110000",
  23951=>"100111101",
  23952=>"000010111",
  23953=>"011001011",
  23954=>"010011100",
  23955=>"110001000",
  23956=>"001011000",
  23957=>"001111000",
  23958=>"110101011",
  23959=>"110000111",
  23960=>"100001100",
  23961=>"000100011",
  23962=>"100101110",
  23963=>"000000000",
  23964=>"110001001",
  23965=>"111010000",
  23966=>"001010010",
  23967=>"010110111",
  23968=>"000011010",
  23969=>"111101000",
  23970=>"110111111",
  23971=>"001001101",
  23972=>"101101000",
  23973=>"101011000",
  23974=>"111101010",
  23975=>"010000101",
  23976=>"101110001",
  23977=>"000100010",
  23978=>"000010011",
  23979=>"101001101",
  23980=>"001111100",
  23981=>"100111010",
  23982=>"000011110",
  23983=>"100001001",
  23984=>"001011000",
  23985=>"010100101",
  23986=>"101111101",
  23987=>"110001010",
  23988=>"111011010",
  23989=>"100000110",
  23990=>"111111111",
  23991=>"001000000",
  23992=>"101010001",
  23993=>"101010001",
  23994=>"101001000",
  23995=>"100001001",
  23996=>"111000110",
  23997=>"110111000",
  23998=>"000111111",
  23999=>"010001000",
  24000=>"010011111",
  24001=>"110111011",
  24002=>"110000001",
  24003=>"010010100",
  24004=>"000010011",
  24005=>"111000010",
  24006=>"001000110",
  24007=>"011001000",
  24008=>"101000011",
  24009=>"010100111",
  24010=>"111011110",
  24011=>"110001010",
  24012=>"000011100",
  24013=>"110011011",
  24014=>"101101010",
  24015=>"010000011",
  24016=>"000111100",
  24017=>"100001110",
  24018=>"100000011",
  24019=>"100110111",
  24020=>"001101111",
  24021=>"101100000",
  24022=>"110001101",
  24023=>"011101000",
  24024=>"001000100",
  24025=>"110111101",
  24026=>"010011001",
  24027=>"010000011",
  24028=>"000010001",
  24029=>"100011101",
  24030=>"101000010",
  24031=>"111100101",
  24032=>"000000010",
  24033=>"100011000",
  24034=>"111110101",
  24035=>"111100101",
  24036=>"000001111",
  24037=>"001001000",
  24038=>"011111101",
  24039=>"101000011",
  24040=>"011101100",
  24041=>"010110111",
  24042=>"010101110",
  24043=>"011101111",
  24044=>"000000000",
  24045=>"010011001",
  24046=>"100110111",
  24047=>"001100101",
  24048=>"001100110",
  24049=>"010001100",
  24050=>"111001010",
  24051=>"010111011",
  24052=>"010111100",
  24053=>"011100011",
  24054=>"111011010",
  24055=>"000101101",
  24056=>"111011100",
  24057=>"101100000",
  24058=>"101011110",
  24059=>"000000111",
  24060=>"000101011",
  24061=>"101000110",
  24062=>"100101100",
  24063=>"111000110",
  24064=>"000010010",
  24065=>"011100101",
  24066=>"110111001",
  24067=>"111001000",
  24068=>"110110010",
  24069=>"100000110",
  24070=>"000000100",
  24071=>"101110000",
  24072=>"011111111",
  24073=>"010101011",
  24074=>"010100101",
  24075=>"000010010",
  24076=>"100000000",
  24077=>"111111111",
  24078=>"001000011",
  24079=>"101001111",
  24080=>"111010000",
  24081=>"101001010",
  24082=>"011100000",
  24083=>"000010100",
  24084=>"011001101",
  24085=>"100100100",
  24086=>"101101011",
  24087=>"001110110",
  24088=>"011100001",
  24089=>"010110101",
  24090=>"111011010",
  24091=>"000100001",
  24092=>"101010110",
  24093=>"100111001",
  24094=>"101101011",
  24095=>"000110100",
  24096=>"001010110",
  24097=>"000000100",
  24098=>"000001101",
  24099=>"010000010",
  24100=>"001101110",
  24101=>"100001011",
  24102=>"011111111",
  24103=>"111101111",
  24104=>"000101101",
  24105=>"111010110",
  24106=>"011000000",
  24107=>"110001001",
  24108=>"111101010",
  24109=>"000101100",
  24110=>"100000001",
  24111=>"001101110",
  24112=>"001011011",
  24113=>"110101001",
  24114=>"010011110",
  24115=>"110100100",
  24116=>"000000001",
  24117=>"110101101",
  24118=>"001010001",
  24119=>"110000000",
  24120=>"111111101",
  24121=>"111101011",
  24122=>"000010001",
  24123=>"100000111",
  24124=>"000000111",
  24125=>"010101101",
  24126=>"001001010",
  24127=>"111001101",
  24128=>"000010110",
  24129=>"001100001",
  24130=>"010000000",
  24131=>"001111010",
  24132=>"000110001",
  24133=>"111101011",
  24134=>"000000110",
  24135=>"111000001",
  24136=>"110100110",
  24137=>"011001001",
  24138=>"101110110",
  24139=>"001011000",
  24140=>"111111010",
  24141=>"001111011",
  24142=>"111011011",
  24143=>"110101111",
  24144=>"100101001",
  24145=>"000000101",
  24146=>"001000110",
  24147=>"010100010",
  24148=>"000101011",
  24149=>"000011101",
  24150=>"001100110",
  24151=>"000101010",
  24152=>"101101001",
  24153=>"110011010",
  24154=>"001110000",
  24155=>"010010010",
  24156=>"011000010",
  24157=>"010001010",
  24158=>"010111000",
  24159=>"001111011",
  24160=>"101100101",
  24161=>"110000011",
  24162=>"110011100",
  24163=>"000000000",
  24164=>"010100010",
  24165=>"110110111",
  24166=>"000101100",
  24167=>"101111100",
  24168=>"000100111",
  24169=>"010010011",
  24170=>"111111010",
  24171=>"100101001",
  24172=>"101100111",
  24173=>"011110110",
  24174=>"101111000",
  24175=>"110100000",
  24176=>"010001110",
  24177=>"000100011",
  24178=>"010101100",
  24179=>"000000101",
  24180=>"010101101",
  24181=>"010000011",
  24182=>"011111100",
  24183=>"010000011",
  24184=>"010111010",
  24185=>"100001011",
  24186=>"010000100",
  24187=>"010110111",
  24188=>"101101010",
  24189=>"001100010",
  24190=>"001110000",
  24191=>"001010110",
  24192=>"111011110",
  24193=>"011100111",
  24194=>"110000100",
  24195=>"101001101",
  24196=>"100000000",
  24197=>"000000000",
  24198=>"111110100",
  24199=>"001111000",
  24200=>"000000110",
  24201=>"101111011",
  24202=>"001011101",
  24203=>"011111100",
  24204=>"111011100",
  24205=>"101001000",
  24206=>"001111000",
  24207=>"101110010",
  24208=>"010000011",
  24209=>"100001111",
  24210=>"101010111",
  24211=>"101100011",
  24212=>"110100011",
  24213=>"100101111",
  24214=>"100100001",
  24215=>"000101010",
  24216=>"111011101",
  24217=>"010111001",
  24218=>"101110110",
  24219=>"111010011",
  24220=>"100000100",
  24221=>"111011001",
  24222=>"000111001",
  24223=>"100110111",
  24224=>"010001100",
  24225=>"001111001",
  24226=>"111001100",
  24227=>"100100110",
  24228=>"101111110",
  24229=>"011010110",
  24230=>"100000100",
  24231=>"111001010",
  24232=>"110111000",
  24233=>"110001001",
  24234=>"001001110",
  24235=>"100010111",
  24236=>"000101100",
  24237=>"011010010",
  24238=>"111001011",
  24239=>"000010000",
  24240=>"001100000",
  24241=>"001100111",
  24242=>"111011001",
  24243=>"011101110",
  24244=>"001010001",
  24245=>"000000100",
  24246=>"111010011",
  24247=>"100011100",
  24248=>"100010100",
  24249=>"011101110",
  24250=>"110111110",
  24251=>"100110000",
  24252=>"010100011",
  24253=>"010101110",
  24254=>"001000000",
  24255=>"111000100",
  24256=>"100011100",
  24257=>"101001000",
  24258=>"011010001",
  24259=>"111011100",
  24260=>"001011010",
  24261=>"011101000",
  24262=>"111000000",
  24263=>"101001111",
  24264=>"110110000",
  24265=>"111010111",
  24266=>"000010110",
  24267=>"011001100",
  24268=>"010101000",
  24269=>"010001010",
  24270=>"000110111",
  24271=>"011110101",
  24272=>"101011011",
  24273=>"110000000",
  24274=>"010001001",
  24275=>"001001011",
  24276=>"100010110",
  24277=>"001100010",
  24278=>"011101001",
  24279=>"010111111",
  24280=>"111001101",
  24281=>"000110001",
  24282=>"011101000",
  24283=>"110000000",
  24284=>"101101001",
  24285=>"111011100",
  24286=>"100101101",
  24287=>"110000111",
  24288=>"001001000",
  24289=>"100101011",
  24290=>"010111001",
  24291=>"011100110",
  24292=>"000010000",
  24293=>"010010111",
  24294=>"010000001",
  24295=>"010000111",
  24296=>"000000000",
  24297=>"110101111",
  24298=>"111011110",
  24299=>"011111000",
  24300=>"111011001",
  24301=>"010111100",
  24302=>"100001001",
  24303=>"001000001",
  24304=>"111111110",
  24305=>"011001111",
  24306=>"011110101",
  24307=>"001010001",
  24308=>"110011000",
  24309=>"110011011",
  24310=>"100101100",
  24311=>"111110000",
  24312=>"000110101",
  24313=>"011101110",
  24314=>"111011110",
  24315=>"010010100",
  24316=>"110101011",
  24317=>"011011000",
  24318=>"011100111",
  24319=>"010011101",
  24320=>"011010000",
  24321=>"110110111",
  24322=>"100111110",
  24323=>"111000000",
  24324=>"110000100",
  24325=>"011101111",
  24326=>"111100010",
  24327=>"101100000",
  24328=>"000100010",
  24329=>"010100010",
  24330=>"001100000",
  24331=>"111100011",
  24332=>"001100010",
  24333=>"000111101",
  24334=>"000111011",
  24335=>"011001111",
  24336=>"101000011",
  24337=>"101010110",
  24338=>"011101101",
  24339=>"001001011",
  24340=>"111000110",
  24341=>"001000100",
  24342=>"011100000",
  24343=>"111001001",
  24344=>"111101011",
  24345=>"000110100",
  24346=>"000010111",
  24347=>"001010101",
  24348=>"010100011",
  24349=>"100001100",
  24350=>"100110010",
  24351=>"111110100",
  24352=>"000111001",
  24353=>"101001001",
  24354=>"111010101",
  24355=>"000101000",
  24356=>"100100101",
  24357=>"000001000",
  24358=>"001010110",
  24359=>"011011110",
  24360=>"101100110",
  24361=>"111010000",
  24362=>"000000111",
  24363=>"110110001",
  24364=>"111111111",
  24365=>"000010001",
  24366=>"001010101",
  24367=>"111101010",
  24368=>"110101101",
  24369=>"011101001",
  24370=>"100011001",
  24371=>"111000001",
  24372=>"001101101",
  24373=>"011001010",
  24374=>"111110111",
  24375=>"000100111",
  24376=>"011011000",
  24377=>"101001010",
  24378=>"010010110",
  24379=>"100101110",
  24380=>"011011000",
  24381=>"100011011",
  24382=>"000010011",
  24383=>"010110101",
  24384=>"000000001",
  24385=>"000001010",
  24386=>"110011011",
  24387=>"001000011",
  24388=>"111010111",
  24389=>"101010111",
  24390=>"011001010",
  24391=>"010000100",
  24392=>"011101110",
  24393=>"100110000",
  24394=>"101111110",
  24395=>"111000111",
  24396=>"000100110",
  24397=>"000000010",
  24398=>"011001101",
  24399=>"001110100",
  24400=>"000000011",
  24401=>"110010100",
  24402=>"101001010",
  24403=>"011001100",
  24404=>"001101110",
  24405=>"111001011",
  24406=>"111000110",
  24407=>"010111001",
  24408=>"101001000",
  24409=>"101101001",
  24410=>"111000000",
  24411=>"110010010",
  24412=>"101110111",
  24413=>"001001010",
  24414=>"010001100",
  24415=>"000000000",
  24416=>"110000000",
  24417=>"110000000",
  24418=>"001000110",
  24419=>"100101010",
  24420=>"011010010",
  24421=>"001001001",
  24422=>"001000110",
  24423=>"000111010",
  24424=>"111000010",
  24425=>"010000110",
  24426=>"000010100",
  24427=>"111000101",
  24428=>"110010010",
  24429=>"001100000",
  24430=>"011011011",
  24431=>"101000110",
  24432=>"111000001",
  24433=>"000110001",
  24434=>"111010010",
  24435=>"100001100",
  24436=>"001010000",
  24437=>"000100010",
  24438=>"110011001",
  24439=>"000111111",
  24440=>"111000011",
  24441=>"101000000",
  24442=>"101100110",
  24443=>"010101111",
  24444=>"011010110",
  24445=>"110000101",
  24446=>"111000011",
  24447=>"010011010",
  24448=>"010101011",
  24449=>"101101111",
  24450=>"101000011",
  24451=>"101110101",
  24452=>"100100011",
  24453=>"011101010",
  24454=>"110100001",
  24455=>"000011001",
  24456=>"111110011",
  24457=>"110000010",
  24458=>"011011001",
  24459=>"111111100",
  24460=>"001001101",
  24461=>"011101101",
  24462=>"010011000",
  24463=>"111100111",
  24464=>"001110111",
  24465=>"001111000",
  24466=>"001000001",
  24467=>"100001001",
  24468=>"100011011",
  24469=>"011011001",
  24470=>"110010110",
  24471=>"000011001",
  24472=>"010000010",
  24473=>"110000111",
  24474=>"101011011",
  24475=>"010000010",
  24476=>"111001101",
  24477=>"010000111",
  24478=>"101110111",
  24479=>"010001010",
  24480=>"010100001",
  24481=>"100111010",
  24482=>"111011000",
  24483=>"010001010",
  24484=>"110011111",
  24485=>"010001101",
  24486=>"001010010",
  24487=>"101111010",
  24488=>"101111111",
  24489=>"111010101",
  24490=>"000111000",
  24491=>"110011000",
  24492=>"001110001",
  24493=>"000000000",
  24494=>"010011110",
  24495=>"011001011",
  24496=>"001010111",
  24497=>"000001010",
  24498=>"000111100",
  24499=>"010010010",
  24500=>"010000011",
  24501=>"001011101",
  24502=>"001100110",
  24503=>"010010010",
  24504=>"100101010",
  24505=>"111101110",
  24506=>"010011000",
  24507=>"001001010",
  24508=>"110111001",
  24509=>"011101110",
  24510=>"010111001",
  24511=>"001000011",
  24512=>"011010100",
  24513=>"001111101",
  24514=>"011000000",
  24515=>"111011110",
  24516=>"111111100",
  24517=>"001011001",
  24518=>"000011011",
  24519=>"111100000",
  24520=>"010101100",
  24521=>"000011000",
  24522=>"000111011",
  24523=>"101001101",
  24524=>"010101000",
  24525=>"000000100",
  24526=>"010000111",
  24527=>"011010000",
  24528=>"010110101",
  24529=>"101110101",
  24530=>"010101001",
  24531=>"010100010",
  24532=>"000011100",
  24533=>"011111101",
  24534=>"000010000",
  24535=>"110100011",
  24536=>"110011111",
  24537=>"000011111",
  24538=>"110110110",
  24539=>"110011110",
  24540=>"110100111",
  24541=>"000110010",
  24542=>"000101100",
  24543=>"100111110",
  24544=>"101101011",
  24545=>"011111111",
  24546=>"110111110",
  24547=>"100100101",
  24548=>"101010100",
  24549=>"100101011",
  24550=>"101110010",
  24551=>"111101010",
  24552=>"111101101",
  24553=>"101011011",
  24554=>"011100010",
  24555=>"011110111",
  24556=>"011101010",
  24557=>"011001111",
  24558=>"110001111",
  24559=>"100000110",
  24560=>"001110110",
  24561=>"010110010",
  24562=>"101001110",
  24563=>"001000000",
  24564=>"110011001",
  24565=>"011100011",
  24566=>"000011000",
  24567=>"100110110",
  24568=>"101110101",
  24569=>"111100010",
  24570=>"010110110",
  24571=>"010110000",
  24572=>"011111111",
  24573=>"110100111",
  24574=>"000011000",
  24575=>"110010010",
  24576=>"101011101",
  24577=>"101010111",
  24578=>"001110010",
  24579=>"010100110",
  24580=>"001011111",
  24581=>"000110000",
  24582=>"111001101",
  24583=>"111101100",
  24584=>"100001001",
  24585=>"000101100",
  24586=>"110001100",
  24587=>"011111111",
  24588=>"111010001",
  24589=>"000011000",
  24590=>"011010110",
  24591=>"111001000",
  24592=>"110010100",
  24593=>"110011101",
  24594=>"000111101",
  24595=>"000000010",
  24596=>"110111101",
  24597=>"001011101",
  24598=>"001010111",
  24599=>"001000011",
  24600=>"000100001",
  24601=>"000010110",
  24602=>"011110010",
  24603=>"100001100",
  24604=>"100010110",
  24605=>"011000001",
  24606=>"011001111",
  24607=>"000011101",
  24608=>"101111101",
  24609=>"000111101",
  24610=>"001101011",
  24611=>"000001011",
  24612=>"110111111",
  24613=>"001110011",
  24614=>"100011111",
  24615=>"000010111",
  24616=>"000010110",
  24617=>"110100111",
  24618=>"111011101",
  24619=>"110101101",
  24620=>"000101000",
  24621=>"100111000",
  24622=>"001110000",
  24623=>"001011000",
  24624=>"011010001",
  24625=>"010110010",
  24626=>"101001111",
  24627=>"011111011",
  24628=>"101101111",
  24629=>"101111001",
  24630=>"010000001",
  24631=>"111001000",
  24632=>"011100001",
  24633=>"011001100",
  24634=>"011100011",
  24635=>"101001010",
  24636=>"000100000",
  24637=>"000000111",
  24638=>"000101111",
  24639=>"001010000",
  24640=>"010000000",
  24641=>"000000000",
  24642=>"101100000",
  24643=>"000010110",
  24644=>"010011000",
  24645=>"000010011",
  24646=>"000010111",
  24647=>"011111000",
  24648=>"010011111",
  24649=>"100101110",
  24650=>"010011101",
  24651=>"110011001",
  24652=>"011101100",
  24653=>"111111111",
  24654=>"010010111",
  24655=>"110001110",
  24656=>"011100111",
  24657=>"000010000",
  24658=>"010000010",
  24659=>"101010101",
  24660=>"100011011",
  24661=>"001011001",
  24662=>"100100001",
  24663=>"110100101",
  24664=>"101010010",
  24665=>"110100110",
  24666=>"001001000",
  24667=>"101100010",
  24668=>"011011000",
  24669=>"001000010",
  24670=>"111011010",
  24671=>"010000011",
  24672=>"100110100",
  24673=>"001011000",
  24674=>"000010110",
  24675=>"110111110",
  24676=>"100010000",
  24677=>"101101111",
  24678=>"100100010",
  24679=>"101000110",
  24680=>"010111011",
  24681=>"001111000",
  24682=>"010011010",
  24683=>"111111001",
  24684=>"000000011",
  24685=>"010100111",
  24686=>"101110111",
  24687=>"010000100",
  24688=>"111101011",
  24689=>"011001001",
  24690=>"011001001",
  24691=>"111000100",
  24692=>"000010101",
  24693=>"101100010",
  24694=>"011001010",
  24695=>"111001001",
  24696=>"101001011",
  24697=>"101010110",
  24698=>"101110110",
  24699=>"000010000",
  24700=>"110100111",
  24701=>"000011100",
  24702=>"101110001",
  24703=>"000010111",
  24704=>"101100011",
  24705=>"010100010",
  24706=>"101111111",
  24707=>"101000100",
  24708=>"001010000",
  24709=>"111001110",
  24710=>"011010111",
  24711=>"110111111",
  24712=>"000000101",
  24713=>"010000000",
  24714=>"110111111",
  24715=>"111011100",
  24716=>"000000010",
  24717=>"101011000",
  24718=>"110011110",
  24719=>"100110011",
  24720=>"100101001",
  24721=>"001101100",
  24722=>"011010111",
  24723=>"101100010",
  24724=>"100011001",
  24725=>"100110101",
  24726=>"001101111",
  24727=>"010111110",
  24728=>"101110111",
  24729=>"110110000",
  24730=>"111001111",
  24731=>"110000100",
  24732=>"111110100",
  24733=>"010111011",
  24734=>"011000011",
  24735=>"111011010",
  24736=>"011010100",
  24737=>"010001100",
  24738=>"010011010",
  24739=>"111000110",
  24740=>"111000001",
  24741=>"011110101",
  24742=>"001110011",
  24743=>"110100000",
  24744=>"110010000",
  24745=>"010010100",
  24746=>"011100001",
  24747=>"010111100",
  24748=>"001011111",
  24749=>"110100100",
  24750=>"001000011",
  24751=>"010010001",
  24752=>"111010101",
  24753=>"101011010",
  24754=>"000001011",
  24755=>"100010001",
  24756=>"000101110",
  24757=>"110110111",
  24758=>"111101111",
  24759=>"100111111",
  24760=>"000011111",
  24761=>"001110100",
  24762=>"101010100",
  24763=>"000000011",
  24764=>"011111110",
  24765=>"011001001",
  24766=>"100011010",
  24767=>"010001111",
  24768=>"010000000",
  24769=>"011001111",
  24770=>"010010010",
  24771=>"100001111",
  24772=>"000000110",
  24773=>"101000011",
  24774=>"000010111",
  24775=>"001001111",
  24776=>"100001100",
  24777=>"101101011",
  24778=>"011111001",
  24779=>"100111101",
  24780=>"001100111",
  24781=>"011000101",
  24782=>"110000010",
  24783=>"110110110",
  24784=>"110000000",
  24785=>"110100110",
  24786=>"000001110",
  24787=>"000010010",
  24788=>"110101001",
  24789=>"010000000",
  24790=>"000100111",
  24791=>"000110010",
  24792=>"101100011",
  24793=>"100010001",
  24794=>"010001100",
  24795=>"000000010",
  24796=>"010001000",
  24797=>"111011001",
  24798=>"111000000",
  24799=>"101101101",
  24800=>"010111000",
  24801=>"010010001",
  24802=>"010011001",
  24803=>"110101100",
  24804=>"001101011",
  24805=>"111001001",
  24806=>"000001010",
  24807=>"010001011",
  24808=>"000100001",
  24809=>"001000100",
  24810=>"111101111",
  24811=>"111011101",
  24812=>"010100101",
  24813=>"110100110",
  24814=>"000010100",
  24815=>"000000100",
  24816=>"111010110",
  24817=>"110101101",
  24818=>"111100111",
  24819=>"110000110",
  24820=>"101001101",
  24821=>"101000001",
  24822=>"011110001",
  24823=>"100111000",
  24824=>"110001110",
  24825=>"001111101",
  24826=>"000111000",
  24827=>"000011010",
  24828=>"010010010",
  24829=>"111100000",
  24830=>"111010111",
  24831=>"001101110",
  24832=>"101110011",
  24833=>"011100101",
  24834=>"111101111",
  24835=>"111001111",
  24836=>"000111110",
  24837=>"001111011",
  24838=>"101100101",
  24839=>"101001100",
  24840=>"101101010",
  24841=>"101100010",
  24842=>"110000111",
  24843=>"101101111",
  24844=>"111001001",
  24845=>"001010001",
  24846=>"101000000",
  24847=>"101001100",
  24848=>"110110100",
  24849=>"000100000",
  24850=>"110000100",
  24851=>"001010010",
  24852=>"100101001",
  24853=>"110000010",
  24854=>"110110000",
  24855=>"100000011",
  24856=>"101010111",
  24857=>"000000100",
  24858=>"110011011",
  24859=>"111011101",
  24860=>"101101110",
  24861=>"011000100",
  24862=>"001011111",
  24863=>"101100000",
  24864=>"110001101",
  24865=>"010001000",
  24866=>"100000111",
  24867=>"111011011",
  24868=>"010110110",
  24869=>"011011000",
  24870=>"110100101",
  24871=>"111010111",
  24872=>"111010100",
  24873=>"110110011",
  24874=>"110101101",
  24875=>"101110110",
  24876=>"001001111",
  24877=>"101101111",
  24878=>"001000000",
  24879=>"010110001",
  24880=>"111011001",
  24881=>"111100011",
  24882=>"111101000",
  24883=>"000001101",
  24884=>"111100011",
  24885=>"010100000",
  24886=>"111100100",
  24887=>"100011110",
  24888=>"111001000",
  24889=>"101001111",
  24890=>"111011101",
  24891=>"000011000",
  24892=>"000111100",
  24893=>"110010011",
  24894=>"101011010",
  24895=>"001101111",
  24896=>"111011010",
  24897=>"010011100",
  24898=>"111011101",
  24899=>"100000000",
  24900=>"110010101",
  24901=>"011010010",
  24902=>"110101011",
  24903=>"001111001",
  24904=>"011001001",
  24905=>"110100000",
  24906=>"000010110",
  24907=>"001000101",
  24908=>"000101101",
  24909=>"111101101",
  24910=>"010111010",
  24911=>"100100000",
  24912=>"100010000",
  24913=>"000111100",
  24914=>"011110001",
  24915=>"000000010",
  24916=>"000100001",
  24917=>"110110101",
  24918=>"010111010",
  24919=>"110001110",
  24920=>"000100010",
  24921=>"011010010",
  24922=>"010101100",
  24923=>"101100100",
  24924=>"000100011",
  24925=>"101011101",
  24926=>"001010010",
  24927=>"111111100",
  24928=>"101100011",
  24929=>"111001001",
  24930=>"010011100",
  24931=>"011000100",
  24932=>"111101100",
  24933=>"111011101",
  24934=>"010110001",
  24935=>"011100111",
  24936=>"111100000",
  24937=>"110101101",
  24938=>"000111101",
  24939=>"001110111",
  24940=>"101011000",
  24941=>"000111100",
  24942=>"111001010",
  24943=>"100001000",
  24944=>"101001000",
  24945=>"100110000",
  24946=>"010110100",
  24947=>"100101010",
  24948=>"110110000",
  24949=>"101000000",
  24950=>"100110010",
  24951=>"111101000",
  24952=>"110011011",
  24953=>"101110010",
  24954=>"110111011",
  24955=>"100111000",
  24956=>"000011010",
  24957=>"110101101",
  24958=>"111100110",
  24959=>"100101001",
  24960=>"110000000",
  24961=>"000111000",
  24962=>"100011111",
  24963=>"011100000",
  24964=>"011111010",
  24965=>"001011100",
  24966=>"110011110",
  24967=>"011110000",
  24968=>"000110000",
  24969=>"000101001",
  24970=>"101011111",
  24971=>"101111100",
  24972=>"010001100",
  24973=>"111100000",
  24974=>"101111110",
  24975=>"010010010",
  24976=>"000001011",
  24977=>"010110010",
  24978=>"101000000",
  24979=>"001110000",
  24980=>"101011000",
  24981=>"001011000",
  24982=>"111010111",
  24983=>"101100100",
  24984=>"010100000",
  24985=>"001000101",
  24986=>"100011011",
  24987=>"000110110",
  24988=>"011000000",
  24989=>"101011101",
  24990=>"111000001",
  24991=>"111111000",
  24992=>"001111001",
  24993=>"111000111",
  24994=>"111111000",
  24995=>"111000110",
  24996=>"100110011",
  24997=>"110010011",
  24998=>"000011110",
  24999=>"010011110",
  25000=>"000100011",
  25001=>"001011110",
  25002=>"010000000",
  25003=>"001000100",
  25004=>"000110010",
  25005=>"100010100",
  25006=>"101001110",
  25007=>"011111101",
  25008=>"101001010",
  25009=>"111010111",
  25010=>"011110001",
  25011=>"111100101",
  25012=>"010100000",
  25013=>"000000100",
  25014=>"000111101",
  25015=>"010111000",
  25016=>"001100100",
  25017=>"000001001",
  25018=>"111110100",
  25019=>"111000010",
  25020=>"011111111",
  25021=>"001101111",
  25022=>"110011100",
  25023=>"101001010",
  25024=>"100000001",
  25025=>"111010110",
  25026=>"010001011",
  25027=>"001100011",
  25028=>"100100110",
  25029=>"000111001",
  25030=>"100110100",
  25031=>"000000000",
  25032=>"111100111",
  25033=>"101001010",
  25034=>"000111000",
  25035=>"000100110",
  25036=>"100100001",
  25037=>"000011110",
  25038=>"011101011",
  25039=>"001110101",
  25040=>"011110000",
  25041=>"011101011",
  25042=>"011100101",
  25043=>"100001001",
  25044=>"011010000",
  25045=>"000010011",
  25046=>"001000001",
  25047=>"001011101",
  25048=>"001000101",
  25049=>"110111101",
  25050=>"100010010",
  25051=>"110000101",
  25052=>"011010110",
  25053=>"010101110",
  25054=>"000001111",
  25055=>"000010011",
  25056=>"001110110",
  25057=>"010100100",
  25058=>"000101111",
  25059=>"100111001",
  25060=>"111100111",
  25061=>"010000000",
  25062=>"001000001",
  25063=>"010101011",
  25064=>"111000000",
  25065=>"111001001",
  25066=>"001000000",
  25067=>"000010111",
  25068=>"001110001",
  25069=>"101000000",
  25070=>"011000000",
  25071=>"110110010",
  25072=>"000000010",
  25073=>"000010010",
  25074=>"001001111",
  25075=>"100111100",
  25076=>"100000110",
  25077=>"110101011",
  25078=>"000101000",
  25079=>"111011000",
  25080=>"111101101",
  25081=>"010010111",
  25082=>"011111011",
  25083=>"110000000",
  25084=>"100111111",
  25085=>"000010011",
  25086=>"111010001",
  25087=>"000000011",
  25088=>"000000000",
  25089=>"101101001",
  25090=>"111110101",
  25091=>"000011010",
  25092=>"101010100",
  25093=>"110000010",
  25094=>"010100000",
  25095=>"100001110",
  25096=>"001010001",
  25097=>"110111110",
  25098=>"010110011",
  25099=>"011011001",
  25100=>"000001000",
  25101=>"000100101",
  25102=>"001000010",
  25103=>"111100100",
  25104=>"011101110",
  25105=>"111101000",
  25106=>"000100010",
  25107=>"001101011",
  25108=>"011111101",
  25109=>"001100100",
  25110=>"111001010",
  25111=>"000101100",
  25112=>"000011010",
  25113=>"101100101",
  25114=>"111111110",
  25115=>"100001100",
  25116=>"010100001",
  25117=>"111001100",
  25118=>"000111101",
  25119=>"010000011",
  25120=>"010110100",
  25121=>"000001110",
  25122=>"010000100",
  25123=>"000010011",
  25124=>"011111110",
  25125=>"010101100",
  25126=>"100001100",
  25127=>"110100111",
  25128=>"101110000",
  25129=>"101101000",
  25130=>"000000100",
  25131=>"110101100",
  25132=>"011110100",
  25133=>"111101010",
  25134=>"110110011",
  25135=>"101001010",
  25136=>"010100011",
  25137=>"000011010",
  25138=>"001111111",
  25139=>"101100111",
  25140=>"111011101",
  25141=>"001111011",
  25142=>"011101110",
  25143=>"001101110",
  25144=>"100010111",
  25145=>"011000100",
  25146=>"110101000",
  25147=>"100001111",
  25148=>"010100111",
  25149=>"000110000",
  25150=>"110011001",
  25151=>"000000000",
  25152=>"111011011",
  25153=>"010010011",
  25154=>"000000010",
  25155=>"111010110",
  25156=>"110100101",
  25157=>"101110000",
  25158=>"010111010",
  25159=>"110010100",
  25160=>"001011010",
  25161=>"011101000",
  25162=>"011101110",
  25163=>"100000010",
  25164=>"110000010",
  25165=>"110101110",
  25166=>"011100010",
  25167=>"001111101",
  25168=>"100010111",
  25169=>"010000001",
  25170=>"000110101",
  25171=>"001101001",
  25172=>"001111001",
  25173=>"001110011",
  25174=>"011110010",
  25175=>"111000101",
  25176=>"000000000",
  25177=>"000101101",
  25178=>"010001100",
  25179=>"100111101",
  25180=>"010110110",
  25181=>"001101011",
  25182=>"010011111",
  25183=>"000111000",
  25184=>"010011110",
  25185=>"100101000",
  25186=>"110110110",
  25187=>"010100100",
  25188=>"001111101",
  25189=>"100001000",
  25190=>"110101000",
  25191=>"010000101",
  25192=>"110000111",
  25193=>"101011010",
  25194=>"010010110",
  25195=>"111100100",
  25196=>"011101111",
  25197=>"000011010",
  25198=>"100001010",
  25199=>"010010110",
  25200=>"100110111",
  25201=>"111100001",
  25202=>"111110010",
  25203=>"010110011",
  25204=>"101010010",
  25205=>"111010010",
  25206=>"111111101",
  25207=>"000011101",
  25208=>"000110000",
  25209=>"111011001",
  25210=>"100000001",
  25211=>"101010100",
  25212=>"010001011",
  25213=>"111110101",
  25214=>"000011100",
  25215=>"011010110",
  25216=>"010111011",
  25217=>"011111001",
  25218=>"100001000",
  25219=>"000110100",
  25220=>"111100101",
  25221=>"101101101",
  25222=>"110110000",
  25223=>"101101110",
  25224=>"000101001",
  25225=>"001111001",
  25226=>"110101101",
  25227=>"110110011",
  25228=>"101101011",
  25229=>"110111100",
  25230=>"010011001",
  25231=>"111001111",
  25232=>"100110101",
  25233=>"111101000",
  25234=>"001010010",
  25235=>"111010100",
  25236=>"010100100",
  25237=>"100011111",
  25238=>"001011101",
  25239=>"001111001",
  25240=>"001101000",
  25241=>"000000100",
  25242=>"100011110",
  25243=>"001110010",
  25244=>"000111110",
  25245=>"100000111",
  25246=>"111110010",
  25247=>"001111000",
  25248=>"101000000",
  25249=>"010111110",
  25250=>"111101010",
  25251=>"010011111",
  25252=>"011100100",
  25253=>"011111001",
  25254=>"010011100",
  25255=>"010100111",
  25256=>"111010101",
  25257=>"010111001",
  25258=>"011000000",
  25259=>"110010011",
  25260=>"111010000",
  25261=>"010101111",
  25262=>"001101010",
  25263=>"001010100",
  25264=>"011000101",
  25265=>"011111111",
  25266=>"010010010",
  25267=>"010010010",
  25268=>"010001101",
  25269=>"010001000",
  25270=>"100100001",
  25271=>"011001001",
  25272=>"011001011",
  25273=>"101001111",
  25274=>"100101011",
  25275=>"100010010",
  25276=>"010010001",
  25277=>"100110110",
  25278=>"101101000",
  25279=>"110010011",
  25280=>"010110000",
  25281=>"111101001",
  25282=>"010100011",
  25283=>"000000010",
  25284=>"001111011",
  25285=>"001011100",
  25286=>"001111000",
  25287=>"000001011",
  25288=>"101001011",
  25289=>"100001100",
  25290=>"111101111",
  25291=>"111001100",
  25292=>"011010011",
  25293=>"110010010",
  25294=>"101111100",
  25295=>"011000010",
  25296=>"111011000",
  25297=>"101001011",
  25298=>"111101100",
  25299=>"100110100",
  25300=>"010111010",
  25301=>"011101101",
  25302=>"110111011",
  25303=>"101000100",
  25304=>"001100001",
  25305=>"000001110",
  25306=>"000100110",
  25307=>"000010001",
  25308=>"110001101",
  25309=>"010101011",
  25310=>"101110100",
  25311=>"000101111",
  25312=>"110100100",
  25313=>"001010100",
  25314=>"000110101",
  25315=>"100100011",
  25316=>"111011001",
  25317=>"110101011",
  25318=>"010101001",
  25319=>"000010100",
  25320=>"100000100",
  25321=>"000001100",
  25322=>"011000011",
  25323=>"101100001",
  25324=>"011001011",
  25325=>"010111111",
  25326=>"110111100",
  25327=>"001100011",
  25328=>"100111101",
  25329=>"100100011",
  25330=>"001000100",
  25331=>"000101011",
  25332=>"111001111",
  25333=>"101000011",
  25334=>"011101101",
  25335=>"110100000",
  25336=>"100111111",
  25337=>"110011111",
  25338=>"010001110",
  25339=>"011111000",
  25340=>"110100000",
  25341=>"001110110",
  25342=>"010100111",
  25343=>"101100001",
  25344=>"000010101",
  25345=>"101111011",
  25346=>"000101000",
  25347=>"110011001",
  25348=>"100100101",
  25349=>"000000001",
  25350=>"010101001",
  25351=>"011111100",
  25352=>"100010100",
  25353=>"101010000",
  25354=>"011110010",
  25355=>"001110001",
  25356=>"111011101",
  25357=>"111110100",
  25358=>"011000100",
  25359=>"100110011",
  25360=>"011111110",
  25361=>"001001100",
  25362=>"001101111",
  25363=>"001000001",
  25364=>"011111000",
  25365=>"001001111",
  25366=>"011010010",
  25367=>"111100000",
  25368=>"100011101",
  25369=>"011000110",
  25370=>"110000111",
  25371=>"010111011",
  25372=>"111111010",
  25373=>"011111011",
  25374=>"010010101",
  25375=>"011100101",
  25376=>"011010001",
  25377=>"101111101",
  25378=>"000011110",
  25379=>"100111000",
  25380=>"001011001",
  25381=>"000101100",
  25382=>"000111110",
  25383=>"010101001",
  25384=>"011010010",
  25385=>"111001001",
  25386=>"100011100",
  25387=>"001111111",
  25388=>"010101011",
  25389=>"010111101",
  25390=>"110001010",
  25391=>"110100110",
  25392=>"100100110",
  25393=>"110101011",
  25394=>"001110000",
  25395=>"000110101",
  25396=>"001010111",
  25397=>"010001100",
  25398=>"101000001",
  25399=>"111111110",
  25400=>"011101000",
  25401=>"110011110",
  25402=>"110101010",
  25403=>"101111111",
  25404=>"111111111",
  25405=>"010000101",
  25406=>"000101000",
  25407=>"010000001",
  25408=>"101001110",
  25409=>"100011111",
  25410=>"001001000",
  25411=>"001001111",
  25412=>"100000010",
  25413=>"011010011",
  25414=>"101010111",
  25415=>"001001000",
  25416=>"010001000",
  25417=>"000100110",
  25418=>"011100111",
  25419=>"011010001",
  25420=>"000101000",
  25421=>"110011111",
  25422=>"011100010",
  25423=>"010101000",
  25424=>"000101011",
  25425=>"100110000",
  25426=>"110110010",
  25427=>"111111111",
  25428=>"111000001",
  25429=>"110100010",
  25430=>"010011100",
  25431=>"001000111",
  25432=>"101110011",
  25433=>"010111110",
  25434=>"100001101",
  25435=>"001001010",
  25436=>"000011100",
  25437=>"001001100",
  25438=>"101100010",
  25439=>"110100001",
  25440=>"000001010",
  25441=>"010000010",
  25442=>"111010010",
  25443=>"111111101",
  25444=>"110101011",
  25445=>"111000000",
  25446=>"010101111",
  25447=>"001100101",
  25448=>"100110110",
  25449=>"111101101",
  25450=>"110101011",
  25451=>"010010001",
  25452=>"110010111",
  25453=>"001001111",
  25454=>"100110100",
  25455=>"000100001",
  25456=>"100111110",
  25457=>"100000110",
  25458=>"010010010",
  25459=>"100001110",
  25460=>"110110100",
  25461=>"010100011",
  25462=>"001110110",
  25463=>"001011000",
  25464=>"101001000",
  25465=>"001001011",
  25466=>"110100111",
  25467=>"110000011",
  25468=>"111110101",
  25469=>"000000000",
  25470=>"110100010",
  25471=>"111110111",
  25472=>"101011111",
  25473=>"101101101",
  25474=>"001010001",
  25475=>"010000011",
  25476=>"001100000",
  25477=>"101101101",
  25478=>"101101100",
  25479=>"011110100",
  25480=>"010110110",
  25481=>"000011000",
  25482=>"000011111",
  25483=>"100000001",
  25484=>"001001011",
  25485=>"100001010",
  25486=>"000101110",
  25487=>"010111111",
  25488=>"011011111",
  25489=>"101100001",
  25490=>"000001000",
  25491=>"111011000",
  25492=>"010010000",
  25493=>"011111101",
  25494=>"000101110",
  25495=>"010110101",
  25496=>"000111011",
  25497=>"111000000",
  25498=>"100000001",
  25499=>"100001011",
  25500=>"000010001",
  25501=>"111111111",
  25502=>"110100000",
  25503=>"110100010",
  25504=>"011110111",
  25505=>"000111101",
  25506=>"100000111",
  25507=>"010001101",
  25508=>"110001111",
  25509=>"100000100",
  25510=>"010011000",
  25511=>"010110001",
  25512=>"110111101",
  25513=>"100010001",
  25514=>"010011001",
  25515=>"101000010",
  25516=>"000100100",
  25517=>"111110101",
  25518=>"110001101",
  25519=>"011110011",
  25520=>"100100110",
  25521=>"110111110",
  25522=>"111000011",
  25523=>"110111111",
  25524=>"101011001",
  25525=>"000010100",
  25526=>"110100010",
  25527=>"111111110",
  25528=>"101101000",
  25529=>"001111011",
  25530=>"111110000",
  25531=>"001111001",
  25532=>"100000100",
  25533=>"001001010",
  25534=>"001010011",
  25535=>"011010011",
  25536=>"100011001",
  25537=>"101010101",
  25538=>"000010111",
  25539=>"100011110",
  25540=>"110011111",
  25541=>"011010000",
  25542=>"111010101",
  25543=>"101111110",
  25544=>"101000000",
  25545=>"110101110",
  25546=>"111011011",
  25547=>"000001100",
  25548=>"101111111",
  25549=>"001000110",
  25550=>"101101011",
  25551=>"110110000",
  25552=>"101100101",
  25553=>"000111010",
  25554=>"110101100",
  25555=>"001000100",
  25556=>"010001010",
  25557=>"111110111",
  25558=>"001100111",
  25559=>"001011111",
  25560=>"111100110",
  25561=>"001000001",
  25562=>"110011011",
  25563=>"111001100",
  25564=>"100000100",
  25565=>"110000111",
  25566=>"011100111",
  25567=>"011000100",
  25568=>"100110001",
  25569=>"110100011",
  25570=>"011110111",
  25571=>"110001000",
  25572=>"001001000",
  25573=>"111111010",
  25574=>"001000111",
  25575=>"001110111",
  25576=>"101111000",
  25577=>"001011001",
  25578=>"110001000",
  25579=>"100000010",
  25580=>"000110101",
  25581=>"100110101",
  25582=>"001010100",
  25583=>"010011000",
  25584=>"011011001",
  25585=>"101001010",
  25586=>"001011100",
  25587=>"001001001",
  25588=>"111101101",
  25589=>"010111010",
  25590=>"001100010",
  25591=>"011110101",
  25592=>"101110001",
  25593=>"001100111",
  25594=>"100000000",
  25595=>"111001001",
  25596=>"010010010",
  25597=>"000101011",
  25598=>"110001000",
  25599=>"110010011",
  25600=>"000101100",
  25601=>"110001100",
  25602=>"001110110",
  25603=>"110110010",
  25604=>"010000111",
  25605=>"100100011",
  25606=>"110111001",
  25607=>"111110000",
  25608=>"011101110",
  25609=>"001111100",
  25610=>"111101000",
  25611=>"001110011",
  25612=>"010010001",
  25613=>"100001001",
  25614=>"101010000",
  25615=>"011010011",
  25616=>"100111111",
  25617=>"001010001",
  25618=>"001111011",
  25619=>"001001111",
  25620=>"000011011",
  25621=>"111101110",
  25622=>"110101001",
  25623=>"001101011",
  25624=>"101000001",
  25625=>"011010101",
  25626=>"010010101",
  25627=>"101011100",
  25628=>"010100101",
  25629=>"010101101",
  25630=>"011101011",
  25631=>"001111111",
  25632=>"010101010",
  25633=>"010110011",
  25634=>"010001011",
  25635=>"110111111",
  25636=>"111101011",
  25637=>"000110011",
  25638=>"010110001",
  25639=>"101101111",
  25640=>"010001110",
  25641=>"111001111",
  25642=>"011110000",
  25643=>"000110000",
  25644=>"110101101",
  25645=>"010010110",
  25646=>"001101101",
  25647=>"001000000",
  25648=>"010001101",
  25649=>"001111000",
  25650=>"101001111",
  25651=>"010001101",
  25652=>"001010100",
  25653=>"000101001",
  25654=>"000100100",
  25655=>"111011010",
  25656=>"111000101",
  25657=>"011010110",
  25658=>"111110100",
  25659=>"100001000",
  25660=>"010111111",
  25661=>"100100111",
  25662=>"111010000",
  25663=>"100100000",
  25664=>"010111010",
  25665=>"001101100",
  25666=>"101000000",
  25667=>"101101100",
  25668=>"111111010",
  25669=>"110101101",
  25670=>"111010011",
  25671=>"110101111",
  25672=>"111100111",
  25673=>"000000011",
  25674=>"000000110",
  25675=>"000001010",
  25676=>"111010000",
  25677=>"101010100",
  25678=>"100010000",
  25679=>"010001011",
  25680=>"001110110",
  25681=>"110011111",
  25682=>"100011100",
  25683=>"000110111",
  25684=>"101001110",
  25685=>"010010011",
  25686=>"000000010",
  25687=>"001000000",
  25688=>"110001000",
  25689=>"000110110",
  25690=>"100011101",
  25691=>"000000000",
  25692=>"000000000",
  25693=>"010010011",
  25694=>"110110100",
  25695=>"011001101",
  25696=>"100001101",
  25697=>"010010011",
  25698=>"000001010",
  25699=>"111011000",
  25700=>"001101000",
  25701=>"011000000",
  25702=>"001111001",
  25703=>"101001000",
  25704=>"010100111",
  25705=>"001000101",
  25706=>"101000101",
  25707=>"010110011",
  25708=>"000100101",
  25709=>"101111111",
  25710=>"100110111",
  25711=>"110000010",
  25712=>"001001100",
  25713=>"110111001",
  25714=>"000001001",
  25715=>"111000011",
  25716=>"000101110",
  25717=>"111011100",
  25718=>"011110001",
  25719=>"100101001",
  25720=>"001111101",
  25721=>"111100101",
  25722=>"001100011",
  25723=>"100110110",
  25724=>"110001100",
  25725=>"110001010",
  25726=>"101110101",
  25727=>"110101010",
  25728=>"000000101",
  25729=>"111111100",
  25730=>"011010011",
  25731=>"010100000",
  25732=>"000000011",
  25733=>"010100010",
  25734=>"111101001",
  25735=>"000111011",
  25736=>"011010001",
  25737=>"101111110",
  25738=>"010011010",
  25739=>"010100101",
  25740=>"111000010",
  25741=>"001010100",
  25742=>"000001000",
  25743=>"111111111",
  25744=>"010011000",
  25745=>"111001000",
  25746=>"011011000",
  25747=>"110010000",
  25748=>"110010100",
  25749=>"111001100",
  25750=>"011101100",
  25751=>"100010001",
  25752=>"100101101",
  25753=>"000110111",
  25754=>"101001001",
  25755=>"011000000",
  25756=>"100111000",
  25757=>"000110010",
  25758=>"100110011",
  25759=>"011110010",
  25760=>"010111100",
  25761=>"110111000",
  25762=>"101011101",
  25763=>"000001000",
  25764=>"001011110",
  25765=>"010001101",
  25766=>"010010011",
  25767=>"001100011",
  25768=>"000001011",
  25769=>"001111101",
  25770=>"000100110",
  25771=>"111101011",
  25772=>"110110100",
  25773=>"100001000",
  25774=>"001100011",
  25775=>"000000011",
  25776=>"110000110",
  25777=>"111010011",
  25778=>"111011101",
  25779=>"011110101",
  25780=>"011000110",
  25781=>"111011000",
  25782=>"101101001",
  25783=>"100100010",
  25784=>"010101111",
  25785=>"011110000",
  25786=>"010010001",
  25787=>"000101100",
  25788=>"111011000",
  25789=>"001111011",
  25790=>"100010111",
  25791=>"100111101",
  25792=>"010111010",
  25793=>"111000101",
  25794=>"000111101",
  25795=>"111110101",
  25796=>"010001001",
  25797=>"011000111",
  25798=>"011101010",
  25799=>"100010101",
  25800=>"000110000",
  25801=>"011000011",
  25802=>"001001011",
  25803=>"001100000",
  25804=>"000101110",
  25805=>"111110000",
  25806=>"000110001",
  25807=>"110101111",
  25808=>"101100100",
  25809=>"111010001",
  25810=>"010010000",
  25811=>"010011110",
  25812=>"000111110",
  25813=>"101110011",
  25814=>"001111010",
  25815=>"101001000",
  25816=>"010111010",
  25817=>"100110001",
  25818=>"001100001",
  25819=>"100011000",
  25820=>"101100110",
  25821=>"000010101",
  25822=>"001101110",
  25823=>"110001000",
  25824=>"110111011",
  25825=>"001100001",
  25826=>"000110111",
  25827=>"110111101",
  25828=>"000011010",
  25829=>"010110000",
  25830=>"010101000",
  25831=>"100101111",
  25832=>"101010111",
  25833=>"001011100",
  25834=>"111101000",
  25835=>"001110110",
  25836=>"000000101",
  25837=>"010111100",
  25838=>"000110010",
  25839=>"100111100",
  25840=>"101101000",
  25841=>"011100010",
  25842=>"101100000",
  25843=>"110010111",
  25844=>"010101110",
  25845=>"011000000",
  25846=>"000000101",
  25847=>"000000001",
  25848=>"010010011",
  25849=>"011100101",
  25850=>"001010110",
  25851=>"000110011",
  25852=>"000100111",
  25853=>"110000101",
  25854=>"000011010",
  25855=>"111001110",
  25856=>"010101010",
  25857=>"100011011",
  25858=>"001110000",
  25859=>"110001001",
  25860=>"001011001",
  25861=>"000011011",
  25862=>"111111001",
  25863=>"110110010",
  25864=>"000110001",
  25865=>"010110111",
  25866=>"111001110",
  25867=>"100001110",
  25868=>"101000100",
  25869=>"111100011",
  25870=>"101001101",
  25871=>"011001010",
  25872=>"100101000",
  25873=>"001100011",
  25874=>"101110001",
  25875=>"011010000",
  25876=>"010001010",
  25877=>"101000110",
  25878=>"001100010",
  25879=>"001111011",
  25880=>"111101100",
  25881=>"010010110",
  25882=>"001011000",
  25883=>"100001001",
  25884=>"000001011",
  25885=>"111011101",
  25886=>"101110001",
  25887=>"100101011",
  25888=>"101101101",
  25889=>"001011111",
  25890=>"010011110",
  25891=>"010110011",
  25892=>"001110011",
  25893=>"010000000",
  25894=>"101001010",
  25895=>"100010000",
  25896=>"111001101",
  25897=>"100000010",
  25898=>"100010000",
  25899=>"111001001",
  25900=>"100101100",
  25901=>"000000100",
  25902=>"010010010",
  25903=>"111111101",
  25904=>"101100111",
  25905=>"011001111",
  25906=>"010010001",
  25907=>"101111110",
  25908=>"101011001",
  25909=>"100001100",
  25910=>"111101101",
  25911=>"110111001",
  25912=>"000000110",
  25913=>"100000111",
  25914=>"111101011",
  25915=>"001100100",
  25916=>"010101010",
  25917=>"010011001",
  25918=>"100001000",
  25919=>"100010101",
  25920=>"000110111",
  25921=>"010111110",
  25922=>"101111010",
  25923=>"011111000",
  25924=>"111001010",
  25925=>"010000100",
  25926=>"000100110",
  25927=>"011001011",
  25928=>"100000000",
  25929=>"110101100",
  25930=>"010111110",
  25931=>"101000000",
  25932=>"010101000",
  25933=>"111100111",
  25934=>"111001110",
  25935=>"111010010",
  25936=>"010000100",
  25937=>"110001001",
  25938=>"000001101",
  25939=>"010110001",
  25940=>"111110101",
  25941=>"000111000",
  25942=>"011110010",
  25943=>"100010100",
  25944=>"000111011",
  25945=>"111101111",
  25946=>"100111110",
  25947=>"000000100",
  25948=>"011001101",
  25949=>"101011011",
  25950=>"111010011",
  25951=>"100111001",
  25952=>"010100011",
  25953=>"011101011",
  25954=>"100010111",
  25955=>"110001011",
  25956=>"000001100",
  25957=>"110000101",
  25958=>"110100100",
  25959=>"100011000",
  25960=>"010100110",
  25961=>"100101101",
  25962=>"000111001",
  25963=>"111011111",
  25964=>"101000011",
  25965=>"010100110",
  25966=>"101010010",
  25967=>"111011000",
  25968=>"101011001",
  25969=>"101111001",
  25970=>"000010001",
  25971=>"001011001",
  25972=>"101110000",
  25973=>"110001101",
  25974=>"111110010",
  25975=>"110011101",
  25976=>"110101011",
  25977=>"110011000",
  25978=>"000100000",
  25979=>"100000001",
  25980=>"011000110",
  25981=>"000111000",
  25982=>"110001010",
  25983=>"000101000",
  25984=>"100100010",
  25985=>"110000000",
  25986=>"100000101",
  25987=>"000100001",
  25988=>"000001100",
  25989=>"000101100",
  25990=>"010111100",
  25991=>"000111001",
  25992=>"110011010",
  25993=>"101101000",
  25994=>"000001101",
  25995=>"001100101",
  25996=>"110110011",
  25997=>"101101010",
  25998=>"011111110",
  25999=>"001101011",
  26000=>"110010010",
  26001=>"000001100",
  26002=>"111001101",
  26003=>"001110100",
  26004=>"101101000",
  26005=>"100010110",
  26006=>"010000010",
  26007=>"100100101",
  26008=>"101110010",
  26009=>"000111101",
  26010=>"001111111",
  26011=>"001000001",
  26012=>"100111101",
  26013=>"000000100",
  26014=>"110111110",
  26015=>"110111000",
  26016=>"001110101",
  26017=>"001110000",
  26018=>"111111000",
  26019=>"101001001",
  26020=>"000001011",
  26021=>"110011010",
  26022=>"000001001",
  26023=>"011101001",
  26024=>"010111100",
  26025=>"101000111",
  26026=>"010001110",
  26027=>"100000111",
  26028=>"011101010",
  26029=>"101111010",
  26030=>"011000101",
  26031=>"010010111",
  26032=>"110110101",
  26033=>"111110111",
  26034=>"010000110",
  26035=>"000101111",
  26036=>"110111010",
  26037=>"111111100",
  26038=>"011110110",
  26039=>"110001101",
  26040=>"011100010",
  26041=>"000010010",
  26042=>"010000000",
  26043=>"010001000",
  26044=>"111101000",
  26045=>"000010101",
  26046=>"001000100",
  26047=>"100111110",
  26048=>"010110001",
  26049=>"001110001",
  26050=>"101011011",
  26051=>"111010111",
  26052=>"111101111",
  26053=>"001001101",
  26054=>"110010000",
  26055=>"111110111",
  26056=>"111111111",
  26057=>"000010000",
  26058=>"110100100",
  26059=>"011101001",
  26060=>"111100100",
  26061=>"011100101",
  26062=>"010011100",
  26063=>"101001011",
  26064=>"100111100",
  26065=>"000110111",
  26066=>"110010110",
  26067=>"100010111",
  26068=>"000111111",
  26069=>"000101111",
  26070=>"001111101",
  26071=>"111110101",
  26072=>"100100000",
  26073=>"011100000",
  26074=>"011000101",
  26075=>"100010011",
  26076=>"111011001",
  26077=>"101110111",
  26078=>"110110110",
  26079=>"001100101",
  26080=>"111001001",
  26081=>"110000101",
  26082=>"110111011",
  26083=>"110000011",
  26084=>"111111000",
  26085=>"010100100",
  26086=>"011000101",
  26087=>"110001001",
  26088=>"001010111",
  26089=>"110011111",
  26090=>"000010011",
  26091=>"001100111",
  26092=>"101100101",
  26093=>"000010010",
  26094=>"000100100",
  26095=>"111111110",
  26096=>"100011000",
  26097=>"110100101",
  26098=>"011011101",
  26099=>"100011111",
  26100=>"001101111",
  26101=>"010111101",
  26102=>"100001100",
  26103=>"010001011",
  26104=>"110110110",
  26105=>"110001001",
  26106=>"101000000",
  26107=>"100001101",
  26108=>"101010010",
  26109=>"111101000",
  26110=>"111000001",
  26111=>"111111011",
  26112=>"001100111",
  26113=>"111110111",
  26114=>"001111111",
  26115=>"111001000",
  26116=>"011111111",
  26117=>"100000001",
  26118=>"011001110",
  26119=>"010101010",
  26120=>"001001100",
  26121=>"001010011",
  26122=>"100000110",
  26123=>"001001110",
  26124=>"100101010",
  26125=>"111111011",
  26126=>"001001010",
  26127=>"011001101",
  26128=>"000110010",
  26129=>"111100111",
  26130=>"111100100",
  26131=>"001000110",
  26132=>"001001000",
  26133=>"011011111",
  26134=>"100001010",
  26135=>"001110110",
  26136=>"011001011",
  26137=>"101100011",
  26138=>"100100101",
  26139=>"010100011",
  26140=>"100001010",
  26141=>"110111010",
  26142=>"010110000",
  26143=>"011010001",
  26144=>"001001111",
  26145=>"010000010",
  26146=>"001111111",
  26147=>"010010000",
  26148=>"101001001",
  26149=>"011100001",
  26150=>"000100011",
  26151=>"010110000",
  26152=>"001010001",
  26153=>"010110001",
  26154=>"011000000",
  26155=>"101100001",
  26156=>"100111111",
  26157=>"010100000",
  26158=>"111010110",
  26159=>"100000101",
  26160=>"111000110",
  26161=>"101000001",
  26162=>"001111111",
  26163=>"001111001",
  26164=>"111011110",
  26165=>"001101111",
  26166=>"110010100",
  26167=>"110010110",
  26168=>"100100000",
  26169=>"111011001",
  26170=>"100100010",
  26171=>"000010111",
  26172=>"000110110",
  26173=>"000011010",
  26174=>"011000011",
  26175=>"011101111",
  26176=>"011011101",
  26177=>"110001110",
  26178=>"000110000",
  26179=>"101010110",
  26180=>"000001000",
  26181=>"101100001",
  26182=>"110000100",
  26183=>"100001111",
  26184=>"000100001",
  26185=>"001101000",
  26186=>"101111100",
  26187=>"000011100",
  26188=>"101101111",
  26189=>"010000010",
  26190=>"000011100",
  26191=>"111111000",
  26192=>"001111001",
  26193=>"101010100",
  26194=>"000110001",
  26195=>"010110111",
  26196=>"001010111",
  26197=>"000000101",
  26198=>"000011011",
  26199=>"100010011",
  26200=>"011011000",
  26201=>"010001010",
  26202=>"000111100",
  26203=>"001001110",
  26204=>"111111001",
  26205=>"110111110",
  26206=>"111111111",
  26207=>"110100111",
  26208=>"001111100",
  26209=>"001110000",
  26210=>"001110010",
  26211=>"000100100",
  26212=>"011100111",
  26213=>"000001100",
  26214=>"010011110",
  26215=>"111011111",
  26216=>"100101000",
  26217=>"001000010",
  26218=>"010011110",
  26219=>"001000101",
  26220=>"001110111",
  26221=>"000100111",
  26222=>"000111101",
  26223=>"101010010",
  26224=>"101000110",
  26225=>"100001101",
  26226=>"011000010",
  26227=>"111111110",
  26228=>"011100111",
  26229=>"011000100",
  26230=>"111111110",
  26231=>"111111111",
  26232=>"001110110",
  26233=>"000000001",
  26234=>"100010000",
  26235=>"100011010",
  26236=>"110011000",
  26237=>"000101010",
  26238=>"111101011",
  26239=>"101010010",
  26240=>"110011111",
  26241=>"000010101",
  26242=>"001011000",
  26243=>"000001001",
  26244=>"010000000",
  26245=>"111001010",
  26246=>"011100111",
  26247=>"100101101",
  26248=>"010110001",
  26249=>"111010011",
  26250=>"010001011",
  26251=>"110110011",
  26252=>"000101011",
  26253=>"110001100",
  26254=>"001000000",
  26255=>"011010011",
  26256=>"101100001",
  26257=>"000011011",
  26258=>"010101001",
  26259=>"101101001",
  26260=>"100101110",
  26261=>"011001011",
  26262=>"001000111",
  26263=>"001011100",
  26264=>"011011001",
  26265=>"011111110",
  26266=>"000110011",
  26267=>"000111011",
  26268=>"001100110",
  26269=>"000011111",
  26270=>"100001110",
  26271=>"001011010",
  26272=>"011100110",
  26273=>"101001110",
  26274=>"100001110",
  26275=>"111101101",
  26276=>"001110000",
  26277=>"001010001",
  26278=>"011010101",
  26279=>"000011001",
  26280=>"111111101",
  26281=>"000101010",
  26282=>"010000110",
  26283=>"110000001",
  26284=>"101100100",
  26285=>"101011001",
  26286=>"111111011",
  26287=>"010010111",
  26288=>"001000010",
  26289=>"010001100",
  26290=>"011000100",
  26291=>"011110101",
  26292=>"001001010",
  26293=>"001101010",
  26294=>"000101101",
  26295=>"101001001",
  26296=>"000000001",
  26297=>"100110001",
  26298=>"010100110",
  26299=>"100101100",
  26300=>"000111001",
  26301=>"111100100",
  26302=>"101001001",
  26303=>"000101000",
  26304=>"001101110",
  26305=>"001000000",
  26306=>"011000011",
  26307=>"001001100",
  26308=>"011010101",
  26309=>"101011111",
  26310=>"111100010",
  26311=>"000000010",
  26312=>"110011010",
  26313=>"111111101",
  26314=>"100000111",
  26315=>"110110010",
  26316=>"110111110",
  26317=>"000101001",
  26318=>"011011001",
  26319=>"110100101",
  26320=>"110001111",
  26321=>"000000100",
  26322=>"011010111",
  26323=>"010000010",
  26324=>"000010011",
  26325=>"110110000",
  26326=>"101100000",
  26327=>"101100110",
  26328=>"101111001",
  26329=>"001000010",
  26330=>"101111110",
  26331=>"011010001",
  26332=>"011111101",
  26333=>"101010011",
  26334=>"110001001",
  26335=>"010011110",
  26336=>"100111011",
  26337=>"100010000",
  26338=>"001101100",
  26339=>"101110011",
  26340=>"101001011",
  26341=>"001100001",
  26342=>"101010000",
  26343=>"011001111",
  26344=>"110101111",
  26345=>"100100111",
  26346=>"100111111",
  26347=>"011011101",
  26348=>"100100101",
  26349=>"011010010",
  26350=>"000111111",
  26351=>"111101001",
  26352=>"101001000",
  26353=>"110111111",
  26354=>"100011000",
  26355=>"111001111",
  26356=>"111001001",
  26357=>"000100001",
  26358=>"110110010",
  26359=>"101000101",
  26360=>"101011101",
  26361=>"010010100",
  26362=>"111010111",
  26363=>"011000111",
  26364=>"110111001",
  26365=>"011100111",
  26366=>"101011000",
  26367=>"010010110",
  26368=>"000001000",
  26369=>"111111001",
  26370=>"101011101",
  26371=>"111011010",
  26372=>"101010111",
  26373=>"011010001",
  26374=>"011110110",
  26375=>"010010010",
  26376=>"111101101",
  26377=>"110111001",
  26378=>"100000000",
  26379=>"110111101",
  26380=>"110010001",
  26381=>"000001100",
  26382=>"000111001",
  26383=>"100110011",
  26384=>"001001100",
  26385=>"100100110",
  26386=>"110010001",
  26387=>"111001100",
  26388=>"101111000",
  26389=>"100010001",
  26390=>"010000111",
  26391=>"110010111",
  26392=>"000101101",
  26393=>"101111110",
  26394=>"101001100",
  26395=>"101110111",
  26396=>"011110111",
  26397=>"010011000",
  26398=>"010001000",
  26399=>"100010001",
  26400=>"101011110",
  26401=>"000100011",
  26402=>"000110000",
  26403=>"001111110",
  26404=>"010010111",
  26405=>"111001011",
  26406=>"011000110",
  26407=>"110011001",
  26408=>"110000100",
  26409=>"111110101",
  26410=>"100000001",
  26411=>"000011101",
  26412=>"000001000",
  26413=>"110011111",
  26414=>"000111010",
  26415=>"101000110",
  26416=>"000000010",
  26417=>"111110111",
  26418=>"011100111",
  26419=>"111110001",
  26420=>"101100110",
  26421=>"110101110",
  26422=>"000101110",
  26423=>"011001100",
  26424=>"111101101",
  26425=>"011110010",
  26426=>"110111001",
  26427=>"011000100",
  26428=>"110000001",
  26429=>"100000010",
  26430=>"010000101",
  26431=>"101011101",
  26432=>"100101000",
  26433=>"111111011",
  26434=>"011111001",
  26435=>"011111011",
  26436=>"100101100",
  26437=>"101110100",
  26438=>"010011111",
  26439=>"000010110",
  26440=>"011011100",
  26441=>"111101101",
  26442=>"101001011",
  26443=>"101010100",
  26444=>"100000010",
  26445=>"010100111",
  26446=>"010011101",
  26447=>"001100101",
  26448=>"111010011",
  26449=>"000000101",
  26450=>"100110110",
  26451=>"111010110",
  26452=>"001111110",
  26453=>"010000001",
  26454=>"011111111",
  26455=>"110111000",
  26456=>"010011111",
  26457=>"101110111",
  26458=>"001101000",
  26459=>"111000000",
  26460=>"111110000",
  26461=>"101110100",
  26462=>"101001001",
  26463=>"010001101",
  26464=>"110101110",
  26465=>"101000010",
  26466=>"111000110",
  26467=>"000000011",
  26468=>"000001100",
  26469=>"111010101",
  26470=>"010001000",
  26471=>"010111011",
  26472=>"000000101",
  26473=>"010011110",
  26474=>"111100110",
  26475=>"000111010",
  26476=>"011000000",
  26477=>"010001010",
  26478=>"101111011",
  26479=>"000010010",
  26480=>"101100111",
  26481=>"011111011",
  26482=>"111111000",
  26483=>"011110000",
  26484=>"010000011",
  26485=>"000111011",
  26486=>"100010010",
  26487=>"000010110",
  26488=>"100100100",
  26489=>"111011010",
  26490=>"001001111",
  26491=>"000011100",
  26492=>"010000100",
  26493=>"110110110",
  26494=>"110111001",
  26495=>"111111011",
  26496=>"010101101",
  26497=>"010110101",
  26498=>"111101110",
  26499=>"010000001",
  26500=>"000000111",
  26501=>"110101101",
  26502=>"010010101",
  26503=>"001011001",
  26504=>"011010100",
  26505=>"011011001",
  26506=>"011000000",
  26507=>"110100011",
  26508=>"101101111",
  26509=>"011111010",
  26510=>"110110011",
  26511=>"010111100",
  26512=>"111011011",
  26513=>"110000101",
  26514=>"010000100",
  26515=>"010100000",
  26516=>"111001110",
  26517=>"101111001",
  26518=>"011001010",
  26519=>"001110000",
  26520=>"110011010",
  26521=>"111100111",
  26522=>"010000110",
  26523=>"101011000",
  26524=>"000111000",
  26525=>"011011100",
  26526=>"011110101",
  26527=>"010110100",
  26528=>"101110110",
  26529=>"000010110",
  26530=>"100101100",
  26531=>"110011000",
  26532=>"010101011",
  26533=>"011011110",
  26534=>"000100011",
  26535=>"110111001",
  26536=>"001110100",
  26537=>"011101100",
  26538=>"001011010",
  26539=>"101100100",
  26540=>"000010001",
  26541=>"011101001",
  26542=>"001101010",
  26543=>"100111000",
  26544=>"111010101",
  26545=>"101111010",
  26546=>"001010000",
  26547=>"111110111",
  26548=>"010101100",
  26549=>"000001010",
  26550=>"110111111",
  26551=>"100111011",
  26552=>"110011110",
  26553=>"110000001",
  26554=>"010101100",
  26555=>"101001110",
  26556=>"000110111",
  26557=>"101101010",
  26558=>"110100000",
  26559=>"000000010",
  26560=>"100000000",
  26561=>"000011111",
  26562=>"000101101",
  26563=>"000111100",
  26564=>"100010000",
  26565=>"111101110",
  26566=>"010011000",
  26567=>"101111110",
  26568=>"000010001",
  26569=>"101110011",
  26570=>"001001011",
  26571=>"011101011",
  26572=>"110011000",
  26573=>"110011101",
  26574=>"111101011",
  26575=>"010111000",
  26576=>"100111111",
  26577=>"010010100",
  26578=>"111111111",
  26579=>"111000000",
  26580=>"000111011",
  26581=>"110101110",
  26582=>"010001100",
  26583=>"010010010",
  26584=>"010101110",
  26585=>"000111111",
  26586=>"110111110",
  26587=>"000001001",
  26588=>"010101100",
  26589=>"101110110",
  26590=>"110010001",
  26591=>"101000100",
  26592=>"100010110",
  26593=>"001000101",
  26594=>"011110000",
  26595=>"000011001",
  26596=>"000000111",
  26597=>"111101101",
  26598=>"001010110",
  26599=>"000000000",
  26600=>"100011110",
  26601=>"100010010",
  26602=>"011100000",
  26603=>"111111000",
  26604=>"110100110",
  26605=>"010000000",
  26606=>"011010000",
  26607=>"100110010",
  26608=>"000000011",
  26609=>"110100100",
  26610=>"111111011",
  26611=>"001110011",
  26612=>"001100001",
  26613=>"110011111",
  26614=>"110100011",
  26615=>"000100000",
  26616=>"100000001",
  26617=>"001111011",
  26618=>"011111010",
  26619=>"000101010",
  26620=>"000011101",
  26621=>"100011001",
  26622=>"101111010",
  26623=>"011011010",
  26624=>"111110101",
  26625=>"111101111",
  26626=>"001000110",
  26627=>"000110011",
  26628=>"001000101",
  26629=>"111101100",
  26630=>"001011001",
  26631=>"011000101",
  26632=>"110000100",
  26633=>"010011001",
  26634=>"000011111",
  26635=>"110000111",
  26636=>"101111100",
  26637=>"001111001",
  26638=>"100110010",
  26639=>"001100101",
  26640=>"011100000",
  26641=>"001001010",
  26642=>"110001111",
  26643=>"000111110",
  26644=>"000111111",
  26645=>"100000000",
  26646=>"000001011",
  26647=>"000011001",
  26648=>"001110100",
  26649=>"000000000",
  26650=>"000001110",
  26651=>"001011111",
  26652=>"111000100",
  26653=>"101001000",
  26654=>"000100011",
  26655=>"011111110",
  26656=>"100110111",
  26657=>"101000001",
  26658=>"110110001",
  26659=>"000001010",
  26660=>"111011010",
  26661=>"001111011",
  26662=>"111011101",
  26663=>"001101001",
  26664=>"101111000",
  26665=>"011110000",
  26666=>"010001011",
  26667=>"010110000",
  26668=>"010111001",
  26669=>"111001111",
  26670=>"101101100",
  26671=>"001011111",
  26672=>"100010000",
  26673=>"010010101",
  26674=>"000111010",
  26675=>"011101111",
  26676=>"011010000",
  26677=>"000010000",
  26678=>"111111111",
  26679=>"010111001",
  26680=>"000010101",
  26681=>"001011001",
  26682=>"010011000",
  26683=>"000000000",
  26684=>"100001010",
  26685=>"111101110",
  26686=>"100000110",
  26687=>"001111000",
  26688=>"011111001",
  26689=>"010001010",
  26690=>"110010010",
  26691=>"110011100",
  26692=>"011010101",
  26693=>"101010000",
  26694=>"001001101",
  26695=>"000101011",
  26696=>"110100000",
  26697=>"000110000",
  26698=>"011101100",
  26699=>"111000101",
  26700=>"000010100",
  26701=>"010110000",
  26702=>"001110001",
  26703=>"101110111",
  26704=>"010000111",
  26705=>"110111010",
  26706=>"101011000",
  26707=>"100000110",
  26708=>"100101011",
  26709=>"100010100",
  26710=>"111001000",
  26711=>"001100100",
  26712=>"000110010",
  26713=>"010111011",
  26714=>"110001110",
  26715=>"100010100",
  26716=>"010001110",
  26717=>"110010010",
  26718=>"110111000",
  26719=>"000000010",
  26720=>"101111001",
  26721=>"010100011",
  26722=>"111011010",
  26723=>"100111111",
  26724=>"110010111",
  26725=>"110000011",
  26726=>"001101110",
  26727=>"110010111",
  26728=>"110011111",
  26729=>"110101011",
  26730=>"111011011",
  26731=>"000000001",
  26732=>"000011100",
  26733=>"111101100",
  26734=>"011111001",
  26735=>"000100110",
  26736=>"111100101",
  26737=>"111100001",
  26738=>"011101010",
  26739=>"100101100",
  26740=>"101011001",
  26741=>"111010110",
  26742=>"011110101",
  26743=>"111011101",
  26744=>"011100110",
  26745=>"101011100",
  26746=>"000110000",
  26747=>"011010111",
  26748=>"011000001",
  26749=>"101001010",
  26750=>"001110110",
  26751=>"110011001",
  26752=>"000000100",
  26753=>"000001110",
  26754=>"000010110",
  26755=>"000011010",
  26756=>"111001100",
  26757=>"001100110",
  26758=>"001110111",
  26759=>"111011101",
  26760=>"110110100",
  26761=>"001000000",
  26762=>"001001101",
  26763=>"001100100",
  26764=>"010010010",
  26765=>"001110101",
  26766=>"100001001",
  26767=>"101011111",
  26768=>"011110000",
  26769=>"100100101",
  26770=>"110011110",
  26771=>"100011010",
  26772=>"010011101",
  26773=>"110100001",
  26774=>"001110011",
  26775=>"000100011",
  26776=>"001101000",
  26777=>"001011100",
  26778=>"100110001",
  26779=>"011101111",
  26780=>"001110111",
  26781=>"100000000",
  26782=>"001101001",
  26783=>"001110101",
  26784=>"100111111",
  26785=>"000000001",
  26786=>"100011000",
  26787=>"010010100",
  26788=>"101101111",
  26789=>"000000111",
  26790=>"011001000",
  26791=>"001001111",
  26792=>"001000001",
  26793=>"111101000",
  26794=>"100001100",
  26795=>"111000011",
  26796=>"010100010",
  26797=>"001101001",
  26798=>"100011100",
  26799=>"111111110",
  26800=>"100100001",
  26801=>"000001100",
  26802=>"110111111",
  26803=>"000010100",
  26804=>"001001001",
  26805=>"000110101",
  26806=>"010000000",
  26807=>"111101111",
  26808=>"110010011",
  26809=>"100110110",
  26810=>"100000001",
  26811=>"011100010",
  26812=>"001010001",
  26813=>"111111010",
  26814=>"000001011",
  26815=>"000000011",
  26816=>"110101111",
  26817=>"110100101",
  26818=>"011001111",
  26819=>"001010000",
  26820=>"001011101",
  26821=>"000111000",
  26822=>"111101000",
  26823=>"000001010",
  26824=>"111110100",
  26825=>"110100111",
  26826=>"010001010",
  26827=>"010110001",
  26828=>"100100000",
  26829=>"010100000",
  26830=>"011101011",
  26831=>"000111101",
  26832=>"011100011",
  26833=>"000010000",
  26834=>"011110111",
  26835=>"010110010",
  26836=>"000101001",
  26837=>"010111001",
  26838=>"010011111",
  26839=>"001101000",
  26840=>"100110100",
  26841=>"010000111",
  26842=>"001011000",
  26843=>"100101110",
  26844=>"011100111",
  26845=>"100111100",
  26846=>"101100001",
  26847=>"001110111",
  26848=>"000000000",
  26849=>"011000011",
  26850=>"010101010",
  26851=>"101010110",
  26852=>"000101101",
  26853=>"011011011",
  26854=>"000001000",
  26855=>"000111001",
  26856=>"100101001",
  26857=>"110011101",
  26858=>"000001100",
  26859=>"000100101",
  26860=>"100011111",
  26861=>"100011100",
  26862=>"110111001",
  26863=>"100000000",
  26864=>"001000010",
  26865=>"000111011",
  26866=>"010000111",
  26867=>"100001001",
  26868=>"010101100",
  26869=>"110001100",
  26870=>"000111101",
  26871=>"110000110",
  26872=>"111110001",
  26873=>"110110010",
  26874=>"101010101",
  26875=>"110100101",
  26876=>"001100000",
  26877=>"001010000",
  26878=>"001110011",
  26879=>"010011101",
  26880=>"011110001",
  26881=>"110010010",
  26882=>"000011000",
  26883=>"001110100",
  26884=>"111110010",
  26885=>"001001000",
  26886=>"111010011",
  26887=>"110100001",
  26888=>"000001000",
  26889=>"011111011",
  26890=>"111110000",
  26891=>"011000110",
  26892=>"101111101",
  26893=>"110111000",
  26894=>"001111110",
  26895=>"100000101",
  26896=>"110111001",
  26897=>"001010000",
  26898=>"011010010",
  26899=>"000000101",
  26900=>"000101110",
  26901=>"001001111",
  26902=>"110101110",
  26903=>"000011001",
  26904=>"001111011",
  26905=>"010010110",
  26906=>"100110110",
  26907=>"011111000",
  26908=>"110111001",
  26909=>"010001010",
  26910=>"111111011",
  26911=>"010111100",
  26912=>"111101000",
  26913=>"110001000",
  26914=>"101111100",
  26915=>"001111011",
  26916=>"111011010",
  26917=>"110011010",
  26918=>"101111111",
  26919=>"010101110",
  26920=>"011011111",
  26921=>"110011100",
  26922=>"001101011",
  26923=>"100111100",
  26924=>"101011110",
  26925=>"010111011",
  26926=>"111101001",
  26927=>"000110000",
  26928=>"111100011",
  26929=>"011011110",
  26930=>"111011111",
  26931=>"010010110",
  26932=>"100100101",
  26933=>"010111100",
  26934=>"110010001",
  26935=>"001001101",
  26936=>"110110011",
  26937=>"111001111",
  26938=>"000000111",
  26939=>"101101100",
  26940=>"101100100",
  26941=>"001001001",
  26942=>"101000111",
  26943=>"111110111",
  26944=>"101111111",
  26945=>"100111011",
  26946=>"010100101",
  26947=>"010101100",
  26948=>"110000010",
  26949=>"110001110",
  26950=>"010110000",
  26951=>"001100100",
  26952=>"111110110",
  26953=>"000101100",
  26954=>"100000101",
  26955=>"001000100",
  26956=>"111101010",
  26957=>"110010101",
  26958=>"011110001",
  26959=>"001010111",
  26960=>"110110101",
  26961=>"011110110",
  26962=>"100101011",
  26963=>"011110000",
  26964=>"000000101",
  26965=>"010111110",
  26966=>"100110101",
  26967=>"100010111",
  26968=>"010000100",
  26969=>"101010000",
  26970=>"110011001",
  26971=>"010100010",
  26972=>"010001100",
  26973=>"111011111",
  26974=>"101001101",
  26975=>"111010111",
  26976=>"000100111",
  26977=>"000011000",
  26978=>"000110000",
  26979=>"110100110",
  26980=>"111001111",
  26981=>"110010110",
  26982=>"000011000",
  26983=>"011111111",
  26984=>"100100100",
  26985=>"000011000",
  26986=>"000001010",
  26987=>"100101011",
  26988=>"110110111",
  26989=>"100100111",
  26990=>"010010001",
  26991=>"101100110",
  26992=>"011001010",
  26993=>"111001000",
  26994=>"101100101",
  26995=>"000110011",
  26996=>"010010010",
  26997=>"011110011",
  26998=>"100000001",
  26999=>"110010101",
  27000=>"101011000",
  27001=>"001000011",
  27002=>"111000110",
  27003=>"100101110",
  27004=>"010100101",
  27005=>"110110001",
  27006=>"111000011",
  27007=>"000000101",
  27008=>"111000000",
  27009=>"100101111",
  27010=>"010110101",
  27011=>"001111000",
  27012=>"100100001",
  27013=>"000111101",
  27014=>"001111101",
  27015=>"101101101",
  27016=>"000000110",
  27017=>"111110011",
  27018=>"001000011",
  27019=>"111111100",
  27020=>"001111000",
  27021=>"010101100",
  27022=>"101010100",
  27023=>"000011001",
  27024=>"100010010",
  27025=>"000000100",
  27026=>"000110000",
  27027=>"000001010",
  27028=>"000100101",
  27029=>"001111100",
  27030=>"001000100",
  27031=>"010100100",
  27032=>"100001000",
  27033=>"101000011",
  27034=>"000111101",
  27035=>"000101001",
  27036=>"000100011",
  27037=>"010010001",
  27038=>"100100011",
  27039=>"101100101",
  27040=>"010101101",
  27041=>"100101100",
  27042=>"010100001",
  27043=>"001010000",
  27044=>"001010101",
  27045=>"001110111",
  27046=>"001011011",
  27047=>"010001101",
  27048=>"110101110",
  27049=>"111101101",
  27050=>"000110011",
  27051=>"011111100",
  27052=>"011001001",
  27053=>"100011100",
  27054=>"011110111",
  27055=>"100001011",
  27056=>"010101000",
  27057=>"101000100",
  27058=>"100011111",
  27059=>"110000100",
  27060=>"001011100",
  27061=>"010101111",
  27062=>"001011101",
  27063=>"010010110",
  27064=>"110110000",
  27065=>"100011010",
  27066=>"000000011",
  27067=>"111101000",
  27068=>"000101010",
  27069=>"100101000",
  27070=>"000011010",
  27071=>"100101000",
  27072=>"010100101",
  27073=>"010000101",
  27074=>"101111010",
  27075=>"001100110",
  27076=>"101010100",
  27077=>"111111101",
  27078=>"010010101",
  27079=>"001111000",
  27080=>"100100011",
  27081=>"001111011",
  27082=>"111001001",
  27083=>"011101111",
  27084=>"001100101",
  27085=>"111000100",
  27086=>"100101011",
  27087=>"011001110",
  27088=>"011100001",
  27089=>"100110001",
  27090=>"011011111",
  27091=>"111010101",
  27092=>"110010010",
  27093=>"001000000",
  27094=>"111101001",
  27095=>"101101110",
  27096=>"111100011",
  27097=>"000011001",
  27098=>"000110101",
  27099=>"001100100",
  27100=>"110100110",
  27101=>"110110100",
  27102=>"011001100",
  27103=>"110001011",
  27104=>"010000011",
  27105=>"011001100",
  27106=>"110101100",
  27107=>"110010011",
  27108=>"001100100",
  27109=>"111100101",
  27110=>"011100110",
  27111=>"101000100",
  27112=>"001111101",
  27113=>"011001110",
  27114=>"010011111",
  27115=>"110100111",
  27116=>"011011111",
  27117=>"110001111",
  27118=>"100110110",
  27119=>"101111110",
  27120=>"011111111",
  27121=>"101000111",
  27122=>"010111101",
  27123=>"011000001",
  27124=>"001001101",
  27125=>"101111000",
  27126=>"001101110",
  27127=>"100100000",
  27128=>"001110111",
  27129=>"010000001",
  27130=>"010100000",
  27131=>"011111111",
  27132=>"100100011",
  27133=>"010000101",
  27134=>"100001101",
  27135=>"100101111",
  27136=>"011100001",
  27137=>"111110111",
  27138=>"110100110",
  27139=>"110110110",
  27140=>"001010010",
  27141=>"011010000",
  27142=>"101010000",
  27143=>"001110110",
  27144=>"011010000",
  27145=>"100101101",
  27146=>"001011000",
  27147=>"011010010",
  27148=>"100111011",
  27149=>"101000111",
  27150=>"100101010",
  27151=>"010100110",
  27152=>"110001010",
  27153=>"010000001",
  27154=>"100011010",
  27155=>"111101010",
  27156=>"110101100",
  27157=>"000101111",
  27158=>"100111110",
  27159=>"111100100",
  27160=>"000101110",
  27161=>"011111110",
  27162=>"000001011",
  27163=>"010100001",
  27164=>"110010100",
  27165=>"101010001",
  27166=>"100110001",
  27167=>"000100000",
  27168=>"101011001",
  27169=>"001101011",
  27170=>"111100111",
  27171=>"101010100",
  27172=>"110000100",
  27173=>"100010110",
  27174=>"000000000",
  27175=>"010011010",
  27176=>"110010010",
  27177=>"010110101",
  27178=>"101110000",
  27179=>"001001000",
  27180=>"101011001",
  27181=>"111010111",
  27182=>"101000010",
  27183=>"011010010",
  27184=>"100100000",
  27185=>"100110001",
  27186=>"110010000",
  27187=>"110100110",
  27188=>"001011101",
  27189=>"110000110",
  27190=>"000000001",
  27191=>"101110111",
  27192=>"000000010",
  27193=>"000011111",
  27194=>"000010111",
  27195=>"100111111",
  27196=>"101110101",
  27197=>"011001000",
  27198=>"011001100",
  27199=>"100100011",
  27200=>"010011111",
  27201=>"011101010",
  27202=>"000100010",
  27203=>"111110101",
  27204=>"010000011",
  27205=>"100001111",
  27206=>"101001101",
  27207=>"010110110",
  27208=>"111111000",
  27209=>"001000100",
  27210=>"001001111",
  27211=>"011010000",
  27212=>"110011101",
  27213=>"010000100",
  27214=>"011001111",
  27215=>"100001001",
  27216=>"101101100",
  27217=>"001101111",
  27218=>"101001001",
  27219=>"010100100",
  27220=>"100101100",
  27221=>"010001110",
  27222=>"100001100",
  27223=>"110000001",
  27224=>"010010111",
  27225=>"111111001",
  27226=>"011001100",
  27227=>"000000000",
  27228=>"000000111",
  27229=>"001000010",
  27230=>"101011110",
  27231=>"001111010",
  27232=>"000110000",
  27233=>"000010001",
  27234=>"001001001",
  27235=>"100011001",
  27236=>"011101101",
  27237=>"011010111",
  27238=>"111010111",
  27239=>"110000000",
  27240=>"100101100",
  27241=>"000011101",
  27242=>"010100011",
  27243=>"011011000",
  27244=>"100010100",
  27245=>"000000100",
  27246=>"000101111",
  27247=>"001110101",
  27248=>"011001100",
  27249=>"010110111",
  27250=>"101011001",
  27251=>"100000010",
  27252=>"110111010",
  27253=>"001001011",
  27254=>"011001000",
  27255=>"111101101",
  27256=>"011010011",
  27257=>"010111000",
  27258=>"000011010",
  27259=>"111111001",
  27260=>"100001001",
  27261=>"000011100",
  27262=>"101100010",
  27263=>"000011000",
  27264=>"100011010",
  27265=>"101000011",
  27266=>"000101000",
  27267=>"100001000",
  27268=>"101010010",
  27269=>"011110001",
  27270=>"111000000",
  27271=>"010011010",
  27272=>"111001100",
  27273=>"001100101",
  27274=>"010011110",
  27275=>"100111100",
  27276=>"010111001",
  27277=>"110011011",
  27278=>"111001000",
  27279=>"000010001",
  27280=>"011001100",
  27281=>"100000101",
  27282=>"100100110",
  27283=>"100110000",
  27284=>"111000010",
  27285=>"001011010",
  27286=>"000100010",
  27287=>"010110011",
  27288=>"000111011",
  27289=>"010101111",
  27290=>"110000010",
  27291=>"000110100",
  27292=>"001111001",
  27293=>"111111011",
  27294=>"000000000",
  27295=>"110101100",
  27296=>"001001110",
  27297=>"100000001",
  27298=>"111111000",
  27299=>"110001000",
  27300=>"101001001",
  27301=>"111000001",
  27302=>"101111001",
  27303=>"100101101",
  27304=>"100001100",
  27305=>"100000010",
  27306=>"100101001",
  27307=>"111010100",
  27308=>"111011011",
  27309=>"111111100",
  27310=>"000000011",
  27311=>"110101111",
  27312=>"000010010",
  27313=>"000010011",
  27314=>"010000000",
  27315=>"011111001",
  27316=>"000110010",
  27317=>"100001100",
  27318=>"111110000",
  27319=>"010100101",
  27320=>"111101101",
  27321=>"100011111",
  27322=>"110001110",
  27323=>"110101110",
  27324=>"000101101",
  27325=>"101000000",
  27326=>"001000101",
  27327=>"100111100",
  27328=>"101010100",
  27329=>"011001011",
  27330=>"100000000",
  27331=>"011111011",
  27332=>"111111101",
  27333=>"101001000",
  27334=>"110100010",
  27335=>"000110101",
  27336=>"001010000",
  27337=>"110000000",
  27338=>"011001111",
  27339=>"100100011",
  27340=>"000001100",
  27341=>"111100100",
  27342=>"110011001",
  27343=>"111110100",
  27344=>"110111110",
  27345=>"100010100",
  27346=>"110101110",
  27347=>"100010011",
  27348=>"000000110",
  27349=>"010001011",
  27350=>"110011101",
  27351=>"100011101",
  27352=>"000001100",
  27353=>"001001111",
  27354=>"000010000",
  27355=>"101110011",
  27356=>"100111010",
  27357=>"000010010",
  27358=>"100001111",
  27359=>"010110011",
  27360=>"001010110",
  27361=>"110011011",
  27362=>"111001010",
  27363=>"100111101",
  27364=>"100010011",
  27365=>"110110000",
  27366=>"110011000",
  27367=>"101011000",
  27368=>"010001101",
  27369=>"010000101",
  27370=>"111011011",
  27371=>"101000001",
  27372=>"000110011",
  27373=>"000001110",
  27374=>"010100000",
  27375=>"101100101",
  27376=>"001100110",
  27377=>"101110101",
  27378=>"111010001",
  27379=>"101100000",
  27380=>"100111111",
  27381=>"011111101",
  27382=>"010100111",
  27383=>"101010000",
  27384=>"000101101",
  27385=>"111010001",
  27386=>"000010010",
  27387=>"000000101",
  27388=>"011000100",
  27389=>"011100011",
  27390=>"110101010",
  27391=>"100010011",
  27392=>"100000011",
  27393=>"001100001",
  27394=>"000000110",
  27395=>"001011111",
  27396=>"101101000",
  27397=>"110011000",
  27398=>"101111111",
  27399=>"111001101",
  27400=>"000101001",
  27401=>"111100100",
  27402=>"111000001",
  27403=>"101110000",
  27404=>"110011011",
  27405=>"011101110",
  27406=>"111111010",
  27407=>"011010010",
  27408=>"001010011",
  27409=>"100000110",
  27410=>"110000011",
  27411=>"101001100",
  27412=>"000000110",
  27413=>"010100110",
  27414=>"110000010",
  27415=>"001100011",
  27416=>"010101010",
  27417=>"001100111",
  27418=>"100001101",
  27419=>"001111111",
  27420=>"000111011",
  27421=>"101001110",
  27422=>"010010001",
  27423=>"100111101",
  27424=>"100111000",
  27425=>"001001010",
  27426=>"111110001",
  27427=>"100011100",
  27428=>"111111110",
  27429=>"110100111",
  27430=>"011010101",
  27431=>"100000011",
  27432=>"011010010",
  27433=>"001011001",
  27434=>"000011100",
  27435=>"101101010",
  27436=>"000010000",
  27437=>"000010110",
  27438=>"111101110",
  27439=>"001000111",
  27440=>"101010001",
  27441=>"011010100",
  27442=>"110010001",
  27443=>"010011011",
  27444=>"001101111",
  27445=>"101111101",
  27446=>"000111011",
  27447=>"010101100",
  27448=>"111000000",
  27449=>"100000010",
  27450=>"011111011",
  27451=>"101100101",
  27452=>"001001000",
  27453=>"101110000",
  27454=>"010110011",
  27455=>"000110110",
  27456=>"001111011",
  27457=>"100001011",
  27458=>"100111111",
  27459=>"100010000",
  27460=>"101101000",
  27461=>"101000110",
  27462=>"101000000",
  27463=>"111101101",
  27464=>"100101111",
  27465=>"010001010",
  27466=>"001111111",
  27467=>"001010010",
  27468=>"100001000",
  27469=>"010000000",
  27470=>"100001001",
  27471=>"011101110",
  27472=>"101010010",
  27473=>"001110110",
  27474=>"101101000",
  27475=>"010010111",
  27476=>"011110010",
  27477=>"010111000",
  27478=>"010010101",
  27479=>"100110100",
  27480=>"110100010",
  27481=>"011000100",
  27482=>"111110110",
  27483=>"000000101",
  27484=>"111101001",
  27485=>"010011001",
  27486=>"011111000",
  27487=>"101111111",
  27488=>"100010111",
  27489=>"010000010",
  27490=>"001101011",
  27491=>"101011100",
  27492=>"010000011",
  27493=>"110101000",
  27494=>"011100000",
  27495=>"010100101",
  27496=>"010100001",
  27497=>"010011011",
  27498=>"000010101",
  27499=>"101101001",
  27500=>"000001100",
  27501=>"010110011",
  27502=>"111010001",
  27503=>"001010011",
  27504=>"110001001",
  27505=>"111100011",
  27506=>"101001100",
  27507=>"101011101",
  27508=>"101010001",
  27509=>"010000100",
  27510=>"000101110",
  27511=>"000101000",
  27512=>"110110100",
  27513=>"101010110",
  27514=>"001000101",
  27515=>"010010000",
  27516=>"011111101",
  27517=>"010010001",
  27518=>"111111110",
  27519=>"100110111",
  27520=>"000101110",
  27521=>"100010101",
  27522=>"000001000",
  27523=>"011010011",
  27524=>"001001101",
  27525=>"000000101",
  27526=>"011110000",
  27527=>"111010110",
  27528=>"011101100",
  27529=>"110100010",
  27530=>"101100111",
  27531=>"000110010",
  27532=>"111101111",
  27533=>"001111010",
  27534=>"111011100",
  27535=>"110001111",
  27536=>"101101101",
  27537=>"000010000",
  27538=>"000110111",
  27539=>"111001100",
  27540=>"111010110",
  27541=>"000011100",
  27542=>"100010001",
  27543=>"011110000",
  27544=>"000000001",
  27545=>"111001111",
  27546=>"101000100",
  27547=>"010100100",
  27548=>"001000100",
  27549=>"010100100",
  27550=>"000010000",
  27551=>"100001111",
  27552=>"010101100",
  27553=>"011011110",
  27554=>"101100000",
  27555=>"101100100",
  27556=>"110010101",
  27557=>"011010010",
  27558=>"011011101",
  27559=>"001111011",
  27560=>"011001100",
  27561=>"000000000",
  27562=>"011101101",
  27563=>"000110110",
  27564=>"011110101",
  27565=>"011101100",
  27566=>"110001100",
  27567=>"110011100",
  27568=>"011001111",
  27569=>"111101010",
  27570=>"100000001",
  27571=>"101101000",
  27572=>"000111110",
  27573=>"101100000",
  27574=>"101001010",
  27575=>"000001001",
  27576=>"011111001",
  27577=>"010100001",
  27578=>"011011111",
  27579=>"001101001",
  27580=>"000111111",
  27581=>"000000000",
  27582=>"000001000",
  27583=>"000001100",
  27584=>"000011001",
  27585=>"100000011",
  27586=>"111010001",
  27587=>"000111010",
  27588=>"101110011",
  27589=>"100001001",
  27590=>"010010001",
  27591=>"001101101",
  27592=>"000111000",
  27593=>"000111111",
  27594=>"111100001",
  27595=>"001111001",
  27596=>"011010101",
  27597=>"000101110",
  27598=>"101000011",
  27599=>"100111111",
  27600=>"110010110",
  27601=>"100010100",
  27602=>"000100010",
  27603=>"011111101",
  27604=>"000110110",
  27605=>"111011011",
  27606=>"111111000",
  27607=>"001111001",
  27608=>"111010000",
  27609=>"110001001",
  27610=>"000101000",
  27611=>"001101001",
  27612=>"001010000",
  27613=>"110010001",
  27614=>"001100101",
  27615=>"010110101",
  27616=>"011000001",
  27617=>"110100011",
  27618=>"100011001",
  27619=>"100000011",
  27620=>"100111100",
  27621=>"010111010",
  27622=>"001111001",
  27623=>"000111110",
  27624=>"100000001",
  27625=>"101000101",
  27626=>"000010100",
  27627=>"110100001",
  27628=>"111100110",
  27629=>"111110101",
  27630=>"011101100",
  27631=>"011000001",
  27632=>"100011011",
  27633=>"111011110",
  27634=>"110111000",
  27635=>"011111010",
  27636=>"110101011",
  27637=>"100011010",
  27638=>"011001100",
  27639=>"111101101",
  27640=>"110010001",
  27641=>"000000001",
  27642=>"101110100",
  27643=>"001001011",
  27644=>"001000110",
  27645=>"000110011",
  27646=>"000000000",
  27647=>"101101110",
  27648=>"101001011",
  27649=>"001011101",
  27650=>"100110101",
  27651=>"110100111",
  27652=>"101110011",
  27653=>"110010110",
  27654=>"001110111",
  27655=>"000001110",
  27656=>"110111100",
  27657=>"011010010",
  27658=>"010001101",
  27659=>"111111001",
  27660=>"111000010",
  27661=>"011101101",
  27662=>"001001010",
  27663=>"100010001",
  27664=>"110110110",
  27665=>"001010101",
  27666=>"100101010",
  27667=>"001010010",
  27668=>"101010010",
  27669=>"010000010",
  27670=>"011100000",
  27671=>"110111111",
  27672=>"010001011",
  27673=>"001100011",
  27674=>"110010001",
  27675=>"101111010",
  27676=>"101101001",
  27677=>"111101110",
  27678=>"011100001",
  27679=>"001011110",
  27680=>"010011100",
  27681=>"001100110",
  27682=>"100000100",
  27683=>"101111100",
  27684=>"101111001",
  27685=>"011100010",
  27686=>"101000111",
  27687=>"110100001",
  27688=>"101011011",
  27689=>"011100110",
  27690=>"100101100",
  27691=>"000101111",
  27692=>"111110111",
  27693=>"100001001",
  27694=>"001100001",
  27695=>"010110010",
  27696=>"011011010",
  27697=>"100100101",
  27698=>"001001100",
  27699=>"111111000",
  27700=>"001100110",
  27701=>"011110000",
  27702=>"011010010",
  27703=>"110111111",
  27704=>"111110000",
  27705=>"010110001",
  27706=>"100110110",
  27707=>"111010110",
  27708=>"000000010",
  27709=>"100111011",
  27710=>"010100001",
  27711=>"100101010",
  27712=>"101000110",
  27713=>"101000100",
  27714=>"100011100",
  27715=>"001001000",
  27716=>"001110010",
  27717=>"001100101",
  27718=>"000001110",
  27719=>"100111100",
  27720=>"110001100",
  27721=>"111101000",
  27722=>"001000101",
  27723=>"000101111",
  27724=>"111001001",
  27725=>"010011011",
  27726=>"000111101",
  27727=>"100001000",
  27728=>"011110000",
  27729=>"100101100",
  27730=>"010010010",
  27731=>"000100101",
  27732=>"001011000",
  27733=>"010010011",
  27734=>"101011111",
  27735=>"111110000",
  27736=>"011110111",
  27737=>"011100110",
  27738=>"001010001",
  27739=>"011111001",
  27740=>"001001000",
  27741=>"011011011",
  27742=>"010101101",
  27743=>"110010101",
  27744=>"000110100",
  27745=>"100000000",
  27746=>"111001111",
  27747=>"001000000",
  27748=>"110001000",
  27749=>"010111101",
  27750=>"010101011",
  27751=>"101110001",
  27752=>"101100010",
  27753=>"011000101",
  27754=>"010101100",
  27755=>"011100000",
  27756=>"111101001",
  27757=>"011101000",
  27758=>"110010110",
  27759=>"111011111",
  27760=>"011011010",
  27761=>"110100010",
  27762=>"001111101",
  27763=>"000111111",
  27764=>"101111111",
  27765=>"110101010",
  27766=>"001110111",
  27767=>"000011000",
  27768=>"101111011",
  27769=>"100010001",
  27770=>"010101000",
  27771=>"111001101",
  27772=>"101001101",
  27773=>"101111101",
  27774=>"101100101",
  27775=>"000010110",
  27776=>"100001110",
  27777=>"111001000",
  27778=>"110100111",
  27779=>"001010101",
  27780=>"101010110",
  27781=>"100100111",
  27782=>"010011111",
  27783=>"011011100",
  27784=>"011000000",
  27785=>"000001000",
  27786=>"000010010",
  27787=>"110101110",
  27788=>"111101101",
  27789=>"110011101",
  27790=>"110101000",
  27791=>"011010000",
  27792=>"101101011",
  27793=>"111111111",
  27794=>"101111101",
  27795=>"000110010",
  27796=>"011110101",
  27797=>"111111110",
  27798=>"010011111",
  27799=>"110111010",
  27800=>"000100110",
  27801=>"100111100",
  27802=>"111011001",
  27803=>"100110010",
  27804=>"011010000",
  27805=>"000111011",
  27806=>"111010001",
  27807=>"010011000",
  27808=>"001010100",
  27809=>"001111110",
  27810=>"011000001",
  27811=>"000111111",
  27812=>"101111101",
  27813=>"000110110",
  27814=>"100111101",
  27815=>"111011111",
  27816=>"001110111",
  27817=>"011000101",
  27818=>"100011101",
  27819=>"010011001",
  27820=>"000100000",
  27821=>"101011000",
  27822=>"011101000",
  27823=>"000100001",
  27824=>"111100001",
  27825=>"100001000",
  27826=>"000101100",
  27827=>"010101111",
  27828=>"110110111",
  27829=>"111101010",
  27830=>"110010000",
  27831=>"100110111",
  27832=>"110100110",
  27833=>"000001100",
  27834=>"110100110",
  27835=>"100101011",
  27836=>"001101101",
  27837=>"110001000",
  27838=>"101101110",
  27839=>"111011010",
  27840=>"011101011",
  27841=>"100111111",
  27842=>"100011001",
  27843=>"100101000",
  27844=>"101101100",
  27845=>"001110010",
  27846=>"110101010",
  27847=>"001010001",
  27848=>"100000000",
  27849=>"101101010",
  27850=>"100000011",
  27851=>"011011110",
  27852=>"000010001",
  27853=>"011011011",
  27854=>"100000011",
  27855=>"001001111",
  27856=>"000111000",
  27857=>"111101001",
  27858=>"001001010",
  27859=>"010111111",
  27860=>"110010110",
  27861=>"010001010",
  27862=>"010010100",
  27863=>"101000110",
  27864=>"011010101",
  27865=>"100000011",
  27866=>"110100011",
  27867=>"110110100",
  27868=>"000111010",
  27869=>"011111000",
  27870=>"011011100",
  27871=>"001011101",
  27872=>"000011010",
  27873=>"111111110",
  27874=>"011011110",
  27875=>"101111010",
  27876=>"100010110",
  27877=>"010000101",
  27878=>"111010001",
  27879=>"000001000",
  27880=>"110111001",
  27881=>"011111110",
  27882=>"100011111",
  27883=>"100100100",
  27884=>"100000101",
  27885=>"011001111",
  27886=>"011001111",
  27887=>"111000000",
  27888=>"101100011",
  27889=>"011001111",
  27890=>"001100101",
  27891=>"111011000",
  27892=>"101111011",
  27893=>"100100001",
  27894=>"111011010",
  27895=>"100111100",
  27896=>"000100011",
  27897=>"101111100",
  27898=>"100110010",
  27899=>"111001000",
  27900=>"100000000",
  27901=>"000011110",
  27902=>"110010110",
  27903=>"000110001",
  27904=>"110110000",
  27905=>"001101000",
  27906=>"011101101",
  27907=>"000011001",
  27908=>"100110111",
  27909=>"111101110",
  27910=>"010000011",
  27911=>"110100100",
  27912=>"001111110",
  27913=>"000001110",
  27914=>"110100111",
  27915=>"101011101",
  27916=>"101101110",
  27917=>"011110001",
  27918=>"011110110",
  27919=>"011001110",
  27920=>"001111010",
  27921=>"000010101",
  27922=>"101110010",
  27923=>"001010001",
  27924=>"100111011",
  27925=>"110000111",
  27926=>"100000111",
  27927=>"111101101",
  27928=>"000111010",
  27929=>"011001100",
  27930=>"101100001",
  27931=>"011100000",
  27932=>"000011010",
  27933=>"111010100",
  27934=>"000010011",
  27935=>"011010101",
  27936=>"000111101",
  27937=>"010000101",
  27938=>"111010011",
  27939=>"001010110",
  27940=>"110010000",
  27941=>"011000110",
  27942=>"000001010",
  27943=>"011100101",
  27944=>"000111110",
  27945=>"000010101",
  27946=>"011111111",
  27947=>"111100101",
  27948=>"001101101",
  27949=>"001000000",
  27950=>"111011001",
  27951=>"000111111",
  27952=>"110011000",
  27953=>"111110100",
  27954=>"001001001",
  27955=>"110100000",
  27956=>"100010111",
  27957=>"001001100",
  27958=>"110010110",
  27959=>"011111100",
  27960=>"100000101",
  27961=>"100000010",
  27962=>"011000001",
  27963=>"100110101",
  27964=>"001111110",
  27965=>"010000100",
  27966=>"001110100",
  27967=>"000000010",
  27968=>"011101101",
  27969=>"000000010",
  27970=>"011011110",
  27971=>"010000110",
  27972=>"111011001",
  27973=>"000110010",
  27974=>"001001000",
  27975=>"001010110",
  27976=>"001011101",
  27977=>"100011111",
  27978=>"110111100",
  27979=>"100000001",
  27980=>"000010101",
  27981=>"011110100",
  27982=>"010110001",
  27983=>"110110110",
  27984=>"010010100",
  27985=>"101110000",
  27986=>"000000111",
  27987=>"001000101",
  27988=>"010011110",
  27989=>"010101011",
  27990=>"000000110",
  27991=>"011111011",
  27992=>"010111100",
  27993=>"001000101",
  27994=>"100001101",
  27995=>"111010000",
  27996=>"001110110",
  27997=>"101101111",
  27998=>"101100000",
  27999=>"111100011",
  28000=>"111101010",
  28001=>"011110000",
  28002=>"000100110",
  28003=>"101110111",
  28004=>"001001000",
  28005=>"111101100",
  28006=>"010011010",
  28007=>"000000001",
  28008=>"010011101",
  28009=>"001101111",
  28010=>"010101111",
  28011=>"100101111",
  28012=>"110101110",
  28013=>"011111100",
  28014=>"001110011",
  28015=>"110001011",
  28016=>"001000010",
  28017=>"011011101",
  28018=>"011100111",
  28019=>"101011110",
  28020=>"011010100",
  28021=>"000001111",
  28022=>"100011010",
  28023=>"011011011",
  28024=>"001101001",
  28025=>"111111011",
  28026=>"010010001",
  28027=>"101000000",
  28028=>"000000110",
  28029=>"101001100",
  28030=>"111001100",
  28031=>"101000000",
  28032=>"100010100",
  28033=>"010111010",
  28034=>"010011010",
  28035=>"010111100",
  28036=>"100110101",
  28037=>"010100100",
  28038=>"010101010",
  28039=>"100001110",
  28040=>"100110001",
  28041=>"100010000",
  28042=>"011000111",
  28043=>"101111001",
  28044=>"000000000",
  28045=>"001111101",
  28046=>"110010100",
  28047=>"111100101",
  28048=>"000110110",
  28049=>"010011101",
  28050=>"010011001",
  28051=>"001000000",
  28052=>"111101101",
  28053=>"010000010",
  28054=>"100000000",
  28055=>"111000100",
  28056=>"001100001",
  28057=>"110101001",
  28058=>"100010110",
  28059=>"111101001",
  28060=>"111011010",
  28061=>"111001111",
  28062=>"100110111",
  28063=>"111011110",
  28064=>"001110011",
  28065=>"000110011",
  28066=>"111001110",
  28067=>"000111010",
  28068=>"001100000",
  28069=>"101010111",
  28070=>"110101011",
  28071=>"110100101",
  28072=>"101111100",
  28073=>"010011011",
  28074=>"001000111",
  28075=>"001100000",
  28076=>"010000001",
  28077=>"010011101",
  28078=>"010101100",
  28079=>"010001001",
  28080=>"111110101",
  28081=>"011001100",
  28082=>"000001000",
  28083=>"010100111",
  28084=>"010111110",
  28085=>"100110100",
  28086=>"101010111",
  28087=>"000010000",
  28088=>"001110100",
  28089=>"010001100",
  28090=>"000101110",
  28091=>"101110100",
  28092=>"000001111",
  28093=>"011110111",
  28094=>"000101111",
  28095=>"110110001",
  28096=>"010111111",
  28097=>"000111011",
  28098=>"001001010",
  28099=>"100100000",
  28100=>"111110010",
  28101=>"101111110",
  28102=>"011110101",
  28103=>"001001111",
  28104=>"110100000",
  28105=>"101100111",
  28106=>"110010011",
  28107=>"000100001",
  28108=>"010110001",
  28109=>"000101100",
  28110=>"010101011",
  28111=>"011001010",
  28112=>"101011110",
  28113=>"011110010",
  28114=>"011011000",
  28115=>"110010001",
  28116=>"011000101",
  28117=>"101010010",
  28118=>"110010011",
  28119=>"011100001",
  28120=>"111110001",
  28121=>"101100101",
  28122=>"110000001",
  28123=>"111001001",
  28124=>"101010100",
  28125=>"111110000",
  28126=>"101100011",
  28127=>"001011110",
  28128=>"111011000",
  28129=>"110101101",
  28130=>"111010110",
  28131=>"110010101",
  28132=>"000010111",
  28133=>"101010100",
  28134=>"010001011",
  28135=>"111111100",
  28136=>"001001111",
  28137=>"001110000",
  28138=>"111011111",
  28139=>"111101100",
  28140=>"101000010",
  28141=>"101110110",
  28142=>"010101011",
  28143=>"101001000",
  28144=>"110001100",
  28145=>"010101101",
  28146=>"001100110",
  28147=>"100101000",
  28148=>"110100010",
  28149=>"100111111",
  28150=>"100111010",
  28151=>"010000001",
  28152=>"110111000",
  28153=>"101101001",
  28154=>"011100111",
  28155=>"001111100",
  28156=>"110001100",
  28157=>"110010100",
  28158=>"001101110",
  28159=>"011000001",
  28160=>"000101011",
  28161=>"010010000",
  28162=>"110011100",
  28163=>"111000000",
  28164=>"001110111",
  28165=>"001111111",
  28166=>"011101010",
  28167=>"000000001",
  28168=>"001000101",
  28169=>"111000011",
  28170=>"101101110",
  28171=>"011001000",
  28172=>"011111101",
  28173=>"000001100",
  28174=>"101101100",
  28175=>"011111011",
  28176=>"110010111",
  28177=>"001101101",
  28178=>"011101010",
  28179=>"001110010",
  28180=>"110001011",
  28181=>"001111100",
  28182=>"011011010",
  28183=>"011100111",
  28184=>"111001011",
  28185=>"101100110",
  28186=>"111001110",
  28187=>"011111001",
  28188=>"000100101",
  28189=>"000010011",
  28190=>"100111101",
  28191=>"011000011",
  28192=>"000001011",
  28193=>"111010001",
  28194=>"100000000",
  28195=>"011100001",
  28196=>"011110101",
  28197=>"010101010",
  28198=>"001010000",
  28199=>"010000111",
  28200=>"100110011",
  28201=>"110110101",
  28202=>"110000010",
  28203=>"000001101",
  28204=>"100011111",
  28205=>"010111000",
  28206=>"101110001",
  28207=>"110111110",
  28208=>"000000100",
  28209=>"011101101",
  28210=>"000000011",
  28211=>"111101000",
  28212=>"111000101",
  28213=>"010110101",
  28214=>"101000110",
  28215=>"101000111",
  28216=>"001111011",
  28217=>"001011001",
  28218=>"101000101",
  28219=>"100000000",
  28220=>"101010000",
  28221=>"011101101",
  28222=>"000100111",
  28223=>"000111110",
  28224=>"111110010",
  28225=>"001110001",
  28226=>"001011101",
  28227=>"110011111",
  28228=>"100001100",
  28229=>"101110001",
  28230=>"110000101",
  28231=>"010000011",
  28232=>"011110101",
  28233=>"100101110",
  28234=>"100110011",
  28235=>"001100001",
  28236=>"111110100",
  28237=>"101001111",
  28238=>"001001101",
  28239=>"011011111",
  28240=>"100010100",
  28241=>"110000001",
  28242=>"100010101",
  28243=>"010011000",
  28244=>"000100110",
  28245=>"011101010",
  28246=>"011010101",
  28247=>"100010001",
  28248=>"010011110",
  28249=>"010101111",
  28250=>"101000101",
  28251=>"101011010",
  28252=>"010010000",
  28253=>"111100110",
  28254=>"000001000",
  28255=>"110011010",
  28256=>"000100011",
  28257=>"101111000",
  28258=>"100110111",
  28259=>"101000000",
  28260=>"111100110",
  28261=>"110110100",
  28262=>"000100101",
  28263=>"110010010",
  28264=>"000010001",
  28265=>"100101101",
  28266=>"110010011",
  28267=>"010110000",
  28268=>"000010111",
  28269=>"101001110",
  28270=>"011001100",
  28271=>"001010110",
  28272=>"011100110",
  28273=>"000010000",
  28274=>"110011000",
  28275=>"100101100",
  28276=>"111111000",
  28277=>"100100110",
  28278=>"011010101",
  28279=>"101111010",
  28280=>"011011100",
  28281=>"111111000",
  28282=>"110101100",
  28283=>"100001110",
  28284=>"111101000",
  28285=>"010000010",
  28286=>"110011000",
  28287=>"000111110",
  28288=>"000000100",
  28289=>"010111001",
  28290=>"100010010",
  28291=>"001010100",
  28292=>"100100111",
  28293=>"111110100",
  28294=>"010011010",
  28295=>"001000101",
  28296=>"000100110",
  28297=>"010001101",
  28298=>"011110000",
  28299=>"000101101",
  28300=>"010010000",
  28301=>"000001100",
  28302=>"111011111",
  28303=>"011111011",
  28304=>"100010011",
  28305=>"001100100",
  28306=>"011011000",
  28307=>"111111101",
  28308=>"101110010",
  28309=>"010100100",
  28310=>"001100011",
  28311=>"101001110",
  28312=>"111001101",
  28313=>"010001101",
  28314=>"011000010",
  28315=>"100000100",
  28316=>"000000000",
  28317=>"000000111",
  28318=>"110111011",
  28319=>"010100000",
  28320=>"010001000",
  28321=>"111011010",
  28322=>"010010001",
  28323=>"000100000",
  28324=>"110100000",
  28325=>"001111100",
  28326=>"000110111",
  28327=>"100000001",
  28328=>"110001111",
  28329=>"000011001",
  28330=>"100101100",
  28331=>"110010010",
  28332=>"000111010",
  28333=>"001110110",
  28334=>"110100010",
  28335=>"110111100",
  28336=>"110010000",
  28337=>"001010110",
  28338=>"000111101",
  28339=>"101000001",
  28340=>"000110011",
  28341=>"111001111",
  28342=>"010100101",
  28343=>"000010000",
  28344=>"010001100",
  28345=>"011000000",
  28346=>"101111111",
  28347=>"111001001",
  28348=>"011000101",
  28349=>"011100010",
  28350=>"001000001",
  28351=>"010111011",
  28352=>"011110101",
  28353=>"111010000",
  28354=>"111010001",
  28355=>"110011010",
  28356=>"011000011",
  28357=>"000111001",
  28358=>"110101111",
  28359=>"111000011",
  28360=>"001001111",
  28361=>"000111000",
  28362=>"101110011",
  28363=>"110100110",
  28364=>"001010010",
  28365=>"111011001",
  28366=>"010100001",
  28367=>"111101111",
  28368=>"010110111",
  28369=>"010110011",
  28370=>"000000010",
  28371=>"001110000",
  28372=>"010011100",
  28373=>"100010110",
  28374=>"100000101",
  28375=>"010101100",
  28376=>"001110101",
  28377=>"011110111",
  28378=>"010100100",
  28379=>"110101111",
  28380=>"101101100",
  28381=>"111111011",
  28382=>"011001101",
  28383=>"111010001",
  28384=>"010011111",
  28385=>"111110101",
  28386=>"000011101",
  28387=>"101111100",
  28388=>"111110100",
  28389=>"101101011",
  28390=>"000000000",
  28391=>"110011010",
  28392=>"100010111",
  28393=>"010000011",
  28394=>"011000110",
  28395=>"101011111",
  28396=>"000010111",
  28397=>"100011100",
  28398=>"110010010",
  28399=>"001110000",
  28400=>"001010010",
  28401=>"000100111",
  28402=>"011010110",
  28403=>"000011010",
  28404=>"000111100",
  28405=>"101100100",
  28406=>"101010111",
  28407=>"010110011",
  28408=>"101011100",
  28409=>"000000000",
  28410=>"011001101",
  28411=>"100000100",
  28412=>"001101111",
  28413=>"100100010",
  28414=>"011111010",
  28415=>"000010001",
  28416=>"111111110",
  28417=>"101000011",
  28418=>"111000110",
  28419=>"000001111",
  28420=>"011111011",
  28421=>"101111101",
  28422=>"111000100",
  28423=>"100101010",
  28424=>"110111100",
  28425=>"010010110",
  28426=>"111001000",
  28427=>"101001000",
  28428=>"111010100",
  28429=>"100011000",
  28430=>"000001001",
  28431=>"010011010",
  28432=>"001101111",
  28433=>"101100010",
  28434=>"101101110",
  28435=>"110001000",
  28436=>"101110111",
  28437=>"100110101",
  28438=>"011100011",
  28439=>"111001001",
  28440=>"010010110",
  28441=>"000011101",
  28442=>"000100111",
  28443=>"111011000",
  28444=>"101000001",
  28445=>"100101101",
  28446=>"110110100",
  28447=>"000110011",
  28448=>"000110000",
  28449=>"001101110",
  28450=>"001011111",
  28451=>"101001000",
  28452=>"001000110",
  28453=>"011000001",
  28454=>"011101010",
  28455=>"010101000",
  28456=>"000111110",
  28457=>"010101100",
  28458=>"001011100",
  28459=>"011010000",
  28460=>"000000101",
  28461=>"000110111",
  28462=>"100010011",
  28463=>"000011110",
  28464=>"110001101",
  28465=>"110101011",
  28466=>"011011000",
  28467=>"000011110",
  28468=>"110101000",
  28469=>"001111010",
  28470=>"011010101",
  28471=>"111100101",
  28472=>"100011010",
  28473=>"110001000",
  28474=>"101110000",
  28475=>"001110001",
  28476=>"110000110",
  28477=>"001111001",
  28478=>"111000101",
  28479=>"110101010",
  28480=>"100001101",
  28481=>"100001010",
  28482=>"010010101",
  28483=>"110100001",
  28484=>"101000011",
  28485=>"000001010",
  28486=>"111000100",
  28487=>"011101111",
  28488=>"100000111",
  28489=>"000100010",
  28490=>"100101011",
  28491=>"100010101",
  28492=>"111100010",
  28493=>"101111010",
  28494=>"110000010",
  28495=>"100000000",
  28496=>"011010010",
  28497=>"111001011",
  28498=>"101110000",
  28499=>"011000000",
  28500=>"101111010",
  28501=>"111101101",
  28502=>"000110110",
  28503=>"101110111",
  28504=>"100111110",
  28505=>"110010110",
  28506=>"000010010",
  28507=>"001100000",
  28508=>"111100010",
  28509=>"111011001",
  28510=>"010011010",
  28511=>"111111110",
  28512=>"000001011",
  28513=>"111111011",
  28514=>"001010101",
  28515=>"110111111",
  28516=>"100101100",
  28517=>"100010010",
  28518=>"100111111",
  28519=>"001111000",
  28520=>"100111110",
  28521=>"000000110",
  28522=>"101000101",
  28523=>"000010111",
  28524=>"011101111",
  28525=>"111011000",
  28526=>"010010000",
  28527=>"010001111",
  28528=>"110111000",
  28529=>"100110010",
  28530=>"100110101",
  28531=>"110110001",
  28532=>"110011110",
  28533=>"111001011",
  28534=>"110001000",
  28535=>"111111110",
  28536=>"011011111",
  28537=>"001001010",
  28538=>"000111100",
  28539=>"000001011",
  28540=>"111111000",
  28541=>"010110110",
  28542=>"010110001",
  28543=>"011110000",
  28544=>"010110110",
  28545=>"101110001",
  28546=>"100101000",
  28547=>"011010110",
  28548=>"100110111",
  28549=>"100111000",
  28550=>"110001111",
  28551=>"000000100",
  28552=>"011111111",
  28553=>"010000010",
  28554=>"000110011",
  28555=>"011001010",
  28556=>"011101000",
  28557=>"011011010",
  28558=>"100101110",
  28559=>"011000111",
  28560=>"101000010",
  28561=>"100100001",
  28562=>"011000100",
  28563=>"010110001",
  28564=>"100011011",
  28565=>"111011110",
  28566=>"011111100",
  28567=>"000101000",
  28568=>"110111111",
  28569=>"011100010",
  28570=>"110111110",
  28571=>"110001010",
  28572=>"010010100",
  28573=>"011000000",
  28574=>"011010011",
  28575=>"101110010",
  28576=>"001001011",
  28577=>"110100111",
  28578=>"111100001",
  28579=>"000001000",
  28580=>"111111010",
  28581=>"000000111",
  28582=>"111100010",
  28583=>"110010011",
  28584=>"110010100",
  28585=>"011010001",
  28586=>"000100011",
  28587=>"010011011",
  28588=>"101011001",
  28589=>"101110111",
  28590=>"110001100",
  28591=>"001001001",
  28592=>"101000010",
  28593=>"111000101",
  28594=>"011100010",
  28595=>"011111101",
  28596=>"001000010",
  28597=>"101011100",
  28598=>"111011001",
  28599=>"001000000",
  28600=>"000000101",
  28601=>"000000010",
  28602=>"010000011",
  28603=>"110011101",
  28604=>"101110101",
  28605=>"110101110",
  28606=>"001010000",
  28607=>"100001101",
  28608=>"001100010",
  28609=>"010000000",
  28610=>"100001001",
  28611=>"100010001",
  28612=>"101111111",
  28613=>"001010000",
  28614=>"001101010",
  28615=>"011111000",
  28616=>"100100100",
  28617=>"110111111",
  28618=>"010110011",
  28619=>"000110100",
  28620=>"001010110",
  28621=>"000111001",
  28622=>"010010000",
  28623=>"011100011",
  28624=>"101001010",
  28625=>"111110101",
  28626=>"001011011",
  28627=>"000000001",
  28628=>"110000011",
  28629=>"110100110",
  28630=>"000010101",
  28631=>"001000111",
  28632=>"100010111",
  28633=>"010110100",
  28634=>"000100011",
  28635=>"100010100",
  28636=>"011010100",
  28637=>"111101010",
  28638=>"001101001",
  28639=>"000100111",
  28640=>"001001110",
  28641=>"000000000",
  28642=>"001111011",
  28643=>"000001111",
  28644=>"111001010",
  28645=>"011110001",
  28646=>"010011100",
  28647=>"010011111",
  28648=>"101000100",
  28649=>"101101010",
  28650=>"001010110",
  28651=>"010100011",
  28652=>"001111000",
  28653=>"011111000",
  28654=>"010011110",
  28655=>"101110001",
  28656=>"111010100",
  28657=>"110100101",
  28658=>"101000001",
  28659=>"000001111",
  28660=>"100111010",
  28661=>"000001101",
  28662=>"101100101",
  28663=>"010010011",
  28664=>"000011111",
  28665=>"110010001",
  28666=>"001001011",
  28667=>"100111001",
  28668=>"100100110",
  28669=>"111011010",
  28670=>"000111111",
  28671=>"110111111",
  28672=>"000001000",
  28673=>"110000010",
  28674=>"011111000",
  28675=>"001000000",
  28676=>"001101101",
  28677=>"011000000",
  28678=>"000111110",
  28679=>"010100100",
  28680=>"101000011",
  28681=>"101001001",
  28682=>"000010011",
  28683=>"001111000",
  28684=>"100000000",
  28685=>"011111011",
  28686=>"000000000",
  28687=>"010111010",
  28688=>"100100101",
  28689=>"100001110",
  28690=>"111110001",
  28691=>"011001000",
  28692=>"001010000",
  28693=>"101001101",
  28694=>"100011101",
  28695=>"111101111",
  28696=>"111000011",
  28697=>"001010001",
  28698=>"010111110",
  28699=>"101110011",
  28700=>"110010110",
  28701=>"010101110",
  28702=>"001100001",
  28703=>"111001000",
  28704=>"101101111",
  28705=>"101010000",
  28706=>"011000100",
  28707=>"001011011",
  28708=>"001001111",
  28709=>"010101100",
  28710=>"001101011",
  28711=>"100101000",
  28712=>"001011011",
  28713=>"000000000",
  28714=>"010111001",
  28715=>"100011010",
  28716=>"101110101",
  28717=>"110111101",
  28718=>"000001101",
  28719=>"001101111",
  28720=>"100111110",
  28721=>"010001101",
  28722=>"000101101",
  28723=>"011110101",
  28724=>"101100011",
  28725=>"101100000",
  28726=>"110100011",
  28727=>"100111101",
  28728=>"101001000",
  28729=>"101111010",
  28730=>"010001100",
  28731=>"011111100",
  28732=>"001010011",
  28733=>"000010100",
  28734=>"010110111",
  28735=>"101010000",
  28736=>"011010111",
  28737=>"001000110",
  28738=>"101000111",
  28739=>"110101100",
  28740=>"100101001",
  28741=>"110011110",
  28742=>"001111111",
  28743=>"100100010",
  28744=>"101101000",
  28745=>"100001010",
  28746=>"111100001",
  28747=>"111111100",
  28748=>"000000010",
  28749=>"010100101",
  28750=>"110111010",
  28751=>"011000001",
  28752=>"110111001",
  28753=>"010111011",
  28754=>"111010111",
  28755=>"101011010",
  28756=>"111110010",
  28757=>"110011111",
  28758=>"101011001",
  28759=>"000101001",
  28760=>"110100011",
  28761=>"100100010",
  28762=>"101000111",
  28763=>"000101001",
  28764=>"110011010",
  28765=>"110010100",
  28766=>"000110001",
  28767=>"110000101",
  28768=>"001100100",
  28769=>"101001010",
  28770=>"001010101",
  28771=>"101100000",
  28772=>"111011001",
  28773=>"011101101",
  28774=>"111011000",
  28775=>"000110000",
  28776=>"000011101",
  28777=>"110010001",
  28778=>"000001100",
  28779=>"011010111",
  28780=>"010000110",
  28781=>"110100100",
  28782=>"000111111",
  28783=>"101000101",
  28784=>"000010000",
  28785=>"101110010",
  28786=>"101111011",
  28787=>"000100100",
  28788=>"111001001",
  28789=>"000010010",
  28790=>"111011110",
  28791=>"101110011",
  28792=>"011101111",
  28793=>"010011001",
  28794=>"000010110",
  28795=>"011100011",
  28796=>"100000100",
  28797=>"000001000",
  28798=>"110110000",
  28799=>"100101110",
  28800=>"110001101",
  28801=>"010111100",
  28802=>"011000000",
  28803=>"110000010",
  28804=>"001110101",
  28805=>"101100011",
  28806=>"001101011",
  28807=>"000100110",
  28808=>"011100100",
  28809=>"010000001",
  28810=>"100010010",
  28811=>"110111110",
  28812=>"000000000",
  28813=>"111001001",
  28814=>"111110111",
  28815=>"100111011",
  28816=>"000111000",
  28817=>"011101110",
  28818=>"011000101",
  28819=>"001100011",
  28820=>"011010010",
  28821=>"100110011",
  28822=>"101001001",
  28823=>"111010000",
  28824=>"101000110",
  28825=>"011100000",
  28826=>"011100111",
  28827=>"101110101",
  28828=>"001001000",
  28829=>"010110110",
  28830=>"100010011",
  28831=>"110111011",
  28832=>"101000101",
  28833=>"000110100",
  28834=>"010110000",
  28835=>"110000101",
  28836=>"011110000",
  28837=>"001100101",
  28838=>"000101000",
  28839=>"001001110",
  28840=>"011001110",
  28841=>"000111001",
  28842=>"010000000",
  28843=>"000101010",
  28844=>"011010111",
  28845=>"010011000",
  28846=>"000111100",
  28847=>"111111110",
  28848=>"011011000",
  28849=>"011010111",
  28850=>"100111110",
  28851=>"000000011",
  28852=>"111100010",
  28853=>"011000010",
  28854=>"101110011",
  28855=>"110001000",
  28856=>"010101111",
  28857=>"000000100",
  28858=>"001101100",
  28859=>"101010011",
  28860=>"010111110",
  28861=>"011110100",
  28862=>"000111011",
  28863=>"100001011",
  28864=>"011110010",
  28865=>"000110000",
  28866=>"100000100",
  28867=>"010110100",
  28868=>"111100011",
  28869=>"110010011",
  28870=>"001111010",
  28871=>"000011011",
  28872=>"011010010",
  28873=>"111000000",
  28874=>"001000111",
  28875=>"101101010",
  28876=>"111111111",
  28877=>"100100111",
  28878=>"101101010",
  28879=>"101100111",
  28880=>"010001101",
  28881=>"100111010",
  28882=>"010000100",
  28883=>"000111000",
  28884=>"111001110",
  28885=>"001101100",
  28886=>"101000010",
  28887=>"011010011",
  28888=>"100010100",
  28889=>"111111111",
  28890=>"001011110",
  28891=>"111010111",
  28892=>"010100011",
  28893=>"010011110",
  28894=>"010110001",
  28895=>"111000100",
  28896=>"110101000",
  28897=>"110000011",
  28898=>"111011101",
  28899=>"010010100",
  28900=>"100000100",
  28901=>"101011000",
  28902=>"000100011",
  28903=>"000100001",
  28904=>"010000010",
  28905=>"101001001",
  28906=>"011001101",
  28907=>"100111100",
  28908=>"010110011",
  28909=>"000011101",
  28910=>"110001101",
  28911=>"011111010",
  28912=>"100111110",
  28913=>"000011010",
  28914=>"100001001",
  28915=>"001101011",
  28916=>"100110011",
  28917=>"011110111",
  28918=>"110101000",
  28919=>"011100001",
  28920=>"010000010",
  28921=>"111001100",
  28922=>"111110011",
  28923=>"110001101",
  28924=>"110101110",
  28925=>"000111111",
  28926=>"000110100",
  28927=>"111011111",
  28928=>"110001001",
  28929=>"010110010",
  28930=>"010100011",
  28931=>"101100001",
  28932=>"111011111",
  28933=>"110000110",
  28934=>"101000010",
  28935=>"110000011",
  28936=>"000100001",
  28937=>"001001001",
  28938=>"011100011",
  28939=>"001001001",
  28940=>"101010000",
  28941=>"111101000",
  28942=>"100000000",
  28943=>"100110110",
  28944=>"011010011",
  28945=>"011010000",
  28946=>"110010100",
  28947=>"111110001",
  28948=>"110111001",
  28949=>"011100101",
  28950=>"100111111",
  28951=>"100111111",
  28952=>"110010000",
  28953=>"001001001",
  28954=>"010011000",
  28955=>"000010101",
  28956=>"100111111",
  28957=>"101001010",
  28958=>"111101011",
  28959=>"001011010",
  28960=>"100100111",
  28961=>"111111101",
  28962=>"111011000",
  28963=>"001100001",
  28964=>"111000101",
  28965=>"010000000",
  28966=>"010011000",
  28967=>"100010100",
  28968=>"001100101",
  28969=>"010101000",
  28970=>"011001101",
  28971=>"111011110",
  28972=>"011101011",
  28973=>"100101111",
  28974=>"011111111",
  28975=>"111011011",
  28976=>"100110100",
  28977=>"111011010",
  28978=>"010011111",
  28979=>"010111101",
  28980=>"000001000",
  28981=>"000110011",
  28982=>"110110000",
  28983=>"101100100",
  28984=>"001101000",
  28985=>"000101011",
  28986=>"100101110",
  28987=>"011111111",
  28988=>"011101011",
  28989=>"001111010",
  28990=>"101100001",
  28991=>"111110111",
  28992=>"110011011",
  28993=>"110001100",
  28994=>"100111001",
  28995=>"011110010",
  28996=>"101000001",
  28997=>"011011010",
  28998=>"010100011",
  28999=>"101111001",
  29000=>"101011110",
  29001=>"001100011",
  29002=>"101011000",
  29003=>"111100111",
  29004=>"011001001",
  29005=>"101011011",
  29006=>"100001010",
  29007=>"000010010",
  29008=>"100111001",
  29009=>"000101100",
  29010=>"100010101",
  29011=>"101001111",
  29012=>"001010010",
  29013=>"001000010",
  29014=>"000000010",
  29015=>"000111100",
  29016=>"110010101",
  29017=>"001010001",
  29018=>"110011011",
  29019=>"001101101",
  29020=>"001000110",
  29021=>"111010110",
  29022=>"001100100",
  29023=>"011000100",
  29024=>"110011100",
  29025=>"010010011",
  29026=>"011101001",
  29027=>"001101100",
  29028=>"110010000",
  29029=>"101101001",
  29030=>"000110110",
  29031=>"010110001",
  29032=>"001010000",
  29033=>"000111101",
  29034=>"010000111",
  29035=>"101100111",
  29036=>"101001100",
  29037=>"100100110",
  29038=>"100000001",
  29039=>"101101110",
  29040=>"000000111",
  29041=>"010110100",
  29042=>"010000101",
  29043=>"110111010",
  29044=>"110111001",
  29045=>"001111110",
  29046=>"010001100",
  29047=>"110110001",
  29048=>"100101100",
  29049=>"010010100",
  29050=>"001011110",
  29051=>"110111000",
  29052=>"100001011",
  29053=>"000110100",
  29054=>"000101111",
  29055=>"100110111",
  29056=>"100101000",
  29057=>"100000001",
  29058=>"001010000",
  29059=>"100000111",
  29060=>"010110111",
  29061=>"011100001",
  29062=>"110001011",
  29063=>"001000011",
  29064=>"111001001",
  29065=>"011000110",
  29066=>"011001100",
  29067=>"100010100",
  29068=>"000110101",
  29069=>"110011001",
  29070=>"100001110",
  29071=>"101010100",
  29072=>"100110100",
  29073=>"100000001",
  29074=>"001101010",
  29075=>"001101011",
  29076=>"001011101",
  29077=>"000100110",
  29078=>"111100111",
  29079=>"010001101",
  29080=>"110110100",
  29081=>"000011010",
  29082=>"000010010",
  29083=>"011001010",
  29084=>"000100110",
  29085=>"110001010",
  29086=>"000101001",
  29087=>"100110001",
  29088=>"100010010",
  29089=>"100010000",
  29090=>"000000101",
  29091=>"000100011",
  29092=>"011111110",
  29093=>"000000001",
  29094=>"001010011",
  29095=>"111000101",
  29096=>"111100110",
  29097=>"111000000",
  29098=>"101001110",
  29099=>"010100110",
  29100=>"011001011",
  29101=>"111100111",
  29102=>"000111100",
  29103=>"101000101",
  29104=>"110001100",
  29105=>"010100000",
  29106=>"101101100",
  29107=>"001110000",
  29108=>"100000011",
  29109=>"110110010",
  29110=>"011110111",
  29111=>"110010110",
  29112=>"100010010",
  29113=>"101011010",
  29114=>"001011000",
  29115=>"000000110",
  29116=>"100000000",
  29117=>"001100111",
  29118=>"010011101",
  29119=>"111011001",
  29120=>"110101110",
  29121=>"001000110",
  29122=>"011001110",
  29123=>"110110110",
  29124=>"101010111",
  29125=>"000000100",
  29126=>"000011101",
  29127=>"100100101",
  29128=>"100011111",
  29129=>"110000000",
  29130=>"001110100",
  29131=>"101110001",
  29132=>"011011111",
  29133=>"110000000",
  29134=>"001100111",
  29135=>"110101111",
  29136=>"100000100",
  29137=>"001010010",
  29138=>"000000011",
  29139=>"010111001",
  29140=>"011110101",
  29141=>"100001011",
  29142=>"111010110",
  29143=>"110000011",
  29144=>"011000111",
  29145=>"100010100",
  29146=>"011010101",
  29147=>"000000011",
  29148=>"100000110",
  29149=>"111101100",
  29150=>"010111001",
  29151=>"000100001",
  29152=>"111111111",
  29153=>"001101001",
  29154=>"101110110",
  29155=>"011001100",
  29156=>"011101110",
  29157=>"000011100",
  29158=>"101100100",
  29159=>"101001101",
  29160=>"111101001",
  29161=>"101110111",
  29162=>"000100001",
  29163=>"100000010",
  29164=>"101011010",
  29165=>"100001011",
  29166=>"000110000",
  29167=>"000111000",
  29168=>"110000001",
  29169=>"111101110",
  29170=>"001101110",
  29171=>"001110101",
  29172=>"010010101",
  29173=>"010110001",
  29174=>"101011110",
  29175=>"010010111",
  29176=>"101110000",
  29177=>"011010110",
  29178=>"000110001",
  29179=>"001101101",
  29180=>"000110011",
  29181=>"101110000",
  29182=>"100011111",
  29183=>"101010101",
  29184=>"011001100",
  29185=>"011010100",
  29186=>"011000001",
  29187=>"110001110",
  29188=>"000100110",
  29189=>"111110101",
  29190=>"011101000",
  29191=>"110101110",
  29192=>"011100000",
  29193=>"011010010",
  29194=>"110111110",
  29195=>"000011011",
  29196=>"110001011",
  29197=>"111110001",
  29198=>"010001000",
  29199=>"010101010",
  29200=>"100111010",
  29201=>"111111101",
  29202=>"100011000",
  29203=>"011100111",
  29204=>"001110100",
  29205=>"000111010",
  29206=>"101011010",
  29207=>"110010111",
  29208=>"000100101",
  29209=>"001101010",
  29210=>"010000010",
  29211=>"111010001",
  29212=>"101010001",
  29213=>"000000010",
  29214=>"100011001",
  29215=>"010100110",
  29216=>"111010101",
  29217=>"011111111",
  29218=>"011000010",
  29219=>"101111001",
  29220=>"001101010",
  29221=>"011101101",
  29222=>"101001011",
  29223=>"111000010",
  29224=>"100100100",
  29225=>"111110010",
  29226=>"100010000",
  29227=>"101100000",
  29228=>"000110011",
  29229=>"010010000",
  29230=>"011000000",
  29231=>"000111001",
  29232=>"000100101",
  29233=>"000010000",
  29234=>"001101000",
  29235=>"100011011",
  29236=>"100101110",
  29237=>"100000100",
  29238=>"111100011",
  29239=>"001010000",
  29240=>"100100101",
  29241=>"001010101",
  29242=>"111111010",
  29243=>"100011000",
  29244=>"101100111",
  29245=>"000101011",
  29246=>"000101000",
  29247=>"111000000",
  29248=>"011110100",
  29249=>"010011101",
  29250=>"001100101",
  29251=>"101000100",
  29252=>"010000010",
  29253=>"000111100",
  29254=>"010101101",
  29255=>"001001110",
  29256=>"101010101",
  29257=>"111101110",
  29258=>"011110101",
  29259=>"011110111",
  29260=>"101111101",
  29261=>"001101001",
  29262=>"101111000",
  29263=>"100000010",
  29264=>"001010111",
  29265=>"111010001",
  29266=>"110010011",
  29267=>"010101001",
  29268=>"000110101",
  29269=>"000110101",
  29270=>"001101001",
  29271=>"001100001",
  29272=>"010011110",
  29273=>"000111000",
  29274=>"000101001",
  29275=>"101011101",
  29276=>"010111110",
  29277=>"000000010",
  29278=>"011000111",
  29279=>"010011001",
  29280=>"001011000",
  29281=>"000101001",
  29282=>"101110110",
  29283=>"100101011",
  29284=>"010000011",
  29285=>"100100100",
  29286=>"101010100",
  29287=>"010010010",
  29288=>"100010010",
  29289=>"100100100",
  29290=>"101011000",
  29291=>"010100110",
  29292=>"100111111",
  29293=>"110101000",
  29294=>"111001111",
  29295=>"111010001",
  29296=>"110011100",
  29297=>"000010010",
  29298=>"111101000",
  29299=>"001001101",
  29300=>"101101010",
  29301=>"011000000",
  29302=>"001010010",
  29303=>"111011001",
  29304=>"011001100",
  29305=>"110001000",
  29306=>"010100010",
  29307=>"010011101",
  29308=>"011010100",
  29309=>"001111111",
  29310=>"100010010",
  29311=>"010010101",
  29312=>"111000011",
  29313=>"110101011",
  29314=>"110001000",
  29315=>"111001001",
  29316=>"001110100",
  29317=>"000100010",
  29318=>"100000100",
  29319=>"100100000",
  29320=>"001110111",
  29321=>"000000100",
  29322=>"101110001",
  29323=>"111101111",
  29324=>"100101010",
  29325=>"100100100",
  29326=>"101110001",
  29327=>"010100001",
  29328=>"000001101",
  29329=>"011010111",
  29330=>"010100101",
  29331=>"001110011",
  29332=>"101110101",
  29333=>"100100000",
  29334=>"010001010",
  29335=>"100001111",
  29336=>"000000000",
  29337=>"101011101",
  29338=>"000101011",
  29339=>"011110111",
  29340=>"001010010",
  29341=>"100011110",
  29342=>"010011010",
  29343=>"010010100",
  29344=>"110000010",
  29345=>"011101110",
  29346=>"010101101",
  29347=>"000001000",
  29348=>"110111111",
  29349=>"000111100",
  29350=>"100001111",
  29351=>"100101000",
  29352=>"010001010",
  29353=>"001000101",
  29354=>"001010010",
  29355=>"101111111",
  29356=>"100001001",
  29357=>"000011011",
  29358=>"111011100",
  29359=>"011101000",
  29360=>"000011101",
  29361=>"011101000",
  29362=>"100101101",
  29363=>"100111001",
  29364=>"110101011",
  29365=>"110010011",
  29366=>"001100010",
  29367=>"010100000",
  29368=>"101001001",
  29369=>"010111110",
  29370=>"101101100",
  29371=>"000010001",
  29372=>"010000111",
  29373=>"001001010",
  29374=>"100111000",
  29375=>"111000010",
  29376=>"000011101",
  29377=>"111011110",
  29378=>"011101101",
  29379=>"110011000",
  29380=>"101111100",
  29381=>"101010011",
  29382=>"100101001",
  29383=>"001101001",
  29384=>"110110000",
  29385=>"100100110",
  29386=>"011001000",
  29387=>"100100111",
  29388=>"000000110",
  29389=>"100011110",
  29390=>"010110011",
  29391=>"010001001",
  29392=>"110101110",
  29393=>"100111111",
  29394=>"011000101",
  29395=>"101100111",
  29396=>"010011011",
  29397=>"000010110",
  29398=>"000101111",
  29399=>"001101010",
  29400=>"000101001",
  29401=>"001001100",
  29402=>"110010000",
  29403=>"011111110",
  29404=>"101000111",
  29405=>"111000011",
  29406=>"101010000",
  29407=>"000110010",
  29408=>"110101000",
  29409=>"100010100",
  29410=>"011001010",
  29411=>"011110101",
  29412=>"111110101",
  29413=>"100100010",
  29414=>"001101000",
  29415=>"100010111",
  29416=>"100100011",
  29417=>"010001110",
  29418=>"000011100",
  29419=>"001000010",
  29420=>"100001110",
  29421=>"000010100",
  29422=>"001111011",
  29423=>"110011011",
  29424=>"010101100",
  29425=>"001101010",
  29426=>"001101000",
  29427=>"110101110",
  29428=>"111101010",
  29429=>"000000001",
  29430=>"111101101",
  29431=>"101111011",
  29432=>"001001110",
  29433=>"011110001",
  29434=>"001101101",
  29435=>"110011101",
  29436=>"011110001",
  29437=>"010111111",
  29438=>"101010110",
  29439=>"011100110",
  29440=>"101110010",
  29441=>"101100010",
  29442=>"100001001",
  29443=>"111011111",
  29444=>"110001101",
  29445=>"010010011",
  29446=>"000001100",
  29447=>"101111111",
  29448=>"010111000",
  29449=>"100000011",
  29450=>"000100110",
  29451=>"000001001",
  29452=>"111000011",
  29453=>"110001111",
  29454=>"100100011",
  29455=>"011100101",
  29456=>"100000100",
  29457=>"010111010",
  29458=>"010110110",
  29459=>"001110100",
  29460=>"111011010",
  29461=>"111100010",
  29462=>"111111101",
  29463=>"111010110",
  29464=>"001001001",
  29465=>"000010011",
  29466=>"001001111",
  29467=>"010010010",
  29468=>"001100111",
  29469=>"100011010",
  29470=>"110011011",
  29471=>"000000001",
  29472=>"000001010",
  29473=>"011100111",
  29474=>"110000001",
  29475=>"001010110",
  29476=>"000111110",
  29477=>"001101001",
  29478=>"100001011",
  29479=>"000111100",
  29480=>"110011011",
  29481=>"101010000",
  29482=>"001111101",
  29483=>"101011011",
  29484=>"011011001",
  29485=>"011110111",
  29486=>"110000010",
  29487=>"110000001",
  29488=>"101011010",
  29489=>"000010101",
  29490=>"100000010",
  29491=>"011111111",
  29492=>"000000010",
  29493=>"101001101",
  29494=>"101010001",
  29495=>"001111110",
  29496=>"011110000",
  29497=>"010011100",
  29498=>"001101111",
  29499=>"011100110",
  29500=>"100000101",
  29501=>"001100011",
  29502=>"000010100",
  29503=>"010010011",
  29504=>"010001011",
  29505=>"000111010",
  29506=>"110110000",
  29507=>"010111101",
  29508=>"001010110",
  29509=>"001111010",
  29510=>"010100110",
  29511=>"010001011",
  29512=>"100110110",
  29513=>"011101011",
  29514=>"000001111",
  29515=>"010101001",
  29516=>"110110110",
  29517=>"010101011",
  29518=>"100011110",
  29519=>"110000101",
  29520=>"111001000",
  29521=>"001100011",
  29522=>"001000101",
  29523=>"101101101",
  29524=>"011010111",
  29525=>"010011100",
  29526=>"110111001",
  29527=>"110101000",
  29528=>"100101111",
  29529=>"101101110",
  29530=>"001011011",
  29531=>"001101010",
  29532=>"011111011",
  29533=>"100100100",
  29534=>"010101011",
  29535=>"000100011",
  29536=>"010011111",
  29537=>"000100110",
  29538=>"000000100",
  29539=>"110110011",
  29540=>"101101010",
  29541=>"110100000",
  29542=>"010111101",
  29543=>"110110000",
  29544=>"110100010",
  29545=>"000000111",
  29546=>"010100111",
  29547=>"000111011",
  29548=>"011001110",
  29549=>"100111010",
  29550=>"110010010",
  29551=>"011111110",
  29552=>"111110110",
  29553=>"011100100",
  29554=>"111110100",
  29555=>"100101110",
  29556=>"111011101",
  29557=>"010101101",
  29558=>"000010101",
  29559=>"001101000",
  29560=>"000110001",
  29561=>"100010100",
  29562=>"011111001",
  29563=>"111110011",
  29564=>"010011000",
  29565=>"111111000",
  29566=>"010110111",
  29567=>"111101100",
  29568=>"111101100",
  29569=>"010010011",
  29570=>"100100010",
  29571=>"100000001",
  29572=>"110001011",
  29573=>"010101000",
  29574=>"001101110",
  29575=>"010100100",
  29576=>"111111110",
  29577=>"110101101",
  29578=>"001011111",
  29579=>"010101011",
  29580=>"100001011",
  29581=>"101111101",
  29582=>"000001011",
  29583=>"001100100",
  29584=>"101100001",
  29585=>"010100101",
  29586=>"000000100",
  29587=>"000000110",
  29588=>"001001011",
  29589=>"111000110",
  29590=>"000111111",
  29591=>"111101101",
  29592=>"011001111",
  29593=>"001010110",
  29594=>"010001111",
  29595=>"100011011",
  29596=>"110111001",
  29597=>"111101100",
  29598=>"100110101",
  29599=>"000011111",
  29600=>"111000001",
  29601=>"110001011",
  29602=>"111001111",
  29603=>"000000101",
  29604=>"000000100",
  29605=>"010010110",
  29606=>"101010100",
  29607=>"011001101",
  29608=>"110001000",
  29609=>"000111101",
  29610=>"011111111",
  29611=>"010100100",
  29612=>"111001101",
  29613=>"110111101",
  29614=>"101110101",
  29615=>"100001110",
  29616=>"110110010",
  29617=>"010111111",
  29618=>"100111100",
  29619=>"011111101",
  29620=>"110111000",
  29621=>"111110000",
  29622=>"110101111",
  29623=>"111010011",
  29624=>"010000101",
  29625=>"000001001",
  29626=>"011100101",
  29627=>"111110111",
  29628=>"110111101",
  29629=>"101101000",
  29630=>"100100000",
  29631=>"110111111",
  29632=>"011000001",
  29633=>"111101100",
  29634=>"100100011",
  29635=>"111100000",
  29636=>"101000001",
  29637=>"111000100",
  29638=>"111101111",
  29639=>"101000100",
  29640=>"000001010",
  29641=>"000011101",
  29642=>"001100010",
  29643=>"011010100",
  29644=>"101000100",
  29645=>"000000001",
  29646=>"000110001",
  29647=>"111100110",
  29648=>"111001100",
  29649=>"000111010",
  29650=>"001011111",
  29651=>"101000000",
  29652=>"010010110",
  29653=>"101001100",
  29654=>"100001101",
  29655=>"111001100",
  29656=>"000010000",
  29657=>"000110110",
  29658=>"011010011",
  29659=>"110000010",
  29660=>"000100000",
  29661=>"101111110",
  29662=>"010111110",
  29663=>"010000101",
  29664=>"000001000",
  29665=>"111001110",
  29666=>"011010010",
  29667=>"110110101",
  29668=>"000011000",
  29669=>"011100011",
  29670=>"101011110",
  29671=>"010000010",
  29672=>"001000000",
  29673=>"011001011",
  29674=>"101100000",
  29675=>"111100101",
  29676=>"001010110",
  29677=>"111001100",
  29678=>"011110000",
  29679=>"111000101",
  29680=>"001011001",
  29681=>"000000101",
  29682=>"001101001",
  29683=>"100000010",
  29684=>"101101100",
  29685=>"000110110",
  29686=>"111010011",
  29687=>"101111100",
  29688=>"001100101",
  29689=>"110000100",
  29690=>"010100100",
  29691=>"111100000",
  29692=>"111000100",
  29693=>"101000101",
  29694=>"101101000",
  29695=>"110011100",
  29696=>"111010101",
  29697=>"000010111",
  29698=>"100111101",
  29699=>"111001010",
  29700=>"111000001",
  29701=>"000011001",
  29702=>"001100011",
  29703=>"011101001",
  29704=>"011001101",
  29705=>"110001111",
  29706=>"000000000",
  29707=>"101010011",
  29708=>"110001100",
  29709=>"101000010",
  29710=>"001110101",
  29711=>"101100111",
  29712=>"101101110",
  29713=>"110100010",
  29714=>"000000010",
  29715=>"110100000",
  29716=>"000011111",
  29717=>"001011001",
  29718=>"011110101",
  29719=>"001101111",
  29720=>"100111000",
  29721=>"111010000",
  29722=>"000100100",
  29723=>"110000110",
  29724=>"010011000",
  29725=>"101110000",
  29726=>"000100111",
  29727=>"000010101",
  29728=>"100011000",
  29729=>"010100010",
  29730=>"101110001",
  29731=>"010010110",
  29732=>"010011111",
  29733=>"001010000",
  29734=>"000010001",
  29735=>"111000010",
  29736=>"000010101",
  29737=>"100011101",
  29738=>"111111011",
  29739=>"000111110",
  29740=>"101110000",
  29741=>"010000010",
  29742=>"110100001",
  29743=>"110011011",
  29744=>"011110001",
  29745=>"001101100",
  29746=>"100000100",
  29747=>"111111001",
  29748=>"111111100",
  29749=>"101111100",
  29750=>"010000010",
  29751=>"111010100",
  29752=>"110000110",
  29753=>"011011100",
  29754=>"001011101",
  29755=>"111111011",
  29756=>"101010100",
  29757=>"000000000",
  29758=>"100010011",
  29759=>"110110010",
  29760=>"000110000",
  29761=>"001001100",
  29762=>"110000111",
  29763=>"011001100",
  29764=>"100000101",
  29765=>"010010000",
  29766=>"000011011",
  29767=>"100111011",
  29768=>"110000101",
  29769=>"111001111",
  29770=>"010101000",
  29771=>"000110000",
  29772=>"111111011",
  29773=>"100001100",
  29774=>"100010110",
  29775=>"110000110",
  29776=>"000000001",
  29777=>"010011000",
  29778=>"011101010",
  29779=>"000010000",
  29780=>"100000100",
  29781=>"110100101",
  29782=>"100111111",
  29783=>"111100111",
  29784=>"110011100",
  29785=>"100000001",
  29786=>"111011111",
  29787=>"010010000",
  29788=>"010100111",
  29789=>"001010001",
  29790=>"110000110",
  29791=>"000110001",
  29792=>"001101010",
  29793=>"111111011",
  29794=>"110110011",
  29795=>"000000010",
  29796=>"000110011",
  29797=>"111000000",
  29798=>"100100100",
  29799=>"110110110",
  29800=>"100011100",
  29801=>"011011100",
  29802=>"100001011",
  29803=>"000110000",
  29804=>"101000101",
  29805=>"011011111",
  29806=>"010101001",
  29807=>"111100001",
  29808=>"011111100",
  29809=>"111101000",
  29810=>"100111101",
  29811=>"000101001",
  29812=>"000010010",
  29813=>"010011100",
  29814=>"000001010",
  29815=>"101001111",
  29816=>"000000011",
  29817=>"001111000",
  29818=>"011110000",
  29819=>"011000100",
  29820=>"100101110",
  29821=>"111011001",
  29822=>"010001010",
  29823=>"001001000",
  29824=>"111001001",
  29825=>"000110101",
  29826=>"100001100",
  29827=>"101100100",
  29828=>"011110011",
  29829=>"011111111",
  29830=>"110111000",
  29831=>"101000100",
  29832=>"001001100",
  29833=>"001010011",
  29834=>"110010110",
  29835=>"110111111",
  29836=>"010100011",
  29837=>"100010010",
  29838=>"111101001",
  29839=>"101111101",
  29840=>"010101100",
  29841=>"111100111",
  29842=>"101000111",
  29843=>"110110011",
  29844=>"001101101",
  29845=>"010100111",
  29846=>"111110100",
  29847=>"011100100",
  29848=>"000100000",
  29849=>"100101011",
  29850=>"010011010",
  29851=>"111011110",
  29852=>"101001110",
  29853=>"011101111",
  29854=>"100111011",
  29855=>"000001011",
  29856=>"000000000",
  29857=>"101111101",
  29858=>"101110001",
  29859=>"000101011",
  29860=>"011111000",
  29861=>"001000111",
  29862=>"000101001",
  29863=>"101010000",
  29864=>"111001100",
  29865=>"011011010",
  29866=>"110111001",
  29867=>"001100000",
  29868=>"101110010",
  29869=>"010111101",
  29870=>"001110010",
  29871=>"111010110",
  29872=>"010100111",
  29873=>"111011000",
  29874=>"010000010",
  29875=>"010101110",
  29876=>"110111111",
  29877=>"011111010",
  29878=>"110111001",
  29879=>"001101100",
  29880=>"011111111",
  29881=>"000011001",
  29882=>"000001100",
  29883=>"101010111",
  29884=>"111111101",
  29885=>"100010111",
  29886=>"000101001",
  29887=>"000000100",
  29888=>"000101100",
  29889=>"011001001",
  29890=>"011011000",
  29891=>"010001001",
  29892=>"111001000",
  29893=>"110011101",
  29894=>"111111011",
  29895=>"001101100",
  29896=>"100111001",
  29897=>"000010000",
  29898=>"100100101",
  29899=>"111100100",
  29900=>"110100100",
  29901=>"101100100",
  29902=>"011100111",
  29903=>"111011111",
  29904=>"100100101",
  29905=>"111001111",
  29906=>"000101101",
  29907=>"001000000",
  29908=>"100110100",
  29909=>"010111011",
  29910=>"001011111",
  29911=>"111000000",
  29912=>"110000010",
  29913=>"001110111",
  29914=>"000101110",
  29915=>"011001011",
  29916=>"000001011",
  29917=>"101010111",
  29918=>"011010011",
  29919=>"100100000",
  29920=>"000111110",
  29921=>"100111001",
  29922=>"000001000",
  29923=>"000010000",
  29924=>"000110000",
  29925=>"010101100",
  29926=>"100011000",
  29927=>"101110101",
  29928=>"011010000",
  29929=>"010011110",
  29930=>"111001000",
  29931=>"011010000",
  29932=>"000110001",
  29933=>"001111110",
  29934=>"110000000",
  29935=>"111111111",
  29936=>"011000111",
  29937=>"001101001",
  29938=>"011100101",
  29939=>"111010010",
  29940=>"010001000",
  29941=>"101010010",
  29942=>"000001000",
  29943=>"110111000",
  29944=>"101000110",
  29945=>"001110100",
  29946=>"001110110",
  29947=>"010101111",
  29948=>"100010110",
  29949=>"000111001",
  29950=>"111101000",
  29951=>"111110010",
  29952=>"010111100",
  29953=>"000010010",
  29954=>"101110111",
  29955=>"110011111",
  29956=>"001110010",
  29957=>"010000111",
  29958=>"100100001",
  29959=>"101111001",
  29960=>"101110010",
  29961=>"011010101",
  29962=>"101100011",
  29963=>"000111110",
  29964=>"011101000",
  29965=>"110000011",
  29966=>"011001011",
  29967=>"001011001",
  29968=>"111100000",
  29969=>"110110010",
  29970=>"101100011",
  29971=>"111010111",
  29972=>"110011101",
  29973=>"110100101",
  29974=>"111000000",
  29975=>"111011000",
  29976=>"111001110",
  29977=>"100101011",
  29978=>"011001000",
  29979=>"011110111",
  29980=>"000011000",
  29981=>"110110100",
  29982=>"010110010",
  29983=>"111101011",
  29984=>"010011000",
  29985=>"010100010",
  29986=>"001000110",
  29987=>"101101111",
  29988=>"000001000",
  29989=>"011010000",
  29990=>"110111001",
  29991=>"011111100",
  29992=>"101110111",
  29993=>"100010111",
  29994=>"001001110",
  29995=>"011100101",
  29996=>"111111101",
  29997=>"110111111",
  29998=>"011100000",
  29999=>"111010000",
  30000=>"000001110",
  30001=>"000010110",
  30002=>"001110101",
  30003=>"100001001",
  30004=>"001100011",
  30005=>"000010110",
  30006=>"000001100",
  30007=>"011011110",
  30008=>"101000010",
  30009=>"111001100",
  30010=>"000011011",
  30011=>"111011100",
  30012=>"001101111",
  30013=>"011000000",
  30014=>"011000111",
  30015=>"010011011",
  30016=>"000101101",
  30017=>"011000000",
  30018=>"110001010",
  30019=>"100100100",
  30020=>"101101011",
  30021=>"010101110",
  30022=>"001001010",
  30023=>"010000100",
  30024=>"100001100",
  30025=>"100100110",
  30026=>"100010111",
  30027=>"101110111",
  30028=>"010100101",
  30029=>"001011100",
  30030=>"101000001",
  30031=>"011000001",
  30032=>"000000110",
  30033=>"000111101",
  30034=>"110110111",
  30035=>"001000010",
  30036=>"011110100",
  30037=>"110011111",
  30038=>"110111001",
  30039=>"111100110",
  30040=>"111100010",
  30041=>"000000101",
  30042=>"011100100",
  30043=>"000111010",
  30044=>"101000010",
  30045=>"101001100",
  30046=>"001011011",
  30047=>"001001010",
  30048=>"101010001",
  30049=>"000000010",
  30050=>"001100110",
  30051=>"100110011",
  30052=>"110101101",
  30053=>"011011011",
  30054=>"011101110",
  30055=>"110110100",
  30056=>"001000110",
  30057=>"111000111",
  30058=>"111111101",
  30059=>"100111011",
  30060=>"111100111",
  30061=>"010001000",
  30062=>"111011000",
  30063=>"100111010",
  30064=>"100100010",
  30065=>"001110010",
  30066=>"001001111",
  30067=>"010100100",
  30068=>"100000110",
  30069=>"000000111",
  30070=>"000100101",
  30071=>"001110001",
  30072=>"110000001",
  30073=>"110000001",
  30074=>"101001011",
  30075=>"100000100",
  30076=>"010100000",
  30077=>"011001011",
  30078=>"011101011",
  30079=>"000001001",
  30080=>"111111101",
  30081=>"101100001",
  30082=>"001011010",
  30083=>"100010010",
  30084=>"010110111",
  30085=>"100101100",
  30086=>"011100011",
  30087=>"011000100",
  30088=>"111011110",
  30089=>"001000000",
  30090=>"111011111",
  30091=>"001000010",
  30092=>"001101110",
  30093=>"010101100",
  30094=>"011111101",
  30095=>"100011100",
  30096=>"110001000",
  30097=>"000001111",
  30098=>"000000100",
  30099=>"100110010",
  30100=>"001001001",
  30101=>"101010011",
  30102=>"111100101",
  30103=>"101101001",
  30104=>"111111101",
  30105=>"100010000",
  30106=>"010010101",
  30107=>"100001010",
  30108=>"011101011",
  30109=>"011000001",
  30110=>"100100110",
  30111=>"000011110",
  30112=>"111001101",
  30113=>"001101011",
  30114=>"110100000",
  30115=>"111111010",
  30116=>"111001101",
  30117=>"011000000",
  30118=>"000101100",
  30119=>"000101011",
  30120=>"000000111",
  30121=>"010101000",
  30122=>"111101100",
  30123=>"111010101",
  30124=>"001111000",
  30125=>"110000101",
  30126=>"101111101",
  30127=>"001100001",
  30128=>"000010010",
  30129=>"011010110",
  30130=>"101001101",
  30131=>"010010010",
  30132=>"101011111",
  30133=>"010000110",
  30134=>"000000101",
  30135=>"111100110",
  30136=>"011101100",
  30137=>"111000111",
  30138=>"101111111",
  30139=>"100110100",
  30140=>"001000111",
  30141=>"100110010",
  30142=>"101110111",
  30143=>"100110010",
  30144=>"111010001",
  30145=>"000101111",
  30146=>"100011110",
  30147=>"010101111",
  30148=>"111111011",
  30149=>"101010101",
  30150=>"011110100",
  30151=>"101010000",
  30152=>"101101011",
  30153=>"000010110",
  30154=>"001111100",
  30155=>"000111001",
  30156=>"000011011",
  30157=>"010001111",
  30158=>"011101111",
  30159=>"011000001",
  30160=>"001111011",
  30161=>"110000110",
  30162=>"111101101",
  30163=>"100100000",
  30164=>"101001101",
  30165=>"111000110",
  30166=>"100011110",
  30167=>"111010100",
  30168=>"001000001",
  30169=>"001111101",
  30170=>"110110110",
  30171=>"111001010",
  30172=>"111000110",
  30173=>"100000110",
  30174=>"000000000",
  30175=>"000110001",
  30176=>"110111000",
  30177=>"000110101",
  30178=>"101100110",
  30179=>"010000011",
  30180=>"110100100",
  30181=>"000110101",
  30182=>"000010000",
  30183=>"110000011",
  30184=>"001111101",
  30185=>"010111011",
  30186=>"111000010",
  30187=>"100101010",
  30188=>"001110011",
  30189=>"101110010",
  30190=>"001101010",
  30191=>"101100000",
  30192=>"100000011",
  30193=>"001111010",
  30194=>"001001011",
  30195=>"100010001",
  30196=>"101001010",
  30197=>"001000100",
  30198=>"110110110",
  30199=>"010001111",
  30200=>"101101110",
  30201=>"100111110",
  30202=>"001001101",
  30203=>"001010000",
  30204=>"111010110",
  30205=>"001111010",
  30206=>"010010110",
  30207=>"011110011",
  30208=>"000111010",
  30209=>"001001100",
  30210=>"100110110",
  30211=>"110101001",
  30212=>"111101111",
  30213=>"010110011",
  30214=>"100100011",
  30215=>"110001100",
  30216=>"001001010",
  30217=>"110001011",
  30218=>"011110001",
  30219=>"000011001",
  30220=>"100010010",
  30221=>"100000000",
  30222=>"111001111",
  30223=>"011010110",
  30224=>"111010101",
  30225=>"001110001",
  30226=>"010100101",
  30227=>"110110100",
  30228=>"110101011",
  30229=>"000101111",
  30230=>"011101001",
  30231=>"111111011",
  30232=>"100101110",
  30233=>"111010011",
  30234=>"101010101",
  30235=>"001001000",
  30236=>"001111101",
  30237=>"101001100",
  30238=>"011010010",
  30239=>"100001100",
  30240=>"010000110",
  30241=>"010101000",
  30242=>"101100001",
  30243=>"100011110",
  30244=>"110011001",
  30245=>"110000010",
  30246=>"011100100",
  30247=>"111111111",
  30248=>"110001101",
  30249=>"101001100",
  30250=>"001000001",
  30251=>"110101110",
  30252=>"100111100",
  30253=>"000101111",
  30254=>"000110110",
  30255=>"011100000",
  30256=>"110100001",
  30257=>"111111111",
  30258=>"111000011",
  30259=>"001011100",
  30260=>"110101011",
  30261=>"111100001",
  30262=>"000100111",
  30263=>"000001100",
  30264=>"111110000",
  30265=>"101100011",
  30266=>"100111101",
  30267=>"100111110",
  30268=>"010110100",
  30269=>"110001010",
  30270=>"111010011",
  30271=>"010010010",
  30272=>"101000111",
  30273=>"001101100",
  30274=>"110101000",
  30275=>"110110000",
  30276=>"110100010",
  30277=>"011111100",
  30278=>"000000001",
  30279=>"101001001",
  30280=>"111010001",
  30281=>"010011101",
  30282=>"111110111",
  30283=>"001001100",
  30284=>"011010110",
  30285=>"000101100",
  30286=>"010100000",
  30287=>"101010111",
  30288=>"001000000",
  30289=>"000000111",
  30290=>"000101000",
  30291=>"100000001",
  30292=>"000010111",
  30293=>"000000100",
  30294=>"111101010",
  30295=>"110101001",
  30296=>"000000101",
  30297=>"001010010",
  30298=>"001011111",
  30299=>"010000011",
  30300=>"110011001",
  30301=>"001101001",
  30302=>"011100000",
  30303=>"010111000",
  30304=>"101111000",
  30305=>"011110011",
  30306=>"110001110",
  30307=>"000001110",
  30308=>"101000100",
  30309=>"001100100",
  30310=>"101011001",
  30311=>"110011111",
  30312=>"000011010",
  30313=>"111010100",
  30314=>"110010101",
  30315=>"011000010",
  30316=>"011000111",
  30317=>"010000000",
  30318=>"100010000",
  30319=>"010011010",
  30320=>"110101001",
  30321=>"000100010",
  30322=>"111001110",
  30323=>"000010000",
  30324=>"000100000",
  30325=>"100000001",
  30326=>"110000000",
  30327=>"001100010",
  30328=>"110111111",
  30329=>"000111000",
  30330=>"101011111",
  30331=>"001000000",
  30332=>"110101110",
  30333=>"100011111",
  30334=>"110011000",
  30335=>"100001001",
  30336=>"101001001",
  30337=>"111110011",
  30338=>"100101000",
  30339=>"010010000",
  30340=>"010111000",
  30341=>"110001111",
  30342=>"011010101",
  30343=>"100011010",
  30344=>"001100110",
  30345=>"001101101",
  30346=>"111010100",
  30347=>"001011000",
  30348=>"001000000",
  30349=>"010111111",
  30350=>"111101111",
  30351=>"000000100",
  30352=>"010000011",
  30353=>"001111110",
  30354=>"100010010",
  30355=>"010001100",
  30356=>"011110110",
  30357=>"111100010",
  30358=>"000101011",
  30359=>"000001101",
  30360=>"111000111",
  30361=>"110100101",
  30362=>"000100001",
  30363=>"101101101",
  30364=>"100011101",
  30365=>"101101111",
  30366=>"010100000",
  30367=>"111001010",
  30368=>"000010011",
  30369=>"110111101",
  30370=>"010101110",
  30371=>"011111101",
  30372=>"111011111",
  30373=>"001100010",
  30374=>"111110000",
  30375=>"001110010",
  30376=>"110010111",
  30377=>"011011111",
  30378=>"101111101",
  30379=>"011011001",
  30380=>"100100010",
  30381=>"001110011",
  30382=>"100100101",
  30383=>"011110010",
  30384=>"011010010",
  30385=>"011000000",
  30386=>"111011010",
  30387=>"100111110",
  30388=>"100001000",
  30389=>"010110110",
  30390=>"101111111",
  30391=>"100000001",
  30392=>"101001100",
  30393=>"100011011",
  30394=>"101000100",
  30395=>"000000101",
  30396=>"100000101",
  30397=>"100000010",
  30398=>"000011010",
  30399=>"110101111",
  30400=>"000100100",
  30401=>"011110010",
  30402=>"001001110",
  30403=>"111111111",
  30404=>"100011001",
  30405=>"111110000",
  30406=>"100010001",
  30407=>"100101010",
  30408=>"011110110",
  30409=>"100110001",
  30410=>"000001010",
  30411=>"000001111",
  30412=>"000011011",
  30413=>"011001101",
  30414=>"001011010",
  30415=>"111110010",
  30416=>"101001000",
  30417=>"011010101",
  30418=>"101111111",
  30419=>"011011001",
  30420=>"100001000",
  30421=>"010001111",
  30422=>"110010010",
  30423=>"000100011",
  30424=>"011100000",
  30425=>"000000111",
  30426=>"001001110",
  30427=>"101110001",
  30428=>"011111000",
  30429=>"010100100",
  30430=>"100100110",
  30431=>"111100000",
  30432=>"000000000",
  30433=>"000001100",
  30434=>"011111010",
  30435=>"010010001",
  30436=>"000010111",
  30437=>"110110110",
  30438=>"111111111",
  30439=>"001100111",
  30440=>"000000001",
  30441=>"111100111",
  30442=>"011111110",
  30443=>"110111011",
  30444=>"000001111",
  30445=>"111110111",
  30446=>"000111101",
  30447=>"110111011",
  30448=>"011100000",
  30449=>"011001001",
  30450=>"000110000",
  30451=>"011110111",
  30452=>"100111110",
  30453=>"100010111",
  30454=>"000001001",
  30455=>"110111111",
  30456=>"111101111",
  30457=>"000001001",
  30458=>"100001100",
  30459=>"110001011",
  30460=>"010010101",
  30461=>"000011000",
  30462=>"010100110",
  30463=>"001010010",
  30464=>"100100100",
  30465=>"110010111",
  30466=>"011111000",
  30467=>"111110000",
  30468=>"101111001",
  30469=>"100101001",
  30470=>"001100101",
  30471=>"101000001",
  30472=>"100000111",
  30473=>"111111101",
  30474=>"011110111",
  30475=>"111110010",
  30476=>"010001010",
  30477=>"100000000",
  30478=>"101001100",
  30479=>"000111100",
  30480=>"000011100",
  30481=>"000000100",
  30482=>"101110001",
  30483=>"111000011",
  30484=>"100001101",
  30485=>"100110011",
  30486=>"011111111",
  30487=>"100101100",
  30488=>"101001011",
  30489=>"000010000",
  30490=>"000101011",
  30491=>"010000000",
  30492=>"011000110",
  30493=>"001100100",
  30494=>"000001000",
  30495=>"111101100",
  30496=>"111100110",
  30497=>"100001000",
  30498=>"001111011",
  30499=>"100101110",
  30500=>"101000100",
  30501=>"001011101",
  30502=>"000101110",
  30503=>"111110110",
  30504=>"111010011",
  30505=>"010111011",
  30506=>"110011011",
  30507=>"001101000",
  30508=>"010011111",
  30509=>"010010010",
  30510=>"001100010",
  30511=>"001110100",
  30512=>"101101000",
  30513=>"100110010",
  30514=>"000101100",
  30515=>"100000010",
  30516=>"101010010",
  30517=>"111110011",
  30518=>"100001110",
  30519=>"111010110",
  30520=>"101000111",
  30521=>"011100011",
  30522=>"001011010",
  30523=>"011010000",
  30524=>"000011111",
  30525=>"111000001",
  30526=>"111100101",
  30527=>"000100011",
  30528=>"100001000",
  30529=>"111100001",
  30530=>"111100001",
  30531=>"101001110",
  30532=>"001010101",
  30533=>"011110001",
  30534=>"110110011",
  30535=>"000000011",
  30536=>"110011000",
  30537=>"111111110",
  30538=>"111011000",
  30539=>"101100100",
  30540=>"100110001",
  30541=>"010001101",
  30542=>"110011101",
  30543=>"000011110",
  30544=>"111100100",
  30545=>"101100100",
  30546=>"100111110",
  30547=>"000100011",
  30548=>"000010101",
  30549=>"000110101",
  30550=>"000100110",
  30551=>"010110100",
  30552=>"111000111",
  30553=>"110001011",
  30554=>"110000110",
  30555=>"110000011",
  30556=>"100011110",
  30557=>"100101011",
  30558=>"101100011",
  30559=>"000000100",
  30560=>"110101100",
  30561=>"111110011",
  30562=>"100111001",
  30563=>"110011100",
  30564=>"011001011",
  30565=>"011111101",
  30566=>"101100101",
  30567=>"111000101",
  30568=>"111101000",
  30569=>"110010010",
  30570=>"001011011",
  30571=>"110101110",
  30572=>"011110011",
  30573=>"110100000",
  30574=>"010101101",
  30575=>"100101000",
  30576=>"010001000",
  30577=>"111111100",
  30578=>"100100001",
  30579=>"100011011",
  30580=>"010010100",
  30581=>"101011100",
  30582=>"010110111",
  30583=>"100100100",
  30584=>"000011001",
  30585=>"000001001",
  30586=>"101111111",
  30587=>"000001000",
  30588=>"111010101",
  30589=>"110100110",
  30590=>"111000111",
  30591=>"010101010",
  30592=>"000001010",
  30593=>"110100100",
  30594=>"011110101",
  30595=>"011110000",
  30596=>"000000000",
  30597=>"111111011",
  30598=>"110101111",
  30599=>"101000011",
  30600=>"101111101",
  30601=>"010010000",
  30602=>"000000011",
  30603=>"110010101",
  30604=>"010100001",
  30605=>"010100000",
  30606=>"011010000",
  30607=>"010001000",
  30608=>"111000011",
  30609=>"001110000",
  30610=>"111000011",
  30611=>"111000100",
  30612=>"110000010",
  30613=>"100000100",
  30614=>"011010001",
  30615=>"110111000",
  30616=>"111110010",
  30617=>"111011100",
  30618=>"000000010",
  30619=>"000000001",
  30620=>"011110111",
  30621=>"100011111",
  30622=>"100101010",
  30623=>"010011110",
  30624=>"001110011",
  30625=>"111001000",
  30626=>"011010100",
  30627=>"011110111",
  30628=>"101110001",
  30629=>"011111010",
  30630=>"001010010",
  30631=>"010010010",
  30632=>"010000011",
  30633=>"111001101",
  30634=>"100010011",
  30635=>"100100010",
  30636=>"100110010",
  30637=>"101000100",
  30638=>"010100001",
  30639=>"001011001",
  30640=>"100001011",
  30641=>"110101000",
  30642=>"000010010",
  30643=>"000101100",
  30644=>"010000000",
  30645=>"100001010",
  30646=>"000100101",
  30647=>"101110111",
  30648=>"101111001",
  30649=>"110110001",
  30650=>"000110101",
  30651=>"011111111",
  30652=>"011101000",
  30653=>"000011010",
  30654=>"110110111",
  30655=>"000000100",
  30656=>"101111011",
  30657=>"111111000",
  30658=>"111010111",
  30659=>"110001010",
  30660=>"111100101",
  30661=>"000111101",
  30662=>"001100001",
  30663=>"010110111",
  30664=>"010001011",
  30665=>"101111111",
  30666=>"001000110",
  30667=>"011110010",
  30668=>"110010010",
  30669=>"111010110",
  30670=>"011010110",
  30671=>"011111101",
  30672=>"001010011",
  30673=>"011010001",
  30674=>"101100111",
  30675=>"100110001",
  30676=>"001010100",
  30677=>"010100111",
  30678=>"110101100",
  30679=>"011000101",
  30680=>"001000100",
  30681=>"111110011",
  30682=>"011111111",
  30683=>"110000011",
  30684=>"110010010",
  30685=>"001001000",
  30686=>"010000010",
  30687=>"100111001",
  30688=>"100110101",
  30689=>"000111001",
  30690=>"001001101",
  30691=>"000111111",
  30692=>"011001001",
  30693=>"101100010",
  30694=>"000001001",
  30695=>"011110101",
  30696=>"001001011",
  30697=>"011111110",
  30698=>"000000100",
  30699=>"011101111",
  30700=>"001000110",
  30701=>"110100011",
  30702=>"111001100",
  30703=>"010010101",
  30704=>"010000001",
  30705=>"110110000",
  30706=>"111100000",
  30707=>"100011110",
  30708=>"001100010",
  30709=>"100010110",
  30710=>"011010001",
  30711=>"000001000",
  30712=>"110111010",
  30713=>"011111001",
  30714=>"001001110",
  30715=>"111100100",
  30716=>"010011001",
  30717=>"011000101",
  30718=>"101110101",
  30719=>"000011101",
  30720=>"110011000",
  30721=>"101011100",
  30722=>"110101110",
  30723=>"100001111",
  30724=>"001111011",
  30725=>"101101010",
  30726=>"011111001",
  30727=>"000110101",
  30728=>"100111110",
  30729=>"100100101",
  30730=>"101000100",
  30731=>"100101011",
  30732=>"111101101",
  30733=>"100110001",
  30734=>"111111001",
  30735=>"001100011",
  30736=>"011000000",
  30737=>"010100001",
  30738=>"001011110",
  30739=>"001000000",
  30740=>"000000101",
  30741=>"110111010",
  30742=>"111111110",
  30743=>"000101101",
  30744=>"011010001",
  30745=>"101101100",
  30746=>"110100010",
  30747=>"111011011",
  30748=>"100110011",
  30749=>"110101001",
  30750=>"001011110",
  30751=>"000010001",
  30752=>"101010111",
  30753=>"011011010",
  30754=>"110110010",
  30755=>"000000001",
  30756=>"001101110",
  30757=>"000010110",
  30758=>"010001011",
  30759=>"110110111",
  30760=>"100100000",
  30761=>"010010100",
  30762=>"000111111",
  30763=>"010101111",
  30764=>"010111101",
  30765=>"011000111",
  30766=>"111001110",
  30767=>"001010000",
  30768=>"000100110",
  30769=>"110000000",
  30770=>"011000001",
  30771=>"111111110",
  30772=>"100111111",
  30773=>"111011101",
  30774=>"001100100",
  30775=>"101101111",
  30776=>"111011011",
  30777=>"100000000",
  30778=>"111111010",
  30779=>"100011010",
  30780=>"110001100",
  30781=>"111111010",
  30782=>"010000100",
  30783=>"000001000",
  30784=>"001110011",
  30785=>"100100010",
  30786=>"100001000",
  30787=>"011101010",
  30788=>"111010100",
  30789=>"010111111",
  30790=>"101001101",
  30791=>"010101000",
  30792=>"101101010",
  30793=>"100000111",
  30794=>"000011010",
  30795=>"101011110",
  30796=>"011010100",
  30797=>"111100101",
  30798=>"111011110",
  30799=>"101001010",
  30800=>"001100000",
  30801=>"000001100",
  30802=>"011001010",
  30803=>"111100110",
  30804=>"100010010",
  30805=>"010100010",
  30806=>"010110110",
  30807=>"110100001",
  30808=>"101111001",
  30809=>"011100101",
  30810=>"100011000",
  30811=>"010001100",
  30812=>"001000111",
  30813=>"100101101",
  30814=>"000001000",
  30815=>"001111110",
  30816=>"001000100",
  30817=>"111000001",
  30818=>"011101001",
  30819=>"101010110",
  30820=>"111101010",
  30821=>"100010111",
  30822=>"001100000",
  30823=>"100011000",
  30824=>"011001101",
  30825=>"111000100",
  30826=>"010110111",
  30827=>"010101000",
  30828=>"101101101",
  30829=>"010101011",
  30830=>"100011111",
  30831=>"001101010",
  30832=>"110111101",
  30833=>"101011101",
  30834=>"011101110",
  30835=>"101010001",
  30836=>"001011110",
  30837=>"111001011",
  30838=>"111100101",
  30839=>"100110110",
  30840=>"000111100",
  30841=>"000001000",
  30842=>"011000101",
  30843=>"001011011",
  30844=>"001001110",
  30845=>"000001110",
  30846=>"110100011",
  30847=>"101011001",
  30848=>"010001010",
  30849=>"001000011",
  30850=>"111011001",
  30851=>"111100111",
  30852=>"111101100",
  30853=>"011001110",
  30854=>"111010000",
  30855=>"100111010",
  30856=>"010010010",
  30857=>"110000111",
  30858=>"010100100",
  30859=>"011011011",
  30860=>"010110111",
  30861=>"100001100",
  30862=>"111100101",
  30863=>"101001010",
  30864=>"101111110",
  30865=>"010010011",
  30866=>"011001101",
  30867=>"101111001",
  30868=>"000010001",
  30869=>"111000111",
  30870=>"101010110",
  30871=>"100011011",
  30872=>"011001111",
  30873=>"011010000",
  30874=>"100110111",
  30875=>"101000000",
  30876=>"101010010",
  30877=>"001011000",
  30878=>"000000100",
  30879=>"001010001",
  30880=>"101101011",
  30881=>"000001111",
  30882=>"011100110",
  30883=>"100110011",
  30884=>"001101000",
  30885=>"110011110",
  30886=>"000101000",
  30887=>"111111011",
  30888=>"011000111",
  30889=>"110011011",
  30890=>"110100000",
  30891=>"101101100",
  30892=>"001011110",
  30893=>"101100110",
  30894=>"000111000",
  30895=>"011011101",
  30896=>"111100010",
  30897=>"101000110",
  30898=>"101100101",
  30899=>"000011110",
  30900=>"001001000",
  30901=>"111010110",
  30902=>"011111011",
  30903=>"110010001",
  30904=>"000010010",
  30905=>"011111011",
  30906=>"011100000",
  30907=>"111101011",
  30908=>"111000111",
  30909=>"101000001",
  30910=>"111000000",
  30911=>"111011101",
  30912=>"100111011",
  30913=>"111111001",
  30914=>"000101110",
  30915=>"111111101",
  30916=>"011001110",
  30917=>"001001000",
  30918=>"001000001",
  30919=>"011000101",
  30920=>"111011010",
  30921=>"000001110",
  30922=>"110110001",
  30923=>"001000110",
  30924=>"101111010",
  30925=>"101101011",
  30926=>"000101111",
  30927=>"010001101",
  30928=>"110111100",
  30929=>"001010101",
  30930=>"000001000",
  30931=>"001101011",
  30932=>"111011011",
  30933=>"000111101",
  30934=>"001000000",
  30935=>"110011010",
  30936=>"100101000",
  30937=>"001001010",
  30938=>"001110100",
  30939=>"010100001",
  30940=>"000010011",
  30941=>"011101010",
  30942=>"111101101",
  30943=>"111011011",
  30944=>"100000100",
  30945=>"010010101",
  30946=>"101010011",
  30947=>"001001011",
  30948=>"011101100",
  30949=>"101000011",
  30950=>"011010010",
  30951=>"111101001",
  30952=>"111001110",
  30953=>"110111011",
  30954=>"001000011",
  30955=>"100001000",
  30956=>"111011000",
  30957=>"110010001",
  30958=>"100101101",
  30959=>"001000000",
  30960=>"001110111",
  30961=>"001111010",
  30962=>"101000001",
  30963=>"010101010",
  30964=>"110001111",
  30965=>"110010111",
  30966=>"100001000",
  30967=>"111100000",
  30968=>"001001101",
  30969=>"011111000",
  30970=>"000011110",
  30971=>"001101011",
  30972=>"111111010",
  30973=>"011111111",
  30974=>"111101110",
  30975=>"000111110",
  30976=>"101101010",
  30977=>"000110000",
  30978=>"110010011",
  30979=>"011110000",
  30980=>"011111111",
  30981=>"101000001",
  30982=>"000011000",
  30983=>"110111101",
  30984=>"101001101",
  30985=>"111111111",
  30986=>"011110110",
  30987=>"100110100",
  30988=>"001000011",
  30989=>"110000000",
  30990=>"111111111",
  30991=>"001011100",
  30992=>"010001011",
  30993=>"111101011",
  30994=>"010001000",
  30995=>"000100110",
  30996=>"110111111",
  30997=>"001000101",
  30998=>"110000001",
  30999=>"101011010",
  31000=>"101111110",
  31001=>"111111100",
  31002=>"110100010",
  31003=>"111111001",
  31004=>"010000110",
  31005=>"000100110",
  31006=>"110110011",
  31007=>"101001101",
  31008=>"100000000",
  31009=>"100011011",
  31010=>"100000000",
  31011=>"101010101",
  31012=>"010100001",
  31013=>"101010100",
  31014=>"001001110",
  31015=>"011000101",
  31016=>"000000110",
  31017=>"010001110",
  31018=>"110101000",
  31019=>"100000101",
  31020=>"001001001",
  31021=>"000000000",
  31022=>"010100110",
  31023=>"100000010",
  31024=>"011001100",
  31025=>"110011000",
  31026=>"101100011",
  31027=>"100010000",
  31028=>"011010100",
  31029=>"011000000",
  31030=>"111001010",
  31031=>"111100000",
  31032=>"001011001",
  31033=>"111000001",
  31034=>"000010010",
  31035=>"001100010",
  31036=>"111110110",
  31037=>"010110110",
  31038=>"011010000",
  31039=>"111111010",
  31040=>"000000001",
  31041=>"011100001",
  31042=>"111111010",
  31043=>"010101110",
  31044=>"000100110",
  31045=>"110100010",
  31046=>"110001011",
  31047=>"101110101",
  31048=>"000010010",
  31049=>"000010110",
  31050=>"001010011",
  31051=>"010110110",
  31052=>"010110111",
  31053=>"011001111",
  31054=>"100110010",
  31055=>"100011000",
  31056=>"110111101",
  31057=>"000001101",
  31058=>"000001000",
  31059=>"001110101",
  31060=>"011000011",
  31061=>"010011000",
  31062=>"101101110",
  31063=>"101111110",
  31064=>"100111011",
  31065=>"010010101",
  31066=>"110001110",
  31067=>"110000001",
  31068=>"001101010",
  31069=>"001100001",
  31070=>"111010010",
  31071=>"000001010",
  31072=>"111000110",
  31073=>"000110001",
  31074=>"000111001",
  31075=>"011001101",
  31076=>"101101111",
  31077=>"111100011",
  31078=>"000101000",
  31079=>"100010001",
  31080=>"001101111",
  31081=>"001000101",
  31082=>"111110101",
  31083=>"100100001",
  31084=>"000101101",
  31085=>"001000011",
  31086=>"111000011",
  31087=>"000100000",
  31088=>"111011000",
  31089=>"000010000",
  31090=>"010110000",
  31091=>"110100110",
  31092=>"101111011",
  31093=>"010000111",
  31094=>"100000111",
  31095=>"111000101",
  31096=>"101000100",
  31097=>"100101101",
  31098=>"011110010",
  31099=>"110111001",
  31100=>"100100010",
  31101=>"101001000",
  31102=>"000100010",
  31103=>"110000001",
  31104=>"000001010",
  31105=>"110001101",
  31106=>"001001011",
  31107=>"000101010",
  31108=>"101101101",
  31109=>"110110010",
  31110=>"010001000",
  31111=>"000000010",
  31112=>"111101000",
  31113=>"111011111",
  31114=>"011000100",
  31115=>"100011100",
  31116=>"000110101",
  31117=>"110100010",
  31118=>"000100101",
  31119=>"100011010",
  31120=>"010000111",
  31121=>"101101000",
  31122=>"111010111",
  31123=>"001111011",
  31124=>"000001101",
  31125=>"100110001",
  31126=>"000010000",
  31127=>"110000101",
  31128=>"100011101",
  31129=>"100000000",
  31130=>"101000011",
  31131=>"011001010",
  31132=>"111011010",
  31133=>"101000101",
  31134=>"101111010",
  31135=>"110110000",
  31136=>"011001011",
  31137=>"011000110",
  31138=>"101111111",
  31139=>"111000001",
  31140=>"011100101",
  31141=>"100110100",
  31142=>"010111001",
  31143=>"011101011",
  31144=>"110101001",
  31145=>"100001111",
  31146=>"000000100",
  31147=>"111000101",
  31148=>"000000010",
  31149=>"110000110",
  31150=>"111100110",
  31151=>"110111001",
  31152=>"011101111",
  31153=>"011110000",
  31154=>"101110000",
  31155=>"101010011",
  31156=>"011010111",
  31157=>"110110110",
  31158=>"110001101",
  31159=>"111010110",
  31160=>"001110100",
  31161=>"001001000",
  31162=>"000010101",
  31163=>"001011101",
  31164=>"000011011",
  31165=>"110000010",
  31166=>"011001110",
  31167=>"100111010",
  31168=>"111111111",
  31169=>"001110010",
  31170=>"011100001",
  31171=>"101011010",
  31172=>"011110011",
  31173=>"110111110",
  31174=>"110110110",
  31175=>"111001010",
  31176=>"001111011",
  31177=>"000001010",
  31178=>"100101110",
  31179=>"010100100",
  31180=>"000101010",
  31181=>"101011010",
  31182=>"001111101",
  31183=>"001100100",
  31184=>"110100111",
  31185=>"001010001",
  31186=>"110010011",
  31187=>"000010011",
  31188=>"001001000",
  31189=>"000111011",
  31190=>"000001001",
  31191=>"110001011",
  31192=>"010110110",
  31193=>"100110011",
  31194=>"010110001",
  31195=>"101110000",
  31196=>"100000011",
  31197=>"111001110",
  31198=>"000110001",
  31199=>"010101111",
  31200=>"000001000",
  31201=>"000001110",
  31202=>"111111000",
  31203=>"101000011",
  31204=>"011001001",
  31205=>"011011100",
  31206=>"010100001",
  31207=>"111011000",
  31208=>"111111111",
  31209=>"011011010",
  31210=>"100100100",
  31211=>"101100011",
  31212=>"001100110",
  31213=>"011010110",
  31214=>"000000011",
  31215=>"001001100",
  31216=>"111001111",
  31217=>"100101011",
  31218=>"111101100",
  31219=>"000011010",
  31220=>"010110111",
  31221=>"110010010",
  31222=>"100010000",
  31223=>"010100011",
  31224=>"110000110",
  31225=>"111110000",
  31226=>"101101000",
  31227=>"000100000",
  31228=>"000110100",
  31229=>"110000101",
  31230=>"101010111",
  31231=>"111101001",
  31232=>"011101111",
  31233=>"111100111",
  31234=>"001110011",
  31235=>"011101001",
  31236=>"011110111",
  31237=>"100001011",
  31238=>"101010000",
  31239=>"101001000",
  31240=>"001101011",
  31241=>"101110101",
  31242=>"000001010",
  31243=>"010100111",
  31244=>"000001011",
  31245=>"010101011",
  31246=>"010010000",
  31247=>"110110001",
  31248=>"101011101",
  31249=>"110100010",
  31250=>"111010100",
  31251=>"100001010",
  31252=>"111010000",
  31253=>"111111011",
  31254=>"000011000",
  31255=>"101011100",
  31256=>"001001011",
  31257=>"001011000",
  31258=>"111101011",
  31259=>"010111101",
  31260=>"111010010",
  31261=>"110011000",
  31262=>"010011001",
  31263=>"101100110",
  31264=>"011011111",
  31265=>"111011000",
  31266=>"101101001",
  31267=>"010010001",
  31268=>"011000110",
  31269=>"010110101",
  31270=>"101011000",
  31271=>"011011101",
  31272=>"000111100",
  31273=>"010111010",
  31274=>"111000000",
  31275=>"000000010",
  31276=>"100010001",
  31277=>"101101001",
  31278=>"001101100",
  31279=>"001000100",
  31280=>"010101000",
  31281=>"011111101",
  31282=>"100111011",
  31283=>"000101000",
  31284=>"001000011",
  31285=>"110110100",
  31286=>"010101000",
  31287=>"101001111",
  31288=>"011110100",
  31289=>"011000101",
  31290=>"100001100",
  31291=>"110110111",
  31292=>"110110100",
  31293=>"100110010",
  31294=>"001001111",
  31295=>"001101010",
  31296=>"001001001",
  31297=>"010010001",
  31298=>"001101100",
  31299=>"001000011",
  31300=>"010010100",
  31301=>"000100001",
  31302=>"000001010",
  31303=>"101011010",
  31304=>"000000100",
  31305=>"001110111",
  31306=>"100111110",
  31307=>"001100011",
  31308=>"111110001",
  31309=>"101001000",
  31310=>"001011101",
  31311=>"011100111",
  31312=>"011010111",
  31313=>"100101100",
  31314=>"101100001",
  31315=>"001001100",
  31316=>"001000110",
  31317=>"000101100",
  31318=>"011101110",
  31319=>"001011001",
  31320=>"010000100",
  31321=>"011100001",
  31322=>"100111001",
  31323=>"001001100",
  31324=>"111110100",
  31325=>"000100011",
  31326=>"001101100",
  31327=>"111101001",
  31328=>"100001111",
  31329=>"010110111",
  31330=>"111101000",
  31331=>"011001011",
  31332=>"111110011",
  31333=>"100111111",
  31334=>"110001000",
  31335=>"010110101",
  31336=>"000100111",
  31337=>"101101101",
  31338=>"100110011",
  31339=>"001000100",
  31340=>"100110010",
  31341=>"000100001",
  31342=>"000101100",
  31343=>"000100000",
  31344=>"011110000",
  31345=>"000000111",
  31346=>"110101111",
  31347=>"011000101",
  31348=>"001010110",
  31349=>"010000000",
  31350=>"111011000",
  31351=>"110100001",
  31352=>"001010110",
  31353=>"101101111",
  31354=>"111110101",
  31355=>"000011110",
  31356=>"000010010",
  31357=>"111011100",
  31358=>"001110111",
  31359=>"010110100",
  31360=>"110011010",
  31361=>"101011110",
  31362=>"101110000",
  31363=>"100100101",
  31364=>"111000100",
  31365=>"111110101",
  31366=>"100110000",
  31367=>"101100100",
  31368=>"001010000",
  31369=>"011010100",
  31370=>"100011100",
  31371=>"110010100",
  31372=>"101111010",
  31373=>"100111001",
  31374=>"011011011",
  31375=>"100000111",
  31376=>"000101111",
  31377=>"101101100",
  31378=>"011010001",
  31379=>"111101100",
  31380=>"000111000",
  31381=>"110000111",
  31382=>"011111010",
  31383=>"010010001",
  31384=>"000000011",
  31385=>"110111111",
  31386=>"011110000",
  31387=>"000001100",
  31388=>"011011001",
  31389=>"001010000",
  31390=>"111110110",
  31391=>"101011010",
  31392=>"010101111",
  31393=>"001100010",
  31394=>"111000100",
  31395=>"101111001",
  31396=>"111000011",
  31397=>"000011000",
  31398=>"110101100",
  31399=>"100000001",
  31400=>"111100010",
  31401=>"000000001",
  31402=>"110011010",
  31403=>"111011001",
  31404=>"011111100",
  31405=>"100000101",
  31406=>"111100110",
  31407=>"010001110",
  31408=>"100100011",
  31409=>"000010011",
  31410=>"111010011",
  31411=>"111011001",
  31412=>"000110110",
  31413=>"001000000",
  31414=>"110011010",
  31415=>"101110100",
  31416=>"101000000",
  31417=>"111100010",
  31418=>"101010001",
  31419=>"010110100",
  31420=>"101010111",
  31421=>"011011001",
  31422=>"001001001",
  31423=>"011000010",
  31424=>"111111000",
  31425=>"101000011",
  31426=>"011111100",
  31427=>"101000100",
  31428=>"110111010",
  31429=>"001100000",
  31430=>"111100001",
  31431=>"010101010",
  31432=>"110011011",
  31433=>"000110010",
  31434=>"100110110",
  31435=>"101101101",
  31436=>"010111100",
  31437=>"010110101",
  31438=>"011011001",
  31439=>"011011001",
  31440=>"111011000",
  31441=>"000000110",
  31442=>"110011011",
  31443=>"111000111",
  31444=>"101011110",
  31445=>"111000100",
  31446=>"001000110",
  31447=>"111010010",
  31448=>"010001011",
  31449=>"110111111",
  31450=>"101110100",
  31451=>"101101011",
  31452=>"100111101",
  31453=>"000101001",
  31454=>"100100111",
  31455=>"000100010",
  31456=>"101001010",
  31457=>"110001000",
  31458=>"101001100",
  31459=>"101101100",
  31460=>"000000111",
  31461=>"110100011",
  31462=>"010000000",
  31463=>"010001010",
  31464=>"001011110",
  31465=>"111100111",
  31466=>"010010110",
  31467=>"010000011",
  31468=>"000000000",
  31469=>"100001111",
  31470=>"101111110",
  31471=>"001110100",
  31472=>"000110110",
  31473=>"110111000",
  31474=>"110100100",
  31475=>"100000000",
  31476=>"100111010",
  31477=>"110100001",
  31478=>"011110111",
  31479=>"001011001",
  31480=>"010101000",
  31481=>"101011010",
  31482=>"110010111",
  31483=>"100110100",
  31484=>"110001101",
  31485=>"011011010",
  31486=>"110110100",
  31487=>"001001101",
  31488=>"100011101",
  31489=>"111100000",
  31490=>"000101000",
  31491=>"101110000",
  31492=>"011100011",
  31493=>"110110001",
  31494=>"000100000",
  31495=>"001100010",
  31496=>"100010100",
  31497=>"010011010",
  31498=>"110111010",
  31499=>"000010011",
  31500=>"110111011",
  31501=>"000110110",
  31502=>"111101101",
  31503=>"100111111",
  31504=>"111111000",
  31505=>"000010100",
  31506=>"110011101",
  31507=>"100001011",
  31508=>"011101100",
  31509=>"101010000",
  31510=>"011111100",
  31511=>"110010100",
  31512=>"101001110",
  31513=>"010110011",
  31514=>"000100000",
  31515=>"000100101",
  31516=>"001010100",
  31517=>"011010010",
  31518=>"001001000",
  31519=>"111111001",
  31520=>"110100101",
  31521=>"111101101",
  31522=>"101111011",
  31523=>"011101101",
  31524=>"011000100",
  31525=>"111001011",
  31526=>"100001111",
  31527=>"011111111",
  31528=>"010011000",
  31529=>"000100011",
  31530=>"101011111",
  31531=>"101001010",
  31532=>"000101101",
  31533=>"000001110",
  31534=>"101101000",
  31535=>"111000000",
  31536=>"000101001",
  31537=>"010011100",
  31538=>"111111011",
  31539=>"100101001",
  31540=>"010011001",
  31541=>"010000000",
  31542=>"011100001",
  31543=>"110110101",
  31544=>"101111000",
  31545=>"001011011",
  31546=>"110000100",
  31547=>"110011000",
  31548=>"111110000",
  31549=>"000010110",
  31550=>"110110000",
  31551=>"000101011",
  31552=>"111100111",
  31553=>"001000100",
  31554=>"100110001",
  31555=>"011101001",
  31556=>"001001010",
  31557=>"100100001",
  31558=>"100000001",
  31559=>"010000100",
  31560=>"111000000",
  31561=>"000010100",
  31562=>"000010001",
  31563=>"100001000",
  31564=>"000011100",
  31565=>"010011101",
  31566=>"010111000",
  31567=>"110011001",
  31568=>"001101011",
  31569=>"001110001",
  31570=>"011110011",
  31571=>"000100101",
  31572=>"101000001",
  31573=>"101110001",
  31574=>"000001101",
  31575=>"110110010",
  31576=>"100111000",
  31577=>"000110010",
  31578=>"110110100",
  31579=>"010000011",
  31580=>"110011011",
  31581=>"000100000",
  31582=>"101000000",
  31583=>"101100100",
  31584=>"010001101",
  31585=>"011010011",
  31586=>"100001010",
  31587=>"111011100",
  31588=>"011000001",
  31589=>"001010010",
  31590=>"111110110",
  31591=>"001111101",
  31592=>"011011001",
  31593=>"000110111",
  31594=>"000111001",
  31595=>"111100100",
  31596=>"000001011",
  31597=>"011001001",
  31598=>"001101111",
  31599=>"111011100",
  31600=>"110011100",
  31601=>"100011011",
  31602=>"001001011",
  31603=>"011001100",
  31604=>"000011011",
  31605=>"000010000",
  31606=>"000101110",
  31607=>"011111001",
  31608=>"010001110",
  31609=>"100010011",
  31610=>"001010011",
  31611=>"100100111",
  31612=>"011011010",
  31613=>"101000100",
  31614=>"001100000",
  31615=>"010101110",
  31616=>"000111000",
  31617=>"110101101",
  31618=>"100010101",
  31619=>"010010001",
  31620=>"111000101",
  31621=>"000110111",
  31622=>"001001000",
  31623=>"001000100",
  31624=>"100100101",
  31625=>"011100100",
  31626=>"000001011",
  31627=>"110001001",
  31628=>"101000111",
  31629=>"010110111",
  31630=>"100110110",
  31631=>"000111100",
  31632=>"000101111",
  31633=>"010000110",
  31634=>"111010000",
  31635=>"011011010",
  31636=>"111101110",
  31637=>"000001011",
  31638=>"001001101",
  31639=>"111110100",
  31640=>"011100111",
  31641=>"111001101",
  31642=>"000011110",
  31643=>"000000000",
  31644=>"001110011",
  31645=>"111010011",
  31646=>"010010001",
  31647=>"000100110",
  31648=>"010011101",
  31649=>"011110111",
  31650=>"001010011",
  31651=>"110100100",
  31652=>"100000000",
  31653=>"110111111",
  31654=>"001001101",
  31655=>"011000110",
  31656=>"111010011",
  31657=>"101011000",
  31658=>"110000001",
  31659=>"011011010",
  31660=>"000111100",
  31661=>"011001101",
  31662=>"101001010",
  31663=>"110010110",
  31664=>"011110010",
  31665=>"111011000",
  31666=>"100101011",
  31667=>"111100101",
  31668=>"011100110",
  31669=>"110110101",
  31670=>"000010010",
  31671=>"011100010",
  31672=>"101111000",
  31673=>"010001011",
  31674=>"011000010",
  31675=>"000100100",
  31676=>"100110011",
  31677=>"111111011",
  31678=>"010101100",
  31679=>"011001010",
  31680=>"101111011",
  31681=>"111000101",
  31682=>"101101011",
  31683=>"000000011",
  31684=>"100110010",
  31685=>"111111100",
  31686=>"001110000",
  31687=>"010000000",
  31688=>"001101100",
  31689=>"011100100",
  31690=>"111100001",
  31691=>"000111110",
  31692=>"111111101",
  31693=>"001000101",
  31694=>"001000010",
  31695=>"010101101",
  31696=>"110011001",
  31697=>"101110110",
  31698=>"100101111",
  31699=>"111111111",
  31700=>"001100101",
  31701=>"110010001",
  31702=>"110101011",
  31703=>"000011110",
  31704=>"010101101",
  31705=>"001101010",
  31706=>"000111010",
  31707=>"110011000",
  31708=>"101010100",
  31709=>"001100101",
  31710=>"000100001",
  31711=>"010001101",
  31712=>"001000001",
  31713=>"011001100",
  31714=>"110110000",
  31715=>"101001000",
  31716=>"011111001",
  31717=>"010011000",
  31718=>"000000010",
  31719=>"111100100",
  31720=>"010010000",
  31721=>"100011010",
  31722=>"000111000",
  31723=>"101110000",
  31724=>"111111110",
  31725=>"110000010",
  31726=>"010111000",
  31727=>"000100001",
  31728=>"001010100",
  31729=>"101101000",
  31730=>"101000111",
  31731=>"001001111",
  31732=>"101010011",
  31733=>"101001000",
  31734=>"000111111",
  31735=>"000000010",
  31736=>"010110100",
  31737=>"101110000",
  31738=>"101010111",
  31739=>"111001001",
  31740=>"011001100",
  31741=>"010000011",
  31742=>"101101101",
  31743=>"110001000",
  31744=>"101000010",
  31745=>"100100110",
  31746=>"101000010",
  31747=>"011011101",
  31748=>"010101101",
  31749=>"011100011",
  31750=>"110000100",
  31751=>"100000101",
  31752=>"000001010",
  31753=>"001111011",
  31754=>"000111100",
  31755=>"011111101",
  31756=>"100010101",
  31757=>"101101011",
  31758=>"101011101",
  31759=>"000011010",
  31760=>"111110100",
  31761=>"001001011",
  31762=>"100010010",
  31763=>"101000100",
  31764=>"100010011",
  31765=>"000000110",
  31766=>"111110110",
  31767=>"000001011",
  31768=>"000111100",
  31769=>"010010101",
  31770=>"000000001",
  31771=>"000111100",
  31772=>"000101100",
  31773=>"101001010",
  31774=>"010100010",
  31775=>"111001011",
  31776=>"100001110",
  31777=>"011001101",
  31778=>"001000110",
  31779=>"011000011",
  31780=>"000010100",
  31781=>"100101110",
  31782=>"111010010",
  31783=>"100001100",
  31784=>"101011100",
  31785=>"011110001",
  31786=>"001111011",
  31787=>"100000110",
  31788=>"100000010",
  31789=>"100000100",
  31790=>"100010001",
  31791=>"111111001",
  31792=>"011111100",
  31793=>"010001011",
  31794=>"101111011",
  31795=>"011000111",
  31796=>"001101010",
  31797=>"001100100",
  31798=>"011111111",
  31799=>"111001001",
  31800=>"001001000",
  31801=>"010011010",
  31802=>"100110001",
  31803=>"001110011",
  31804=>"001001110",
  31805=>"110110000",
  31806=>"000111110",
  31807=>"100100110",
  31808=>"000101001",
  31809=>"001010110",
  31810=>"000000100",
  31811=>"110001001",
  31812=>"101010111",
  31813=>"111110101",
  31814=>"011010101",
  31815=>"010000101",
  31816=>"001010110",
  31817=>"110010010",
  31818=>"100011010",
  31819=>"110100001",
  31820=>"100001000",
  31821=>"100001001",
  31822=>"011000000",
  31823=>"111111011",
  31824=>"101001000",
  31825=>"100010011",
  31826=>"000101111",
  31827=>"101101000",
  31828=>"011001100",
  31829=>"001011010",
  31830=>"001110110",
  31831=>"000110111",
  31832=>"111001111",
  31833=>"001010110",
  31834=>"101110100",
  31835=>"011010101",
  31836=>"110000001",
  31837=>"001001010",
  31838=>"111110011",
  31839=>"110001100",
  31840=>"101111010",
  31841=>"011001000",
  31842=>"110111101",
  31843=>"100001001",
  31844=>"010110101",
  31845=>"010101101",
  31846=>"100101011",
  31847=>"011110000",
  31848=>"110001000",
  31849=>"001111101",
  31850=>"011000100",
  31851=>"011000001",
  31852=>"010100010",
  31853=>"010001100",
  31854=>"001000011",
  31855=>"100111101",
  31856=>"001010001",
  31857=>"000110111",
  31858=>"000100111",
  31859=>"101000000",
  31860=>"001110111",
  31861=>"101011001",
  31862=>"101010001",
  31863=>"010001001",
  31864=>"100011010",
  31865=>"100101111",
  31866=>"111011100",
  31867=>"001011000",
  31868=>"000001001",
  31869=>"010100110",
  31870=>"000001000",
  31871=>"111011111",
  31872=>"010111000",
  31873=>"011000111",
  31874=>"001111000",
  31875=>"100111111",
  31876=>"110100100",
  31877=>"000100100",
  31878=>"010101101",
  31879=>"101011110",
  31880=>"000101010",
  31881=>"000001100",
  31882=>"000011100",
  31883=>"111111011",
  31884=>"110000111",
  31885=>"101110001",
  31886=>"111000110",
  31887=>"011011001",
  31888=>"011111101",
  31889=>"101001000",
  31890=>"011011111",
  31891=>"011010100",
  31892=>"100011001",
  31893=>"101011100",
  31894=>"000010010",
  31895=>"001001011",
  31896=>"100101000",
  31897=>"010111110",
  31898=>"101101110",
  31899=>"110000100",
  31900=>"000111111",
  31901=>"010011111",
  31902=>"000010011",
  31903=>"001100111",
  31904=>"001010111",
  31905=>"000100010",
  31906=>"101010100",
  31907=>"011111111",
  31908=>"010010011",
  31909=>"101010111",
  31910=>"110100101",
  31911=>"110101001",
  31912=>"001001001",
  31913=>"001001111",
  31914=>"101001011",
  31915=>"011100010",
  31916=>"111001111",
  31917=>"011011111",
  31918=>"111011110",
  31919=>"001011110",
  31920=>"111111010",
  31921=>"111101101",
  31922=>"101101110",
  31923=>"110111111",
  31924=>"011101001",
  31925=>"010101101",
  31926=>"111101001",
  31927=>"010101100",
  31928=>"011001001",
  31929=>"110111010",
  31930=>"111010100",
  31931=>"100001110",
  31932=>"000001011",
  31933=>"010111001",
  31934=>"100001010",
  31935=>"111011101",
  31936=>"111110000",
  31937=>"011101110",
  31938=>"001000010",
  31939=>"010110110",
  31940=>"110011110",
  31941=>"001011110",
  31942=>"110111111",
  31943=>"010000110",
  31944=>"101101101",
  31945=>"100011011",
  31946=>"011101010",
  31947=>"111000000",
  31948=>"010011010",
  31949=>"111100110",
  31950=>"100011111",
  31951=>"011001100",
  31952=>"111001001",
  31953=>"001111110",
  31954=>"000010101",
  31955=>"000111010",
  31956=>"010000110",
  31957=>"010101001",
  31958=>"010111110",
  31959=>"011101001",
  31960=>"111101101",
  31961=>"101000100",
  31962=>"001111101",
  31963=>"010011100",
  31964=>"000010101",
  31965=>"010100100",
  31966=>"000001001",
  31967=>"001110101",
  31968=>"100100001",
  31969=>"010010100",
  31970=>"101000010",
  31971=>"010010010",
  31972=>"011100000",
  31973=>"010001010",
  31974=>"011111011",
  31975=>"100000101",
  31976=>"001111101",
  31977=>"101111011",
  31978=>"000110001",
  31979=>"010011101",
  31980=>"111101100",
  31981=>"000101001",
  31982=>"101101110",
  31983=>"000100011",
  31984=>"011100111",
  31985=>"100001000",
  31986=>"011100010",
  31987=>"101000110",
  31988=>"100010001",
  31989=>"101011111",
  31990=>"001111001",
  31991=>"011111101",
  31992=>"000100000",
  31993=>"000100110",
  31994=>"010000001",
  31995=>"000001001",
  31996=>"110010010",
  31997=>"110101101",
  31998=>"110111011",
  31999=>"101110110",
  32000=>"100011001",
  32001=>"100110011",
  32002=>"011011000",
  32003=>"110011000",
  32004=>"100101010",
  32005=>"010111111",
  32006=>"011001110",
  32007=>"011011101",
  32008=>"001101101",
  32009=>"110000111",
  32010=>"110111100",
  32011=>"010101010",
  32012=>"011010111",
  32013=>"110111111",
  32014=>"011001111",
  32015=>"001001010",
  32016=>"001110111",
  32017=>"100101111",
  32018=>"011010001",
  32019=>"100000100",
  32020=>"001100010",
  32021=>"000000101",
  32022=>"000010110",
  32023=>"100011011",
  32024=>"010010011",
  32025=>"111110101",
  32026=>"011010010",
  32027=>"000111011",
  32028=>"101101011",
  32029=>"001110101",
  32030=>"110011010",
  32031=>"000011111",
  32032=>"010010111",
  32033=>"100001111",
  32034=>"011011011",
  32035=>"111100100",
  32036=>"101110101",
  32037=>"100011011",
  32038=>"101111011",
  32039=>"100100100",
  32040=>"011101110",
  32041=>"110010110",
  32042=>"011011000",
  32043=>"110010101",
  32044=>"000110001",
  32045=>"011000000",
  32046=>"010011111",
  32047=>"110101010",
  32048=>"001000110",
  32049=>"010010101",
  32050=>"111010100",
  32051=>"000000111",
  32052=>"010100101",
  32053=>"100111101",
  32054=>"011110011",
  32055=>"111010110",
  32056=>"111111101",
  32057=>"101000011",
  32058=>"000110000",
  32059=>"110111010",
  32060=>"010101011",
  32061=>"011111011",
  32062=>"101011001",
  32063=>"110111000",
  32064=>"101000100",
  32065=>"000100110",
  32066=>"010110011",
  32067=>"110001100",
  32068=>"000111110",
  32069=>"001011111",
  32070=>"010110010",
  32071=>"100110101",
  32072=>"101101111",
  32073=>"010110110",
  32074=>"111011000",
  32075=>"101101010",
  32076=>"001110100",
  32077=>"011011001",
  32078=>"100100100",
  32079=>"000001000",
  32080=>"101100100",
  32081=>"110001111",
  32082=>"111010111",
  32083=>"100001100",
  32084=>"111110101",
  32085=>"011001010",
  32086=>"110101101",
  32087=>"111011000",
  32088=>"001110100",
  32089=>"000111000",
  32090=>"000000000",
  32091=>"101001101",
  32092=>"101001001",
  32093=>"001011101",
  32094=>"000000100",
  32095=>"100110011",
  32096=>"000101101",
  32097=>"101010110",
  32098=>"010000100",
  32099=>"000110010",
  32100=>"111000011",
  32101=>"001111011",
  32102=>"111010010",
  32103=>"111010110",
  32104=>"000100001",
  32105=>"111100010",
  32106=>"111111110",
  32107=>"111011010",
  32108=>"110111110",
  32109=>"111110011",
  32110=>"000101100",
  32111=>"011111100",
  32112=>"011011100",
  32113=>"011100110",
  32114=>"111101110",
  32115=>"000110101",
  32116=>"001001000",
  32117=>"000110010",
  32118=>"100111011",
  32119=>"001110100",
  32120=>"001111110",
  32121=>"110000000",
  32122=>"100000000",
  32123=>"010111000",
  32124=>"101011000",
  32125=>"111001010",
  32126=>"110110100",
  32127=>"111111111",
  32128=>"101100000",
  32129=>"001001110",
  32130=>"110001100",
  32131=>"101010010",
  32132=>"010111101",
  32133=>"001101100",
  32134=>"110110110",
  32135=>"001010000",
  32136=>"000011101",
  32137=>"000110011",
  32138=>"011111010",
  32139=>"111011111",
  32140=>"111001101",
  32141=>"001011110",
  32142=>"100011010",
  32143=>"000101000",
  32144=>"010001000",
  32145=>"001101011",
  32146=>"101001001",
  32147=>"100110000",
  32148=>"000111011",
  32149=>"111111110",
  32150=>"110111011",
  32151=>"001110110",
  32152=>"101010010",
  32153=>"111011011",
  32154=>"011111100",
  32155=>"001011100",
  32156=>"010010010",
  32157=>"011000110",
  32158=>"011111011",
  32159=>"110011101",
  32160=>"110110010",
  32161=>"110000111",
  32162=>"111010000",
  32163=>"011110110",
  32164=>"110111011",
  32165=>"010000100",
  32166=>"000011010",
  32167=>"010000000",
  32168=>"010111001",
  32169=>"111100111",
  32170=>"010100111",
  32171=>"111100110",
  32172=>"100010001",
  32173=>"110100111",
  32174=>"001011011",
  32175=>"111101000",
  32176=>"111001111",
  32177=>"101111101",
  32178=>"000011111",
  32179=>"100011000",
  32180=>"111010001",
  32181=>"100110010",
  32182=>"010111011",
  32183=>"011111011",
  32184=>"011010011",
  32185=>"110010111",
  32186=>"000000011",
  32187=>"011101001",
  32188=>"110010011",
  32189=>"011111100",
  32190=>"011011100",
  32191=>"110110001",
  32192=>"001000110",
  32193=>"110011010",
  32194=>"111010001",
  32195=>"101110110",
  32196=>"001010000",
  32197=>"101001101",
  32198=>"101000011",
  32199=>"000011010",
  32200=>"011111101",
  32201=>"100011011",
  32202=>"101010101",
  32203=>"111001100",
  32204=>"101111110",
  32205=>"000011010",
  32206=>"110010110",
  32207=>"011101000",
  32208=>"100010011",
  32209=>"101100001",
  32210=>"000101010",
  32211=>"001011100",
  32212=>"010000110",
  32213=>"001001100",
  32214=>"110110000",
  32215=>"100100101",
  32216=>"100001010",
  32217=>"001010011",
  32218=>"010110110",
  32219=>"111101010",
  32220=>"010110000",
  32221=>"001011000",
  32222=>"100111110",
  32223=>"101001011",
  32224=>"111100100",
  32225=>"111000001",
  32226=>"100110101",
  32227=>"101100001",
  32228=>"110100100",
  32229=>"111100101",
  32230=>"010110011",
  32231=>"101011010",
  32232=>"011101110",
  32233=>"100110111",
  32234=>"011100111",
  32235=>"001000101",
  32236=>"110110011",
  32237=>"110110100",
  32238=>"100100000",
  32239=>"111001100",
  32240=>"110001100",
  32241=>"111001011",
  32242=>"000111100",
  32243=>"010110001",
  32244=>"111100011",
  32245=>"011101101",
  32246=>"111101001",
  32247=>"001100111",
  32248=>"100110001",
  32249=>"001011110",
  32250=>"101011111",
  32251=>"101000110",
  32252=>"101001001",
  32253=>"101001010",
  32254=>"000010000",
  32255=>"010110001",
  32256=>"001100100",
  32257=>"011100100",
  32258=>"001100100",
  32259=>"000011111",
  32260=>"100010100",
  32261=>"100101010",
  32262=>"100111110",
  32263=>"111111110",
  32264=>"101101011",
  32265=>"000011100",
  32266=>"010111101",
  32267=>"000110001",
  32268=>"010011000",
  32269=>"010101110",
  32270=>"101011011",
  32271=>"000110011",
  32272=>"100001010",
  32273=>"110011010",
  32274=>"000101000",
  32275=>"101001000",
  32276=>"010011000",
  32277=>"100011000",
  32278=>"110100110",
  32279=>"111101101",
  32280=>"111010010",
  32281=>"001001000",
  32282=>"111100100",
  32283=>"101011010",
  32284=>"000011011",
  32285=>"011000101",
  32286=>"001100011",
  32287=>"101010111",
  32288=>"011111000",
  32289=>"111000010",
  32290=>"010010101",
  32291=>"010110110",
  32292=>"010010110",
  32293=>"101000000",
  32294=>"101111100",
  32295=>"011011010",
  32296=>"010000011",
  32297=>"110011101",
  32298=>"000100010",
  32299=>"011101110",
  32300=>"011001010",
  32301=>"110110001",
  32302=>"001110010",
  32303=>"011011101",
  32304=>"011011111",
  32305=>"111000000",
  32306=>"111010000",
  32307=>"100100001",
  32308=>"000111001",
  32309=>"100000000",
  32310=>"100110110",
  32311=>"111000110",
  32312=>"001000000",
  32313=>"100110010",
  32314=>"001001111",
  32315=>"001101001",
  32316=>"100110110",
  32317=>"001010000",
  32318=>"010000111",
  32319=>"000011100",
  32320=>"111101110",
  32321=>"001100001",
  32322=>"010000111",
  32323=>"010101000",
  32324=>"101011000",
  32325=>"100011101",
  32326=>"000010001",
  32327=>"010011000",
  32328=>"101011101",
  32329=>"010010011",
  32330=>"111100001",
  32331=>"100000101",
  32332=>"101001100",
  32333=>"110110010",
  32334=>"111111111",
  32335=>"111110101",
  32336=>"000111111",
  32337=>"111111010",
  32338=>"101101000",
  32339=>"101001011",
  32340=>"010100101",
  32341=>"000001000",
  32342=>"110000011",
  32343=>"111000111",
  32344=>"100111011",
  32345=>"010011101",
  32346=>"000000110",
  32347=>"001000001",
  32348=>"011111010",
  32349=>"110111010",
  32350=>"011001010",
  32351=>"101101001",
  32352=>"100000101",
  32353=>"101101111",
  32354=>"001111101",
  32355=>"111010101",
  32356=>"111111110",
  32357=>"000000110",
  32358=>"111011010",
  32359=>"100000101",
  32360=>"110000000",
  32361=>"000111000",
  32362=>"011011110",
  32363=>"010101010",
  32364=>"010101101",
  32365=>"111011110",
  32366=>"011011010",
  32367=>"001011110",
  32368=>"100011000",
  32369=>"111010110",
  32370=>"101110111",
  32371=>"111001101",
  32372=>"111110111",
  32373=>"101100001",
  32374=>"101010100",
  32375=>"011000101",
  32376=>"110101111",
  32377=>"000110010",
  32378=>"110101011",
  32379=>"101100101",
  32380=>"010000011",
  32381=>"001001100",
  32382=>"010000011",
  32383=>"001111000",
  32384=>"111101010",
  32385=>"101010001",
  32386=>"000110110",
  32387=>"011110110",
  32388=>"001100001",
  32389=>"111010011",
  32390=>"100001101",
  32391=>"011010001",
  32392=>"110101111",
  32393=>"100000101",
  32394=>"101100010",
  32395=>"101111100",
  32396=>"011011101",
  32397=>"000100111",
  32398=>"001011000",
  32399=>"101111111",
  32400=>"001000101",
  32401=>"000100011",
  32402=>"111001000",
  32403=>"111100011",
  32404=>"100000011",
  32405=>"001101100",
  32406=>"001101111",
  32407=>"100010010",
  32408=>"101111101",
  32409=>"000001110",
  32410=>"000110000",
  32411=>"110000101",
  32412=>"110111000",
  32413=>"000000000",
  32414=>"110100111",
  32415=>"111110100",
  32416=>"000001010",
  32417=>"101011110",
  32418=>"011111001",
  32419=>"110001110",
  32420=>"100000010",
  32421=>"000011111",
  32422=>"000010100",
  32423=>"000110101",
  32424=>"110111011",
  32425=>"110100110",
  32426=>"000010100",
  32427=>"001010010",
  32428=>"110011100",
  32429=>"101000111",
  32430=>"010111010",
  32431=>"100011010",
  32432=>"000001101",
  32433=>"001101000",
  32434=>"110011010",
  32435=>"010010100",
  32436=>"101001010",
  32437=>"101010001",
  32438=>"111010000",
  32439=>"101011001",
  32440=>"001101001",
  32441=>"010001110",
  32442=>"001010100",
  32443=>"000011100",
  32444=>"000001000",
  32445=>"011111001",
  32446=>"101100011",
  32447=>"010000001",
  32448=>"011011101",
  32449=>"010001100",
  32450=>"000011011",
  32451=>"000100100",
  32452=>"000000101",
  32453=>"101110111",
  32454=>"110011111",
  32455=>"110010111",
  32456=>"010000111",
  32457=>"110000100",
  32458=>"101100101",
  32459=>"001100100",
  32460=>"000011001",
  32461=>"100111011",
  32462=>"111111001",
  32463=>"110000000",
  32464=>"010001011",
  32465=>"000101111",
  32466=>"000010010",
  32467=>"000010110",
  32468=>"101001100",
  32469=>"000010010",
  32470=>"010101000",
  32471=>"100010100",
  32472=>"110100000",
  32473=>"110010000",
  32474=>"011100100",
  32475=>"001000101",
  32476=>"001011111",
  32477=>"000110100",
  32478=>"100101011",
  32479=>"101101011",
  32480=>"111011010",
  32481=>"101000000",
  32482=>"111011110",
  32483=>"001100010",
  32484=>"000100101",
  32485=>"100001000",
  32486=>"111110110",
  32487=>"000100100",
  32488=>"001000010",
  32489=>"011000000",
  32490=>"100100111",
  32491=>"011100000",
  32492=>"000000111",
  32493=>"010000011",
  32494=>"111111100",
  32495=>"110010011",
  32496=>"100100011",
  32497=>"111110011",
  32498=>"100001100",
  32499=>"011100000",
  32500=>"001101010",
  32501=>"111010111",
  32502=>"111011110",
  32503=>"110001100",
  32504=>"101101100",
  32505=>"100010111",
  32506=>"010000000",
  32507=>"011001001",
  32508=>"010101000",
  32509=>"000000101",
  32510=>"101010100",
  32511=>"110010110",
  32512=>"110000001",
  32513=>"000000100",
  32514=>"111000010",
  32515=>"001001001",
  32516=>"100001111",
  32517=>"001101001",
  32518=>"011101000",
  32519=>"000001111",
  32520=>"001011010",
  32521=>"110100010",
  32522=>"011000000",
  32523=>"011000101",
  32524=>"000101101",
  32525=>"011000110",
  32526=>"110000100",
  32527=>"111100011",
  32528=>"011111100",
  32529=>"101001101",
  32530=>"001001010",
  32531=>"011101101",
  32532=>"001101010",
  32533=>"000000010",
  32534=>"110100110",
  32535=>"010011100",
  32536=>"111100000",
  32537=>"100000100",
  32538=>"000000110",
  32539=>"101000001",
  32540=>"011100011",
  32541=>"001001110",
  32542=>"111110110",
  32543=>"011100111",
  32544=>"010110111",
  32545=>"110010111",
  32546=>"001000010",
  32547=>"000111101",
  32548=>"000111010",
  32549=>"000110001",
  32550=>"101100001",
  32551=>"111110011",
  32552=>"111001011",
  32553=>"001010111",
  32554=>"110010010",
  32555=>"001000000",
  32556=>"100011011",
  32557=>"000010000",
  32558=>"000111010",
  32559=>"110000111",
  32560=>"001010101",
  32561=>"110000100",
  32562=>"011111100",
  32563=>"010011111",
  32564=>"101101101",
  32565=>"000010001",
  32566=>"101001100",
  32567=>"000110011",
  32568=>"100100111",
  32569=>"011110110",
  32570=>"111111110",
  32571=>"011101100",
  32572=>"001101100",
  32573=>"110101000",
  32574=>"100101101",
  32575=>"101100111",
  32576=>"010000100",
  32577=>"001101010",
  32578=>"000010101",
  32579=>"101001111",
  32580=>"000111111",
  32581=>"011011111",
  32582=>"100010000",
  32583=>"100001001",
  32584=>"111100010",
  32585=>"010100100",
  32586=>"100010101",
  32587=>"110110001",
  32588=>"110010010",
  32589=>"110101111",
  32590=>"001110000",
  32591=>"000001001",
  32592=>"010101010",
  32593=>"101010001",
  32594=>"010100001",
  32595=>"010111100",
  32596=>"101100111",
  32597=>"111100101",
  32598=>"001101111",
  32599=>"111110100",
  32600=>"111101010",
  32601=>"000110111",
  32602=>"110000001",
  32603=>"011011000",
  32604=>"011011010",
  32605=>"111110001",
  32606=>"011111100",
  32607=>"010100101",
  32608=>"001001000",
  32609=>"001010111",
  32610=>"000111001",
  32611=>"010111101",
  32612=>"100000001",
  32613=>"000010000",
  32614=>"001000000",
  32615=>"001011010",
  32616=>"111000001",
  32617=>"010010101",
  32618=>"001011101",
  32619=>"111111101",
  32620=>"110011001",
  32621=>"011000010",
  32622=>"000100110",
  32623=>"001010100",
  32624=>"000001001",
  32625=>"011110110",
  32626=>"100100010",
  32627=>"101101110",
  32628=>"111100001",
  32629=>"101110000",
  32630=>"111100001",
  32631=>"011111010",
  32632=>"110101111",
  32633=>"000111110",
  32634=>"000010101",
  32635=>"000011011",
  32636=>"110111010",
  32637=>"000011110",
  32638=>"100110111",
  32639=>"111101010",
  32640=>"101000001",
  32641=>"011010011",
  32642=>"001000010",
  32643=>"110100110",
  32644=>"111101000",
  32645=>"000011101",
  32646=>"111001101",
  32647=>"110010100",
  32648=>"100111111",
  32649=>"111100011",
  32650=>"101111100",
  32651=>"000111100",
  32652=>"101000010",
  32653=>"001001011",
  32654=>"110000001",
  32655=>"010000001",
  32656=>"111101000",
  32657=>"001001001",
  32658=>"010001001",
  32659=>"010101001",
  32660=>"011010001",
  32661=>"101011011",
  32662=>"101011000",
  32663=>"110000000",
  32664=>"001000110",
  32665=>"000010111",
  32666=>"100110100",
  32667=>"001110110",
  32668=>"110011000",
  32669=>"000000111",
  32670=>"110001111",
  32671=>"000000000",
  32672=>"011000101",
  32673=>"100110101",
  32674=>"010001100",
  32675=>"011010010",
  32676=>"000100010",
  32677=>"110000101",
  32678=>"111110000",
  32679=>"000110010",
  32680=>"000111010",
  32681=>"100010010",
  32682=>"000111101",
  32683=>"111101000",
  32684=>"100000010",
  32685=>"110100010",
  32686=>"010001011",
  32687=>"011010000",
  32688=>"101001111",
  32689=>"101111011",
  32690=>"001111101",
  32691=>"111010010",
  32692=>"000100100",
  32693=>"011010111",
  32694=>"000001110",
  32695=>"110001000",
  32696=>"110101011",
  32697=>"100011011",
  32698=>"000100000",
  32699=>"111100001",
  32700=>"010100110",
  32701=>"111111010",
  32702=>"100001100",
  32703=>"001100011",
  32704=>"111011001",
  32705=>"000011110",
  32706=>"110111010",
  32707=>"110011111",
  32708=>"111111111",
  32709=>"101010110",
  32710=>"111101111",
  32711=>"000111110",
  32712=>"001100000",
  32713=>"001010001",
  32714=>"000100100",
  32715=>"110110111",
  32716=>"010011000",
  32717=>"100001101",
  32718=>"111000000",
  32719=>"111110100",
  32720=>"001011000",
  32721=>"000100111",
  32722=>"001001011",
  32723=>"001100011",
  32724=>"001100001",
  32725=>"100001000",
  32726=>"101000000",
  32727=>"000010111",
  32728=>"111001100",
  32729=>"100101100",
  32730=>"010001001",
  32731=>"100001010",
  32732=>"011000100",
  32733=>"001001001",
  32734=>"011100101",
  32735=>"111110011",
  32736=>"111111100",
  32737=>"111001010",
  32738=>"011000111",
  32739=>"111001001",
  32740=>"011001001",
  32741=>"101110000",
  32742=>"010000110",
  32743=>"100000001",
  32744=>"000001111",
  32745=>"001110101",
  32746=>"100000101",
  32747=>"011110110",
  32748=>"111110010",
  32749=>"100111001",
  32750=>"010001010",
  32751=>"010010000",
  32752=>"000101111",
  32753=>"111001001",
  32754=>"100000110",
  32755=>"110101000",
  32756=>"100010010",
  32757=>"110111000",
  32758=>"001001000",
  32759=>"111100101",
  32760=>"011010110",
  32761=>"001010000",
  32762=>"111100001",
  32763=>"000001110",
  32764=>"101011000",
  32765=>"000011010",
  32766=>"011001000",
  32767=>"011000010",
  32768=>"010101011",
  32769=>"111011001",
  32770=>"110011100",
  32771=>"100110010",
  32772=>"010110001",
  32773=>"001100100",
  32774=>"101101010",
  32775=>"011101010",
  32776=>"000100100",
  32777=>"011011100",
  32778=>"001111111",
  32779=>"011111010",
  32780=>"010010101",
  32781=>"101101100",
  32782=>"100001011",
  32783=>"111010110",
  32784=>"100101100",
  32785=>"111010110",
  32786=>"011011100",
  32787=>"011000110",
  32788=>"111100011",
  32789=>"101111110",
  32790=>"110101100",
  32791=>"000011101",
  32792=>"011001100",
  32793=>"010100000",
  32794=>"001000110",
  32795=>"010000101",
  32796=>"111101010",
  32797=>"001101100",
  32798=>"101001111",
  32799=>"110101111",
  32800=>"010001101",
  32801=>"010010011",
  32802=>"010101000",
  32803=>"110110001",
  32804=>"101011101",
  32805=>"011110000",
  32806=>"011000010",
  32807=>"000011000",
  32808=>"001101110",
  32809=>"101000111",
  32810=>"011011111",
  32811=>"000100000",
  32812=>"110010011",
  32813=>"111111110",
  32814=>"011000010",
  32815=>"101000001",
  32816=>"101110001",
  32817=>"011001001",
  32818=>"011110010",
  32819=>"001001101",
  32820=>"100101110",
  32821=>"011111100",
  32822=>"100110001",
  32823=>"010010011",
  32824=>"000100100",
  32825=>"111111001",
  32826=>"000010110",
  32827=>"110100100",
  32828=>"100010010",
  32829=>"011100101",
  32830=>"001001001",
  32831=>"110011111",
  32832=>"100000100",
  32833=>"010000110",
  32834=>"110001010",
  32835=>"010010100",
  32836=>"001101101",
  32837=>"001110101",
  32838=>"111011000",
  32839=>"000100011",
  32840=>"011010101",
  32841=>"001000111",
  32842=>"000110000",
  32843=>"100100111",
  32844=>"000010111",
  32845=>"010000011",
  32846=>"100001111",
  32847=>"100111101",
  32848=>"001100010",
  32849=>"110010110",
  32850=>"000010110",
  32851=>"000100001",
  32852=>"100100011",
  32853=>"000010010",
  32854=>"010110111",
  32855=>"000111111",
  32856=>"010001111",
  32857=>"101010000",
  32858=>"100100000",
  32859=>"101101111",
  32860=>"110110001",
  32861=>"000100101",
  32862=>"111000010",
  32863=>"000000100",
  32864=>"001010011",
  32865=>"001000100",
  32866=>"000011001",
  32867=>"101100001",
  32868=>"001110110",
  32869=>"111001100",
  32870=>"000101111",
  32871=>"110000000",
  32872=>"010110010",
  32873=>"100110010",
  32874=>"101100110",
  32875=>"010110001",
  32876=>"011110010",
  32877=>"001100011",
  32878=>"010101011",
  32879=>"110100011",
  32880=>"111101111",
  32881=>"011100101",
  32882=>"100010101",
  32883=>"111000100",
  32884=>"110000110",
  32885=>"011101011",
  32886=>"100010101",
  32887=>"000010101",
  32888=>"101010111",
  32889=>"110110101",
  32890=>"010100111",
  32891=>"000110101",
  32892=>"110111111",
  32893=>"101001011",
  32894=>"000010010",
  32895=>"101100110",
  32896=>"100001111",
  32897=>"101010100",
  32898=>"100101111",
  32899=>"101000100",
  32900=>"101011001",
  32901=>"100011011",
  32902=>"101100000",
  32903=>"010001000",
  32904=>"001100001",
  32905=>"101111110",
  32906=>"110000110",
  32907=>"001111111",
  32908=>"010010110",
  32909=>"101101000",
  32910=>"000000111",
  32911=>"100111111",
  32912=>"010110001",
  32913=>"001100111",
  32914=>"010101100",
  32915=>"000001010",
  32916=>"100000010",
  32917=>"000001000",
  32918=>"001111110",
  32919=>"101011000",
  32920=>"101011110",
  32921=>"100100010",
  32922=>"010010010",
  32923=>"000001111",
  32924=>"110111011",
  32925=>"001000000",
  32926=>"101110010",
  32927=>"000000110",
  32928=>"010000100",
  32929=>"011101100",
  32930=>"110010000",
  32931=>"100000000",
  32932=>"001011000",
  32933=>"011000111",
  32934=>"011001100",
  32935=>"011011010",
  32936=>"100110001",
  32937=>"010011100",
  32938=>"101000110",
  32939=>"111010101",
  32940=>"111100100",
  32941=>"100101101",
  32942=>"000100001",
  32943=>"001101111",
  32944=>"111000100",
  32945=>"010111001",
  32946=>"000100100",
  32947=>"001010000",
  32948=>"000010110",
  32949=>"000010110",
  32950=>"101011111",
  32951=>"001000111",
  32952=>"110100011",
  32953=>"100001011",
  32954=>"101111110",
  32955=>"111101100",
  32956=>"000001110",
  32957=>"111011100",
  32958=>"010111010",
  32959=>"000001010",
  32960=>"101110101",
  32961=>"010100111",
  32962=>"101101000",
  32963=>"101100000",
  32964=>"110110100",
  32965=>"010000110",
  32966=>"010101100",
  32967=>"010101001",
  32968=>"010101101",
  32969=>"110010001",
  32970=>"000101010",
  32971=>"110100010",
  32972=>"100000101",
  32973=>"010100111",
  32974=>"110110010",
  32975=>"010001111",
  32976=>"010011001",
  32977=>"001011010",
  32978=>"110110011",
  32979=>"000000001",
  32980=>"010100100",
  32981=>"011101101",
  32982=>"001000101",
  32983=>"001110111",
  32984=>"000111100",
  32985=>"001110110",
  32986=>"011111011",
  32987=>"011001011",
  32988=>"000010010",
  32989=>"110010100",
  32990=>"011011111",
  32991=>"101100111",
  32992=>"001001110",
  32993=>"100110011",
  32994=>"011101000",
  32995=>"110001011",
  32996=>"000011110",
  32997=>"100101010",
  32998=>"000111111",
  32999=>"010001010",
  33000=>"000000010",
  33001=>"000011010",
  33002=>"001011101",
  33003=>"001000100",
  33004=>"110110010",
  33005=>"111101101",
  33006=>"011011100",
  33007=>"010001000",
  33008=>"101011110",
  33009=>"100010010",
  33010=>"110010000",
  33011=>"010011011",
  33012=>"010101000",
  33013=>"000000100",
  33014=>"110110001",
  33015=>"011100111",
  33016=>"011110101",
  33017=>"110111001",
  33018=>"011000010",
  33019=>"111111100",
  33020=>"010110111",
  33021=>"000011011",
  33022=>"111100111",
  33023=>"001101001",
  33024=>"001011000",
  33025=>"000011011",
  33026=>"000011010",
  33027=>"001110111",
  33028=>"000100011",
  33029=>"110011101",
  33030=>"001101100",
  33031=>"111110111",
  33032=>"000101001",
  33033=>"001000100",
  33034=>"001110100",
  33035=>"101000000",
  33036=>"101110011",
  33037=>"011101010",
  33038=>"100100101",
  33039=>"111000001",
  33040=>"001111101",
  33041=>"101010000",
  33042=>"101010101",
  33043=>"111110111",
  33044=>"010000110",
  33045=>"101001111",
  33046=>"010101001",
  33047=>"101110111",
  33048=>"011010010",
  33049=>"011011011",
  33050=>"100110011",
  33051=>"010010101",
  33052=>"000010010",
  33053=>"001010110",
  33054=>"010100001",
  33055=>"100011010",
  33056=>"110100010",
  33057=>"110110010",
  33058=>"001011011",
  33059=>"000100000",
  33060=>"111101111",
  33061=>"110000001",
  33062=>"010111011",
  33063=>"111100101",
  33064=>"000100101",
  33065=>"011110000",
  33066=>"111010011",
  33067=>"111001001",
  33068=>"100001010",
  33069=>"011001010",
  33070=>"110111010",
  33071=>"000100011",
  33072=>"110000110",
  33073=>"100100010",
  33074=>"100101001",
  33075=>"001100001",
  33076=>"101010010",
  33077=>"010010110",
  33078=>"010001101",
  33079=>"000101001",
  33080=>"111101011",
  33081=>"010110100",
  33082=>"110011010",
  33083=>"111101111",
  33084=>"001100010",
  33085=>"000000110",
  33086=>"011110100",
  33087=>"010010111",
  33088=>"110011001",
  33089=>"010010000",
  33090=>"001110110",
  33091=>"001100111",
  33092=>"010100111",
  33093=>"010101000",
  33094=>"101000111",
  33095=>"000010000",
  33096=>"001101110",
  33097=>"000100000",
  33098=>"100100101",
  33099=>"101110100",
  33100=>"101111111",
  33101=>"110010011",
  33102=>"101110111",
  33103=>"110111110",
  33104=>"101101111",
  33105=>"011110001",
  33106=>"010001101",
  33107=>"000111011",
  33108=>"000101110",
  33109=>"100010011",
  33110=>"000100010",
  33111=>"001100100",
  33112=>"110001100",
  33113=>"100101100",
  33114=>"011010110",
  33115=>"100000100",
  33116=>"011011101",
  33117=>"001000011",
  33118=>"000101111",
  33119=>"000110001",
  33120=>"110101101",
  33121=>"101111000",
  33122=>"001000101",
  33123=>"100101101",
  33124=>"010011100",
  33125=>"101000010",
  33126=>"000001110",
  33127=>"000011100",
  33128=>"011010010",
  33129=>"110000111",
  33130=>"000100110",
  33131=>"100010000",
  33132=>"111001001",
  33133=>"111011010",
  33134=>"100010001",
  33135=>"110101101",
  33136=>"010000011",
  33137=>"111110110",
  33138=>"000010010",
  33139=>"011000111",
  33140=>"110100101",
  33141=>"110101001",
  33142=>"010011000",
  33143=>"011100010",
  33144=>"001010110",
  33145=>"011111001",
  33146=>"011011111",
  33147=>"111000101",
  33148=>"011110010",
  33149=>"111010011",
  33150=>"111101011",
  33151=>"001000110",
  33152=>"100001111",
  33153=>"110101001",
  33154=>"001111010",
  33155=>"100000000",
  33156=>"001101110",
  33157=>"110111000",
  33158=>"011000010",
  33159=>"000111101",
  33160=>"000010111",
  33161=>"011010011",
  33162=>"001000101",
  33163=>"010000110",
  33164=>"111010100",
  33165=>"000010001",
  33166=>"100011011",
  33167=>"001110011",
  33168=>"111100111",
  33169=>"011001000",
  33170=>"110100010",
  33171=>"110000001",
  33172=>"101010011",
  33173=>"010101101",
  33174=>"010100101",
  33175=>"011100001",
  33176=>"110011000",
  33177=>"001000101",
  33178=>"110101011",
  33179=>"000010111",
  33180=>"100000111",
  33181=>"001001011",
  33182=>"101111100",
  33183=>"010000001",
  33184=>"010010110",
  33185=>"001011111",
  33186=>"101101100",
  33187=>"100000101",
  33188=>"011101011",
  33189=>"111001011",
  33190=>"110101100",
  33191=>"111001010",
  33192=>"001010010",
  33193=>"010101000",
  33194=>"101011011",
  33195=>"111001000",
  33196=>"000010011",
  33197=>"010000110",
  33198=>"010010100",
  33199=>"101110000",
  33200=>"000100001",
  33201=>"011001000",
  33202=>"101111111",
  33203=>"101100101",
  33204=>"011000111",
  33205=>"010101101",
  33206=>"011001100",
  33207=>"000100000",
  33208=>"101010010",
  33209=>"111000101",
  33210=>"100100001",
  33211=>"010001100",
  33212=>"010110011",
  33213=>"011101110",
  33214=>"001100100",
  33215=>"001000111",
  33216=>"001001011",
  33217=>"011111110",
  33218=>"100111111",
  33219=>"111111001",
  33220=>"111111110",
  33221=>"101100001",
  33222=>"010000001",
  33223=>"101100100",
  33224=>"010101101",
  33225=>"101101010",
  33226=>"010011101",
  33227=>"001001000",
  33228=>"010111100",
  33229=>"101110111",
  33230=>"010000101",
  33231=>"011111110",
  33232=>"101111001",
  33233=>"000010110",
  33234=>"100010001",
  33235=>"100011111",
  33236=>"110000111",
  33237=>"100101011",
  33238=>"010110000",
  33239=>"111001011",
  33240=>"101110110",
  33241=>"100110010",
  33242=>"110011000",
  33243=>"111100010",
  33244=>"110010001",
  33245=>"000101101",
  33246=>"001000011",
  33247=>"001110111",
  33248=>"101110100",
  33249=>"101010100",
  33250=>"000110000",
  33251=>"110111100",
  33252=>"100010110",
  33253=>"110110010",
  33254=>"100000000",
  33255=>"101101101",
  33256=>"010110111",
  33257=>"010111010",
  33258=>"011111110",
  33259=>"010100010",
  33260=>"011001110",
  33261=>"111111001",
  33262=>"011110110",
  33263=>"000000000",
  33264=>"101010101",
  33265=>"101010110",
  33266=>"111010000",
  33267=>"101101000",
  33268=>"000111000",
  33269=>"001011010",
  33270=>"101110000",
  33271=>"010000010",
  33272=>"111001010",
  33273=>"000100100",
  33274=>"111110010",
  33275=>"100011110",
  33276=>"001110101",
  33277=>"000011011",
  33278=>"000110110",
  33279=>"101011011",
  33280=>"001111011",
  33281=>"111001100",
  33282=>"000111001",
  33283=>"000111101",
  33284=>"100000011",
  33285=>"111011011",
  33286=>"001100101",
  33287=>"101011001",
  33288=>"100000000",
  33289=>"101001100",
  33290=>"010000000",
  33291=>"111000111",
  33292=>"111010101",
  33293=>"011001110",
  33294=>"011100110",
  33295=>"100001111",
  33296=>"000111100",
  33297=>"001111000",
  33298=>"101000011",
  33299=>"000000000",
  33300=>"010000000",
  33301=>"111001110",
  33302=>"101111111",
  33303=>"001001001",
  33304=>"110111011",
  33305=>"001001110",
  33306=>"100000100",
  33307=>"011000000",
  33308=>"111110101",
  33309=>"000110111",
  33310=>"100011011",
  33311=>"110110000",
  33312=>"100001010",
  33313=>"111000011",
  33314=>"010000000",
  33315=>"111011110",
  33316=>"001100011",
  33317=>"100010111",
  33318=>"011011110",
  33319=>"100101111",
  33320=>"110011110",
  33321=>"011111110",
  33322=>"011101000",
  33323=>"111011100",
  33324=>"100100100",
  33325=>"001000001",
  33326=>"000001011",
  33327=>"001000001",
  33328=>"110000111",
  33329=>"010001011",
  33330=>"000111101",
  33331=>"010111110",
  33332=>"011111011",
  33333=>"100011101",
  33334=>"101100101",
  33335=>"101100101",
  33336=>"001111100",
  33337=>"010000001",
  33338=>"000010010",
  33339=>"010111111",
  33340=>"001100000",
  33341=>"100110100",
  33342=>"101001101",
  33343=>"011100100",
  33344=>"001010110",
  33345=>"000101100",
  33346=>"010000001",
  33347=>"011100001",
  33348=>"010001110",
  33349=>"000010101",
  33350=>"001010000",
  33351=>"001001111",
  33352=>"010011100",
  33353=>"001111011",
  33354=>"001000111",
  33355=>"000111011",
  33356=>"111111110",
  33357=>"011101000",
  33358=>"001001100",
  33359=>"100011110",
  33360=>"001001000",
  33361=>"001010000",
  33362=>"011001011",
  33363=>"001001010",
  33364=>"000010000",
  33365=>"010000011",
  33366=>"000000111",
  33367=>"011010101",
  33368=>"010010000",
  33369=>"011011011",
  33370=>"110010010",
  33371=>"101110111",
  33372=>"100111001",
  33373=>"001010000",
  33374=>"000111101",
  33375=>"110111011",
  33376=>"101000001",
  33377=>"110000010",
  33378=>"011111010",
  33379=>"110110000",
  33380=>"111101110",
  33381=>"000001011",
  33382=>"101000011",
  33383=>"000011000",
  33384=>"011001010",
  33385=>"010110010",
  33386=>"101110100",
  33387=>"110110110",
  33388=>"100100111",
  33389=>"001000010",
  33390=>"000100000",
  33391=>"110010110",
  33392=>"110111101",
  33393=>"100111101",
  33394=>"101011001",
  33395=>"010101101",
  33396=>"101001000",
  33397=>"001100100",
  33398=>"111000111",
  33399=>"110001100",
  33400=>"100100100",
  33401=>"000111001",
  33402=>"010000010",
  33403=>"110111101",
  33404=>"101010011",
  33405=>"010101100",
  33406=>"111010001",
  33407=>"101010001",
  33408=>"010010010",
  33409=>"001001111",
  33410=>"001101111",
  33411=>"000001011",
  33412=>"011100100",
  33413=>"110000010",
  33414=>"000010000",
  33415=>"010010110",
  33416=>"100010100",
  33417=>"000110110",
  33418=>"111110111",
  33419=>"100101111",
  33420=>"001000110",
  33421=>"110011100",
  33422=>"001000010",
  33423=>"010111101",
  33424=>"101000010",
  33425=>"110111111",
  33426=>"101000100",
  33427=>"110111110",
  33428=>"001001000",
  33429=>"110110011",
  33430=>"100101101",
  33431=>"011110110",
  33432=>"011111100",
  33433=>"000000011",
  33434=>"011111110",
  33435=>"001111000",
  33436=>"100100100",
  33437=>"000001111",
  33438=>"000011000",
  33439=>"111111101",
  33440=>"101010000",
  33441=>"010001101",
  33442=>"100101100",
  33443=>"011010000",
  33444=>"010111000",
  33445=>"001110111",
  33446=>"101011101",
  33447=>"001010011",
  33448=>"011000011",
  33449=>"111000110",
  33450=>"010010100",
  33451=>"001111101",
  33452=>"111101100",
  33453=>"011000000",
  33454=>"011011011",
  33455=>"111100000",
  33456=>"100100101",
  33457=>"000000110",
  33458=>"010011100",
  33459=>"110101001",
  33460=>"010010001",
  33461=>"100111110",
  33462=>"101100001",
  33463=>"001010100",
  33464=>"101111110",
  33465=>"111010101",
  33466=>"101010000",
  33467=>"110001101",
  33468=>"010100111",
  33469=>"010100110",
  33470=>"000011110",
  33471=>"010100101",
  33472=>"110101101",
  33473=>"011011001",
  33474=>"011100110",
  33475=>"001101101",
  33476=>"111111001",
  33477=>"000110000",
  33478=>"110001111",
  33479=>"010001001",
  33480=>"111000111",
  33481=>"001001101",
  33482=>"101110000",
  33483=>"001001011",
  33484=>"000011000",
  33485=>"011001011",
  33486=>"000101011",
  33487=>"110101011",
  33488=>"001001111",
  33489=>"011101010",
  33490=>"101101011",
  33491=>"110011000",
  33492=>"111100001",
  33493=>"000010100",
  33494=>"110001011",
  33495=>"101101110",
  33496=>"000100000",
  33497=>"101110101",
  33498=>"111101101",
  33499=>"111101101",
  33500=>"000110010",
  33501=>"011100000",
  33502=>"110100010",
  33503=>"110111100",
  33504=>"000101100",
  33505=>"101010100",
  33506=>"100001111",
  33507=>"011101100",
  33508=>"111111011",
  33509=>"001001000",
  33510=>"000111001",
  33511=>"011011000",
  33512=>"100111011",
  33513=>"000010011",
  33514=>"001101010",
  33515=>"111000001",
  33516=>"101001100",
  33517=>"110100010",
  33518=>"011110011",
  33519=>"011000110",
  33520=>"100111101",
  33521=>"111111100",
  33522=>"111111110",
  33523=>"101010000",
  33524=>"011010111",
  33525=>"000000010",
  33526=>"011001000",
  33527=>"011011001",
  33528=>"010001011",
  33529=>"011110001",
  33530=>"001111100",
  33531=>"000000000",
  33532=>"101010000",
  33533=>"000101100",
  33534=>"011101000",
  33535=>"011101000",
  33536=>"101010110",
  33537=>"001111011",
  33538=>"110001010",
  33539=>"110110010",
  33540=>"011110100",
  33541=>"001101101",
  33542=>"110100010",
  33543=>"100111110",
  33544=>"001001000",
  33545=>"100010110",
  33546=>"010000001",
  33547=>"001001100",
  33548=>"111101011",
  33549=>"111111111",
  33550=>"000000101",
  33551=>"100101010",
  33552=>"001110001",
  33553=>"100100100",
  33554=>"001010000",
  33555=>"110100111",
  33556=>"100100111",
  33557=>"010100101",
  33558=>"101001011",
  33559=>"111111100",
  33560=>"010100111",
  33561=>"011001101",
  33562=>"001100110",
  33563=>"000000000",
  33564=>"100001000",
  33565=>"000101100",
  33566=>"011000110",
  33567=>"101011001",
  33568=>"100000101",
  33569=>"000010001",
  33570=>"010110010",
  33571=>"111011010",
  33572=>"100111000",
  33573=>"000000000",
  33574=>"101001111",
  33575=>"101110011",
  33576=>"111000101",
  33577=>"011010010",
  33578=>"010011000",
  33579=>"011000111",
  33580=>"001111100",
  33581=>"010100001",
  33582=>"100010110",
  33583=>"011110111",
  33584=>"100010000",
  33585=>"111010010",
  33586=>"110011101",
  33587=>"100100100",
  33588=>"100000101",
  33589=>"011010010",
  33590=>"001100010",
  33591=>"010001101",
  33592=>"000001110",
  33593=>"000000000",
  33594=>"000111000",
  33595=>"000000001",
  33596=>"101101100",
  33597=>"011100111",
  33598=>"001000100",
  33599=>"011011011",
  33600=>"100001011",
  33601=>"011001011",
  33602=>"011111011",
  33603=>"110111100",
  33604=>"101111011",
  33605=>"110110111",
  33606=>"111111000",
  33607=>"101100101",
  33608=>"110000001",
  33609=>"101110011",
  33610=>"110011101",
  33611=>"100001110",
  33612=>"110100010",
  33613=>"001011100",
  33614=>"000110100",
  33615=>"101100101",
  33616=>"111001100",
  33617=>"101101001",
  33618=>"010000001",
  33619=>"011111011",
  33620=>"110001010",
  33621=>"010100111",
  33622=>"001100100",
  33623=>"010011100",
  33624=>"000110100",
  33625=>"000101001",
  33626=>"100110110",
  33627=>"110000001",
  33628=>"000100011",
  33629=>"110100001",
  33630=>"001011100",
  33631=>"100111101",
  33632=>"110000000",
  33633=>"001011011",
  33634=>"011110011",
  33635=>"101011111",
  33636=>"111000111",
  33637=>"100000100",
  33638=>"100011010",
  33639=>"101010001",
  33640=>"000011100",
  33641=>"000010011",
  33642=>"101010100",
  33643=>"100110010",
  33644=>"101111010",
  33645=>"010011010",
  33646=>"010101100",
  33647=>"001000001",
  33648=>"100011101",
  33649=>"011100011",
  33650=>"010110000",
  33651=>"000101111",
  33652=>"111011010",
  33653=>"110111111",
  33654=>"011101011",
  33655=>"110000010",
  33656=>"111101000",
  33657=>"100100000",
  33658=>"100111000",
  33659=>"000001101",
  33660=>"001101000",
  33661=>"000011001",
  33662=>"001000111",
  33663=>"101110110",
  33664=>"111001010",
  33665=>"001101010",
  33666=>"000001111",
  33667=>"010001101",
  33668=>"010110011",
  33669=>"110100000",
  33670=>"010010101",
  33671=>"001001010",
  33672=>"101111110",
  33673=>"010111001",
  33674=>"010000101",
  33675=>"110010000",
  33676=>"101001001",
  33677=>"011001001",
  33678=>"101101000",
  33679=>"101010101",
  33680=>"111001001",
  33681=>"100111111",
  33682=>"011001101",
  33683=>"000101100",
  33684=>"110011101",
  33685=>"110001011",
  33686=>"001010010",
  33687=>"001010101",
  33688=>"100010010",
  33689=>"010101100",
  33690=>"011010010",
  33691=>"111001110",
  33692=>"000110100",
  33693=>"100101010",
  33694=>"010001110",
  33695=>"001111100",
  33696=>"001011100",
  33697=>"001011000",
  33698=>"001011000",
  33699=>"001110011",
  33700=>"010010000",
  33701=>"000010000",
  33702=>"111111100",
  33703=>"000001010",
  33704=>"011010100",
  33705=>"000000111",
  33706=>"001101100",
  33707=>"001111111",
  33708=>"100010101",
  33709=>"100010010",
  33710=>"100001010",
  33711=>"000101101",
  33712=>"000010100",
  33713=>"011010110",
  33714=>"010111110",
  33715=>"000011111",
  33716=>"100001111",
  33717=>"000100110",
  33718=>"011000101",
  33719=>"101001000",
  33720=>"111100100",
  33721=>"010001011",
  33722=>"010000010",
  33723=>"011001011",
  33724=>"010101000",
  33725=>"101111101",
  33726=>"000101010",
  33727=>"000010000",
  33728=>"001000110",
  33729=>"011111011",
  33730=>"011111110",
  33731=>"001011001",
  33732=>"011110010",
  33733=>"110111100",
  33734=>"010110101",
  33735=>"000001101",
  33736=>"000001000",
  33737=>"111001010",
  33738=>"011010010",
  33739=>"010111010",
  33740=>"010110110",
  33741=>"010101111",
  33742=>"100000101",
  33743=>"101011110",
  33744=>"101001000",
  33745=>"011111010",
  33746=>"110011011",
  33747=>"000010111",
  33748=>"100101110",
  33749=>"100011100",
  33750=>"000110111",
  33751=>"001111111",
  33752=>"111111110",
  33753=>"111000011",
  33754=>"010011000",
  33755=>"100111111",
  33756=>"000110110",
  33757=>"000001110",
  33758=>"010101001",
  33759=>"010110100",
  33760=>"110000011",
  33761=>"110101010",
  33762=>"001101111",
  33763=>"010101100",
  33764=>"101001101",
  33765=>"011111011",
  33766=>"111100110",
  33767=>"101100100",
  33768=>"000100101",
  33769=>"011011101",
  33770=>"100011111",
  33771=>"000000001",
  33772=>"011001100",
  33773=>"011111111",
  33774=>"011010011",
  33775=>"110011110",
  33776=>"010010011",
  33777=>"110000000",
  33778=>"101010010",
  33779=>"110001011",
  33780=>"001010001",
  33781=>"101110110",
  33782=>"010010010",
  33783=>"000010110",
  33784=>"000111111",
  33785=>"101001100",
  33786=>"111101000",
  33787=>"110010111",
  33788=>"000001101",
  33789=>"010100000",
  33790=>"101000010",
  33791=>"111000100",
  33792=>"001111111",
  33793=>"111010111",
  33794=>"011100111",
  33795=>"101001110",
  33796=>"000000011",
  33797=>"001111101",
  33798=>"001110010",
  33799=>"011110111",
  33800=>"110000000",
  33801=>"101011001",
  33802=>"011100111",
  33803=>"011101111",
  33804=>"001110000",
  33805=>"000100000",
  33806=>"010011001",
  33807=>"111111000",
  33808=>"111001110",
  33809=>"110000001",
  33810=>"111100100",
  33811=>"110011110",
  33812=>"001101010",
  33813=>"011011110",
  33814=>"010100111",
  33815=>"111110000",
  33816=>"010001001",
  33817=>"101010101",
  33818=>"100100010",
  33819=>"001111100",
  33820=>"111111111",
  33821=>"101000110",
  33822=>"110001000",
  33823=>"001000111",
  33824=>"100011001",
  33825=>"100100101",
  33826=>"011100000",
  33827=>"101100101",
  33828=>"010101101",
  33829=>"110000100",
  33830=>"100100100",
  33831=>"111111010",
  33832=>"100010101",
  33833=>"001100001",
  33834=>"111110011",
  33835=>"010000010",
  33836=>"100010111",
  33837=>"010110111",
  33838=>"100011110",
  33839=>"111000000",
  33840=>"001101011",
  33841=>"000001010",
  33842=>"000100101",
  33843=>"111111110",
  33844=>"111100001",
  33845=>"111001111",
  33846=>"000110000",
  33847=>"101011101",
  33848=>"010110010",
  33849=>"001100001",
  33850=>"110111110",
  33851=>"001011100",
  33852=>"111011110",
  33853=>"001100011",
  33854=>"100010001",
  33855=>"110010000",
  33856=>"111111001",
  33857=>"111110000",
  33858=>"001000000",
  33859=>"111000100",
  33860=>"110010010",
  33861=>"110101101",
  33862=>"101101110",
  33863=>"001000101",
  33864=>"110010001",
  33865=>"111011111",
  33866=>"100111011",
  33867=>"000000101",
  33868=>"110101101",
  33869=>"000111011",
  33870=>"010100001",
  33871=>"010011000",
  33872=>"110101111",
  33873=>"000100101",
  33874=>"001011011",
  33875=>"110110010",
  33876=>"001110110",
  33877=>"010100100",
  33878=>"000001001",
  33879=>"111001011",
  33880=>"000100011",
  33881=>"100010011",
  33882=>"001100111",
  33883=>"000110000",
  33884=>"111001000",
  33885=>"100100001",
  33886=>"101011110",
  33887=>"001110000",
  33888=>"110011100",
  33889=>"111100010",
  33890=>"001010111",
  33891=>"100011000",
  33892=>"010110101",
  33893=>"000001001",
  33894=>"101001101",
  33895=>"111001100",
  33896=>"000001100",
  33897=>"110001111",
  33898=>"110000001",
  33899=>"001000110",
  33900=>"111101000",
  33901=>"100101011",
  33902=>"000101100",
  33903=>"110011100",
  33904=>"101110010",
  33905=>"111011011",
  33906=>"100000011",
  33907=>"011111101",
  33908=>"000001011",
  33909=>"111111011",
  33910=>"100000010",
  33911=>"110010100",
  33912=>"100100101",
  33913=>"001010101",
  33914=>"101001110",
  33915=>"000001101",
  33916=>"111011001",
  33917=>"010100000",
  33918=>"100011111",
  33919=>"110111001",
  33920=>"111010011",
  33921=>"000101000",
  33922=>"010101111",
  33923=>"000010001",
  33924=>"111001100",
  33925=>"000010110",
  33926=>"100011101",
  33927=>"101100110",
  33928=>"111101111",
  33929=>"000000000",
  33930=>"101000101",
  33931=>"111011100",
  33932=>"010110001",
  33933=>"100101101",
  33934=>"011111100",
  33935=>"010100100",
  33936=>"000011001",
  33937=>"101101001",
  33938=>"111111111",
  33939=>"001011101",
  33940=>"100100111",
  33941=>"001011101",
  33942=>"000101001",
  33943=>"011110110",
  33944=>"100111100",
  33945=>"010101110",
  33946=>"100011111",
  33947=>"010111111",
  33948=>"111111011",
  33949=>"011000101",
  33950=>"100000110",
  33951=>"111000110",
  33952=>"001100000",
  33953=>"000000101",
  33954=>"101110110",
  33955=>"011010110",
  33956=>"011001111",
  33957=>"001100101",
  33958=>"011111100",
  33959=>"101001000",
  33960=>"011110111",
  33961=>"111100010",
  33962=>"101000100",
  33963=>"101111111",
  33964=>"101100011",
  33965=>"100001001",
  33966=>"000100010",
  33967=>"011110011",
  33968=>"100010101",
  33969=>"010011001",
  33970=>"010111100",
  33971=>"000011101",
  33972=>"011100101",
  33973=>"001110001",
  33974=>"000100010",
  33975=>"111010000",
  33976=>"001101001",
  33977=>"100001000",
  33978=>"000001100",
  33979=>"011110011",
  33980=>"001110011",
  33981=>"100001001",
  33982=>"110011101",
  33983=>"011111011",
  33984=>"100101101",
  33985=>"001011010",
  33986=>"011110010",
  33987=>"101011011",
  33988=>"101110111",
  33989=>"011010100",
  33990=>"010000110",
  33991=>"101101111",
  33992=>"101100010",
  33993=>"001111111",
  33994=>"000011100",
  33995=>"110011101",
  33996=>"010010000",
  33997=>"101100011",
  33998=>"100000011",
  33999=>"110011000",
  34000=>"011011100",
  34001=>"100011100",
  34002=>"101101110",
  34003=>"111011110",
  34004=>"000111111",
  34005=>"000101100",
  34006=>"000110100",
  34007=>"110101000",
  34008=>"000101010",
  34009=>"100000000",
  34010=>"010010110",
  34011=>"010100000",
  34012=>"111111001",
  34013=>"110011101",
  34014=>"110001000",
  34015=>"101011011",
  34016=>"011100011",
  34017=>"000001000",
  34018=>"110100000",
  34019=>"110100011",
  34020=>"001000110",
  34021=>"001010111",
  34022=>"010010010",
  34023=>"000000110",
  34024=>"101001111",
  34025=>"011111100",
  34026=>"010000011",
  34027=>"111101011",
  34028=>"001111010",
  34029=>"101000011",
  34030=>"110101000",
  34031=>"111010111",
  34032=>"110111100",
  34033=>"010010000",
  34034=>"011010111",
  34035=>"110111110",
  34036=>"110000011",
  34037=>"000010000",
  34038=>"011011000",
  34039=>"101110001",
  34040=>"001011100",
  34041=>"000000001",
  34042=>"010000110",
  34043=>"010000000",
  34044=>"000000110",
  34045=>"101100111",
  34046=>"100111011",
  34047=>"010100101",
  34048=>"111111110",
  34049=>"011110001",
  34050=>"001011000",
  34051=>"000000100",
  34052=>"111010110",
  34053=>"011000101",
  34054=>"000111011",
  34055=>"110101111",
  34056=>"101001111",
  34057=>"011101000",
  34058=>"101110111",
  34059=>"110010001",
  34060=>"111011100",
  34061=>"010001001",
  34062=>"100010101",
  34063=>"010000001",
  34064=>"000000110",
  34065=>"000010000",
  34066=>"000001100",
  34067=>"111001110",
  34068=>"110001110",
  34069=>"011111001",
  34070=>"000101111",
  34071=>"000000101",
  34072=>"111000110",
  34073=>"000010100",
  34074=>"101010100",
  34075=>"000000011",
  34076=>"100000110",
  34077=>"110100010",
  34078=>"110111000",
  34079=>"000100001",
  34080=>"010101100",
  34081=>"011001100",
  34082=>"110101111",
  34083=>"000010101",
  34084=>"000011001",
  34085=>"101010100",
  34086=>"100110111",
  34087=>"001000011",
  34088=>"010100011",
  34089=>"111100011",
  34090=>"110010001",
  34091=>"100001111",
  34092=>"110001111",
  34093=>"011111010",
  34094=>"000011001",
  34095=>"101101011",
  34096=>"111101101",
  34097=>"101010011",
  34098=>"000001110",
  34099=>"111001001",
  34100=>"111100100",
  34101=>"111101100",
  34102=>"111101110",
  34103=>"011000001",
  34104=>"110111001",
  34105=>"000110011",
  34106=>"100000101",
  34107=>"011101100",
  34108=>"111101110",
  34109=>"110011001",
  34110=>"110001011",
  34111=>"110100011",
  34112=>"010100100",
  34113=>"110110110",
  34114=>"010011111",
  34115=>"100000111",
  34116=>"010010101",
  34117=>"111000010",
  34118=>"100000000",
  34119=>"110100001",
  34120=>"001101000",
  34121=>"000001011",
  34122=>"010000101",
  34123=>"100100101",
  34124=>"001110000",
  34125=>"100111000",
  34126=>"010011001",
  34127=>"110000111",
  34128=>"110011000",
  34129=>"000010101",
  34130=>"001000011",
  34131=>"001011010",
  34132=>"000101011",
  34133=>"001010001",
  34134=>"111000011",
  34135=>"001101000",
  34136=>"000101110",
  34137=>"001010100",
  34138=>"101111111",
  34139=>"111011001",
  34140=>"100010110",
  34141=>"100011101",
  34142=>"100011010",
  34143=>"001110001",
  34144=>"101100001",
  34145=>"110011010",
  34146=>"010110010",
  34147=>"000000110",
  34148=>"101000110",
  34149=>"001101111",
  34150=>"110000100",
  34151=>"100110111",
  34152=>"100110100",
  34153=>"100001100",
  34154=>"000010011",
  34155=>"101011010",
  34156=>"001111101",
  34157=>"110110000",
  34158=>"001011111",
  34159=>"101011111",
  34160=>"100100101",
  34161=>"001111010",
  34162=>"000011100",
  34163=>"011010011",
  34164=>"011111101",
  34165=>"010101101",
  34166=>"010101000",
  34167=>"110011011",
  34168=>"110110110",
  34169=>"010110100",
  34170=>"011111111",
  34171=>"111011101",
  34172=>"110100001",
  34173=>"011111000",
  34174=>"001111100",
  34175=>"010100000",
  34176=>"101010001",
  34177=>"111100110",
  34178=>"000010111",
  34179=>"001000111",
  34180=>"100111011",
  34181=>"101110000",
  34182=>"110010001",
  34183=>"001001010",
  34184=>"000101010",
  34185=>"000000010",
  34186=>"010001010",
  34187=>"000100000",
  34188=>"101101101",
  34189=>"011011111",
  34190=>"101000100",
  34191=>"000010111",
  34192=>"001011010",
  34193=>"001010000",
  34194=>"011011001",
  34195=>"100110001",
  34196=>"000011000",
  34197=>"001111000",
  34198=>"001001111",
  34199=>"100001000",
  34200=>"001100100",
  34201=>"011100001",
  34202=>"011001111",
  34203=>"000101000",
  34204=>"001010000",
  34205=>"011010111",
  34206=>"101000011",
  34207=>"111010111",
  34208=>"010100000",
  34209=>"110000110",
  34210=>"010101111",
  34211=>"011111001",
  34212=>"011101110",
  34213=>"011111000",
  34214=>"011101000",
  34215=>"000111101",
  34216=>"101001000",
  34217=>"100111000",
  34218=>"000111111",
  34219=>"111111100",
  34220=>"100001010",
  34221=>"001101110",
  34222=>"101001000",
  34223=>"011010100",
  34224=>"110010000",
  34225=>"100101100",
  34226=>"111110001",
  34227=>"111111010",
  34228=>"101000100",
  34229=>"011000000",
  34230=>"000000101",
  34231=>"111100100",
  34232=>"010000000",
  34233=>"011100101",
  34234=>"011111000",
  34235=>"111111111",
  34236=>"110001011",
  34237=>"110010111",
  34238=>"000001001",
  34239=>"001000011",
  34240=>"111001110",
  34241=>"001001110",
  34242=>"010001100",
  34243=>"011100111",
  34244=>"101111000",
  34245=>"010100000",
  34246=>"001001101",
  34247=>"001101000",
  34248=>"011010110",
  34249=>"011111101",
  34250=>"000001111",
  34251=>"001001111",
  34252=>"011111010",
  34253=>"001000011",
  34254=>"001011010",
  34255=>"011110111",
  34256=>"011111100",
  34257=>"000111000",
  34258=>"010010111",
  34259=>"000000000",
  34260=>"100101110",
  34261=>"001110010",
  34262=>"011001100",
  34263=>"011001111",
  34264=>"011001001",
  34265=>"100011100",
  34266=>"101000111",
  34267=>"000000100",
  34268=>"101000101",
  34269=>"000100000",
  34270=>"101101000",
  34271=>"100001110",
  34272=>"100111011",
  34273=>"011101000",
  34274=>"111111011",
  34275=>"100100000",
  34276=>"111000011",
  34277=>"101101100",
  34278=>"001100111",
  34279=>"000100010",
  34280=>"001011100",
  34281=>"000001001",
  34282=>"110101111",
  34283=>"011001100",
  34284=>"001110001",
  34285=>"111011001",
  34286=>"101110100",
  34287=>"000111010",
  34288=>"001001111",
  34289=>"110011011",
  34290=>"000101101",
  34291=>"010101000",
  34292=>"000010001",
  34293=>"100100100",
  34294=>"010111001",
  34295=>"111001000",
  34296=>"111011000",
  34297=>"111110100",
  34298=>"001001101",
  34299=>"101010101",
  34300=>"111011110",
  34301=>"011000100",
  34302=>"000000100",
  34303=>"010010100",
  34304=>"110010110",
  34305=>"011100100",
  34306=>"100101001",
  34307=>"101000100",
  34308=>"110011000",
  34309=>"000011110",
  34310=>"001000010",
  34311=>"100101010",
  34312=>"010011101",
  34313=>"110011111",
  34314=>"010111110",
  34315=>"111110000",
  34316=>"101011110",
  34317=>"011011111",
  34318=>"010001001",
  34319=>"110110111",
  34320=>"011001011",
  34321=>"100110101",
  34322=>"001010101",
  34323=>"101101001",
  34324=>"011011001",
  34325=>"010101100",
  34326=>"010000100",
  34327=>"111010100",
  34328=>"100000100",
  34329=>"001101010",
  34330=>"100101111",
  34331=>"101101000",
  34332=>"001111010",
  34333=>"011010110",
  34334=>"101011110",
  34335=>"100000110",
  34336=>"001101011",
  34337=>"000110000",
  34338=>"001011100",
  34339=>"000000000",
  34340=>"010101111",
  34341=>"011001001",
  34342=>"000000011",
  34343=>"110110101",
  34344=>"000000110",
  34345=>"101001000",
  34346=>"111110000",
  34347=>"010101000",
  34348=>"000111101",
  34349=>"010001100",
  34350=>"000000110",
  34351=>"111001001",
  34352=>"111000100",
  34353=>"000111010",
  34354=>"101000101",
  34355=>"101001011",
  34356=>"110101001",
  34357=>"111101001",
  34358=>"101010001",
  34359=>"101000100",
  34360=>"100101101",
  34361=>"100000000",
  34362=>"010101011",
  34363=>"110010101",
  34364=>"001000100",
  34365=>"010011111",
  34366=>"001001001",
  34367=>"001111101",
  34368=>"110011001",
  34369=>"111100110",
  34370=>"101001001",
  34371=>"001101111",
  34372=>"100100010",
  34373=>"010101011",
  34374=>"100001110",
  34375=>"101101111",
  34376=>"101011110",
  34377=>"010010001",
  34378=>"100110001",
  34379=>"011000101",
  34380=>"100100100",
  34381=>"101101111",
  34382=>"000111000",
  34383=>"111111001",
  34384=>"111111101",
  34385=>"001100000",
  34386=>"110010101",
  34387=>"101011110",
  34388=>"111101101",
  34389=>"100100011",
  34390=>"000111000",
  34391=>"011011000",
  34392=>"100100100",
  34393=>"010111110",
  34394=>"010010001",
  34395=>"001000010",
  34396=>"010100001",
  34397=>"111101111",
  34398=>"101011000",
  34399=>"001001101",
  34400=>"101000011",
  34401=>"111111001",
  34402=>"010010010",
  34403=>"010000111",
  34404=>"001000000",
  34405=>"110100111",
  34406=>"101000101",
  34407=>"100100000",
  34408=>"011011110",
  34409=>"001000110",
  34410=>"001001111",
  34411=>"101110001",
  34412=>"011001000",
  34413=>"011101011",
  34414=>"101010001",
  34415=>"011011101",
  34416=>"001101001",
  34417=>"101110000",
  34418=>"000001111",
  34419=>"111001111",
  34420=>"101101110",
  34421=>"110101000",
  34422=>"000111011",
  34423=>"011101011",
  34424=>"100010111",
  34425=>"101001001",
  34426=>"110000100",
  34427=>"110100110",
  34428=>"000000001",
  34429=>"001111001",
  34430=>"101010000",
  34431=>"010111101",
  34432=>"101111011",
  34433=>"100010000",
  34434=>"001010001",
  34435=>"010010100",
  34436=>"010110010",
  34437=>"110100000",
  34438=>"100110110",
  34439=>"000100000",
  34440=>"111110010",
  34441=>"010001100",
  34442=>"000001000",
  34443=>"110011111",
  34444=>"001100001",
  34445=>"101001110",
  34446=>"101010010",
  34447=>"001110100",
  34448=>"010011001",
  34449=>"000010100",
  34450=>"000011000",
  34451=>"000010111",
  34452=>"100110100",
  34453=>"000001110",
  34454=>"011110111",
  34455=>"000011000",
  34456=>"111111101",
  34457=>"111100111",
  34458=>"111011011",
  34459=>"000001101",
  34460=>"000010110",
  34461=>"111110000",
  34462=>"110100110",
  34463=>"100101110",
  34464=>"011110100",
  34465=>"001000111",
  34466=>"110000001",
  34467=>"110010100",
  34468=>"101101011",
  34469=>"111111110",
  34470=>"000100000",
  34471=>"111010111",
  34472=>"000010101",
  34473=>"111100100",
  34474=>"100110000",
  34475=>"101001110",
  34476=>"111100111",
  34477=>"111010110",
  34478=>"111101100",
  34479=>"110001100",
  34480=>"111000001",
  34481=>"100010011",
  34482=>"111001101",
  34483=>"000011010",
  34484=>"101111011",
  34485=>"011000100",
  34486=>"011001111",
  34487=>"100110110",
  34488=>"110001001",
  34489=>"110011001",
  34490=>"100010100",
  34491=>"001111100",
  34492=>"111000110",
  34493=>"011001010",
  34494=>"111001001",
  34495=>"010001011",
  34496=>"110101000",
  34497=>"110111101",
  34498=>"111110100",
  34499=>"100011011",
  34500=>"000011111",
  34501=>"100101011",
  34502=>"010001011",
  34503=>"011111101",
  34504=>"111100110",
  34505=>"000100001",
  34506=>"010110111",
  34507=>"010011100",
  34508=>"000100010",
  34509=>"001001001",
  34510=>"010010011",
  34511=>"011010110",
  34512=>"010101111",
  34513=>"110000111",
  34514=>"001001111",
  34515=>"111110001",
  34516=>"101101110",
  34517=>"101001000",
  34518=>"001110011",
  34519=>"001110100",
  34520=>"001000011",
  34521=>"000000000",
  34522=>"100100100",
  34523=>"111001000",
  34524=>"110011101",
  34525=>"010100101",
  34526=>"011000111",
  34527=>"001100010",
  34528=>"111111100",
  34529=>"000100110",
  34530=>"011010011",
  34531=>"110011000",
  34532=>"101101001",
  34533=>"111100100",
  34534=>"101001000",
  34535=>"101000110",
  34536=>"000000000",
  34537=>"000000000",
  34538=>"011100010",
  34539=>"111110101",
  34540=>"111011111",
  34541=>"010100111",
  34542=>"100010010",
  34543=>"101111111",
  34544=>"110110000",
  34545=>"010111111",
  34546=>"101111000",
  34547=>"010010001",
  34548=>"000101001",
  34549=>"100010001",
  34550=>"000111111",
  34551=>"111101001",
  34552=>"001110101",
  34553=>"011010001",
  34554=>"001100111",
  34555=>"110000010",
  34556=>"000000001",
  34557=>"010000110",
  34558=>"010010010",
  34559=>"001110000",
  34560=>"100011111",
  34561=>"111101110",
  34562=>"010000100",
  34563=>"111101100",
  34564=>"000011000",
  34565=>"110010010",
  34566=>"111010100",
  34567=>"101010011",
  34568=>"100010101",
  34569=>"100010101",
  34570=>"110010001",
  34571=>"011011101",
  34572=>"111110100",
  34573=>"000100000",
  34574=>"000001101",
  34575=>"101111000",
  34576=>"011011111",
  34577=>"110000001",
  34578=>"010110000",
  34579=>"010001111",
  34580=>"101111101",
  34581=>"001001000",
  34582=>"111111011",
  34583=>"011110000",
  34584=>"000101010",
  34585=>"011100001",
  34586=>"011000110",
  34587=>"100101011",
  34588=>"110111001",
  34589=>"100111110",
  34590=>"011001101",
  34591=>"001110110",
  34592=>"000001011",
  34593=>"000111011",
  34594=>"111100110",
  34595=>"001010000",
  34596=>"010111100",
  34597=>"110010000",
  34598=>"000001110",
  34599=>"110011111",
  34600=>"001010001",
  34601=>"111101011",
  34602=>"110011011",
  34603=>"010111110",
  34604=>"101100010",
  34605=>"111111101",
  34606=>"001010101",
  34607=>"010110110",
  34608=>"110000011",
  34609=>"010100110",
  34610=>"111100000",
  34611=>"110100011",
  34612=>"010011010",
  34613=>"101100010",
  34614=>"100111110",
  34615=>"011111100",
  34616=>"001110100",
  34617=>"010001111",
  34618=>"100111101",
  34619=>"101110001",
  34620=>"101010100",
  34621=>"110011011",
  34622=>"111010000",
  34623=>"001000110",
  34624=>"000001000",
  34625=>"001111000",
  34626=>"001010000",
  34627=>"001100010",
  34628=>"101101010",
  34629=>"100101010",
  34630=>"001011000",
  34631=>"111000110",
  34632=>"110000111",
  34633=>"001100011",
  34634=>"110101111",
  34635=>"011101010",
  34636=>"110100111",
  34637=>"011000010",
  34638=>"000011110",
  34639=>"111100110",
  34640=>"100101010",
  34641=>"000001100",
  34642=>"101111110",
  34643=>"101000001",
  34644=>"111101110",
  34645=>"100101100",
  34646=>"111101111",
  34647=>"010100100",
  34648=>"101111001",
  34649=>"111000101",
  34650=>"010000101",
  34651=>"111110101",
  34652=>"000001000",
  34653=>"010000110",
  34654=>"101100111",
  34655=>"101000110",
  34656=>"110100001",
  34657=>"010111001",
  34658=>"100010111",
  34659=>"010000100",
  34660=>"011101000",
  34661=>"111101001",
  34662=>"001111011",
  34663=>"010111010",
  34664=>"110111011",
  34665=>"010100001",
  34666=>"110000000",
  34667=>"111111011",
  34668=>"001111011",
  34669=>"011100101",
  34670=>"000101100",
  34671=>"001111111",
  34672=>"001011000",
  34673=>"010000111",
  34674=>"001010111",
  34675=>"000101110",
  34676=>"111100011",
  34677=>"111111000",
  34678=>"110101010",
  34679=>"010100001",
  34680=>"100000000",
  34681=>"110011101",
  34682=>"001111101",
  34683=>"001101111",
  34684=>"111010010",
  34685=>"010011010",
  34686=>"101111100",
  34687=>"011110011",
  34688=>"011010100",
  34689=>"000011111",
  34690=>"101001110",
  34691=>"011110110",
  34692=>"100010000",
  34693=>"001100100",
  34694=>"011111010",
  34695=>"000101100",
  34696=>"010111111",
  34697=>"011010100",
  34698=>"101110000",
  34699=>"101010010",
  34700=>"111110010",
  34701=>"010001001",
  34702=>"100101000",
  34703=>"101100100",
  34704=>"000010111",
  34705=>"000011001",
  34706=>"100000011",
  34707=>"111011111",
  34708=>"101111100",
  34709=>"111101101",
  34710=>"001100101",
  34711=>"011000010",
  34712=>"010011010",
  34713=>"000101011",
  34714=>"000111010",
  34715=>"110110100",
  34716=>"110001101",
  34717=>"111000111",
  34718=>"001100000",
  34719=>"010100011",
  34720=>"110111111",
  34721=>"111100011",
  34722=>"100011110",
  34723=>"100101100",
  34724=>"111000000",
  34725=>"100101100",
  34726=>"100101110",
  34727=>"110110111",
  34728=>"000001101",
  34729=>"001100001",
  34730=>"000001111",
  34731=>"011101011",
  34732=>"111000000",
  34733=>"110110000",
  34734=>"100110000",
  34735=>"101110000",
  34736=>"110110111",
  34737=>"010010001",
  34738=>"000000000",
  34739=>"011111101",
  34740=>"110101111",
  34741=>"111101110",
  34742=>"110011000",
  34743=>"110010000",
  34744=>"001110111",
  34745=>"001010001",
  34746=>"001011000",
  34747=>"011110000",
  34748=>"000010000",
  34749=>"111110011",
  34750=>"010011101",
  34751=>"100100110",
  34752=>"010101010",
  34753=>"000001111",
  34754=>"001010011",
  34755=>"011000101",
  34756=>"000001011",
  34757=>"001111101",
  34758=>"001110001",
  34759=>"000001110",
  34760=>"111001010",
  34761=>"101011101",
  34762=>"000100101",
  34763=>"111101000",
  34764=>"001110100",
  34765=>"101001110",
  34766=>"010110101",
  34767=>"111100101",
  34768=>"010011011",
  34769=>"111101001",
  34770=>"111011001",
  34771=>"010001000",
  34772=>"111001000",
  34773=>"010001010",
  34774=>"011001001",
  34775=>"000001011",
  34776=>"010011000",
  34777=>"011110011",
  34778=>"111110100",
  34779=>"011010010",
  34780=>"000101011",
  34781=>"000110100",
  34782=>"111110101",
  34783=>"000010000",
  34784=>"101011000",
  34785=>"111010110",
  34786=>"100101001",
  34787=>"011001000",
  34788=>"101001000",
  34789=>"100000111",
  34790=>"110100110",
  34791=>"010110111",
  34792=>"101000000",
  34793=>"001111111",
  34794=>"000110111",
  34795=>"100010001",
  34796=>"000001000",
  34797=>"011101111",
  34798=>"100001111",
  34799=>"011111010",
  34800=>"001100010",
  34801=>"000011101",
  34802=>"000001001",
  34803=>"001011001",
  34804=>"011101101",
  34805=>"010000010",
  34806=>"111011100",
  34807=>"000000110",
  34808=>"111001000",
  34809=>"111100000",
  34810=>"000110111",
  34811=>"000100111",
  34812=>"011001011",
  34813=>"010010010",
  34814=>"110111000",
  34815=>"111011000",
  34816=>"101100010",
  34817=>"000001110",
  34818=>"001100010",
  34819=>"110010011",
  34820=>"011011100",
  34821=>"010100001",
  34822=>"111110010",
  34823=>"101001111",
  34824=>"101011000",
  34825=>"101011110",
  34826=>"001011110",
  34827=>"111010011",
  34828=>"011111101",
  34829=>"110011100",
  34830=>"101100100",
  34831=>"000101000",
  34832=>"101100100",
  34833=>"011011010",
  34834=>"000000000",
  34835=>"010110101",
  34836=>"101011000",
  34837=>"101000011",
  34838=>"110000001",
  34839=>"100000011",
  34840=>"111010111",
  34841=>"000000001",
  34842=>"011010001",
  34843=>"111101001",
  34844=>"101000110",
  34845=>"001111000",
  34846=>"011010001",
  34847=>"110010001",
  34848=>"001100010",
  34849=>"001111110",
  34850=>"011111100",
  34851=>"011000111",
  34852=>"011001101",
  34853=>"100100110",
  34854=>"011111000",
  34855=>"110000111",
  34856=>"110000010",
  34857=>"100111111",
  34858=>"111101101",
  34859=>"100001100",
  34860=>"110101100",
  34861=>"101000110",
  34862=>"111011101",
  34863=>"100110100",
  34864=>"001101001",
  34865=>"100110000",
  34866=>"111111111",
  34867=>"001110011",
  34868=>"111101010",
  34869=>"010010101",
  34870=>"000010011",
  34871=>"010110010",
  34872=>"110010001",
  34873=>"110001011",
  34874=>"101111110",
  34875=>"110011011",
  34876=>"011001111",
  34877=>"011001110",
  34878=>"111100111",
  34879=>"001011101",
  34880=>"111101011",
  34881=>"000110011",
  34882=>"011001001",
  34883=>"011101011",
  34884=>"000010010",
  34885=>"001000011",
  34886=>"100101000",
  34887=>"111100010",
  34888=>"111010011",
  34889=>"101010101",
  34890=>"010011010",
  34891=>"101001010",
  34892=>"010010000",
  34893=>"111101110",
  34894=>"100100000",
  34895=>"010100111",
  34896=>"011001111",
  34897=>"010110010",
  34898=>"010101010",
  34899=>"011000101",
  34900=>"001010110",
  34901=>"010000000",
  34902=>"100110110",
  34903=>"100111110",
  34904=>"100010100",
  34905=>"101111011",
  34906=>"000001010",
  34907=>"000110010",
  34908=>"000010010",
  34909=>"110110110",
  34910=>"001110111",
  34911=>"001010100",
  34912=>"000101110",
  34913=>"100001010",
  34914=>"001000011",
  34915=>"010000011",
  34916=>"110100011",
  34917=>"110011000",
  34918=>"100100110",
  34919=>"010100101",
  34920=>"100000111",
  34921=>"111010100",
  34922=>"110001010",
  34923=>"001010101",
  34924=>"100110101",
  34925=>"111000010",
  34926=>"001001001",
  34927=>"001100010",
  34928=>"000000000",
  34929=>"010101011",
  34930=>"111000000",
  34931=>"101110011",
  34932=>"011111111",
  34933=>"011100101",
  34934=>"101011100",
  34935=>"000111101",
  34936=>"100011100",
  34937=>"001101100",
  34938=>"001010101",
  34939=>"000010000",
  34940=>"001000101",
  34941=>"000011100",
  34942=>"011000001",
  34943=>"011010000",
  34944=>"010010111",
  34945=>"110010000",
  34946=>"111010001",
  34947=>"000100111",
  34948=>"011010000",
  34949=>"111101010",
  34950=>"111001110",
  34951=>"111111010",
  34952=>"000101010",
  34953=>"101010110",
  34954=>"100110111",
  34955=>"011101100",
  34956=>"101101000",
  34957=>"111111101",
  34958=>"110101011",
  34959=>"001000101",
  34960=>"110010101",
  34961=>"111011001",
  34962=>"111110111",
  34963=>"010111111",
  34964=>"011000001",
  34965=>"110101001",
  34966=>"100000111",
  34967=>"001111001",
  34968=>"111101100",
  34969=>"111001111",
  34970=>"110111111",
  34971=>"011100011",
  34972=>"011101010",
  34973=>"111100110",
  34974=>"111001101",
  34975=>"111011011",
  34976=>"000000111",
  34977=>"011100111",
  34978=>"001000110",
  34979=>"000010010",
  34980=>"011101100",
  34981=>"010111101",
  34982=>"001100111",
  34983=>"000000010",
  34984=>"101010010",
  34985=>"110110001",
  34986=>"001111011",
  34987=>"011110001",
  34988=>"001000110",
  34989=>"011001110",
  34990=>"000110000",
  34991=>"000011111",
  34992=>"000010010",
  34993=>"000110101",
  34994=>"101101000",
  34995=>"000000010",
  34996=>"001000110",
  34997=>"100101000",
  34998=>"000011110",
  34999=>"010000010",
  35000=>"000101000",
  35001=>"110110110",
  35002=>"000000110",
  35003=>"110101110",
  35004=>"110110000",
  35005=>"111100000",
  35006=>"001010011",
  35007=>"100100011",
  35008=>"100010011",
  35009=>"011011001",
  35010=>"100001101",
  35011=>"111111011",
  35012=>"100000001",
  35013=>"001100111",
  35014=>"010001000",
  35015=>"101100111",
  35016=>"111111000",
  35017=>"111000001",
  35018=>"010011011",
  35019=>"011110001",
  35020=>"100000110",
  35021=>"011100001",
  35022=>"101111010",
  35023=>"010111001",
  35024=>"010100000",
  35025=>"000111111",
  35026=>"011101101",
  35027=>"001111010",
  35028=>"000000100",
  35029=>"010001011",
  35030=>"000000001",
  35031=>"000011001",
  35032=>"101011100",
  35033=>"001011010",
  35034=>"001000001",
  35035=>"111111100",
  35036=>"011110001",
  35037=>"011101001",
  35038=>"000001000",
  35039=>"001000000",
  35040=>"001111111",
  35041=>"000001000",
  35042=>"111111101",
  35043=>"000000000",
  35044=>"001111100",
  35045=>"111100001",
  35046=>"010100001",
  35047=>"000110111",
  35048=>"000111001",
  35049=>"110111101",
  35050=>"001110001",
  35051=>"010000010",
  35052=>"001010001",
  35053=>"100100010",
  35054=>"111101111",
  35055=>"000000000",
  35056=>"010001001",
  35057=>"110000011",
  35058=>"110110111",
  35059=>"001111000",
  35060=>"000100010",
  35061=>"010001001",
  35062=>"010101110",
  35063=>"101100001",
  35064=>"000111101",
  35065=>"101110110",
  35066=>"010011001",
  35067=>"001100110",
  35068=>"110111000",
  35069=>"000011000",
  35070=>"100111111",
  35071=>"101000001",
  35072=>"110010001",
  35073=>"010000110",
  35074=>"111100000",
  35075=>"111101100",
  35076=>"110111110",
  35077=>"011000111",
  35078=>"100011011",
  35079=>"100011100",
  35080=>"000000001",
  35081=>"101001111",
  35082=>"010100010",
  35083=>"101011111",
  35084=>"000010110",
  35085=>"000001000",
  35086=>"111100011",
  35087=>"000100000",
  35088=>"100011011",
  35089=>"101011111",
  35090=>"000001101",
  35091=>"001011010",
  35092=>"111011011",
  35093=>"110101011",
  35094=>"011010000",
  35095=>"101001101",
  35096=>"111000001",
  35097=>"111110111",
  35098=>"101100100",
  35099=>"101001010",
  35100=>"110001100",
  35101=>"011111100",
  35102=>"001010010",
  35103=>"110100011",
  35104=>"010110010",
  35105=>"010110000",
  35106=>"100001100",
  35107=>"101101011",
  35108=>"010101011",
  35109=>"000110101",
  35110=>"111111010",
  35111=>"101011111",
  35112=>"001001011",
  35113=>"111101011",
  35114=>"010011001",
  35115=>"010001111",
  35116=>"001010001",
  35117=>"010111111",
  35118=>"110011110",
  35119=>"010000100",
  35120=>"000101101",
  35121=>"110110100",
  35122=>"110111100",
  35123=>"010001001",
  35124=>"011011011",
  35125=>"101011111",
  35126=>"110110101",
  35127=>"000010000",
  35128=>"111110110",
  35129=>"000010010",
  35130=>"000111010",
  35131=>"011010000",
  35132=>"000100111",
  35133=>"111111001",
  35134=>"011011101",
  35135=>"100010010",
  35136=>"000100010",
  35137=>"111101101",
  35138=>"001000000",
  35139=>"111000100",
  35140=>"011110001",
  35141=>"110000100",
  35142=>"111100101",
  35143=>"011001000",
  35144=>"110011010",
  35145=>"011110001",
  35146=>"100000011",
  35147=>"010000101",
  35148=>"100111111",
  35149=>"000110001",
  35150=>"001101001",
  35151=>"010101001",
  35152=>"010110110",
  35153=>"010101110",
  35154=>"010001100",
  35155=>"000010111",
  35156=>"001000110",
  35157=>"110100101",
  35158=>"011000000",
  35159=>"101111010",
  35160=>"001101011",
  35161=>"001111001",
  35162=>"110111001",
  35163=>"001010011",
  35164=>"010101100",
  35165=>"011001010",
  35166=>"101101111",
  35167=>"111001101",
  35168=>"110100101",
  35169=>"100001111",
  35170=>"100101111",
  35171=>"111001010",
  35172=>"101100101",
  35173=>"100111111",
  35174=>"110110010",
  35175=>"000110111",
  35176=>"101001010",
  35177=>"100001011",
  35178=>"101111101",
  35179=>"011111011",
  35180=>"011110001",
  35181=>"111100001",
  35182=>"111100001",
  35183=>"110110111",
  35184=>"111111001",
  35185=>"100101101",
  35186=>"010000010",
  35187=>"001000001",
  35188=>"000010010",
  35189=>"011110011",
  35190=>"000011010",
  35191=>"010001001",
  35192=>"111110010",
  35193=>"101000111",
  35194=>"010000011",
  35195=>"001101010",
  35196=>"011010010",
  35197=>"000010010",
  35198=>"000010100",
  35199=>"001011100",
  35200=>"000111010",
  35201=>"000011110",
  35202=>"111001011",
  35203=>"001010100",
  35204=>"110011111",
  35205=>"101100001",
  35206=>"011011001",
  35207=>"110110011",
  35208=>"100111111",
  35209=>"010110000",
  35210=>"010000000",
  35211=>"110101110",
  35212=>"011011011",
  35213=>"110111101",
  35214=>"101100111",
  35215=>"001010001",
  35216=>"101011111",
  35217=>"011110101",
  35218=>"011010000",
  35219=>"100010100",
  35220=>"111101000",
  35221=>"000100100",
  35222=>"100010010",
  35223=>"110010000",
  35224=>"011001100",
  35225=>"101101001",
  35226=>"000110001",
  35227=>"010011000",
  35228=>"011111001",
  35229=>"010010110",
  35230=>"111110000",
  35231=>"111000111",
  35232=>"100000000",
  35233=>"101000111",
  35234=>"000001100",
  35235=>"001111101",
  35236=>"010111010",
  35237=>"110010101",
  35238=>"101100000",
  35239=>"001010100",
  35240=>"011010100",
  35241=>"110001011",
  35242=>"100110010",
  35243=>"100110101",
  35244=>"010011100",
  35245=>"010000001",
  35246=>"000011010",
  35247=>"001001010",
  35248=>"000000000",
  35249=>"111000110",
  35250=>"101010101",
  35251=>"010000010",
  35252=>"111000110",
  35253=>"011010011",
  35254=>"001111001",
  35255=>"000111010",
  35256=>"110100101",
  35257=>"010100101",
  35258=>"000100100",
  35259=>"110010000",
  35260=>"101101110",
  35261=>"000101110",
  35262=>"010100101",
  35263=>"010100010",
  35264=>"011111011",
  35265=>"101111000",
  35266=>"001011011",
  35267=>"110000111",
  35268=>"010000000",
  35269=>"101000101",
  35270=>"010000101",
  35271=>"111000101",
  35272=>"111101110",
  35273=>"111011011",
  35274=>"100000100",
  35275=>"011101100",
  35276=>"111111111",
  35277=>"001101010",
  35278=>"000000000",
  35279=>"111001000",
  35280=>"101011111",
  35281=>"110111000",
  35282=>"010110010",
  35283=>"000010001",
  35284=>"010111011",
  35285=>"110010011",
  35286=>"001101010",
  35287=>"010010010",
  35288=>"001000000",
  35289=>"011010110",
  35290=>"100000100",
  35291=>"011010110",
  35292=>"101011111",
  35293=>"011001110",
  35294=>"100101111",
  35295=>"001111101",
  35296=>"100101110",
  35297=>"001001000",
  35298=>"000001110",
  35299=>"101000011",
  35300=>"000010111",
  35301=>"110101011",
  35302=>"100001100",
  35303=>"011010100",
  35304=>"001101010",
  35305=>"101110010",
  35306=>"010000000",
  35307=>"010111101",
  35308=>"110111110",
  35309=>"110101000",
  35310=>"011010100",
  35311=>"111000100",
  35312=>"111111010",
  35313=>"110011101",
  35314=>"101010101",
  35315=>"000010001",
  35316=>"110111011",
  35317=>"001101001",
  35318=>"110101110",
  35319=>"101111110",
  35320=>"101100010",
  35321=>"100110000",
  35322=>"000001001",
  35323=>"000010011",
  35324=>"010010110",
  35325=>"111010100",
  35326=>"010110010",
  35327=>"101101010",
  35328=>"101101111",
  35329=>"101001001",
  35330=>"101011011",
  35331=>"100011110",
  35332=>"001100101",
  35333=>"111010110",
  35334=>"011011101",
  35335=>"110101101",
  35336=>"010110111",
  35337=>"011010000",
  35338=>"000110010",
  35339=>"100110010",
  35340=>"011100000",
  35341=>"111101010",
  35342=>"010011010",
  35343=>"110110110",
  35344=>"101011111",
  35345=>"111101110",
  35346=>"111101011",
  35347=>"101111111",
  35348=>"010100111",
  35349=>"100011000",
  35350=>"111101010",
  35351=>"011110010",
  35352=>"011010101",
  35353=>"101100010",
  35354=>"100101000",
  35355=>"001001001",
  35356=>"010001111",
  35357=>"110010001",
  35358=>"101110110",
  35359=>"001110001",
  35360=>"100100100",
  35361=>"001000101",
  35362=>"111011111",
  35363=>"001000110",
  35364=>"110100000",
  35365=>"101000110",
  35366=>"100010000",
  35367=>"100110111",
  35368=>"001011010",
  35369=>"011010100",
  35370=>"111101111",
  35371=>"110010101",
  35372=>"101001110",
  35373=>"110010000",
  35374=>"011111011",
  35375=>"000000010",
  35376=>"100001101",
  35377=>"111100101",
  35378=>"001011010",
  35379=>"011110100",
  35380=>"111011111",
  35381=>"001100001",
  35382=>"000010001",
  35383=>"001011000",
  35384=>"101100111",
  35385=>"111010001",
  35386=>"000000000",
  35387=>"011111100",
  35388=>"101011001",
  35389=>"111101110",
  35390=>"111000111",
  35391=>"100100101",
  35392=>"010001111",
  35393=>"110000100",
  35394=>"010110010",
  35395=>"000010011",
  35396=>"110101101",
  35397=>"100000101",
  35398=>"001001111",
  35399=>"111011100",
  35400=>"010011110",
  35401=>"110111110",
  35402=>"111001100",
  35403=>"110011010",
  35404=>"000001100",
  35405=>"000011001",
  35406=>"101100000",
  35407=>"010111100",
  35408=>"010101111",
  35409=>"011100100",
  35410=>"000101010",
  35411=>"111100011",
  35412=>"001010011",
  35413=>"100110011",
  35414=>"001111001",
  35415=>"010111111",
  35416=>"000010010",
  35417=>"101100111",
  35418=>"000100101",
  35419=>"111011110",
  35420=>"000010000",
  35421=>"000100011",
  35422=>"011011101",
  35423=>"100000000",
  35424=>"101110110",
  35425=>"010010011",
  35426=>"101000100",
  35427=>"011000011",
  35428=>"010100101",
  35429=>"011101111",
  35430=>"110111101",
  35431=>"000010110",
  35432=>"100110001",
  35433=>"011011010",
  35434=>"000111001",
  35435=>"000101011",
  35436=>"001011111",
  35437=>"000100101",
  35438=>"100100011",
  35439=>"000111110",
  35440=>"110000011",
  35441=>"000001100",
  35442=>"101001001",
  35443=>"110001000",
  35444=>"001010011",
  35445=>"001100111",
  35446=>"101001001",
  35447=>"001010001",
  35448=>"001010001",
  35449=>"010000100",
  35450=>"010011001",
  35451=>"101001011",
  35452=>"111000001",
  35453=>"100011011",
  35454=>"001111100",
  35455=>"111001011",
  35456=>"110010111",
  35457=>"101011111",
  35458=>"101100111",
  35459=>"100100111",
  35460=>"101110011",
  35461=>"010010000",
  35462=>"101010000",
  35463=>"111010001",
  35464=>"001100010",
  35465=>"100111100",
  35466=>"101110100",
  35467=>"100110101",
  35468=>"011101101",
  35469=>"011101001",
  35470=>"100111110",
  35471=>"010011101",
  35472=>"101101011",
  35473=>"100110100",
  35474=>"000001010",
  35475=>"101111011",
  35476=>"101101100",
  35477=>"011001000",
  35478=>"001100011",
  35479=>"100110100",
  35480=>"000101100",
  35481=>"111110101",
  35482=>"010100001",
  35483=>"110100111",
  35484=>"111001111",
  35485=>"111000001",
  35486=>"100100111",
  35487=>"010101011",
  35488=>"011101111",
  35489=>"001100010",
  35490=>"010101011",
  35491=>"010011110",
  35492=>"100100100",
  35493=>"000010110",
  35494=>"111010110",
  35495=>"011011110",
  35496=>"000111000",
  35497=>"011001011",
  35498=>"100110000",
  35499=>"011000111",
  35500=>"001000001",
  35501=>"000101000",
  35502=>"110000000",
  35503=>"010000111",
  35504=>"010001101",
  35505=>"001000110",
  35506=>"111100101",
  35507=>"001100110",
  35508=>"000111001",
  35509=>"010000011",
  35510=>"010010101",
  35511=>"111011011",
  35512=>"010100010",
  35513=>"110000001",
  35514=>"101000101",
  35515=>"110010111",
  35516=>"110100010",
  35517=>"000011100",
  35518=>"100011110",
  35519=>"001111110",
  35520=>"011010011",
  35521=>"100100011",
  35522=>"100011000",
  35523=>"101000000",
  35524=>"011010010",
  35525=>"010011010",
  35526=>"110011111",
  35527=>"000001100",
  35528=>"011010000",
  35529=>"001101111",
  35530=>"001001011",
  35531=>"010111111",
  35532=>"011111011",
  35533=>"101101001",
  35534=>"110100111",
  35535=>"011011000",
  35536=>"101000110",
  35537=>"111111101",
  35538=>"111110110",
  35539=>"010100101",
  35540=>"100010001",
  35541=>"100000100",
  35542=>"010000010",
  35543=>"100100010",
  35544=>"010001111",
  35545=>"111011110",
  35546=>"101010011",
  35547=>"110100110",
  35548=>"100011000",
  35549=>"011001011",
  35550=>"000001100",
  35551=>"010100000",
  35552=>"000110101",
  35553=>"000111110",
  35554=>"000111111",
  35555=>"010011101",
  35556=>"100011000",
  35557=>"101011001",
  35558=>"100100011",
  35559=>"110001110",
  35560=>"011111010",
  35561=>"101101110",
  35562=>"110111010",
  35563=>"011101111",
  35564=>"010000000",
  35565=>"010110111",
  35566=>"111110000",
  35567=>"011110011",
  35568=>"111111000",
  35569=>"001001110",
  35570=>"001101011",
  35571=>"001001111",
  35572=>"010110101",
  35573=>"010100111",
  35574=>"101001100",
  35575=>"001010010",
  35576=>"011110011",
  35577=>"111001000",
  35578=>"111000001",
  35579=>"001100000",
  35580=>"100011100",
  35581=>"101100000",
  35582=>"111100001",
  35583=>"010101110",
  35584=>"111001100",
  35585=>"011100010",
  35586=>"000101100",
  35587=>"101111101",
  35588=>"001001111",
  35589=>"111001111",
  35590=>"011101101",
  35591=>"010100110",
  35592=>"110110010",
  35593=>"000111000",
  35594=>"001000001",
  35595=>"101010101",
  35596=>"110111100",
  35597=>"111100100",
  35598=>"110100010",
  35599=>"101110000",
  35600=>"100110011",
  35601=>"000101010",
  35602=>"001101001",
  35603=>"001000010",
  35604=>"100011001",
  35605=>"011000010",
  35606=>"111101110",
  35607=>"000100000",
  35608=>"101000110",
  35609=>"110011100",
  35610=>"101000010",
  35611=>"110000101",
  35612=>"011100110",
  35613=>"100111011",
  35614=>"000111000",
  35615=>"011100001",
  35616=>"111111001",
  35617=>"111101011",
  35618=>"001001101",
  35619=>"011011110",
  35620=>"010110000",
  35621=>"000000010",
  35622=>"010000001",
  35623=>"110010111",
  35624=>"001101101",
  35625=>"111101111",
  35626=>"111111011",
  35627=>"011011101",
  35628=>"011111001",
  35629=>"100010110",
  35630=>"010100000",
  35631=>"101110100",
  35632=>"000000110",
  35633=>"111011011",
  35634=>"010100000",
  35635=>"100111011",
  35636=>"001100000",
  35637=>"001010011",
  35638=>"100100000",
  35639=>"100010100",
  35640=>"001000001",
  35641=>"000010010",
  35642=>"101101110",
  35643=>"011101100",
  35644=>"101001001",
  35645=>"111001100",
  35646=>"100010000",
  35647=>"100001101",
  35648=>"110111101",
  35649=>"000000100",
  35650=>"000101101",
  35651=>"001001011",
  35652=>"000000000",
  35653=>"111011110",
  35654=>"011101110",
  35655=>"101010111",
  35656=>"011110000",
  35657=>"010011010",
  35658=>"111000111",
  35659=>"111110110",
  35660=>"010000110",
  35661=>"000101101",
  35662=>"001000100",
  35663=>"001001111",
  35664=>"001001000",
  35665=>"100110001",
  35666=>"110110000",
  35667=>"101101111",
  35668=>"110011011",
  35669=>"101011011",
  35670=>"011100000",
  35671=>"010101111",
  35672=>"111011010",
  35673=>"100011001",
  35674=>"011101111",
  35675=>"111001000",
  35676=>"100000001",
  35677=>"000110100",
  35678=>"101010001",
  35679=>"000000001",
  35680=>"100100100",
  35681=>"011011000",
  35682=>"111010010",
  35683=>"100111100",
  35684=>"011010111",
  35685=>"101100111",
  35686=>"101011011",
  35687=>"001110001",
  35688=>"101000000",
  35689=>"110010010",
  35690=>"101110001",
  35691=>"000010101",
  35692=>"010100111",
  35693=>"111010001",
  35694=>"111101100",
  35695=>"001100101",
  35696=>"011000100",
  35697=>"111001001",
  35698=>"100000101",
  35699=>"001100000",
  35700=>"000110011",
  35701=>"010010011",
  35702=>"110110111",
  35703=>"001011111",
  35704=>"110110100",
  35705=>"011011001",
  35706=>"111001100",
  35707=>"110110000",
  35708=>"110110010",
  35709=>"001101001",
  35710=>"100101011",
  35711=>"001111100",
  35712=>"110000001",
  35713=>"100100101",
  35714=>"101111101",
  35715=>"011011101",
  35716=>"111011001",
  35717=>"111000101",
  35718=>"111001111",
  35719=>"011100111",
  35720=>"001101110",
  35721=>"100001001",
  35722=>"111000000",
  35723=>"101001001",
  35724=>"110001111",
  35725=>"110100110",
  35726=>"000101111",
  35727=>"111011101",
  35728=>"010010011",
  35729=>"011011101",
  35730=>"001011011",
  35731=>"101011111",
  35732=>"110101100",
  35733=>"001011010",
  35734=>"110111010",
  35735=>"010010100",
  35736=>"001111110",
  35737=>"111110100",
  35738=>"100011011",
  35739=>"001101010",
  35740=>"110001111",
  35741=>"111110111",
  35742=>"101011100",
  35743=>"110011010",
  35744=>"111001001",
  35745=>"010001111",
  35746=>"110111111",
  35747=>"111111100",
  35748=>"100011000",
  35749=>"101000011",
  35750=>"010110011",
  35751=>"001001001",
  35752=>"010100100",
  35753=>"111100111",
  35754=>"001101111",
  35755=>"110010010",
  35756=>"001110010",
  35757=>"010001000",
  35758=>"011110010",
  35759=>"011101011",
  35760=>"111001100",
  35761=>"010010001",
  35762=>"011110101",
  35763=>"010011111",
  35764=>"011010001",
  35765=>"100010000",
  35766=>"101101010",
  35767=>"000001111",
  35768=>"101100010",
  35769=>"001011011",
  35770=>"111001000",
  35771=>"011101100",
  35772=>"001011101",
  35773=>"000000010",
  35774=>"101000101",
  35775=>"110110001",
  35776=>"010011110",
  35777=>"001100001",
  35778=>"111101101",
  35779=>"011101000",
  35780=>"110110100",
  35781=>"010100111",
  35782=>"000101101",
  35783=>"111101000",
  35784=>"000100010",
  35785=>"000001000",
  35786=>"111100101",
  35787=>"001010100",
  35788=>"110010011",
  35789=>"010110001",
  35790=>"011000101",
  35791=>"100001010",
  35792=>"100110101",
  35793=>"000010110",
  35794=>"111111111",
  35795=>"000110100",
  35796=>"100110000",
  35797=>"111111100",
  35798=>"001000100",
  35799=>"101100111",
  35800=>"001011111",
  35801=>"001101111",
  35802=>"100100110",
  35803=>"110010011",
  35804=>"010001111",
  35805=>"111100101",
  35806=>"110011001",
  35807=>"110100001",
  35808=>"001110001",
  35809=>"011111111",
  35810=>"000010110",
  35811=>"010001110",
  35812=>"001011000",
  35813=>"101100110",
  35814=>"101111010",
  35815=>"011110101",
  35816=>"101101011",
  35817=>"101100101",
  35818=>"000010010",
  35819=>"010110110",
  35820=>"111000100",
  35821=>"010101101",
  35822=>"010111111",
  35823=>"110100111",
  35824=>"111011011",
  35825=>"100011010",
  35826=>"100000100",
  35827=>"110001001",
  35828=>"011111100",
  35829=>"100001111",
  35830=>"101011001",
  35831=>"010010111",
  35832=>"011100101",
  35833=>"110010010",
  35834=>"101111011",
  35835=>"010101010",
  35836=>"110010110",
  35837=>"001100011",
  35838=>"111110110",
  35839=>"100110001",
  35840=>"110111111",
  35841=>"100010101",
  35842=>"011011111",
  35843=>"000110011",
  35844=>"110011110",
  35845=>"011010000",
  35846=>"111100100",
  35847=>"101110000",
  35848=>"010101011",
  35849=>"100001001",
  35850=>"001000000",
  35851=>"100101101",
  35852=>"100100101",
  35853=>"001010010",
  35854=>"100111111",
  35855=>"110110111",
  35856=>"101010001",
  35857=>"111101010",
  35858=>"110101110",
  35859=>"001001011",
  35860=>"000001110",
  35861=>"001011101",
  35862=>"001110000",
  35863=>"001010010",
  35864=>"000010000",
  35865=>"111000011",
  35866=>"000111000",
  35867=>"100111111",
  35868=>"101010101",
  35869=>"011011010",
  35870=>"001100001",
  35871=>"010111010",
  35872=>"101010010",
  35873=>"101111000",
  35874=>"010111000",
  35875=>"011010000",
  35876=>"101100011",
  35877=>"110010010",
  35878=>"000100111",
  35879=>"111100110",
  35880=>"001000000",
  35881=>"111011100",
  35882=>"111010111",
  35883=>"111101111",
  35884=>"110001100",
  35885=>"111100100",
  35886=>"000101110",
  35887=>"110111110",
  35888=>"011111000",
  35889=>"100001001",
  35890=>"010000010",
  35891=>"110111000",
  35892=>"111111110",
  35893=>"010001110",
  35894=>"100001101",
  35895=>"100011010",
  35896=>"001001101",
  35897=>"011111101",
  35898=>"011010100",
  35899=>"001100010",
  35900=>"001010111",
  35901=>"001001011",
  35902=>"001110001",
  35903=>"000110010",
  35904=>"000010010",
  35905=>"111000001",
  35906=>"011100000",
  35907=>"100111010",
  35908=>"110110100",
  35909=>"111011011",
  35910=>"111111101",
  35911=>"011100100",
  35912=>"100010100",
  35913=>"001011100",
  35914=>"101010100",
  35915=>"001001101",
  35916=>"111100100",
  35917=>"101010000",
  35918=>"100101011",
  35919=>"101001000",
  35920=>"010110010",
  35921=>"000110001",
  35922=>"100101110",
  35923=>"111101010",
  35924=>"100110011",
  35925=>"110111001",
  35926=>"101010100",
  35927=>"000010010",
  35928=>"111011010",
  35929=>"101101000",
  35930=>"100001000",
  35931=>"101011001",
  35932=>"001000101",
  35933=>"000100000",
  35934=>"110010011",
  35935=>"011100000",
  35936=>"100111100",
  35937=>"011110101",
  35938=>"101011011",
  35939=>"010110010",
  35940=>"101011101",
  35941=>"011011111",
  35942=>"011001110",
  35943=>"000011000",
  35944=>"010110010",
  35945=>"011111011",
  35946=>"111011001",
  35947=>"001001100",
  35948=>"000101011",
  35949=>"111110111",
  35950=>"101100011",
  35951=>"101011000",
  35952=>"011111010",
  35953=>"000011101",
  35954=>"010111000",
  35955=>"101010101",
  35956=>"010100000",
  35957=>"101101011",
  35958=>"011110110",
  35959=>"111100101",
  35960=>"000100110",
  35961=>"100000000",
  35962=>"110111100",
  35963=>"010101110",
  35964=>"110010001",
  35965=>"101110111",
  35966=>"100101110",
  35967=>"011000011",
  35968=>"011100111",
  35969=>"011001001",
  35970=>"101111110",
  35971=>"100101101",
  35972=>"011111011",
  35973=>"001001100",
  35974=>"110111111",
  35975=>"101111010",
  35976=>"110000000",
  35977=>"000010101",
  35978=>"001000101",
  35979=>"010100010",
  35980=>"100000111",
  35981=>"000011011",
  35982=>"010100001",
  35983=>"010000001",
  35984=>"110000111",
  35985=>"111110111",
  35986=>"011010100",
  35987=>"110100011",
  35988=>"010011101",
  35989=>"101000110",
  35990=>"111000010",
  35991=>"000000000",
  35992=>"011010100",
  35993=>"111010111",
  35994=>"001011100",
  35995=>"100010010",
  35996=>"110010011",
  35997=>"100111001",
  35998=>"111110000",
  35999=>"100011111",
  36000=>"101110000",
  36001=>"001111111",
  36002=>"000010000",
  36003=>"010100101",
  36004=>"110010100",
  36005=>"110000110",
  36006=>"100101100",
  36007=>"011010111",
  36008=>"111111100",
  36009=>"101111111",
  36010=>"110001010",
  36011=>"000010000",
  36012=>"101100010",
  36013=>"011011000",
  36014=>"001110101",
  36015=>"100000000",
  36016=>"010011001",
  36017=>"111110000",
  36018=>"110011110",
  36019=>"110110000",
  36020=>"000101111",
  36021=>"000000100",
  36022=>"110110010",
  36023=>"010011001",
  36024=>"010000100",
  36025=>"101110101",
  36026=>"001000111",
  36027=>"000100111",
  36028=>"110010000",
  36029=>"101100010",
  36030=>"010110011",
  36031=>"001000000",
  36032=>"000101100",
  36033=>"110101011",
  36034=>"000010001",
  36035=>"100110111",
  36036=>"111100100",
  36037=>"101000100",
  36038=>"000110011",
  36039=>"110000101",
  36040=>"110001111",
  36041=>"100011110",
  36042=>"110111011",
  36043=>"011011010",
  36044=>"101100111",
  36045=>"001100110",
  36046=>"110100111",
  36047=>"011110011",
  36048=>"001000100",
  36049=>"000110110",
  36050=>"101111101",
  36051=>"101110011",
  36052=>"011100110",
  36053=>"111011000",
  36054=>"101001011",
  36055=>"100010000",
  36056=>"000001010",
  36057=>"011110000",
  36058=>"000101000",
  36059=>"001110101",
  36060=>"110000010",
  36061=>"000101100",
  36062=>"110111111",
  36063=>"000101101",
  36064=>"001010001",
  36065=>"011000000",
  36066=>"001100010",
  36067=>"110111010",
  36068=>"100000011",
  36069=>"001000000",
  36070=>"000101001",
  36071=>"001110101",
  36072=>"001001010",
  36073=>"111100101",
  36074=>"101100001",
  36075=>"111011101",
  36076=>"111101011",
  36077=>"011010000",
  36078=>"000011010",
  36079=>"000011001",
  36080=>"011001100",
  36081=>"001001000",
  36082=>"010111110",
  36083=>"001011010",
  36084=>"111101010",
  36085=>"000010001",
  36086=>"111001011",
  36087=>"101000111",
  36088=>"100011110",
  36089=>"111000111",
  36090=>"110011011",
  36091=>"110001000",
  36092=>"010000000",
  36093=>"010010001",
  36094=>"101111101",
  36095=>"110010101",
  36096=>"110101000",
  36097=>"110111001",
  36098=>"111101011",
  36099=>"000011100",
  36100=>"011110001",
  36101=>"101001001",
  36102=>"100000001",
  36103=>"101110000",
  36104=>"110011000",
  36105=>"100110000",
  36106=>"100001001",
  36107=>"111101110",
  36108=>"110110010",
  36109=>"100101101",
  36110=>"111000101",
  36111=>"110111000",
  36112=>"101110000",
  36113=>"011000101",
  36114=>"111111110",
  36115=>"110100100",
  36116=>"101010111",
  36117=>"111100001",
  36118=>"100111001",
  36119=>"111010111",
  36120=>"101100111",
  36121=>"111001001",
  36122=>"010001100",
  36123=>"000010111",
  36124=>"011001100",
  36125=>"101001010",
  36126=>"111010011",
  36127=>"111111111",
  36128=>"010111101",
  36129=>"010000101",
  36130=>"110111000",
  36131=>"000100010",
  36132=>"101100001",
  36133=>"000001011",
  36134=>"100100000",
  36135=>"100110001",
  36136=>"101010010",
  36137=>"001110110",
  36138=>"000100110",
  36139=>"001111100",
  36140=>"110111100",
  36141=>"100101011",
  36142=>"111110111",
  36143=>"110001001",
  36144=>"010110010",
  36145=>"110111111",
  36146=>"001000000",
  36147=>"110110111",
  36148=>"010001111",
  36149=>"000001100",
  36150=>"111101001",
  36151=>"010111000",
  36152=>"101001110",
  36153=>"101001001",
  36154=>"001111011",
  36155=>"110100101",
  36156=>"100011101",
  36157=>"001000000",
  36158=>"001100001",
  36159=>"000110000",
  36160=>"110101110",
  36161=>"100011110",
  36162=>"010010010",
  36163=>"100010101",
  36164=>"101100000",
  36165=>"100101001",
  36166=>"100010100",
  36167=>"000000111",
  36168=>"111001001",
  36169=>"110010000",
  36170=>"101001001",
  36171=>"100010101",
  36172=>"110110101",
  36173=>"100010011",
  36174=>"111001111",
  36175=>"100111100",
  36176=>"100111000",
  36177=>"011101110",
  36178=>"110110100",
  36179=>"001101011",
  36180=>"101100101",
  36181=>"110010001",
  36182=>"100010110",
  36183=>"110000101",
  36184=>"000101011",
  36185=>"011010011",
  36186=>"010000111",
  36187=>"000111100",
  36188=>"101011010",
  36189=>"001000011",
  36190=>"111110101",
  36191=>"100011000",
  36192=>"000110011",
  36193=>"100111010",
  36194=>"000011000",
  36195=>"001010010",
  36196=>"010110001",
  36197=>"101011111",
  36198=>"011101000",
  36199=>"011101100",
  36200=>"000100001",
  36201=>"001110011",
  36202=>"110000010",
  36203=>"110011011",
  36204=>"100000101",
  36205=>"000100010",
  36206=>"010011110",
  36207=>"000110001",
  36208=>"001000100",
  36209=>"111011100",
  36210=>"011110111",
  36211=>"010000111",
  36212=>"001100010",
  36213=>"100111101",
  36214=>"100100100",
  36215=>"101100111",
  36216=>"010001000",
  36217=>"001001110",
  36218=>"000001011",
  36219=>"100000110",
  36220=>"001110010",
  36221=>"110111000",
  36222=>"100100101",
  36223=>"010001010",
  36224=>"010011000",
  36225=>"001010000",
  36226=>"111111001",
  36227=>"110000001",
  36228=>"001111111",
  36229=>"000111111",
  36230=>"111100110",
  36231=>"011000101",
  36232=>"010001110",
  36233=>"111000001",
  36234=>"000110011",
  36235=>"011000111",
  36236=>"011100100",
  36237=>"101110001",
  36238=>"111011111",
  36239=>"001010110",
  36240=>"000000001",
  36241=>"010100000",
  36242=>"111100000",
  36243=>"010011100",
  36244=>"100111001",
  36245=>"011010101",
  36246=>"111111101",
  36247=>"001000111",
  36248=>"010100110",
  36249=>"000100111",
  36250=>"000100110",
  36251=>"100000000",
  36252=>"110110010",
  36253=>"001001110",
  36254=>"101011101",
  36255=>"111000000",
  36256=>"111101110",
  36257=>"001110000",
  36258=>"010010011",
  36259=>"000110110",
  36260=>"111101001",
  36261=>"111110000",
  36262=>"101110011",
  36263=>"010000101",
  36264=>"110011111",
  36265=>"011010000",
  36266=>"000001000",
  36267=>"100010111",
  36268=>"000000110",
  36269=>"010000001",
  36270=>"010011001",
  36271=>"011100100",
  36272=>"000010111",
  36273=>"001011000",
  36274=>"001100011",
  36275=>"010000001",
  36276=>"101011010",
  36277=>"110001110",
  36278=>"001011001",
  36279=>"000001100",
  36280=>"111111111",
  36281=>"101011010",
  36282=>"110111011",
  36283=>"010101001",
  36284=>"100100111",
  36285=>"010110101",
  36286=>"011011011",
  36287=>"010011000",
  36288=>"100111000",
  36289=>"001011011",
  36290=>"111111110",
  36291=>"001101100",
  36292=>"001110101",
  36293=>"001101110",
  36294=>"000111001",
  36295=>"000111100",
  36296=>"111000110",
  36297=>"011110111",
  36298=>"000010001",
  36299=>"101011110",
  36300=>"111011101",
  36301=>"000100111",
  36302=>"110000010",
  36303=>"011010010",
  36304=>"111011000",
  36305=>"101000101",
  36306=>"010110011",
  36307=>"011010011",
  36308=>"110001111",
  36309=>"101100010",
  36310=>"010001111",
  36311=>"011110010",
  36312=>"101110001",
  36313=>"100110101",
  36314=>"100100001",
  36315=>"000000000",
  36316=>"111110100",
  36317=>"000100011",
  36318=>"001011000",
  36319=>"010110001",
  36320=>"000101100",
  36321=>"101110101",
  36322=>"100110001",
  36323=>"010001010",
  36324=>"010001000",
  36325=>"111000011",
  36326=>"010001101",
  36327=>"011000100",
  36328=>"010100000",
  36329=>"010000011",
  36330=>"010000110",
  36331=>"001110000",
  36332=>"001100011",
  36333=>"111001101",
  36334=>"110101111",
  36335=>"010100001",
  36336=>"111101100",
  36337=>"111000110",
  36338=>"100000100",
  36339=>"001100000",
  36340=>"111001010",
  36341=>"011000011",
  36342=>"111111100",
  36343=>"110010001",
  36344=>"001110011",
  36345=>"101010111",
  36346=>"101101111",
  36347=>"001001111",
  36348=>"001111110",
  36349=>"000010011",
  36350=>"100000111",
  36351=>"100000100",
  36352=>"011100100",
  36353=>"001001101",
  36354=>"100100101",
  36355=>"000011010",
  36356=>"111101111",
  36357=>"010011011",
  36358=>"100110100",
  36359=>"110101000",
  36360=>"101101100",
  36361=>"001100110",
  36362=>"011101111",
  36363=>"111111100",
  36364=>"110001001",
  36365=>"010100010",
  36366=>"101101100",
  36367=>"010110000",
  36368=>"000110001",
  36369=>"010010011",
  36370=>"001000000",
  36371=>"111010011",
  36372=>"110000011",
  36373=>"000001110",
  36374=>"101011110",
  36375=>"111011010",
  36376=>"000010000",
  36377=>"010100110",
  36378=>"010001100",
  36379=>"110100101",
  36380=>"100101000",
  36381=>"111111000",
  36382=>"011000101",
  36383=>"010111011",
  36384=>"011111011",
  36385=>"001010001",
  36386=>"011011110",
  36387=>"011100110",
  36388=>"110000110",
  36389=>"010000011",
  36390=>"111010001",
  36391=>"000110110",
  36392=>"001010101",
  36393=>"100101010",
  36394=>"111001100",
  36395=>"100010000",
  36396=>"010000101",
  36397=>"000100110",
  36398=>"000100010",
  36399=>"010001100",
  36400=>"001110000",
  36401=>"000101000",
  36402=>"101101111",
  36403=>"100011010",
  36404=>"011101011",
  36405=>"100011011",
  36406=>"111100111",
  36407=>"010000110",
  36408=>"110110110",
  36409=>"101111001",
  36410=>"001011011",
  36411=>"110100010",
  36412=>"110100110",
  36413=>"001001010",
  36414=>"000000100",
  36415=>"011101100",
  36416=>"100110101",
  36417=>"001111100",
  36418=>"010001010",
  36419=>"110001100",
  36420=>"110100010",
  36421=>"010110111",
  36422=>"000100011",
  36423=>"100011110",
  36424=>"001001111",
  36425=>"100010010",
  36426=>"111011101",
  36427=>"000010101",
  36428=>"011011111",
  36429=>"000011001",
  36430=>"111100010",
  36431=>"100111110",
  36432=>"110010001",
  36433=>"001000010",
  36434=>"000000110",
  36435=>"011000100",
  36436=>"111101101",
  36437=>"100101111",
  36438=>"111110100",
  36439=>"110100110",
  36440=>"111101011",
  36441=>"011011101",
  36442=>"000111111",
  36443=>"000101101",
  36444=>"010010100",
  36445=>"110010100",
  36446=>"001010010",
  36447=>"001110000",
  36448=>"100000010",
  36449=>"101011010",
  36450=>"000110110",
  36451=>"100001101",
  36452=>"000101101",
  36453=>"001101100",
  36454=>"011011101",
  36455=>"011000101",
  36456=>"010101010",
  36457=>"111000010",
  36458=>"000000111",
  36459=>"001110010",
  36460=>"110110010",
  36461=>"100000000",
  36462=>"100011110",
  36463=>"001001100",
  36464=>"110110111",
  36465=>"111011010",
  36466=>"011010000",
  36467=>"100001000",
  36468=>"101011100",
  36469=>"111111010",
  36470=>"001101011",
  36471=>"110010000",
  36472=>"100111100",
  36473=>"010110001",
  36474=>"111010110",
  36475=>"110010011",
  36476=>"010001110",
  36477=>"010111000",
  36478=>"000000001",
  36479=>"111010100",
  36480=>"010111011",
  36481=>"111000010",
  36482=>"101010000",
  36483=>"000000100",
  36484=>"001001000",
  36485=>"011101001",
  36486=>"110100010",
  36487=>"011000010",
  36488=>"011011010",
  36489=>"001110010",
  36490=>"110111111",
  36491=>"100001011",
  36492=>"010010110",
  36493=>"010100100",
  36494=>"010000010",
  36495=>"000111011",
  36496=>"101011001",
  36497=>"001110111",
  36498=>"101000000",
  36499=>"010001110",
  36500=>"011000011",
  36501=>"011001010",
  36502=>"000110111",
  36503=>"010101001",
  36504=>"100110001",
  36505=>"011000111",
  36506=>"111001111",
  36507=>"000011111",
  36508=>"101011011",
  36509=>"011110101",
  36510=>"111000100",
  36511=>"011110101",
  36512=>"001101000",
  36513=>"100110110",
  36514=>"000000101",
  36515=>"111101000",
  36516=>"000000101",
  36517=>"001010111",
  36518=>"110000000",
  36519=>"000001010",
  36520=>"100101010",
  36521=>"001110111",
  36522=>"111010110",
  36523=>"101101010",
  36524=>"001011100",
  36525=>"010010111",
  36526=>"001100010",
  36527=>"100100001",
  36528=>"000101111",
  36529=>"000111101",
  36530=>"111001000",
  36531=>"011001001",
  36532=>"001100110",
  36533=>"110001011",
  36534=>"011001101",
  36535=>"000000110",
  36536=>"010001010",
  36537=>"001101111",
  36538=>"001011010",
  36539=>"001001011",
  36540=>"001001000",
  36541=>"110010011",
  36542=>"001000011",
  36543=>"100101110",
  36544=>"100110111",
  36545=>"011011100",
  36546=>"011010110",
  36547=>"000110000",
  36548=>"001011000",
  36549=>"001000001",
  36550=>"000110100",
  36551=>"011000001",
  36552=>"110000001",
  36553=>"100110101",
  36554=>"000100110",
  36555=>"110001000",
  36556=>"100001111",
  36557=>"101100010",
  36558=>"000011110",
  36559=>"101110110",
  36560=>"001110010",
  36561=>"110001000",
  36562=>"001101001",
  36563=>"010100100",
  36564=>"111011011",
  36565=>"010111111",
  36566=>"000010000",
  36567=>"110110101",
  36568=>"010100010",
  36569=>"000010010",
  36570=>"010101000",
  36571=>"000110010",
  36572=>"010110011",
  36573=>"010100011",
  36574=>"110111010",
  36575=>"110011000",
  36576=>"001000100",
  36577=>"010000000",
  36578=>"101001000",
  36579=>"011100000",
  36580=>"101000111",
  36581=>"111110100",
  36582=>"011100010",
  36583=>"001111100",
  36584=>"010110000",
  36585=>"100111000",
  36586=>"001111011",
  36587=>"001101100",
  36588=>"011010111",
  36589=>"001010001",
  36590=>"111000001",
  36591=>"100001000",
  36592=>"110010101",
  36593=>"101100111",
  36594=>"111011001",
  36595=>"000011010",
  36596=>"111100001",
  36597=>"110010111",
  36598=>"111110110",
  36599=>"001110101",
  36600=>"010011100",
  36601=>"010011000",
  36602=>"010001000",
  36603=>"101001110",
  36604=>"110100011",
  36605=>"010000111",
  36606=>"011101010",
  36607=>"011101101",
  36608=>"001001011",
  36609=>"110010010",
  36610=>"000101001",
  36611=>"000110111",
  36612=>"001000101",
  36613=>"100000110",
  36614=>"101010000",
  36615=>"101110010",
  36616=>"001000011",
  36617=>"101100111",
  36618=>"000001010",
  36619=>"101010100",
  36620=>"010111111",
  36621=>"110100100",
  36622=>"100101001",
  36623=>"111000011",
  36624=>"001001001",
  36625=>"000101011",
  36626=>"011101101",
  36627=>"001100110",
  36628=>"111100100",
  36629=>"010010010",
  36630=>"100100001",
  36631=>"100010101",
  36632=>"011110100",
  36633=>"000101110",
  36634=>"111101001",
  36635=>"110001001",
  36636=>"111010110",
  36637=>"010111011",
  36638=>"000110101",
  36639=>"101001011",
  36640=>"000001101",
  36641=>"111111000",
  36642=>"101011010",
  36643=>"111100111",
  36644=>"100101001",
  36645=>"000101010",
  36646=>"011011101",
  36647=>"010001100",
  36648=>"000001100",
  36649=>"001110101",
  36650=>"011011110",
  36651=>"000110011",
  36652=>"001010111",
  36653=>"001101100",
  36654=>"011000011",
  36655=>"101011011",
  36656=>"001111100",
  36657=>"000100111",
  36658=>"000010011",
  36659=>"101110101",
  36660=>"110100011",
  36661=>"001011110",
  36662=>"011000001",
  36663=>"111001100",
  36664=>"000100111",
  36665=>"011111101",
  36666=>"100011010",
  36667=>"000100100",
  36668=>"011001001",
  36669=>"111111100",
  36670=>"110100111",
  36671=>"010100100",
  36672=>"100100001",
  36673=>"111000000",
  36674=>"101100111",
  36675=>"011010001",
  36676=>"101001000",
  36677=>"110010100",
  36678=>"100001000",
  36679=>"111000010",
  36680=>"111011010",
  36681=>"100000010",
  36682=>"011110111",
  36683=>"100000100",
  36684=>"101010011",
  36685=>"101000100",
  36686=>"011010000",
  36687=>"000011111",
  36688=>"001011111",
  36689=>"001011011",
  36690=>"001001101",
  36691=>"001010100",
  36692=>"101000100",
  36693=>"110010001",
  36694=>"001111100",
  36695=>"101011000",
  36696=>"010101111",
  36697=>"011110011",
  36698=>"000100011",
  36699=>"001001000",
  36700=>"111101011",
  36701=>"000000010",
  36702=>"101011001",
  36703=>"000101101",
  36704=>"001101000",
  36705=>"010010111",
  36706=>"101010000",
  36707=>"011010110",
  36708=>"101111110",
  36709=>"010110000",
  36710=>"110111110",
  36711=>"110000100",
  36712=>"010001001",
  36713=>"010001000",
  36714=>"011100111",
  36715=>"101111111",
  36716=>"101010101",
  36717=>"011011010",
  36718=>"011111111",
  36719=>"110101010",
  36720=>"110100100",
  36721=>"010111011",
  36722=>"010001010",
  36723=>"001000011",
  36724=>"011101110",
  36725=>"000001000",
  36726=>"010010000",
  36727=>"111010010",
  36728=>"111000100",
  36729=>"111101100",
  36730=>"000111101",
  36731=>"101100111",
  36732=>"000000010",
  36733=>"011111101",
  36734=>"100010111",
  36735=>"010011101",
  36736=>"001001111",
  36737=>"100000010",
  36738=>"010100010",
  36739=>"000101111",
  36740=>"101000011",
  36741=>"110010000",
  36742=>"011011110",
  36743=>"100101010",
  36744=>"000101000",
  36745=>"001010000",
  36746=>"001010001",
  36747=>"111111111",
  36748=>"001110101",
  36749=>"000000010",
  36750=>"100001110",
  36751=>"101000000",
  36752=>"001000010",
  36753=>"100100010",
  36754=>"001100000",
  36755=>"011101000",
  36756=>"010011001",
  36757=>"110110110",
  36758=>"101000011",
  36759=>"001101110",
  36760=>"010001101",
  36761=>"110110101",
  36762=>"010110100",
  36763=>"001111100",
  36764=>"110000100",
  36765=>"000110001",
  36766=>"010001001",
  36767=>"111111000",
  36768=>"001001100",
  36769=>"110110001",
  36770=>"001111110",
  36771=>"010000001",
  36772=>"000010010",
  36773=>"000001100",
  36774=>"110110101",
  36775=>"011001011",
  36776=>"010001101",
  36777=>"011100010",
  36778=>"010100000",
  36779=>"001010000",
  36780=>"001000111",
  36781=>"011110011",
  36782=>"011010010",
  36783=>"111001110",
  36784=>"101010100",
  36785=>"001000010",
  36786=>"101100111",
  36787=>"101010111",
  36788=>"011010101",
  36789=>"010001001",
  36790=>"110001101",
  36791=>"101010010",
  36792=>"010111000",
  36793=>"100111000",
  36794=>"010101110",
  36795=>"111011110",
  36796=>"111111101",
  36797=>"101000000",
  36798=>"011011001",
  36799=>"110011101",
  36800=>"101110111",
  36801=>"011011001",
  36802=>"101101110",
  36803=>"100000100",
  36804=>"100011000",
  36805=>"100101111",
  36806=>"110101101",
  36807=>"111100100",
  36808=>"010111111",
  36809=>"000001011",
  36810=>"110101110",
  36811=>"111010001",
  36812=>"000110011",
  36813=>"111110100",
  36814=>"100101101",
  36815=>"100101101",
  36816=>"000101000",
  36817=>"101010011",
  36818=>"000000100",
  36819=>"101101000",
  36820=>"010101001",
  36821=>"110001000",
  36822=>"001111010",
  36823=>"010011101",
  36824=>"010000101",
  36825=>"110011110",
  36826=>"010000110",
  36827=>"011001111",
  36828=>"110000010",
  36829=>"001111101",
  36830=>"010001101",
  36831=>"010100111",
  36832=>"111101101",
  36833=>"001000001",
  36834=>"001010111",
  36835=>"100101110",
  36836=>"000001100",
  36837=>"010101101",
  36838=>"110101101",
  36839=>"110001110",
  36840=>"001011110",
  36841=>"110100100",
  36842=>"010110011",
  36843=>"110001011",
  36844=>"100001110",
  36845=>"000100011",
  36846=>"001001001",
  36847=>"100001110",
  36848=>"111111000",
  36849=>"010000000",
  36850=>"111110101",
  36851=>"010101101",
  36852=>"101110101",
  36853=>"101000101",
  36854=>"101011010",
  36855=>"001100001",
  36856=>"101000000",
  36857=>"011011001",
  36858=>"001010111",
  36859=>"101101011",
  36860=>"011101000",
  36861=>"010011101",
  36862=>"010111000",
  36863=>"011101111",
  36864=>"110100001",
  36865=>"001001100",
  36866=>"111110100",
  36867=>"000110010",
  36868=>"011000001",
  36869=>"111000000",
  36870=>"010011110",
  36871=>"111001101",
  36872=>"101101011",
  36873=>"010001101",
  36874=>"101111111",
  36875=>"010011100",
  36876=>"001011100",
  36877=>"101111011",
  36878=>"011010011",
  36879=>"011001111",
  36880=>"101111101",
  36881=>"111011111",
  36882=>"011000100",
  36883=>"001010111",
  36884=>"101110011",
  36885=>"100111011",
  36886=>"110100100",
  36887=>"101100010",
  36888=>"111110100",
  36889=>"010101100",
  36890=>"010011000",
  36891=>"010111011",
  36892=>"100101100",
  36893=>"100101001",
  36894=>"001011100",
  36895=>"000000011",
  36896=>"010000101",
  36897=>"100011000",
  36898=>"111010000",
  36899=>"101000111",
  36900=>"110011100",
  36901=>"000111011",
  36902=>"001010001",
  36903=>"101111101",
  36904=>"011011001",
  36905=>"001111000",
  36906=>"001001111",
  36907=>"000011011",
  36908=>"001100011",
  36909=>"001110010",
  36910=>"010101111",
  36911=>"101001100",
  36912=>"010111100",
  36913=>"010010110",
  36914=>"010001110",
  36915=>"111000000",
  36916=>"101000000",
  36917=>"111010001",
  36918=>"010011110",
  36919=>"000111001",
  36920=>"010000000",
  36921=>"000010100",
  36922=>"111100010",
  36923=>"000111000",
  36924=>"000010111",
  36925=>"001011000",
  36926=>"000010111",
  36927=>"010000110",
  36928=>"111010001",
  36929=>"000011011",
  36930=>"101111101",
  36931=>"001010010",
  36932=>"001001110",
  36933=>"000011111",
  36934=>"001001111",
  36935=>"001111000",
  36936=>"011101001",
  36937=>"110111010",
  36938=>"110100010",
  36939=>"100001101",
  36940=>"001001111",
  36941=>"101110100",
  36942=>"010101101",
  36943=>"101001010",
  36944=>"001100000",
  36945=>"110001110",
  36946=>"001110100",
  36947=>"001110101",
  36948=>"111111000",
  36949=>"001100000",
  36950=>"011100111",
  36951=>"011100001",
  36952=>"010000010",
  36953=>"100010110",
  36954=>"100101100",
  36955=>"111100111",
  36956=>"010111111",
  36957=>"001101101",
  36958=>"001101011",
  36959=>"010000011",
  36960=>"101110010",
  36961=>"111001001",
  36962=>"011011101",
  36963=>"100101100",
  36964=>"100010100",
  36965=>"010010110",
  36966=>"000100010",
  36967=>"101001000",
  36968=>"111100011",
  36969=>"101111000",
  36970=>"001100010",
  36971=>"011001100",
  36972=>"011101010",
  36973=>"001100001",
  36974=>"111000111",
  36975=>"010111111",
  36976=>"001101100",
  36977=>"000001100",
  36978=>"010000010",
  36979=>"001010011",
  36980=>"001010101",
  36981=>"001100000",
  36982=>"000001010",
  36983=>"011110100",
  36984=>"110000011",
  36985=>"011100100",
  36986=>"001001000",
  36987=>"010001111",
  36988=>"111001011",
  36989=>"111110000",
  36990=>"011000000",
  36991=>"011011001",
  36992=>"111000100",
  36993=>"010010000",
  36994=>"111101100",
  36995=>"001000101",
  36996=>"101101010",
  36997=>"101100110",
  36998=>"011100111",
  36999=>"101011010",
  37000=>"100010110",
  37001=>"110010100",
  37002=>"001001111",
  37003=>"100111001",
  37004=>"001110001",
  37005=>"010110001",
  37006=>"000111011",
  37007=>"101111001",
  37008=>"011011011",
  37009=>"111110011",
  37010=>"101011010",
  37011=>"011000100",
  37012=>"101101101",
  37013=>"100100110",
  37014=>"011111011",
  37015=>"111110101",
  37016=>"011111101",
  37017=>"110000110",
  37018=>"000100101",
  37019=>"111111000",
  37020=>"010010110",
  37021=>"110110000",
  37022=>"011101110",
  37023=>"100100000",
  37024=>"100111111",
  37025=>"111000110",
  37026=>"010000110",
  37027=>"001011101",
  37028=>"000010111",
  37029=>"100011111",
  37030=>"001011110",
  37031=>"000111010",
  37032=>"111101010",
  37033=>"100101010",
  37034=>"000001000",
  37035=>"100100001",
  37036=>"000000111",
  37037=>"000100111",
  37038=>"010101000",
  37039=>"111011100",
  37040=>"011100010",
  37041=>"000010111",
  37042=>"101010111",
  37043=>"100001001",
  37044=>"111001011",
  37045=>"010011110",
  37046=>"001010001",
  37047=>"110101011",
  37048=>"111000101",
  37049=>"001000001",
  37050=>"000000111",
  37051=>"110010111",
  37052=>"111100010",
  37053=>"011011101",
  37054=>"111100001",
  37055=>"101011011",
  37056=>"001111010",
  37057=>"000001100",
  37058=>"011011111",
  37059=>"100100011",
  37060=>"101100101",
  37061=>"100101011",
  37062=>"111101111",
  37063=>"101111100",
  37064=>"100111110",
  37065=>"101000110",
  37066=>"010100001",
  37067=>"010010100",
  37068=>"000111011",
  37069=>"001110100",
  37070=>"001001010",
  37071=>"111101011",
  37072=>"110101000",
  37073=>"101001000",
  37074=>"110000101",
  37075=>"010000101",
  37076=>"010110001",
  37077=>"000110101",
  37078=>"010101010",
  37079=>"010111001",
  37080=>"001100000",
  37081=>"010100011",
  37082=>"101010010",
  37083=>"001101100",
  37084=>"100111110",
  37085=>"010110011",
  37086=>"000000001",
  37087=>"111011010",
  37088=>"001001000",
  37089=>"011000100",
  37090=>"011100000",
  37091=>"110001000",
  37092=>"111001011",
  37093=>"010111010",
  37094=>"110000010",
  37095=>"111111110",
  37096=>"001011001",
  37097=>"101110011",
  37098=>"101010111",
  37099=>"101100101",
  37100=>"000100100",
  37101=>"000100001",
  37102=>"101111001",
  37103=>"000000000",
  37104=>"011111110",
  37105=>"000000110",
  37106=>"011000001",
  37107=>"100011111",
  37108=>"110011011",
  37109=>"110000001",
  37110=>"011000010",
  37111=>"010110010",
  37112=>"100011101",
  37113=>"000100101",
  37114=>"011110100",
  37115=>"011001001",
  37116=>"110001101",
  37117=>"010101010",
  37118=>"101111101",
  37119=>"111101111",
  37120=>"011011011",
  37121=>"100011010",
  37122=>"110111010",
  37123=>"011101000",
  37124=>"111111111",
  37125=>"010010001",
  37126=>"011010110",
  37127=>"000001000",
  37128=>"001001001",
  37129=>"111111011",
  37130=>"110101011",
  37131=>"000000001",
  37132=>"111000000",
  37133=>"010100001",
  37134=>"110011000",
  37135=>"001011111",
  37136=>"000000111",
  37137=>"111011011",
  37138=>"000011110",
  37139=>"011010000",
  37140=>"010000101",
  37141=>"010011000",
  37142=>"111100100",
  37143=>"010100101",
  37144=>"100111001",
  37145=>"101101101",
  37146=>"000001111",
  37147=>"100000010",
  37148=>"000110011",
  37149=>"110000000",
  37150=>"011010100",
  37151=>"100001000",
  37152=>"101100100",
  37153=>"111001000",
  37154=>"010111010",
  37155=>"000101101",
  37156=>"001100000",
  37157=>"101101100",
  37158=>"101011100",
  37159=>"100000011",
  37160=>"001101100",
  37161=>"001011100",
  37162=>"001101010",
  37163=>"110000001",
  37164=>"110001000",
  37165=>"110101000",
  37166=>"001101110",
  37167=>"000011101",
  37168=>"001100111",
  37169=>"101100111",
  37170=>"110111100",
  37171=>"011111000",
  37172=>"011101010",
  37173=>"100011111",
  37174=>"000101000",
  37175=>"100101111",
  37176=>"001100111",
  37177=>"101110101",
  37178=>"010110110",
  37179=>"000011111",
  37180=>"101011000",
  37181=>"001011000",
  37182=>"011000000",
  37183=>"111101011",
  37184=>"000111110",
  37185=>"010110101",
  37186=>"111110111",
  37187=>"011001111",
  37188=>"010100110",
  37189=>"101000010",
  37190=>"000010101",
  37191=>"101010101",
  37192=>"000101001",
  37193=>"101100000",
  37194=>"110011100",
  37195=>"001101101",
  37196=>"110101001",
  37197=>"001101001",
  37198=>"101001110",
  37199=>"110101111",
  37200=>"110000011",
  37201=>"011111110",
  37202=>"111011001",
  37203=>"000100001",
  37204=>"000000110",
  37205=>"101001110",
  37206=>"000000100",
  37207=>"000110011",
  37208=>"100110111",
  37209=>"010000101",
  37210=>"100101100",
  37211=>"111000100",
  37212=>"111100101",
  37213=>"110110011",
  37214=>"101000101",
  37215=>"000001010",
  37216=>"110001010",
  37217=>"000101101",
  37218=>"001101011",
  37219=>"011001011",
  37220=>"011111010",
  37221=>"110110010",
  37222=>"110010011",
  37223=>"001000101",
  37224=>"100101001",
  37225=>"111111110",
  37226=>"101000001",
  37227=>"101010100",
  37228=>"101010111",
  37229=>"100101111",
  37230=>"010100110",
  37231=>"110001001",
  37232=>"000000000",
  37233=>"101100111",
  37234=>"101000000",
  37235=>"011000100",
  37236=>"110011001",
  37237=>"110011010",
  37238=>"001110100",
  37239=>"010011101",
  37240=>"001011100",
  37241=>"000011110",
  37242=>"010000110",
  37243=>"111001100",
  37244=>"010101111",
  37245=>"010011010",
  37246=>"100000100",
  37247=>"011001110",
  37248=>"111111000",
  37249=>"110011001",
  37250=>"010110100",
  37251=>"010000001",
  37252=>"100000111",
  37253=>"011001010",
  37254=>"111110011",
  37255=>"010011011",
  37256=>"000000010",
  37257=>"100010110",
  37258=>"101110111",
  37259=>"011000101",
  37260=>"111010110",
  37261=>"101110001",
  37262=>"101100010",
  37263=>"101000011",
  37264=>"000000000",
  37265=>"000000001",
  37266=>"110001011",
  37267=>"100111010",
  37268=>"000011010",
  37269=>"001110001",
  37270=>"101111001",
  37271=>"101101000",
  37272=>"001111001",
  37273=>"011111101",
  37274=>"100001101",
  37275=>"001111100",
  37276=>"101001000",
  37277=>"001111000",
  37278=>"111100101",
  37279=>"111111101",
  37280=>"001001101",
  37281=>"111001101",
  37282=>"110010011",
  37283=>"000100010",
  37284=>"111000111",
  37285=>"001000110",
  37286=>"101101110",
  37287=>"001011110",
  37288=>"011101111",
  37289=>"011001000",
  37290=>"011100001",
  37291=>"000001100",
  37292=>"011010101",
  37293=>"110110000",
  37294=>"001010010",
  37295=>"111100110",
  37296=>"011000001",
  37297=>"010101101",
  37298=>"001111001",
  37299=>"011100001",
  37300=>"011011011",
  37301=>"011111100",
  37302=>"001011001",
  37303=>"111100000",
  37304=>"101111010",
  37305=>"100011110",
  37306=>"000101000",
  37307=>"110111101",
  37308=>"001001100",
  37309=>"010100010",
  37310=>"001001000",
  37311=>"000011111",
  37312=>"110000000",
  37313=>"000000001",
  37314=>"010000101",
  37315=>"101111111",
  37316=>"011000010",
  37317=>"101101110",
  37318=>"010001101",
  37319=>"000000000",
  37320=>"010100000",
  37321=>"010001101",
  37322=>"000010011",
  37323=>"101001111",
  37324=>"101001100",
  37325=>"010001000",
  37326=>"111011001",
  37327=>"101110000",
  37328=>"011011111",
  37329=>"000110000",
  37330=>"011001111",
  37331=>"101001000",
  37332=>"110001111",
  37333=>"000001100",
  37334=>"001100000",
  37335=>"011100010",
  37336=>"000101111",
  37337=>"100111101",
  37338=>"100100000",
  37339=>"101100000",
  37340=>"100101110",
  37341=>"001011101",
  37342=>"110001100",
  37343=>"001100110",
  37344=>"010100110",
  37345=>"001101100",
  37346=>"101101010",
  37347=>"011101100",
  37348=>"011000010",
  37349=>"101011001",
  37350=>"001111101",
  37351=>"010011001",
  37352=>"001000001",
  37353=>"110101110",
  37354=>"001100010",
  37355=>"100001010",
  37356=>"010110100",
  37357=>"101100001",
  37358=>"000001010",
  37359=>"111001000",
  37360=>"000100001",
  37361=>"110111101",
  37362=>"101100101",
  37363=>"000001001",
  37364=>"101110101",
  37365=>"000111001",
  37366=>"000011011",
  37367=>"110000010",
  37368=>"000000000",
  37369=>"011101100",
  37370=>"011001010",
  37371=>"111000000",
  37372=>"101101010",
  37373=>"111000001",
  37374=>"110110110",
  37375=>"111000010",
  37376=>"101011001",
  37377=>"101011010",
  37378=>"011001000",
  37379=>"000000000",
  37380=>"100010010",
  37381=>"100011111",
  37382=>"100101001",
  37383=>"010011010",
  37384=>"110100100",
  37385=>"000000111",
  37386=>"110001110",
  37387=>"010000111",
  37388=>"000101011",
  37389=>"101001011",
  37390=>"100010001",
  37391=>"100111001",
  37392=>"110101111",
  37393=>"111111101",
  37394=>"101100011",
  37395=>"011111001",
  37396=>"000000010",
  37397=>"100000010",
  37398=>"010111111",
  37399=>"100000101",
  37400=>"111011011",
  37401=>"110100010",
  37402=>"110100101",
  37403=>"011111110",
  37404=>"010100000",
  37405=>"110011001",
  37406=>"010110110",
  37407=>"001101100",
  37408=>"101000000",
  37409=>"100110001",
  37410=>"000101111",
  37411=>"001100101",
  37412=>"111110001",
  37413=>"011001111",
  37414=>"100111100",
  37415=>"111111001",
  37416=>"001110111",
  37417=>"111001111",
  37418=>"101100111",
  37419=>"100111101",
  37420=>"000110101",
  37421=>"010100101",
  37422=>"011101000",
  37423=>"010110010",
  37424=>"100110101",
  37425=>"110011110",
  37426=>"110011011",
  37427=>"110101000",
  37428=>"011000011",
  37429=>"100000000",
  37430=>"101100110",
  37431=>"000110110",
  37432=>"111110010",
  37433=>"001011100",
  37434=>"001110001",
  37435=>"001111111",
  37436=>"111101101",
  37437=>"100110110",
  37438=>"100100010",
  37439=>"000000000",
  37440=>"111001001",
  37441=>"111111011",
  37442=>"001101110",
  37443=>"011010101",
  37444=>"001101101",
  37445=>"110010110",
  37446=>"100100111",
  37447=>"101010111",
  37448=>"001000000",
  37449=>"101000001",
  37450=>"011011111",
  37451=>"010111001",
  37452=>"100011111",
  37453=>"000001000",
  37454=>"000100100",
  37455=>"101001101",
  37456=>"001000011",
  37457=>"010111110",
  37458=>"000001101",
  37459=>"001001010",
  37460=>"001011001",
  37461=>"000011111",
  37462=>"000100010",
  37463=>"001010001",
  37464=>"000011001",
  37465=>"011000101",
  37466=>"000011000",
  37467=>"001010100",
  37468=>"101010101",
  37469=>"001000000",
  37470=>"101010000",
  37471=>"110001101",
  37472=>"001101111",
  37473=>"011110000",
  37474=>"101010111",
  37475=>"110011010",
  37476=>"000010001",
  37477=>"111110100",
  37478=>"000111001",
  37479=>"000011011",
  37480=>"000010110",
  37481=>"000001001",
  37482=>"011110110",
  37483=>"100010111",
  37484=>"110010101",
  37485=>"001101011",
  37486=>"111100111",
  37487=>"100001000",
  37488=>"101010000",
  37489=>"000001011",
  37490=>"010101011",
  37491=>"001100011",
  37492=>"010101110",
  37493=>"100101001",
  37494=>"101010001",
  37495=>"010010000",
  37496=>"110100101",
  37497=>"001000011",
  37498=>"011100000",
  37499=>"011100101",
  37500=>"010101101",
  37501=>"100110110",
  37502=>"110000010",
  37503=>"111111111",
  37504=>"001110001",
  37505=>"011000110",
  37506=>"110101001",
  37507=>"000001111",
  37508=>"101100001",
  37509=>"000101110",
  37510=>"100000111",
  37511=>"001101010",
  37512=>"111000111",
  37513=>"011111000",
  37514=>"011000110",
  37515=>"100110111",
  37516=>"000110000",
  37517=>"010010000",
  37518=>"010110011",
  37519=>"001111000",
  37520=>"011110111",
  37521=>"001110110",
  37522=>"111100101",
  37523=>"010101111",
  37524=>"000101010",
  37525=>"111111001",
  37526=>"111000110",
  37527=>"011110111",
  37528=>"011100011",
  37529=>"100011001",
  37530=>"011000010",
  37531=>"101010001",
  37532=>"011010000",
  37533=>"100111011",
  37534=>"101000100",
  37535=>"011011010",
  37536=>"000000111",
  37537=>"011000100",
  37538=>"001000011",
  37539=>"111101001",
  37540=>"111100001",
  37541=>"000100011",
  37542=>"001000000",
  37543=>"001111101",
  37544=>"010110001",
  37545=>"000010100",
  37546=>"000101101",
  37547=>"001000000",
  37548=>"101010010",
  37549=>"010011100",
  37550=>"110001001",
  37551=>"110100000",
  37552=>"001001110",
  37553=>"001111001",
  37554=>"100111101",
  37555=>"010000111",
  37556=>"111100101",
  37557=>"001100111",
  37558=>"100101100",
  37559=>"001111110",
  37560=>"100101011",
  37561=>"010001010",
  37562=>"010011011",
  37563=>"000011001",
  37564=>"011100000",
  37565=>"111010001",
  37566=>"001001110",
  37567=>"001100101",
  37568=>"111000100",
  37569=>"101110011",
  37570=>"101011110",
  37571=>"010110000",
  37572=>"110010111",
  37573=>"111101000",
  37574=>"111011110",
  37575=>"100000100",
  37576=>"101110001",
  37577=>"000000000",
  37578=>"000110001",
  37579=>"110110001",
  37580=>"110011001",
  37581=>"100010011",
  37582=>"010011011",
  37583=>"000011010",
  37584=>"111111110",
  37585=>"111101101",
  37586=>"110010011",
  37587=>"001111010",
  37588=>"100010011",
  37589=>"000101110",
  37590=>"010110110",
  37591=>"000001111",
  37592=>"110011000",
  37593=>"000001001",
  37594=>"111101011",
  37595=>"100001110",
  37596=>"101101100",
  37597=>"111001011",
  37598=>"100111100",
  37599=>"001111001",
  37600=>"000100011",
  37601=>"101011101",
  37602=>"100110101",
  37603=>"010001010",
  37604=>"000010101",
  37605=>"000010011",
  37606=>"000001100",
  37607=>"110100010",
  37608=>"001001001",
  37609=>"111101110",
  37610=>"101101000",
  37611=>"001000001",
  37612=>"010011100",
  37613=>"110001101",
  37614=>"101010100",
  37615=>"001111100",
  37616=>"110010111",
  37617=>"111000000",
  37618=>"001000000",
  37619=>"001010011",
  37620=>"110011000",
  37621=>"100101110",
  37622=>"000100000",
  37623=>"100011101",
  37624=>"011101000",
  37625=>"110000010",
  37626=>"110100010",
  37627=>"100011100",
  37628=>"100100100",
  37629=>"011101101",
  37630=>"100111000",
  37631=>"001010010",
  37632=>"111110010",
  37633=>"001001000",
  37634=>"000011010",
  37635=>"010001001",
  37636=>"100010110",
  37637=>"001110001",
  37638=>"000010101",
  37639=>"101111010",
  37640=>"010001000",
  37641=>"010111000",
  37642=>"110001110",
  37643=>"010001010",
  37644=>"110011110",
  37645=>"111110101",
  37646=>"000100110",
  37647=>"100001001",
  37648=>"011101010",
  37649=>"110101011",
  37650=>"110110010",
  37651=>"101100101",
  37652=>"011001101",
  37653=>"001011111",
  37654=>"110010111",
  37655=>"000001111",
  37656=>"111010010",
  37657=>"101001001",
  37658=>"000111001",
  37659=>"100101110",
  37660=>"110111010",
  37661=>"001000111",
  37662=>"010010101",
  37663=>"010100100",
  37664=>"011000100",
  37665=>"110110101",
  37666=>"100111010",
  37667=>"100000010",
  37668=>"110111011",
  37669=>"000000101",
  37670=>"101111001",
  37671=>"011000101",
  37672=>"100011010",
  37673=>"111111110",
  37674=>"010001110",
  37675=>"100110111",
  37676=>"101010110",
  37677=>"001111110",
  37678=>"101101011",
  37679=>"010000010",
  37680=>"001100110",
  37681=>"011000001",
  37682=>"000010100",
  37683=>"000111100",
  37684=>"110100110",
  37685=>"001101011",
  37686=>"011100010",
  37687=>"101001111",
  37688=>"001110110",
  37689=>"010000010",
  37690=>"001100000",
  37691=>"110101001",
  37692=>"100100011",
  37693=>"010101111",
  37694=>"111001000",
  37695=>"101101100",
  37696=>"001111011",
  37697=>"100011010",
  37698=>"100101110",
  37699=>"110011111",
  37700=>"010111100",
  37701=>"100000101",
  37702=>"010101001",
  37703=>"101101000",
  37704=>"101001100",
  37705=>"010111111",
  37706=>"110110101",
  37707=>"010100000",
  37708=>"011010110",
  37709=>"001100101",
  37710=>"000011000",
  37711=>"111011111",
  37712=>"100100101",
  37713=>"101100101",
  37714=>"010001000",
  37715=>"100011110",
  37716=>"101111100",
  37717=>"101110000",
  37718=>"100000111",
  37719=>"010011010",
  37720=>"000000000",
  37721=>"000001010",
  37722=>"001010100",
  37723=>"100000011",
  37724=>"111101000",
  37725=>"101100111",
  37726=>"101010001",
  37727=>"000001111",
  37728=>"111011010",
  37729=>"011010001",
  37730=>"000111101",
  37731=>"110111010",
  37732=>"011101001",
  37733=>"101100100",
  37734=>"000100111",
  37735=>"111000010",
  37736=>"111101110",
  37737=>"100111001",
  37738=>"000000000",
  37739=>"110011111",
  37740=>"000001101",
  37741=>"001100000",
  37742=>"001100100",
  37743=>"011110000",
  37744=>"010110110",
  37745=>"101011100",
  37746=>"010001001",
  37747=>"001011100",
  37748=>"011000001",
  37749=>"000000000",
  37750=>"010101000",
  37751=>"000100011",
  37752=>"111110110",
  37753=>"100000100",
  37754=>"011111000",
  37755=>"111111010",
  37756=>"000000101",
  37757=>"110111001",
  37758=>"010000011",
  37759=>"110000110",
  37760=>"101110110",
  37761=>"111001000",
  37762=>"001011001",
  37763=>"000000110",
  37764=>"011001001",
  37765=>"110110111",
  37766=>"101011010",
  37767=>"010111010",
  37768=>"000010011",
  37769=>"100101111",
  37770=>"011010001",
  37771=>"011001101",
  37772=>"101110010",
  37773=>"100001110",
  37774=>"111111001",
  37775=>"011010101",
  37776=>"001101000",
  37777=>"111001010",
  37778=>"101110010",
  37779=>"110111111",
  37780=>"011010010",
  37781=>"000001100",
  37782=>"011010111",
  37783=>"010000111",
  37784=>"111000000",
  37785=>"010001001",
  37786=>"110000100",
  37787=>"101001001",
  37788=>"010011100",
  37789=>"100000001",
  37790=>"011001011",
  37791=>"000000011",
  37792=>"000011001",
  37793=>"110010111",
  37794=>"101101011",
  37795=>"001000011",
  37796=>"100110101",
  37797=>"100110011",
  37798=>"111100000",
  37799=>"011011001",
  37800=>"011111101",
  37801=>"101001011",
  37802=>"111011111",
  37803=>"001001011",
  37804=>"111100000",
  37805=>"010110111",
  37806=>"100111101",
  37807=>"001000010",
  37808=>"010101101",
  37809=>"111111101",
  37810=>"011001001",
  37811=>"101010101",
  37812=>"011010011",
  37813=>"110011100",
  37814=>"110001000",
  37815=>"011000101",
  37816=>"001001000",
  37817=>"010001111",
  37818=>"010001101",
  37819=>"101101100",
  37820=>"010010101",
  37821=>"101010010",
  37822=>"101111000",
  37823=>"001001111",
  37824=>"111001000",
  37825=>"100001111",
  37826=>"100100010",
  37827=>"100000100",
  37828=>"100010110",
  37829=>"111101010",
  37830=>"001110000",
  37831=>"010111110",
  37832=>"100010111",
  37833=>"110001111",
  37834=>"001001101",
  37835=>"010010110",
  37836=>"111111011",
  37837=>"100100110",
  37838=>"010100100",
  37839=>"101001110",
  37840=>"110011100",
  37841=>"110101010",
  37842=>"011011011",
  37843=>"010100111",
  37844=>"010100100",
  37845=>"100001101",
  37846=>"010010001",
  37847=>"010001111",
  37848=>"101000000",
  37849=>"011100000",
  37850=>"010000010",
  37851=>"011000000",
  37852=>"011001000",
  37853=>"101110011",
  37854=>"011110111",
  37855=>"000100111",
  37856=>"111101001",
  37857=>"000001100",
  37858=>"110110011",
  37859=>"000010100",
  37860=>"010111010",
  37861=>"010000101",
  37862=>"000011010",
  37863=>"001100000",
  37864=>"101101010",
  37865=>"010100100",
  37866=>"001110111",
  37867=>"110111111",
  37868=>"001010111",
  37869=>"111100100",
  37870=>"111001000",
  37871=>"110110000",
  37872=>"000000111",
  37873=>"011000010",
  37874=>"101000000",
  37875=>"000101101",
  37876=>"011110101",
  37877=>"001111110",
  37878=>"110101110",
  37879=>"011011111",
  37880=>"111101011",
  37881=>"001011011",
  37882=>"100011010",
  37883=>"110010100",
  37884=>"110001000",
  37885=>"110111100",
  37886=>"001110111",
  37887=>"010011001",
  37888=>"100000001",
  37889=>"110010000",
  37890=>"000001010",
  37891=>"011010010",
  37892=>"101101111",
  37893=>"010010011",
  37894=>"011001001",
  37895=>"111101111",
  37896=>"010111110",
  37897=>"010011000",
  37898=>"010001100",
  37899=>"111111110",
  37900=>"101011011",
  37901=>"001011011",
  37902=>"001000011",
  37903=>"100000100",
  37904=>"111010011",
  37905=>"101000011",
  37906=>"010011110",
  37907=>"010101011",
  37908=>"000000011",
  37909=>"111001011",
  37910=>"100010111",
  37911=>"111001010",
  37912=>"001111010",
  37913=>"011110111",
  37914=>"111101101",
  37915=>"111101000",
  37916=>"000010001",
  37917=>"011101001",
  37918=>"011000111",
  37919=>"000000011",
  37920=>"010000011",
  37921=>"110000101",
  37922=>"100011111",
  37923=>"011001101",
  37924=>"110000101",
  37925=>"001101010",
  37926=>"100111111",
  37927=>"000111001",
  37928=>"110010100",
  37929=>"000000010",
  37930=>"001110011",
  37931=>"100001001",
  37932=>"100001101",
  37933=>"101000001",
  37934=>"110001111",
  37935=>"000111101",
  37936=>"011111000",
  37937=>"111100100",
  37938=>"111110110",
  37939=>"110001111",
  37940=>"011010001",
  37941=>"001010000",
  37942=>"000010010",
  37943=>"011001110",
  37944=>"011000011",
  37945=>"110001111",
  37946=>"111001101",
  37947=>"101011011",
  37948=>"000011100",
  37949=>"001001101",
  37950=>"000110100",
  37951=>"000100110",
  37952=>"101101010",
  37953=>"000001001",
  37954=>"111000111",
  37955=>"010000001",
  37956=>"010010111",
  37957=>"100000010",
  37958=>"010111100",
  37959=>"111010001",
  37960=>"001111111",
  37961=>"011001011",
  37962=>"011000100",
  37963=>"011111110",
  37964=>"000000110",
  37965=>"100001111",
  37966=>"001110001",
  37967=>"100111000",
  37968=>"000111101",
  37969=>"100001110",
  37970=>"110110110",
  37971=>"100010100",
  37972=>"001001000",
  37973=>"010000001",
  37974=>"110011101",
  37975=>"000111111",
  37976=>"100101001",
  37977=>"010111010",
  37978=>"101101100",
  37979=>"111011100",
  37980=>"100010111",
  37981=>"010010011",
  37982=>"000000011",
  37983=>"000011100",
  37984=>"101011100",
  37985=>"001000011",
  37986=>"010001000",
  37987=>"100010001",
  37988=>"101000011",
  37989=>"010001010",
  37990=>"101001101",
  37991=>"000100101",
  37992=>"101011010",
  37993=>"001100000",
  37994=>"000101001",
  37995=>"001110101",
  37996=>"011001011",
  37997=>"010011110",
  37998=>"010000110",
  37999=>"101100000",
  38000=>"100010101",
  38001=>"101111011",
  38002=>"110111010",
  38003=>"101011101",
  38004=>"100111010",
  38005=>"101011101",
  38006=>"000010111",
  38007=>"100010110",
  38008=>"011001011",
  38009=>"111110001",
  38010=>"111010110",
  38011=>"111101111",
  38012=>"001000100",
  38013=>"000010011",
  38014=>"111101001",
  38015=>"110111010",
  38016=>"110000001",
  38017=>"110010111",
  38018=>"000111011",
  38019=>"001001001",
  38020=>"100011001",
  38021=>"011011011",
  38022=>"110010100",
  38023=>"100001101",
  38024=>"011001101",
  38025=>"010100000",
  38026=>"000111011",
  38027=>"010101100",
  38028=>"000110100",
  38029=>"010010010",
  38030=>"010001011",
  38031=>"100011100",
  38032=>"101001101",
  38033=>"010010000",
  38034=>"100101100",
  38035=>"111111111",
  38036=>"000101101",
  38037=>"101001010",
  38038=>"110000111",
  38039=>"011011000",
  38040=>"011111100",
  38041=>"110101100",
  38042=>"010001100",
  38043=>"100100000",
  38044=>"000011001",
  38045=>"000010010",
  38046=>"101000101",
  38047=>"111110001",
  38048=>"110111000",
  38049=>"011101011",
  38050=>"010101100",
  38051=>"111110101",
  38052=>"000000101",
  38053=>"100011101",
  38054=>"001100111",
  38055=>"110101000",
  38056=>"000100111",
  38057=>"100001101",
  38058=>"011111101",
  38059=>"011110111",
  38060=>"011001010",
  38061=>"100010011",
  38062=>"001111101",
  38063=>"001100101",
  38064=>"010100010",
  38065=>"010001100",
  38066=>"001100010",
  38067=>"001100101",
  38068=>"000000011",
  38069=>"000100101",
  38070=>"100010111",
  38071=>"011100011",
  38072=>"100101101",
  38073=>"010101110",
  38074=>"010110110",
  38075=>"011011110",
  38076=>"010010011",
  38077=>"100010110",
  38078=>"101010110",
  38079=>"101010110",
  38080=>"000010001",
  38081=>"100101000",
  38082=>"101100101",
  38083=>"101111001",
  38084=>"000001011",
  38085=>"101110110",
  38086=>"011001101",
  38087=>"101110010",
  38088=>"100000111",
  38089=>"010000001",
  38090=>"101101011",
  38091=>"101111111",
  38092=>"010110000",
  38093=>"000101011",
  38094=>"001111111",
  38095=>"111110110",
  38096=>"110111111",
  38097=>"111001101",
  38098=>"000100010",
  38099=>"010011101",
  38100=>"001111101",
  38101=>"011001101",
  38102=>"001111111",
  38103=>"100011110",
  38104=>"000000100",
  38105=>"101111101",
  38106=>"011000011",
  38107=>"111011111",
  38108=>"110001110",
  38109=>"100010010",
  38110=>"001010000",
  38111=>"010111000",
  38112=>"100111110",
  38113=>"011010000",
  38114=>"110010011",
  38115=>"001111111",
  38116=>"010010010",
  38117=>"000011101",
  38118=>"101101111",
  38119=>"100100011",
  38120=>"011001011",
  38121=>"001001110",
  38122=>"111100011",
  38123=>"010100001",
  38124=>"010111111",
  38125=>"111110100",
  38126=>"000100000",
  38127=>"101000101",
  38128=>"001011110",
  38129=>"111110011",
  38130=>"001111000",
  38131=>"111011010",
  38132=>"100111011",
  38133=>"010001001",
  38134=>"100011100",
  38135=>"000100010",
  38136=>"000010101",
  38137=>"111011111",
  38138=>"000111110",
  38139=>"011111011",
  38140=>"001110000",
  38141=>"011100011",
  38142=>"010001011",
  38143=>"100101001",
  38144=>"110000100",
  38145=>"010110000",
  38146=>"111111101",
  38147=>"101101111",
  38148=>"111000100",
  38149=>"101000111",
  38150=>"011100111",
  38151=>"000000000",
  38152=>"100111100",
  38153=>"101000001",
  38154=>"011100110",
  38155=>"010001101",
  38156=>"110110100",
  38157=>"000110111",
  38158=>"111110101",
  38159=>"000010001",
  38160=>"000101010",
  38161=>"110101101",
  38162=>"010000011",
  38163=>"111000010",
  38164=>"110001010",
  38165=>"000111110",
  38166=>"100110011",
  38167=>"000110001",
  38168=>"011010001",
  38169=>"001000111",
  38170=>"010000100",
  38171=>"001001100",
  38172=>"101111111",
  38173=>"111001100",
  38174=>"000101111",
  38175=>"101000011",
  38176=>"100100000",
  38177=>"001000010",
  38178=>"010011011",
  38179=>"011011110",
  38180=>"101101010",
  38181=>"000000001",
  38182=>"110000000",
  38183=>"100000111",
  38184=>"101011001",
  38185=>"110011100",
  38186=>"001001100",
  38187=>"110100001",
  38188=>"011100111",
  38189=>"100001111",
  38190=>"101001011",
  38191=>"101010011",
  38192=>"000100110",
  38193=>"001000100",
  38194=>"000000001",
  38195=>"101000001",
  38196=>"100011111",
  38197=>"111000010",
  38198=>"010001111",
  38199=>"000111011",
  38200=>"110010111",
  38201=>"000110010",
  38202=>"000110011",
  38203=>"011010100",
  38204=>"110000011",
  38205=>"101010001",
  38206=>"110010001",
  38207=>"101111101",
  38208=>"110001110",
  38209=>"111101010",
  38210=>"011001111",
  38211=>"000001110",
  38212=>"110110101",
  38213=>"010111010",
  38214=>"011101001",
  38215=>"100011100",
  38216=>"100000011",
  38217=>"101000101",
  38218=>"000000011",
  38219=>"000010011",
  38220=>"001011010",
  38221=>"110001100",
  38222=>"111101011",
  38223=>"101001111",
  38224=>"111101010",
  38225=>"000000100",
  38226=>"101111101",
  38227=>"001010011",
  38228=>"101101000",
  38229=>"000010011",
  38230=>"000000010",
  38231=>"111110000",
  38232=>"111000010",
  38233=>"001001010",
  38234=>"111111100",
  38235=>"001100001",
  38236=>"000010001",
  38237=>"100001000",
  38238=>"101101111",
  38239=>"000110010",
  38240=>"110010011",
  38241=>"011100000",
  38242=>"110100111",
  38243=>"010000001",
  38244=>"111110101",
  38245=>"001001101",
  38246=>"111011010",
  38247=>"011110010",
  38248=>"111010001",
  38249=>"010111111",
  38250=>"010000100",
  38251=>"001001111",
  38252=>"011111010",
  38253=>"001011110",
  38254=>"111110100",
  38255=>"101011100",
  38256=>"111110111",
  38257=>"101110010",
  38258=>"101011110",
  38259=>"010100101",
  38260=>"101010011",
  38261=>"001110011",
  38262=>"011001101",
  38263=>"010001001",
  38264=>"000011100",
  38265=>"110110110",
  38266=>"101110001",
  38267=>"101100011",
  38268=>"101000111",
  38269=>"111001111",
  38270=>"010110110",
  38271=>"111010000",
  38272=>"110111001",
  38273=>"011010000",
  38274=>"011111100",
  38275=>"100000010",
  38276=>"100101111",
  38277=>"000010100",
  38278=>"000001100",
  38279=>"011001010",
  38280=>"010101111",
  38281=>"011010100",
  38282=>"111010100",
  38283=>"100101111",
  38284=>"110010001",
  38285=>"101100000",
  38286=>"000000001",
  38287=>"101111101",
  38288=>"111101000",
  38289=>"000100000",
  38290=>"110100010",
  38291=>"111010110",
  38292=>"110001101",
  38293=>"000000001",
  38294=>"100100001",
  38295=>"101100001",
  38296=>"111101100",
  38297=>"010011111",
  38298=>"101110010",
  38299=>"110010100",
  38300=>"001111010",
  38301=>"101011001",
  38302=>"000111010",
  38303=>"001100111",
  38304=>"000111101",
  38305=>"000011111",
  38306=>"000010010",
  38307=>"010000100",
  38308=>"000011001",
  38309=>"010101011",
  38310=>"001110010",
  38311=>"111101101",
  38312=>"100101100",
  38313=>"100110010",
  38314=>"011001111",
  38315=>"111010111",
  38316=>"001000110",
  38317=>"101111111",
  38318=>"111101111",
  38319=>"010100100",
  38320=>"100110010",
  38321=>"010000000",
  38322=>"100010010",
  38323=>"100101101",
  38324=>"010100001",
  38325=>"000001010",
  38326=>"000001111",
  38327=>"010100000",
  38328=>"000111011",
  38329=>"110000011",
  38330=>"000010010",
  38331=>"000001101",
  38332=>"000000011",
  38333=>"100001101",
  38334=>"101001110",
  38335=>"111011110",
  38336=>"001001011",
  38337=>"010100111",
  38338=>"101100001",
  38339=>"111111111",
  38340=>"010011010",
  38341=>"001010000",
  38342=>"001001101",
  38343=>"110101001",
  38344=>"100000110",
  38345=>"011000001",
  38346=>"101111101",
  38347=>"100001001",
  38348=>"100000110",
  38349=>"101011000",
  38350=>"101110110",
  38351=>"011011110",
  38352=>"010100010",
  38353=>"111001110",
  38354=>"101011101",
  38355=>"010111111",
  38356=>"000001111",
  38357=>"100101101",
  38358=>"101011111",
  38359=>"000001010",
  38360=>"100111011",
  38361=>"010100101",
  38362=>"110100100",
  38363=>"111010100",
  38364=>"001010111",
  38365=>"001001011",
  38366=>"100111100",
  38367=>"111100111",
  38368=>"111011011",
  38369=>"010011000",
  38370=>"000010111",
  38371=>"000100011",
  38372=>"101101000",
  38373=>"010010100",
  38374=>"100100001",
  38375=>"011001100",
  38376=>"001000110",
  38377=>"001101110",
  38378=>"000000101",
  38379=>"001110111",
  38380=>"000010000",
  38381=>"110110001",
  38382=>"110000011",
  38383=>"000111001",
  38384=>"000011111",
  38385=>"011101100",
  38386=>"000110010",
  38387=>"000010110",
  38388=>"101000000",
  38389=>"001001001",
  38390=>"111110001",
  38391=>"010101011",
  38392=>"011101000",
  38393=>"100010010",
  38394=>"010101000",
  38395=>"111011011",
  38396=>"001000110",
  38397=>"101101000",
  38398=>"100111001",
  38399=>"000101010",
  38400=>"001101100",
  38401=>"101101011",
  38402=>"110111000",
  38403=>"001000011",
  38404=>"011001010",
  38405=>"011110001",
  38406=>"111110110",
  38407=>"100001010",
  38408=>"011011011",
  38409=>"111011011",
  38410=>"000100111",
  38411=>"100101111",
  38412=>"110000101",
  38413=>"111011111",
  38414=>"001101101",
  38415=>"101110000",
  38416=>"001000100",
  38417=>"101100011",
  38418=>"111111011",
  38419=>"101110101",
  38420=>"000000010",
  38421=>"010111110",
  38422=>"110001011",
  38423=>"101000010",
  38424=>"001111100",
  38425=>"100111110",
  38426=>"001111010",
  38427=>"110000111",
  38428=>"110010010",
  38429=>"010010010",
  38430=>"011100101",
  38431=>"000001111",
  38432=>"010011101",
  38433=>"010011110",
  38434=>"000000001",
  38435=>"010110001",
  38436=>"100001001",
  38437=>"110101011",
  38438=>"011011111",
  38439=>"111001100",
  38440=>"100001110",
  38441=>"000101100",
  38442=>"010000101",
  38443=>"110100110",
  38444=>"100011111",
  38445=>"000100110",
  38446=>"100100101",
  38447=>"000000001",
  38448=>"011000011",
  38449=>"110111000",
  38450=>"101101010",
  38451=>"111101011",
  38452=>"100010110",
  38453=>"101111011",
  38454=>"101011101",
  38455=>"111001100",
  38456=>"001011101",
  38457=>"111001101",
  38458=>"000011010",
  38459=>"011001101",
  38460=>"111000101",
  38461=>"011101101",
  38462=>"111111100",
  38463=>"011100111",
  38464=>"001101101",
  38465=>"101011110",
  38466=>"111010110",
  38467=>"000000001",
  38468=>"110101000",
  38469=>"000111001",
  38470=>"010011100",
  38471=>"001101011",
  38472=>"100110000",
  38473=>"110110111",
  38474=>"100100001",
  38475=>"111010101",
  38476=>"100101010",
  38477=>"000011000",
  38478=>"110100001",
  38479=>"011011011",
  38480=>"011000111",
  38481=>"010011101",
  38482=>"010100001",
  38483=>"000000010",
  38484=>"011011000",
  38485=>"101101001",
  38486=>"001000101",
  38487=>"011100101",
  38488=>"010110101",
  38489=>"011100110",
  38490=>"011110001",
  38491=>"011000111",
  38492=>"000100000",
  38493=>"000101100",
  38494=>"000110100",
  38495=>"010110111",
  38496=>"111101110",
  38497=>"000011000",
  38498=>"001100110",
  38499=>"101110000",
  38500=>"000011111",
  38501=>"000110001",
  38502=>"010111011",
  38503=>"100010110",
  38504=>"000010000",
  38505=>"110001000",
  38506=>"010100111",
  38507=>"001011111",
  38508=>"000001011",
  38509=>"001001010",
  38510=>"101111110",
  38511=>"111010000",
  38512=>"001101110",
  38513=>"011100011",
  38514=>"001000011",
  38515=>"001010011",
  38516=>"000011110",
  38517=>"100101001",
  38518=>"000111110",
  38519=>"111111101",
  38520=>"010010111",
  38521=>"001010111",
  38522=>"000000110",
  38523=>"100100110",
  38524=>"011100111",
  38525=>"100010101",
  38526=>"000010101",
  38527=>"011010110",
  38528=>"111100110",
  38529=>"111111011",
  38530=>"010111001",
  38531=>"010011110",
  38532=>"011111110",
  38533=>"000001001",
  38534=>"111001101",
  38535=>"100111001",
  38536=>"000011100",
  38537=>"010000010",
  38538=>"111010001",
  38539=>"100000101",
  38540=>"111110001",
  38541=>"101111101",
  38542=>"101100111",
  38543=>"100100111",
  38544=>"011101101",
  38545=>"001100110",
  38546=>"011010000",
  38547=>"001001000",
  38548=>"001101101",
  38549=>"111100100",
  38550=>"110011010",
  38551=>"110010111",
  38552=>"100000000",
  38553=>"010010110",
  38554=>"111011101",
  38555=>"110011000",
  38556=>"101110100",
  38557=>"001010000",
  38558=>"100000101",
  38559=>"110000010",
  38560=>"101101111",
  38561=>"000100011",
  38562=>"010111110",
  38563=>"101110010",
  38564=>"011000011",
  38565=>"110000111",
  38566=>"110101101",
  38567=>"100010010",
  38568=>"010111000",
  38569=>"000001111",
  38570=>"001000111",
  38571=>"111111110",
  38572=>"101000110",
  38573=>"111000001",
  38574=>"110111000",
  38575=>"000000001",
  38576=>"000000011",
  38577=>"101001100",
  38578=>"001110100",
  38579=>"011100111",
  38580=>"011101111",
  38581=>"001111101",
  38582=>"101111111",
  38583=>"010010111",
  38584=>"100011010",
  38585=>"011111010",
  38586=>"000111111",
  38587=>"110001111",
  38588=>"111110101",
  38589=>"110111110",
  38590=>"000111101",
  38591=>"001000111",
  38592=>"000110110",
  38593=>"001111101",
  38594=>"001011100",
  38595=>"101100000",
  38596=>"011000011",
  38597=>"010010000",
  38598=>"111011011",
  38599=>"010001011",
  38600=>"101000000",
  38601=>"010010111",
  38602=>"110100100",
  38603=>"010000100",
  38604=>"010110111",
  38605=>"100110110",
  38606=>"101001010",
  38607=>"100010001",
  38608=>"000001101",
  38609=>"011001000",
  38610=>"011110110",
  38611=>"101101001",
  38612=>"000001011",
  38613=>"000010000",
  38614=>"100100011",
  38615=>"010011011",
  38616=>"011011101",
  38617=>"101000110",
  38618=>"000101011",
  38619=>"110111101",
  38620=>"111000110",
  38621=>"111100101",
  38622=>"100010101",
  38623=>"000100111",
  38624=>"001110111",
  38625=>"000100111",
  38626=>"001110000",
  38627=>"101110111",
  38628=>"000000101",
  38629=>"101101111",
  38630=>"111101111",
  38631=>"100101000",
  38632=>"100011111",
  38633=>"101100001",
  38634=>"010111000",
  38635=>"001110001",
  38636=>"100111100",
  38637=>"011111111",
  38638=>"000000110",
  38639=>"111111110",
  38640=>"011110110",
  38641=>"011111010",
  38642=>"110110111",
  38643=>"001001101",
  38644=>"101001001",
  38645=>"101010000",
  38646=>"010001101",
  38647=>"000000101",
  38648=>"000001100",
  38649=>"011010110",
  38650=>"111101110",
  38651=>"000110100",
  38652=>"110001101",
  38653=>"000100111",
  38654=>"110111101",
  38655=>"001001001",
  38656=>"100011111",
  38657=>"110010111",
  38658=>"010101001",
  38659=>"000001000",
  38660=>"000001101",
  38661=>"101111000",
  38662=>"111100101",
  38663=>"010101001",
  38664=>"111110110",
  38665=>"110110010",
  38666=>"110100001",
  38667=>"000001011",
  38668=>"100001110",
  38669=>"000000110",
  38670=>"011110010",
  38671=>"001111110",
  38672=>"101101010",
  38673=>"011001010",
  38674=>"000100011",
  38675=>"000001111",
  38676=>"101100110",
  38677=>"000000101",
  38678=>"100111111",
  38679=>"011001101",
  38680=>"011011100",
  38681=>"100011000",
  38682=>"001100111",
  38683=>"000000110",
  38684=>"100001100",
  38685=>"111110111",
  38686=>"010101000",
  38687=>"001010000",
  38688=>"111111111",
  38689=>"111111101",
  38690=>"000000011",
  38691=>"110000001",
  38692=>"100001010",
  38693=>"010100110",
  38694=>"010000011",
  38695=>"001101001",
  38696=>"011110110",
  38697=>"111101100",
  38698=>"111010010",
  38699=>"011000110",
  38700=>"111010001",
  38701=>"110110101",
  38702=>"000001000",
  38703=>"000001001",
  38704=>"011011110",
  38705=>"010100111",
  38706=>"010110110",
  38707=>"011000110",
  38708=>"101110000",
  38709=>"010000010",
  38710=>"001111011",
  38711=>"000101000",
  38712=>"001100011",
  38713=>"010001001",
  38714=>"111111010",
  38715=>"000111110",
  38716=>"010010111",
  38717=>"000111001",
  38718=>"010000111",
  38719=>"000110011",
  38720=>"000111010",
  38721=>"000001010",
  38722=>"111101110",
  38723=>"000001100",
  38724=>"110010011",
  38725=>"001011011",
  38726=>"111101010",
  38727=>"110001001",
  38728=>"111011001",
  38729=>"101100110",
  38730=>"100011100",
  38731=>"111000010",
  38732=>"001101011",
  38733=>"011111111",
  38734=>"111100011",
  38735=>"111101011",
  38736=>"101111000",
  38737=>"000110000",
  38738=>"010100111",
  38739=>"100100110",
  38740=>"111101101",
  38741=>"011110010",
  38742=>"010010101",
  38743=>"010011100",
  38744=>"110100010",
  38745=>"010100001",
  38746=>"101001100",
  38747=>"000000111",
  38748=>"010100010",
  38749=>"001111111",
  38750=>"100011101",
  38751=>"010000000",
  38752=>"011101010",
  38753=>"010101010",
  38754=>"100010100",
  38755=>"001111101",
  38756=>"011110111",
  38757=>"011111111",
  38758=>"011110111",
  38759=>"101111010",
  38760=>"111001110",
  38761=>"010010111",
  38762=>"101011010",
  38763=>"000010000",
  38764=>"100011111",
  38765=>"101101011",
  38766=>"011101001",
  38767=>"010110111",
  38768=>"110001110",
  38769=>"101001100",
  38770=>"101110011",
  38771=>"001000110",
  38772=>"010010001",
  38773=>"001110001",
  38774=>"010001010",
  38775=>"000001111",
  38776=>"010101110",
  38777=>"111001101",
  38778=>"001110100",
  38779=>"111011111",
  38780=>"000000010",
  38781=>"111101001",
  38782=>"101111000",
  38783=>"001110000",
  38784=>"001010111",
  38785=>"111111101",
  38786=>"010110010",
  38787=>"110100110",
  38788=>"011111100",
  38789=>"110001000",
  38790=>"110110100",
  38791=>"000000101",
  38792=>"001011001",
  38793=>"100001010",
  38794=>"011110001",
  38795=>"101111111",
  38796=>"110000100",
  38797=>"100011011",
  38798=>"011100110",
  38799=>"110001111",
  38800=>"110101100",
  38801=>"101111111",
  38802=>"001010000",
  38803=>"011000000",
  38804=>"101110110",
  38805=>"101110010",
  38806=>"100101110",
  38807=>"010110000",
  38808=>"001001010",
  38809=>"010010011",
  38810=>"011010101",
  38811=>"110001111",
  38812=>"110000100",
  38813=>"010011011",
  38814=>"111101100",
  38815=>"001101011",
  38816=>"101110000",
  38817=>"100111100",
  38818=>"110111101",
  38819=>"001111111",
  38820=>"001000001",
  38821=>"000010111",
  38822=>"001000001",
  38823=>"110101100",
  38824=>"101101110",
  38825=>"111001111",
  38826=>"110110100",
  38827=>"111011110",
  38828=>"000101011",
  38829=>"101110100",
  38830=>"000000000",
  38831=>"001100001",
  38832=>"011101011",
  38833=>"000011101",
  38834=>"110001001",
  38835=>"100000100",
  38836=>"110100100",
  38837=>"010010110",
  38838=>"010001111",
  38839=>"000100110",
  38840=>"000110001",
  38841=>"010000101",
  38842=>"110100010",
  38843=>"000011100",
  38844=>"100000110",
  38845=>"000000100",
  38846=>"111111101",
  38847=>"011110110",
  38848=>"011010101",
  38849=>"011010001",
  38850=>"011001011",
  38851=>"000111110",
  38852=>"010100001",
  38853=>"110010100",
  38854=>"011100000",
  38855=>"110110010",
  38856=>"010000010",
  38857=>"001110011",
  38858=>"111000010",
  38859=>"011001100",
  38860=>"111110001",
  38861=>"111010111",
  38862=>"000100010",
  38863=>"000011001",
  38864=>"110100001",
  38865=>"001011100",
  38866=>"011000110",
  38867=>"100111101",
  38868=>"100111000",
  38869=>"001101100",
  38870=>"101101011",
  38871=>"111100001",
  38872=>"101010000",
  38873=>"011011100",
  38874=>"101010011",
  38875=>"111010001",
  38876=>"000111110",
  38877=>"110100010",
  38878=>"101111111",
  38879=>"100111110",
  38880=>"111010101",
  38881=>"111011010",
  38882=>"000101110",
  38883=>"110111001",
  38884=>"100110001",
  38885=>"001000100",
  38886=>"001110100",
  38887=>"010010000",
  38888=>"011011100",
  38889=>"110111110",
  38890=>"110100001",
  38891=>"001101110",
  38892=>"000000100",
  38893=>"000000111",
  38894=>"111011010",
  38895=>"011100000",
  38896=>"000001100",
  38897=>"011011110",
  38898=>"110001100",
  38899=>"100111011",
  38900=>"110010100",
  38901=>"100111100",
  38902=>"111101100",
  38903=>"010111101",
  38904=>"111000000",
  38905=>"000101001",
  38906=>"110111111",
  38907=>"101101010",
  38908=>"100111110",
  38909=>"110000100",
  38910=>"101010101",
  38911=>"110101000",
  38912=>"000011101",
  38913=>"001010000",
  38914=>"000011100",
  38915=>"010010000",
  38916=>"001111111",
  38917=>"101001010",
  38918=>"001001111",
  38919=>"100000101",
  38920=>"101100000",
  38921=>"100011000",
  38922=>"111111110",
  38923=>"011001011",
  38924=>"001000000",
  38925=>"010011011",
  38926=>"001000011",
  38927=>"111110110",
  38928=>"101100110",
  38929=>"100101010",
  38930=>"101100010",
  38931=>"001110011",
  38932=>"111111001",
  38933=>"111101011",
  38934=>"100110110",
  38935=>"110001111",
  38936=>"011111101",
  38937=>"001111001",
  38938=>"100111000",
  38939=>"011101000",
  38940=>"100111010",
  38941=>"011101001",
  38942=>"101101110",
  38943=>"000101110",
  38944=>"001100000",
  38945=>"001011010",
  38946=>"110000000",
  38947=>"010010101",
  38948=>"011101000",
  38949=>"010111101",
  38950=>"110001100",
  38951=>"001110000",
  38952=>"011110001",
  38953=>"110010000",
  38954=>"001101010",
  38955=>"011010010",
  38956=>"000000000",
  38957=>"111111111",
  38958=>"011101100",
  38959=>"101000111",
  38960=>"010001101",
  38961=>"010011111",
  38962=>"000110101",
  38963=>"011110100",
  38964=>"111000110",
  38965=>"101111111",
  38966=>"010011011",
  38967=>"001101010",
  38968=>"101100100",
  38969=>"001000000",
  38970=>"001110110",
  38971=>"000011010",
  38972=>"000000011",
  38973=>"101110100",
  38974=>"111001001",
  38975=>"100100011",
  38976=>"001110111",
  38977=>"001001000",
  38978=>"000101110",
  38979=>"000000001",
  38980=>"101000010",
  38981=>"110011101",
  38982=>"011111100",
  38983=>"101111110",
  38984=>"111110000",
  38985=>"010100111",
  38986=>"011010001",
  38987=>"100110111",
  38988=>"111101010",
  38989=>"100011000",
  38990=>"110000101",
  38991=>"011011111",
  38992=>"110100111",
  38993=>"110001010",
  38994=>"010010111",
  38995=>"010011110",
  38996=>"100101110",
  38997=>"110100011",
  38998=>"111011010",
  38999=>"001010001",
  39000=>"100110111",
  39001=>"101001010",
  39002=>"010010010",
  39003=>"011001101",
  39004=>"110001010",
  39005=>"101101000",
  39006=>"110001000",
  39007=>"011111001",
  39008=>"011011011",
  39009=>"110011011",
  39010=>"000011011",
  39011=>"011010101",
  39012=>"000010000",
  39013=>"000001001",
  39014=>"010111111",
  39015=>"110101000",
  39016=>"110010111",
  39017=>"001110100",
  39018=>"111010110",
  39019=>"101100000",
  39020=>"110010001",
  39021=>"110100110",
  39022=>"001100100",
  39023=>"100010001",
  39024=>"100101010",
  39025=>"011010000",
  39026=>"011110011",
  39027=>"000100100",
  39028=>"101110101",
  39029=>"000110000",
  39030=>"010010011",
  39031=>"111100011",
  39032=>"010010100",
  39033=>"010000001",
  39034=>"110111101",
  39035=>"101111010",
  39036=>"011011011",
  39037=>"001010100",
  39038=>"010011000",
  39039=>"110001011",
  39040=>"110000010",
  39041=>"100010111",
  39042=>"001111000",
  39043=>"001001100",
  39044=>"011001010",
  39045=>"100000000",
  39046=>"111110111",
  39047=>"010011110",
  39048=>"001110111",
  39049=>"110001111",
  39050=>"001101010",
  39051=>"110000010",
  39052=>"011011011",
  39053=>"110100001",
  39054=>"111011010",
  39055=>"011100000",
  39056=>"001100010",
  39057=>"101110101",
  39058=>"000010001",
  39059=>"111010010",
  39060=>"100110000",
  39061=>"110101010",
  39062=>"101011001",
  39063=>"100010111",
  39064=>"101010101",
  39065=>"001101001",
  39066=>"101000111",
  39067=>"001101000",
  39068=>"001011110",
  39069=>"111001111",
  39070=>"010111111",
  39071=>"000100001",
  39072=>"101111111",
  39073=>"110110110",
  39074=>"001011110",
  39075=>"101001011",
  39076=>"100110000",
  39077=>"000010010",
  39078=>"001011100",
  39079=>"101001110",
  39080=>"000010010",
  39081=>"001101101",
  39082=>"101111001",
  39083=>"001101100",
  39084=>"011010110",
  39085=>"100001101",
  39086=>"100100100",
  39087=>"010111011",
  39088=>"011100011",
  39089=>"000001000",
  39090=>"100110010",
  39091=>"111000011",
  39092=>"111010101",
  39093=>"011110000",
  39094=>"101101101",
  39095=>"001110110",
  39096=>"111000011",
  39097=>"100101010",
  39098=>"000101100",
  39099=>"010011001",
  39100=>"001010100",
  39101=>"010010111",
  39102=>"001111100",
  39103=>"111101001",
  39104=>"111101101",
  39105=>"010110100",
  39106=>"101111001",
  39107=>"010110110",
  39108=>"101010110",
  39109=>"000111001",
  39110=>"011001101",
  39111=>"100011010",
  39112=>"110110101",
  39113=>"000111101",
  39114=>"111111001",
  39115=>"001110100",
  39116=>"111010010",
  39117=>"000011001",
  39118=>"010111000",
  39119=>"011111111",
  39120=>"101001000",
  39121=>"010111111",
  39122=>"011101110",
  39123=>"000100001",
  39124=>"011100000",
  39125=>"111100010",
  39126=>"000001000",
  39127=>"101100101",
  39128=>"101100010",
  39129=>"100001000",
  39130=>"100001100",
  39131=>"010100000",
  39132=>"110100000",
  39133=>"111100101",
  39134=>"000100101",
  39135=>"000001001",
  39136=>"100011100",
  39137=>"110010011",
  39138=>"001010000",
  39139=>"111101000",
  39140=>"011010100",
  39141=>"101010010",
  39142=>"100101101",
  39143=>"000100011",
  39144=>"100100011",
  39145=>"011010000",
  39146=>"001011010",
  39147=>"100011001",
  39148=>"110100110",
  39149=>"101001101",
  39150=>"000110000",
  39151=>"101011111",
  39152=>"001010111",
  39153=>"111000110",
  39154=>"010000010",
  39155=>"010000000",
  39156=>"101100010",
  39157=>"010110011",
  39158=>"100000000",
  39159=>"111011000",
  39160=>"101010100",
  39161=>"100000000",
  39162=>"111010100",
  39163=>"110001110",
  39164=>"001110110",
  39165=>"100001001",
  39166=>"001001000",
  39167=>"100000010",
  39168=>"010001101",
  39169=>"001000000",
  39170=>"101001011",
  39171=>"001100010",
  39172=>"011001011",
  39173=>"110101000",
  39174=>"101100111",
  39175=>"101010010",
  39176=>"010000000",
  39177=>"101100100",
  39178=>"110010111",
  39179=>"101101011",
  39180=>"011110101",
  39181=>"101111000",
  39182=>"010101100",
  39183=>"011100100",
  39184=>"011101101",
  39185=>"101101000",
  39186=>"110110010",
  39187=>"100111001",
  39188=>"010100101",
  39189=>"011101101",
  39190=>"110011000",
  39191=>"011001010",
  39192=>"000111100",
  39193=>"100011101",
  39194=>"100001100",
  39195=>"011010110",
  39196=>"111111010",
  39197=>"011100101",
  39198=>"100101001",
  39199=>"111011100",
  39200=>"000001010",
  39201=>"111100001",
  39202=>"111111111",
  39203=>"010010011",
  39204=>"011100100",
  39205=>"100001000",
  39206=>"101101111",
  39207=>"010110000",
  39208=>"001000110",
  39209=>"100011100",
  39210=>"110011101",
  39211=>"100000111",
  39212=>"110001110",
  39213=>"110000111",
  39214=>"001101110",
  39215=>"001100011",
  39216=>"100011011",
  39217=>"100101111",
  39218=>"110111111",
  39219=>"110100010",
  39220=>"011110011",
  39221=>"110001010",
  39222=>"001000111",
  39223=>"010010011",
  39224=>"010001101",
  39225=>"101010001",
  39226=>"110111000",
  39227=>"001000101",
  39228=>"000101010",
  39229=>"010010010",
  39230=>"011101110",
  39231=>"000011001",
  39232=>"010101001",
  39233=>"100000110",
  39234=>"000101000",
  39235=>"101101101",
  39236=>"001000101",
  39237=>"101010100",
  39238=>"011100100",
  39239=>"011100110",
  39240=>"101000001",
  39241=>"000111100",
  39242=>"101000101",
  39243=>"110011000",
  39244=>"011011010",
  39245=>"001001010",
  39246=>"011111010",
  39247=>"111100100",
  39248=>"011111101",
  39249=>"000100001",
  39250=>"111010111",
  39251=>"101010101",
  39252=>"011000111",
  39253=>"000110011",
  39254=>"010011110",
  39255=>"011111101",
  39256=>"010100010",
  39257=>"010101000",
  39258=>"100101001",
  39259=>"101001010",
  39260=>"100100001",
  39261=>"100010111",
  39262=>"010110110",
  39263=>"000010110",
  39264=>"111111101",
  39265=>"010000001",
  39266=>"111100101",
  39267=>"101001110",
  39268=>"100010101",
  39269=>"001111000",
  39270=>"111011111",
  39271=>"010010101",
  39272=>"000001011",
  39273=>"111011110",
  39274=>"110110011",
  39275=>"011000000",
  39276=>"100000101",
  39277=>"101100011",
  39278=>"001101111",
  39279=>"110010010",
  39280=>"011000100",
  39281=>"010010110",
  39282=>"111111110",
  39283=>"111000001",
  39284=>"010110010",
  39285=>"011000101",
  39286=>"000000111",
  39287=>"101101000",
  39288=>"010010011",
  39289=>"011101010",
  39290=>"111011110",
  39291=>"111001110",
  39292=>"110110101",
  39293=>"010000001",
  39294=>"000100001",
  39295=>"110010110",
  39296=>"100010000",
  39297=>"111000100",
  39298=>"010010001",
  39299=>"111110000",
  39300=>"011111101",
  39301=>"100000111",
  39302=>"111111111",
  39303=>"111111101",
  39304=>"011111110",
  39305=>"111111111",
  39306=>"000111111",
  39307=>"000100000",
  39308=>"001101010",
  39309=>"011110110",
  39310=>"111110111",
  39311=>"011011001",
  39312=>"111010010",
  39313=>"011011010",
  39314=>"000001011",
  39315=>"001011101",
  39316=>"000011011",
  39317=>"010100001",
  39318=>"100000000",
  39319=>"101001000",
  39320=>"001110111",
  39321=>"011010000",
  39322=>"111100010",
  39323=>"110101111",
  39324=>"001111100",
  39325=>"000100110",
  39326=>"101000111",
  39327=>"110111011",
  39328=>"111010010",
  39329=>"100000100",
  39330=>"010100111",
  39331=>"101011011",
  39332=>"000101000",
  39333=>"110000101",
  39334=>"111101111",
  39335=>"010110011",
  39336=>"101010011",
  39337=>"101000011",
  39338=>"101000000",
  39339=>"000000000",
  39340=>"001110101",
  39341=>"001110111",
  39342=>"000011110",
  39343=>"011011011",
  39344=>"101001101",
  39345=>"101101111",
  39346=>"111111001",
  39347=>"011110001",
  39348=>"000000010",
  39349=>"011100010",
  39350=>"000101101",
  39351=>"011101111",
  39352=>"101000101",
  39353=>"010011111",
  39354=>"000000100",
  39355=>"110010000",
  39356=>"001101101",
  39357=>"000011110",
  39358=>"001001011",
  39359=>"001001001",
  39360=>"100010010",
  39361=>"001000011",
  39362=>"101011001",
  39363=>"101111000",
  39364=>"010010000",
  39365=>"110110100",
  39366=>"000001101",
  39367=>"101110000",
  39368=>"011111100",
  39369=>"111110010",
  39370=>"011100100",
  39371=>"100010101",
  39372=>"000011010",
  39373=>"011110110",
  39374=>"100101000",
  39375=>"010101110",
  39376=>"110010010",
  39377=>"101011011",
  39378=>"111011011",
  39379=>"010100110",
  39380=>"111110111",
  39381=>"100010000",
  39382=>"101011100",
  39383=>"001001101",
  39384=>"110100110",
  39385=>"010101100",
  39386=>"001101100",
  39387=>"110010011",
  39388=>"100100111",
  39389=>"011101011",
  39390=>"001001101",
  39391=>"010001011",
  39392=>"111010101",
  39393=>"110111110",
  39394=>"110010101",
  39395=>"100110000",
  39396=>"110110101",
  39397=>"110100000",
  39398=>"000001011",
  39399=>"001101010",
  39400=>"000100010",
  39401=>"010001010",
  39402=>"001100110",
  39403=>"011110110",
  39404=>"110101000",
  39405=>"011001001",
  39406=>"111111111",
  39407=>"000101011",
  39408=>"010011101",
  39409=>"111010100",
  39410=>"011110010",
  39411=>"111010010",
  39412=>"011000100",
  39413=>"001111110",
  39414=>"111100110",
  39415=>"000101000",
  39416=>"001011011",
  39417=>"110101100",
  39418=>"011101110",
  39419=>"111101011",
  39420=>"010001000",
  39421=>"010101011",
  39422=>"000000110",
  39423=>"100101110",
  39424=>"111101111",
  39425=>"100101011",
  39426=>"011101110",
  39427=>"111100001",
  39428=>"100000111",
  39429=>"101000001",
  39430=>"010000001",
  39431=>"110011101",
  39432=>"111101011",
  39433=>"011011100",
  39434=>"101011100",
  39435=>"011110110",
  39436=>"011000110",
  39437=>"110010101",
  39438=>"000101010",
  39439=>"110100101",
  39440=>"101111111",
  39441=>"010000001",
  39442=>"010010111",
  39443=>"111011011",
  39444=>"111010001",
  39445=>"101001110",
  39446=>"011111010",
  39447=>"000111000",
  39448=>"001111100",
  39449=>"000001010",
  39450=>"000100100",
  39451=>"001111011",
  39452=>"001001000",
  39453=>"011010001",
  39454=>"111111010",
  39455=>"100101000",
  39456=>"000000001",
  39457=>"101001101",
  39458=>"100000111",
  39459=>"010110001",
  39460=>"110000001",
  39461=>"111110010",
  39462=>"110011110",
  39463=>"011100100",
  39464=>"110110001",
  39465=>"001111101",
  39466=>"010100010",
  39467=>"001100011",
  39468=>"100100100",
  39469=>"100110100",
  39470=>"111100101",
  39471=>"000011010",
  39472=>"011011100",
  39473=>"101010111",
  39474=>"001110110",
  39475=>"011101010",
  39476=>"111011101",
  39477=>"000111100",
  39478=>"100101011",
  39479=>"000000001",
  39480=>"011100011",
  39481=>"110100100",
  39482=>"010010001",
  39483=>"001101000",
  39484=>"110011000",
  39485=>"100010000",
  39486=>"000100100",
  39487=>"100110111",
  39488=>"111111111",
  39489=>"000010000",
  39490=>"101001111",
  39491=>"110101000",
  39492=>"111110111",
  39493=>"010001011",
  39494=>"001010100",
  39495=>"101001000",
  39496=>"001000111",
  39497=>"010110000",
  39498=>"000010001",
  39499=>"100011111",
  39500=>"101101101",
  39501=>"001010000",
  39502=>"000001100",
  39503=>"000111101",
  39504=>"101000001",
  39505=>"010000011",
  39506=>"000010101",
  39507=>"010110100",
  39508=>"100100000",
  39509=>"010000011",
  39510=>"000000000",
  39511=>"010011001",
  39512=>"000000100",
  39513=>"000001000",
  39514=>"111011000",
  39515=>"001100000",
  39516=>"110101110",
  39517=>"111110010",
  39518=>"001101100",
  39519=>"000011111",
  39520=>"111001011",
  39521=>"101011110",
  39522=>"110111000",
  39523=>"110011111",
  39524=>"111110111",
  39525=>"001000100",
  39526=>"010100101",
  39527=>"001101010",
  39528=>"010011011",
  39529=>"000110111",
  39530=>"000111101",
  39531=>"100011011",
  39532=>"110100011",
  39533=>"010011011",
  39534=>"101111110",
  39535=>"111011001",
  39536=>"101111010",
  39537=>"010000100",
  39538=>"001010000",
  39539=>"110101100",
  39540=>"010110101",
  39541=>"011001001",
  39542=>"111101011",
  39543=>"111010010",
  39544=>"100010000",
  39545=>"101111110",
  39546=>"111000010",
  39547=>"101110011",
  39548=>"010111000",
  39549=>"110111110",
  39550=>"000000001",
  39551=>"001011110",
  39552=>"001110000",
  39553=>"110011111",
  39554=>"110100010",
  39555=>"101000001",
  39556=>"100101001",
  39557=>"110010000",
  39558=>"111011100",
  39559=>"100100001",
  39560=>"101111101",
  39561=>"111111110",
  39562=>"110111001",
  39563=>"101011001",
  39564=>"010001011",
  39565=>"001100010",
  39566=>"101011010",
  39567=>"000100111",
  39568=>"100110010",
  39569=>"111101111",
  39570=>"011001110",
  39571=>"111110000",
  39572=>"001000000",
  39573=>"010110100",
  39574=>"001101000",
  39575=>"100110010",
  39576=>"001101100",
  39577=>"110011000",
  39578=>"100101110",
  39579=>"000110000",
  39580=>"100001001",
  39581=>"000110001",
  39582=>"100010001",
  39583=>"010111111",
  39584=>"101111101",
  39585=>"111001000",
  39586=>"000110111",
  39587=>"001101000",
  39588=>"011000011",
  39589=>"010011111",
  39590=>"100011110",
  39591=>"000100101",
  39592=>"110110000",
  39593=>"111100011",
  39594=>"110000000",
  39595=>"010011100",
  39596=>"011000101",
  39597=>"001001000",
  39598=>"111111010",
  39599=>"100001000",
  39600=>"101100001",
  39601=>"000010100",
  39602=>"010111100",
  39603=>"101010001",
  39604=>"010010101",
  39605=>"000100001",
  39606=>"111100100",
  39607=>"110000010",
  39608=>"010111011",
  39609=>"111111110",
  39610=>"101101001",
  39611=>"000011100",
  39612=>"010000011",
  39613=>"001100111",
  39614=>"001101101",
  39615=>"100011000",
  39616=>"111110000",
  39617=>"111111000",
  39618=>"000111110",
  39619=>"100111100",
  39620=>"111100110",
  39621=>"010001111",
  39622=>"001001011",
  39623=>"101010100",
  39624=>"100010010",
  39625=>"001100111",
  39626=>"010110100",
  39627=>"011111110",
  39628=>"100110101",
  39629=>"110000000",
  39630=>"100101011",
  39631=>"000000011",
  39632=>"100000111",
  39633=>"011011000",
  39634=>"011110000",
  39635=>"110000001",
  39636=>"100001000",
  39637=>"001000000",
  39638=>"010101101",
  39639=>"000000111",
  39640=>"010000010",
  39641=>"001110001",
  39642=>"100100010",
  39643=>"001011000",
  39644=>"101101101",
  39645=>"110010111",
  39646=>"000111100",
  39647=>"000011110",
  39648=>"101111010",
  39649=>"001010100",
  39650=>"010001110",
  39651=>"011101011",
  39652=>"010000010",
  39653=>"111110001",
  39654=>"101000100",
  39655=>"111101010",
  39656=>"101110110",
  39657=>"111110011",
  39658=>"011110111",
  39659=>"001011011",
  39660=>"110011001",
  39661=>"111101110",
  39662=>"100011101",
  39663=>"000000010",
  39664=>"010100000",
  39665=>"110111101",
  39666=>"000111011",
  39667=>"100100010",
  39668=>"001101000",
  39669=>"101111110",
  39670=>"010100101",
  39671=>"001111001",
  39672=>"001100010",
  39673=>"101011010",
  39674=>"111011100",
  39675=>"110111101",
  39676=>"000011001",
  39677=>"000000100",
  39678=>"001000011",
  39679=>"100100010",
  39680=>"101001001",
  39681=>"010000101",
  39682=>"010111100",
  39683=>"001101010",
  39684=>"100000100",
  39685=>"001001100",
  39686=>"000011000",
  39687=>"011110110",
  39688=>"010011000",
  39689=>"101100011",
  39690=>"000101110",
  39691=>"110001011",
  39692=>"101111010",
  39693=>"100000111",
  39694=>"000011000",
  39695=>"100110010",
  39696=>"111101000",
  39697=>"110011011",
  39698=>"001001011",
  39699=>"111100110",
  39700=>"101010000",
  39701=>"110110010",
  39702=>"001101110",
  39703=>"111100011",
  39704=>"011010000",
  39705=>"001000000",
  39706=>"010001000",
  39707=>"011011001",
  39708=>"111110001",
  39709=>"110010001",
  39710=>"010111100",
  39711=>"000010010",
  39712=>"001010110",
  39713=>"101000010",
  39714=>"000011110",
  39715=>"011010111",
  39716=>"011101000",
  39717=>"010010100",
  39718=>"011101101",
  39719=>"101100010",
  39720=>"011100110",
  39721=>"000100010",
  39722=>"111101010",
  39723=>"000110000",
  39724=>"111001000",
  39725=>"010101010",
  39726=>"001100101",
  39727=>"011100001",
  39728=>"011101111",
  39729=>"101011100",
  39730=>"000111011",
  39731=>"000001001",
  39732=>"101111111",
  39733=>"011011110",
  39734=>"011001010",
  39735=>"000100110",
  39736=>"110110100",
  39737=>"011000001",
  39738=>"000011111",
  39739=>"001110011",
  39740=>"000101011",
  39741=>"110011000",
  39742=>"101111011",
  39743=>"010001010",
  39744=>"001011001",
  39745=>"010000000",
  39746=>"001010111",
  39747=>"100000110",
  39748=>"111010101",
  39749=>"011000101",
  39750=>"001100100",
  39751=>"101010100",
  39752=>"101100011",
  39753=>"101010000",
  39754=>"101100101",
  39755=>"000110011",
  39756=>"110111000",
  39757=>"011100101",
  39758=>"100000011",
  39759=>"000100111",
  39760=>"010000111",
  39761=>"101011000",
  39762=>"011010100",
  39763=>"110110100",
  39764=>"010000000",
  39765=>"011100000",
  39766=>"110010110",
  39767=>"111000001",
  39768=>"100010000",
  39769=>"111101010",
  39770=>"101010101",
  39771=>"101000001",
  39772=>"100011110",
  39773=>"001111011",
  39774=>"011110111",
  39775=>"110000100",
  39776=>"100110000",
  39777=>"010101001",
  39778=>"000000010",
  39779=>"111100111",
  39780=>"010010111",
  39781=>"000100001",
  39782=>"111010110",
  39783=>"001001010",
  39784=>"101000100",
  39785=>"011101000",
  39786=>"111011110",
  39787=>"100100101",
  39788=>"100101000",
  39789=>"011100011",
  39790=>"000111110",
  39791=>"000001011",
  39792=>"000011010",
  39793=>"101010100",
  39794=>"100110010",
  39795=>"100100110",
  39796=>"111110101",
  39797=>"000000001",
  39798=>"101000011",
  39799=>"010101000",
  39800=>"101000011",
  39801=>"101110100",
  39802=>"101111011",
  39803=>"000010100",
  39804=>"010100100",
  39805=>"110100100",
  39806=>"000100110",
  39807=>"110010010",
  39808=>"011000100",
  39809=>"000001110",
  39810=>"100001001",
  39811=>"011100011",
  39812=>"000100011",
  39813=>"110011011",
  39814=>"010000100",
  39815=>"000110111",
  39816=>"011110011",
  39817=>"010010010",
  39818=>"110011011",
  39819=>"110110111",
  39820=>"110110010",
  39821=>"000111011",
  39822=>"001000110",
  39823=>"101101000",
  39824=>"001110100",
  39825=>"111110010",
  39826=>"110000011",
  39827=>"111101111",
  39828=>"001010000",
  39829=>"010011111",
  39830=>"111110001",
  39831=>"000000000",
  39832=>"111110101",
  39833=>"110010111",
  39834=>"101101011",
  39835=>"100101010",
  39836=>"010101010",
  39837=>"100110011",
  39838=>"101110100",
  39839=>"000011110",
  39840=>"101110010",
  39841=>"111111011",
  39842=>"001110101",
  39843=>"101111111",
  39844=>"111111000",
  39845=>"100001111",
  39846=>"111101100",
  39847=>"011010010",
  39848=>"111000100",
  39849=>"111101111",
  39850=>"011101100",
  39851=>"010001011",
  39852=>"110100101",
  39853=>"111111110",
  39854=>"011110100",
  39855=>"011011100",
  39856=>"100111000",
  39857=>"001100100",
  39858=>"001011011",
  39859=>"101110011",
  39860=>"110100101",
  39861=>"110100111",
  39862=>"000100100",
  39863=>"101001101",
  39864=>"110101110",
  39865=>"101011000",
  39866=>"000011001",
  39867=>"111111101",
  39868=>"111111011",
  39869=>"101000011",
  39870=>"000110101",
  39871=>"100100111",
  39872=>"011111110",
  39873=>"101100100",
  39874=>"111000010",
  39875=>"111001110",
  39876=>"110100110",
  39877=>"110110010",
  39878=>"110100100",
  39879=>"000101110",
  39880=>"100011010",
  39881=>"000111101",
  39882=>"000010001",
  39883=>"001000000",
  39884=>"011100101",
  39885=>"101101111",
  39886=>"001110111",
  39887=>"001011001",
  39888=>"001000111",
  39889=>"100011010",
  39890=>"101000011",
  39891=>"000000010",
  39892=>"110011110",
  39893=>"001010011",
  39894=>"011011111",
  39895=>"010100111",
  39896=>"000101111",
  39897=>"110100010",
  39898=>"000100101",
  39899=>"110100001",
  39900=>"110011001",
  39901=>"110101011",
  39902=>"101101110",
  39903=>"010110101",
  39904=>"010000000",
  39905=>"110100011",
  39906=>"001000000",
  39907=>"110101000",
  39908=>"100001000",
  39909=>"010010000",
  39910=>"111010101",
  39911=>"111100000",
  39912=>"111101010",
  39913=>"110010110",
  39914=>"001100000",
  39915=>"111100000",
  39916=>"110011111",
  39917=>"101011100",
  39918=>"111000101",
  39919=>"101001010",
  39920=>"000000000",
  39921=>"001111000",
  39922=>"010000011",
  39923=>"001101100",
  39924=>"100010100",
  39925=>"000100001",
  39926=>"111001110",
  39927=>"100101000",
  39928=>"000110000",
  39929=>"110001000",
  39930=>"001011001",
  39931=>"010100111",
  39932=>"110001011",
  39933=>"110010110",
  39934=>"000000000",
  39935=>"011101011",
  39936=>"100100100",
  39937=>"000010111",
  39938=>"010000001",
  39939=>"000001010",
  39940=>"010011100",
  39941=>"000001010",
  39942=>"101001001",
  39943=>"101100100",
  39944=>"001101010",
  39945=>"010110010",
  39946=>"100101001",
  39947=>"110110001",
  39948=>"110111111",
  39949=>"110110010",
  39950=>"010011111",
  39951=>"111100110",
  39952=>"001110110",
  39953=>"001101100",
  39954=>"111110001",
  39955=>"100110000",
  39956=>"101100000",
  39957=>"010010100",
  39958=>"011101110",
  39959=>"001000001",
  39960=>"011111111",
  39961=>"010111110",
  39962=>"010111111",
  39963=>"001001000",
  39964=>"000000010",
  39965=>"001010001",
  39966=>"111010101",
  39967=>"011100100",
  39968=>"010111110",
  39969=>"101111100",
  39970=>"110001110",
  39971=>"000101110",
  39972=>"100001101",
  39973=>"111011010",
  39974=>"011100110",
  39975=>"000111000",
  39976=>"101111110",
  39977=>"001011011",
  39978=>"110011110",
  39979=>"001101100",
  39980=>"000000011",
  39981=>"101100100",
  39982=>"011100110",
  39983=>"000011000",
  39984=>"100111001",
  39985=>"110101101",
  39986=>"110011000",
  39987=>"001110101",
  39988=>"011010011",
  39989=>"100100000",
  39990=>"100000100",
  39991=>"111101000",
  39992=>"001000111",
  39993=>"110000100",
  39994=>"000100101",
  39995=>"000111110",
  39996=>"101110101",
  39997=>"100010111",
  39998=>"001011111",
  39999=>"100100010",
  40000=>"101100101",
  40001=>"101000010",
  40002=>"001010111",
  40003=>"110111001",
  40004=>"010010001",
  40005=>"011100101",
  40006=>"110000000",
  40007=>"010000001",
  40008=>"000010100",
  40009=>"101101011",
  40010=>"111111101",
  40011=>"100111001",
  40012=>"000010010",
  40013=>"001111111",
  40014=>"111011001",
  40015=>"011101111",
  40016=>"001011011",
  40017=>"111110001",
  40018=>"010111111",
  40019=>"011010111",
  40020=>"110111011",
  40021=>"001101010",
  40022=>"101110001",
  40023=>"001001101",
  40024=>"111001001",
  40025=>"101000111",
  40026=>"000100010",
  40027=>"101101110",
  40028=>"010010010",
  40029=>"100010011",
  40030=>"100101100",
  40031=>"111101010",
  40032=>"110101000",
  40033=>"110001101",
  40034=>"110111110",
  40035=>"001000010",
  40036=>"011100100",
  40037=>"110100100",
  40038=>"011010010",
  40039=>"100010101",
  40040=>"001111011",
  40041=>"101110001",
  40042=>"101100011",
  40043=>"001101001",
  40044=>"100110111",
  40045=>"111110011",
  40046=>"111000111",
  40047=>"101000001",
  40048=>"010000011",
  40049=>"011101111",
  40050=>"001110101",
  40051=>"101000000",
  40052=>"111100001",
  40053=>"010011111",
  40054=>"011001010",
  40055=>"101110010",
  40056=>"100010010",
  40057=>"111011000",
  40058=>"110100011",
  40059=>"111001100",
  40060=>"100001111",
  40061=>"111111011",
  40062=>"000000101",
  40063=>"111010111",
  40064=>"001000100",
  40065=>"001110000",
  40066=>"101001011",
  40067=>"100000110",
  40068=>"001100100",
  40069=>"100000011",
  40070=>"011101111",
  40071=>"111011000",
  40072=>"000001110",
  40073=>"101001000",
  40074=>"101100000",
  40075=>"111010011",
  40076=>"010010101",
  40077=>"101101111",
  40078=>"100101101",
  40079=>"101011010",
  40080=>"111000101",
  40081=>"110111101",
  40082=>"100011000",
  40083=>"011101011",
  40084=>"101101111",
  40085=>"110110110",
  40086=>"000001000",
  40087=>"111101111",
  40088=>"001000010",
  40089=>"100000011",
  40090=>"101101110",
  40091=>"010111001",
  40092=>"110100001",
  40093=>"001011100",
  40094=>"001101110",
  40095=>"000110011",
  40096=>"010000000",
  40097=>"001001010",
  40098=>"110010111",
  40099=>"111000010",
  40100=>"110000101",
  40101=>"111100111",
  40102=>"100100001",
  40103=>"100110010",
  40104=>"111000101",
  40105=>"010011011",
  40106=>"101110111",
  40107=>"010110110",
  40108=>"110010100",
  40109=>"000001110",
  40110=>"011111110",
  40111=>"010011100",
  40112=>"011000111",
  40113=>"101001000",
  40114=>"100001011",
  40115=>"000000011",
  40116=>"110000011",
  40117=>"110010010",
  40118=>"011100001",
  40119=>"010100101",
  40120=>"010000000",
  40121=>"110100110",
  40122=>"001100000",
  40123=>"101111100",
  40124=>"111001101",
  40125=>"111001010",
  40126=>"001111101",
  40127=>"111100000",
  40128=>"001101001",
  40129=>"001111111",
  40130=>"111100011",
  40131=>"000001001",
  40132=>"110011011",
  40133=>"010111001",
  40134=>"001101101",
  40135=>"001100011",
  40136=>"111101100",
  40137=>"110011111",
  40138=>"001010100",
  40139=>"100100110",
  40140=>"010101111",
  40141=>"000011010",
  40142=>"011011000",
  40143=>"101110001",
  40144=>"100111110",
  40145=>"110110011",
  40146=>"100101101",
  40147=>"001101111",
  40148=>"001110000",
  40149=>"010011101",
  40150=>"001101010",
  40151=>"111110101",
  40152=>"101001000",
  40153=>"101001001",
  40154=>"000010011",
  40155=>"110000011",
  40156=>"110000111",
  40157=>"000000111",
  40158=>"111010010",
  40159=>"101100001",
  40160=>"101011110",
  40161=>"011101000",
  40162=>"110110100",
  40163=>"111100100",
  40164=>"110101001",
  40165=>"110000001",
  40166=>"111110101",
  40167=>"111101011",
  40168=>"011110010",
  40169=>"001010101",
  40170=>"010000110",
  40171=>"100101001",
  40172=>"000100000",
  40173=>"010100011",
  40174=>"010000000",
  40175=>"001011110",
  40176=>"011100001",
  40177=>"101000010",
  40178=>"001000000",
  40179=>"100101000",
  40180=>"100110011",
  40181=>"100011011",
  40182=>"111001011",
  40183=>"001000000",
  40184=>"110000101",
  40185=>"001010101",
  40186=>"101111110",
  40187=>"001011010",
  40188=>"000001111",
  40189=>"001100101",
  40190=>"110100100",
  40191=>"001011101",
  40192=>"000101110",
  40193=>"110010110",
  40194=>"010011001",
  40195=>"000000101",
  40196=>"001000110",
  40197=>"101000111",
  40198=>"001100111",
  40199=>"111100001",
  40200=>"100110100",
  40201=>"011010010",
  40202=>"100000110",
  40203=>"001101011",
  40204=>"001110000",
  40205=>"110000110",
  40206=>"110010000",
  40207=>"111100101",
  40208=>"010111011",
  40209=>"011110011",
  40210=>"111110111",
  40211=>"010001010",
  40212=>"110100001",
  40213=>"000000101",
  40214=>"100101111",
  40215=>"111001100",
  40216=>"000011111",
  40217=>"000101000",
  40218=>"000011000",
  40219=>"101000101",
  40220=>"001000111",
  40221=>"101001001",
  40222=>"010111011",
  40223=>"100010000",
  40224=>"000000100",
  40225=>"100111100",
  40226=>"000001011",
  40227=>"111100101",
  40228=>"010101010",
  40229=>"100011001",
  40230=>"110000000",
  40231=>"100110000",
  40232=>"110101011",
  40233=>"110011100",
  40234=>"111000001",
  40235=>"100000011",
  40236=>"000110100",
  40237=>"101101101",
  40238=>"111001111",
  40239=>"011000111",
  40240=>"101110011",
  40241=>"010011010",
  40242=>"101111101",
  40243=>"101001001",
  40244=>"111110101",
  40245=>"001000110",
  40246=>"010011001",
  40247=>"011101100",
  40248=>"001111100",
  40249=>"001011100",
  40250=>"101000000",
  40251=>"101000100",
  40252=>"111101100",
  40253=>"101101100",
  40254=>"101011101",
  40255=>"010000000",
  40256=>"011100000",
  40257=>"110000111",
  40258=>"000010000",
  40259=>"101110101",
  40260=>"101100101",
  40261=>"011100010",
  40262=>"000001100",
  40263=>"011111001",
  40264=>"000010100",
  40265=>"000001000",
  40266=>"110000111",
  40267=>"010010000",
  40268=>"010110000",
  40269=>"010000100",
  40270=>"111101011",
  40271=>"101100000",
  40272=>"000010110",
  40273=>"100001000",
  40274=>"111001010",
  40275=>"011000011",
  40276=>"101011000",
  40277=>"000011001",
  40278=>"000111011",
  40279=>"100001100",
  40280=>"010000100",
  40281=>"000010100",
  40282=>"010101001",
  40283=>"111100001",
  40284=>"101100010",
  40285=>"101000000",
  40286=>"101010010",
  40287=>"101000000",
  40288=>"100100000",
  40289=>"111101111",
  40290=>"101010110",
  40291=>"011101001",
  40292=>"010100001",
  40293=>"010010000",
  40294=>"010111010",
  40295=>"110100010",
  40296=>"001100010",
  40297=>"100000000",
  40298=>"001001111",
  40299=>"001010011",
  40300=>"110110110",
  40301=>"010111001",
  40302=>"100101111",
  40303=>"011111100",
  40304=>"011001110",
  40305=>"000110001",
  40306=>"000100111",
  40307=>"011001011",
  40308=>"100001101",
  40309=>"001010000",
  40310=>"110111000",
  40311=>"111001111",
  40312=>"010110101",
  40313=>"110011011",
  40314=>"001010111",
  40315=>"100000000",
  40316=>"100100100",
  40317=>"100101110",
  40318=>"111100011",
  40319=>"100010010",
  40320=>"000001000",
  40321=>"001010011",
  40322=>"111100101",
  40323=>"111000101",
  40324=>"111110001",
  40325=>"101000110",
  40326=>"000100110",
  40327=>"101111001",
  40328=>"111001001",
  40329=>"000101101",
  40330=>"010010001",
  40331=>"110001101",
  40332=>"001000010",
  40333=>"110010001",
  40334=>"100101110",
  40335=>"000010010",
  40336=>"001011101",
  40337=>"111101011",
  40338=>"011011010",
  40339=>"000001000",
  40340=>"101111001",
  40341=>"100110001",
  40342=>"111111110",
  40343=>"111111110",
  40344=>"111110000",
  40345=>"001000010",
  40346=>"000011001",
  40347=>"001100010",
  40348=>"101110111",
  40349=>"111111111",
  40350=>"100111000",
  40351=>"010110101",
  40352=>"001101101",
  40353=>"001011100",
  40354=>"011010111",
  40355=>"000101010",
  40356=>"110001100",
  40357=>"011100110",
  40358=>"010011011",
  40359=>"010010100",
  40360=>"001110111",
  40361=>"001001000",
  40362=>"011101010",
  40363=>"001000110",
  40364=>"111011000",
  40365=>"111111111",
  40366=>"000111001",
  40367=>"111101000",
  40368=>"110101000",
  40369=>"000110101",
  40370=>"111101100",
  40371=>"011011111",
  40372=>"010111110",
  40373=>"110100000",
  40374=>"000101111",
  40375=>"010000010",
  40376=>"111100001",
  40377=>"010000110",
  40378=>"001010010",
  40379=>"111000101",
  40380=>"110110110",
  40381=>"100011100",
  40382=>"101011111",
  40383=>"000011101",
  40384=>"100001000",
  40385=>"101010000",
  40386=>"011001011",
  40387=>"011000101",
  40388=>"110000110",
  40389=>"000000011",
  40390=>"110001110",
  40391=>"100011010",
  40392=>"011010000",
  40393=>"101011000",
  40394=>"011000010",
  40395=>"000111101",
  40396=>"111011111",
  40397=>"100000111",
  40398=>"000010000",
  40399=>"000110110",
  40400=>"011010011",
  40401=>"111101111",
  40402=>"101101101",
  40403=>"100100001",
  40404=>"111101001",
  40405=>"000100001",
  40406=>"111001100",
  40407=>"011011101",
  40408=>"000010001",
  40409=>"110011000",
  40410=>"000000001",
  40411=>"000111000",
  40412=>"001001000",
  40413=>"001001110",
  40414=>"101100101",
  40415=>"001010000",
  40416=>"011100111",
  40417=>"100101111",
  40418=>"111111111",
  40419=>"111011011",
  40420=>"001111110",
  40421=>"001110011",
  40422=>"001100111",
  40423=>"100110000",
  40424=>"011001110",
  40425=>"101010110",
  40426=>"001100011",
  40427=>"010011010",
  40428=>"111101110",
  40429=>"101001001",
  40430=>"000010001",
  40431=>"001010001",
  40432=>"100101110",
  40433=>"011100011",
  40434=>"011000111",
  40435=>"000010111",
  40436=>"110001111",
  40437=>"100100101",
  40438=>"101011110",
  40439=>"000000000",
  40440=>"010011101",
  40441=>"010100010",
  40442=>"101110011",
  40443=>"001101001",
  40444=>"101111101",
  40445=>"010001000",
  40446=>"100011010",
  40447=>"001100111",
  40448=>"011001100",
  40449=>"010100010",
  40450=>"111001101",
  40451=>"001101101",
  40452=>"010101101",
  40453=>"010000000",
  40454=>"111101101",
  40455=>"011101110",
  40456=>"001001110",
  40457=>"011110111",
  40458=>"111011011",
  40459=>"100101000",
  40460=>"000001001",
  40461=>"111010011",
  40462=>"010101001",
  40463=>"010011001",
  40464=>"010001110",
  40465=>"110111110",
  40466=>"101100010",
  40467=>"111100110",
  40468=>"101001011",
  40469=>"110110111",
  40470=>"010110110",
  40471=>"010000001",
  40472=>"111000100",
  40473=>"011111001",
  40474=>"001101100",
  40475=>"011100100",
  40476=>"110010010",
  40477=>"010000010",
  40478=>"011010110",
  40479=>"100000110",
  40480=>"111001011",
  40481=>"101001100",
  40482=>"000001000",
  40483=>"001100101",
  40484=>"110100101",
  40485=>"100001011",
  40486=>"100110100",
  40487=>"101111100",
  40488=>"110010100",
  40489=>"001001001",
  40490=>"111110001",
  40491=>"010010101",
  40492=>"010110010",
  40493=>"000010110",
  40494=>"010000011",
  40495=>"010001011",
  40496=>"011111010",
  40497=>"111111010",
  40498=>"001001010",
  40499=>"101000010",
  40500=>"100000010",
  40501=>"110100101",
  40502=>"101100010",
  40503=>"100011101",
  40504=>"101111111",
  40505=>"111010101",
  40506=>"110010000",
  40507=>"010111001",
  40508=>"000100101",
  40509=>"000011111",
  40510=>"101101001",
  40511=>"000000000",
  40512=>"000000000",
  40513=>"010101100",
  40514=>"100111001",
  40515=>"111011010",
  40516=>"100000111",
  40517=>"001000101",
  40518=>"101111110",
  40519=>"101000110",
  40520=>"000111110",
  40521=>"111111000",
  40522=>"010000010",
  40523=>"111011110",
  40524=>"000000010",
  40525=>"101111010",
  40526=>"010011000",
  40527=>"111000010",
  40528=>"110011111",
  40529=>"010100000",
  40530=>"010001000",
  40531=>"000100001",
  40532=>"000110001",
  40533=>"001000001",
  40534=>"000001110",
  40535=>"100101111",
  40536=>"101111001",
  40537=>"100001110",
  40538=>"000000100",
  40539=>"010010100",
  40540=>"010001111",
  40541=>"000110100",
  40542=>"101101100",
  40543=>"001001111",
  40544=>"011100010",
  40545=>"001110110",
  40546=>"001111000",
  40547=>"111111111",
  40548=>"111001111",
  40549=>"001000100",
  40550=>"110111011",
  40551=>"100101001",
  40552=>"000101110",
  40553=>"100110011",
  40554=>"110010110",
  40555=>"000000111",
  40556=>"100000111",
  40557=>"100001101",
  40558=>"111000110",
  40559=>"011101101",
  40560=>"000111100",
  40561=>"000100000",
  40562=>"011111010",
  40563=>"000110100",
  40564=>"100111000",
  40565=>"010000100",
  40566=>"100110000",
  40567=>"101011010",
  40568=>"001100011",
  40569=>"111000001",
  40570=>"010011011",
  40571=>"001111000",
  40572=>"101101000",
  40573=>"101111011",
  40574=>"110101100",
  40575=>"011111100",
  40576=>"110001100",
  40577=>"000001000",
  40578=>"011111100",
  40579=>"100001011",
  40580=>"100001100",
  40581=>"110111110",
  40582=>"011100001",
  40583=>"000111101",
  40584=>"111100111",
  40585=>"000100010",
  40586=>"111011101",
  40587=>"000111010",
  40588=>"110011011",
  40589=>"001111000",
  40590=>"111010010",
  40591=>"011110100",
  40592=>"001001101",
  40593=>"001100111",
  40594=>"110100011",
  40595=>"000110001",
  40596=>"000110001",
  40597=>"100010000",
  40598=>"110001100",
  40599=>"101011100",
  40600=>"111001101",
  40601=>"110000011",
  40602=>"101000100",
  40603=>"101110101",
  40604=>"110101100",
  40605=>"100000001",
  40606=>"000010110",
  40607=>"110001011",
  40608=>"010101111",
  40609=>"010111000",
  40610=>"000111010",
  40611=>"010111101",
  40612=>"110001001",
  40613=>"001010011",
  40614=>"010000100",
  40615=>"000110011",
  40616=>"001000001",
  40617=>"001101010",
  40618=>"101101111",
  40619=>"111111010",
  40620=>"010010011",
  40621=>"111101001",
  40622=>"011101000",
  40623=>"000011101",
  40624=>"101101001",
  40625=>"000101001",
  40626=>"111010000",
  40627=>"011010100",
  40628=>"000001010",
  40629=>"101100000",
  40630=>"101010110",
  40631=>"001010110",
  40632=>"110000111",
  40633=>"001100000",
  40634=>"100001100",
  40635=>"010001010",
  40636=>"111011100",
  40637=>"011001001",
  40638=>"101000100",
  40639=>"111000001",
  40640=>"000011100",
  40641=>"100001110",
  40642=>"001010101",
  40643=>"010010011",
  40644=>"011011111",
  40645=>"000101001",
  40646=>"011110011",
  40647=>"101100001",
  40648=>"001001100",
  40649=>"011000100",
  40650=>"101000011",
  40651=>"011001000",
  40652=>"001111110",
  40653=>"100100110",
  40654=>"010010000",
  40655=>"011101110",
  40656=>"101101100",
  40657=>"101001110",
  40658=>"111000101",
  40659=>"000011001",
  40660=>"000000110",
  40661=>"001101010",
  40662=>"111111111",
  40663=>"010001000",
  40664=>"001110111",
  40665=>"001000011",
  40666=>"100000000",
  40667=>"001010000",
  40668=>"100100011",
  40669=>"010000000",
  40670=>"100000011",
  40671=>"110100110",
  40672=>"011111110",
  40673=>"001000010",
  40674=>"100111110",
  40675=>"001001010",
  40676=>"011011100",
  40677=>"100000111",
  40678=>"010110101",
  40679=>"011110010",
  40680=>"000101111",
  40681=>"100110101",
  40682=>"011110111",
  40683=>"000011000",
  40684=>"010010000",
  40685=>"100101101",
  40686=>"110111100",
  40687=>"110000000",
  40688=>"110011110",
  40689=>"010110000",
  40690=>"101111001",
  40691=>"000000101",
  40692=>"010000100",
  40693=>"110001000",
  40694=>"000000011",
  40695=>"110100110",
  40696=>"001001100",
  40697=>"011111000",
  40698=>"010001011",
  40699=>"010101011",
  40700=>"001011101",
  40701=>"011111101",
  40702=>"101101110",
  40703=>"001000001",
  40704=>"100001001",
  40705=>"001010110",
  40706=>"110100001",
  40707=>"000000101",
  40708=>"111010110",
  40709=>"000100010",
  40710=>"101011001",
  40711=>"101010010",
  40712=>"011001010",
  40713=>"011000100",
  40714=>"111001110",
  40715=>"110100000",
  40716=>"001011000",
  40717=>"101111000",
  40718=>"010111011",
  40719=>"010101111",
  40720=>"111001110",
  40721=>"101001000",
  40722=>"000000000",
  40723=>"011110011",
  40724=>"110010011",
  40725=>"111110011",
  40726=>"000111101",
  40727=>"110000011",
  40728=>"011001001",
  40729=>"010101100",
  40730=>"101000000",
  40731=>"110000100",
  40732=>"111000001",
  40733=>"111010110",
  40734=>"101111111",
  40735=>"010001001",
  40736=>"101011110",
  40737=>"110000001",
  40738=>"011110011",
  40739=>"101101110",
  40740=>"111101011",
  40741=>"111101101",
  40742=>"000011011",
  40743=>"101110011",
  40744=>"110100110",
  40745=>"100011010",
  40746=>"011001100",
  40747=>"111011100",
  40748=>"100111010",
  40749=>"110000000",
  40750=>"101010001",
  40751=>"110101100",
  40752=>"000101110",
  40753=>"111011011",
  40754=>"011011001",
  40755=>"010110001",
  40756=>"100100001",
  40757=>"011111011",
  40758=>"101110110",
  40759=>"000000011",
  40760=>"100001011",
  40761=>"001001100",
  40762=>"000011001",
  40763=>"011000010",
  40764=>"000101111",
  40765=>"010011011",
  40766=>"111100100",
  40767=>"111011110",
  40768=>"100111111",
  40769=>"101010010",
  40770=>"000011101",
  40771=>"100010000",
  40772=>"000100110",
  40773=>"111011111",
  40774=>"111011111",
  40775=>"101000010",
  40776=>"001001010",
  40777=>"000101111",
  40778=>"101000001",
  40779=>"000101001",
  40780=>"011011110",
  40781=>"101011001",
  40782=>"001110010",
  40783=>"101101010",
  40784=>"111000100",
  40785=>"000010110",
  40786=>"110110101",
  40787=>"110001000",
  40788=>"000100111",
  40789=>"000110110",
  40790=>"011101011",
  40791=>"110100010",
  40792=>"110111001",
  40793=>"001100011",
  40794=>"010001000",
  40795=>"001110100",
  40796=>"100011111",
  40797=>"100000011",
  40798=>"010101110",
  40799=>"110100000",
  40800=>"101000111",
  40801=>"111001111",
  40802=>"100010111",
  40803=>"010100110",
  40804=>"101001000",
  40805=>"111111011",
  40806=>"100100100",
  40807=>"011001011",
  40808=>"010001001",
  40809=>"010110000",
  40810=>"010010001",
  40811=>"101110101",
  40812=>"011110011",
  40813=>"001101011",
  40814=>"100000111",
  40815=>"101110011",
  40816=>"011011000",
  40817=>"011101000",
  40818=>"110011110",
  40819=>"010101111",
  40820=>"010011011",
  40821=>"010001101",
  40822=>"000001001",
  40823=>"010100110",
  40824=>"011001001",
  40825=>"110000010",
  40826=>"110111110",
  40827=>"001011101",
  40828=>"110100100",
  40829=>"101100010",
  40830=>"111000110",
  40831=>"110001111",
  40832=>"000110010",
  40833=>"101000010",
  40834=>"001001101",
  40835=>"111101100",
  40836=>"011100111",
  40837=>"010001011",
  40838=>"111101000",
  40839=>"100011101",
  40840=>"010010010",
  40841=>"000000011",
  40842=>"100011000",
  40843=>"101101111",
  40844=>"110010100",
  40845=>"110010110",
  40846=>"000110001",
  40847=>"000100101",
  40848=>"100100011",
  40849=>"011101110",
  40850=>"001011000",
  40851=>"001000100",
  40852=>"100011001",
  40853=>"000110011",
  40854=>"100010000",
  40855=>"011100100",
  40856=>"001010110",
  40857=>"011000010",
  40858=>"000111000",
  40859=>"100111011",
  40860=>"110111010",
  40861=>"000101011",
  40862=>"000010101",
  40863=>"111000111",
  40864=>"001101000",
  40865=>"101100110",
  40866=>"111101011",
  40867=>"000011100",
  40868=>"100100111",
  40869=>"110100011",
  40870=>"101100000",
  40871=>"000000010",
  40872=>"000011000",
  40873=>"110010001",
  40874=>"111110011",
  40875=>"010001100",
  40876=>"111111110",
  40877=>"101000011",
  40878=>"100100010",
  40879=>"000111000",
  40880=>"000100011",
  40881=>"011111011",
  40882=>"010111111",
  40883=>"100100010",
  40884=>"010100111",
  40885=>"010001011",
  40886=>"001111110",
  40887=>"001101101",
  40888=>"001111111",
  40889=>"101110000",
  40890=>"111011110",
  40891=>"100100110",
  40892=>"010000001",
  40893=>"001001011",
  40894=>"001000100",
  40895=>"110000001",
  40896=>"011010001",
  40897=>"100001011",
  40898=>"001101001",
  40899=>"111110110",
  40900=>"100110101",
  40901=>"111100100",
  40902=>"011111010",
  40903=>"110000010",
  40904=>"000000010",
  40905=>"000100010",
  40906=>"001110110",
  40907=>"101011110",
  40908=>"110001000",
  40909=>"101101111",
  40910=>"111111111",
  40911=>"111100101",
  40912=>"011000101",
  40913=>"110010101",
  40914=>"101111000",
  40915=>"100000000",
  40916=>"111000110",
  40917=>"000000111",
  40918=>"111000010",
  40919=>"001000111",
  40920=>"100110000",
  40921=>"100011001",
  40922=>"011101000",
  40923=>"010010110",
  40924=>"010110100",
  40925=>"000010100",
  40926=>"111011011",
  40927=>"100100100",
  40928=>"010101010",
  40929=>"001000000",
  40930=>"010101010",
  40931=>"010010110",
  40932=>"001111101",
  40933=>"011010100",
  40934=>"100011101",
  40935=>"100000011",
  40936=>"000100110",
  40937=>"011111111",
  40938=>"101100010",
  40939=>"010000111",
  40940=>"011110101",
  40941=>"001010010",
  40942=>"011000101",
  40943=>"001010101",
  40944=>"001011001",
  40945=>"001100011",
  40946=>"111001011",
  40947=>"010101100",
  40948=>"111111010",
  40949=>"100000110",
  40950=>"100101101",
  40951=>"010111000",
  40952=>"000010010",
  40953=>"010110101",
  40954=>"100000101",
  40955=>"000011011",
  40956=>"101011100",
  40957=>"010111010",
  40958=>"000111001",
  40959=>"111011110",
  40960=>"000000001",
  40961=>"111010010",
  40962=>"001111100",
  40963=>"000101101",
  40964=>"000000011",
  40965=>"111101101",
  40966=>"011101010",
  40967=>"110111100",
  40968=>"001010111",
  40969=>"111011111",
  40970=>"010111001",
  40971=>"101001101",
  40972=>"000011011",
  40973=>"110100100",
  40974=>"000001100",
  40975=>"110001000",
  40976=>"000111110",
  40977=>"100110011",
  40978=>"011001111",
  40979=>"111100010",
  40980=>"101001011",
  40981=>"101100001",
  40982=>"100010110",
  40983=>"110110110",
  40984=>"000110000",
  40985=>"110001000",
  40986=>"011001100",
  40987=>"111001101",
  40988=>"110001101",
  40989=>"010110100",
  40990=>"011111000",
  40991=>"000001100",
  40992=>"100010110",
  40993=>"000110100",
  40994=>"001001101",
  40995=>"110110010",
  40996=>"010001101",
  40997=>"101101010",
  40998=>"001000110",
  40999=>"111101000",
  41000=>"000111000",
  41001=>"111001001",
  41002=>"110110100",
  41003=>"000001000",
  41004=>"101100111",
  41005=>"010111110",
  41006=>"000011101",
  41007=>"000110011",
  41008=>"000110100",
  41009=>"001000101",
  41010=>"111101011",
  41011=>"000101000",
  41012=>"111100010",
  41013=>"011001100",
  41014=>"111000111",
  41015=>"001111010",
  41016=>"001111110",
  41017=>"010010000",
  41018=>"010010000",
  41019=>"111111111",
  41020=>"001110011",
  41021=>"000010000",
  41022=>"101000000",
  41023=>"111001101",
  41024=>"000011010",
  41025=>"000100011",
  41026=>"111111011",
  41027=>"011100001",
  41028=>"100111001",
  41029=>"110000011",
  41030=>"111101111",
  41031=>"111001000",
  41032=>"111101011",
  41033=>"011001111",
  41034=>"000100000",
  41035=>"000101000",
  41036=>"011100001",
  41037=>"111010110",
  41038=>"110101010",
  41039=>"000001001",
  41040=>"011001111",
  41041=>"100000001",
  41042=>"110001010",
  41043=>"001110101",
  41044=>"111010110",
  41045=>"000101001",
  41046=>"010111011",
  41047=>"000000110",
  41048=>"101010000",
  41049=>"111010101",
  41050=>"100100100",
  41051=>"000001000",
  41052=>"011101110",
  41053=>"000101111",
  41054=>"010110110",
  41055=>"011000010",
  41056=>"011011111",
  41057=>"000010000",
  41058=>"100001110",
  41059=>"101100111",
  41060=>"110011011",
  41061=>"011001100",
  41062=>"100110111",
  41063=>"001110100",
  41064=>"100110101",
  41065=>"110010110",
  41066=>"101100110",
  41067=>"010001100",
  41068=>"001111110",
  41069=>"001001011",
  41070=>"101111001",
  41071=>"100000111",
  41072=>"011111001",
  41073=>"001010111",
  41074=>"011101100",
  41075=>"101100100",
  41076=>"010111111",
  41077=>"111011011",
  41078=>"011011100",
  41079=>"010111111",
  41080=>"000000100",
  41081=>"011011100",
  41082=>"000000101",
  41083=>"100110010",
  41084=>"101111010",
  41085=>"011011100",
  41086=>"100000011",
  41087=>"101011000",
  41088=>"110011110",
  41089=>"000101011",
  41090=>"001001000",
  41091=>"100000001",
  41092=>"111100101",
  41093=>"000011101",
  41094=>"110111011",
  41095=>"100010110",
  41096=>"001111011",
  41097=>"101111111",
  41098=>"111101110",
  41099=>"111011101",
  41100=>"000000110",
  41101=>"011011100",
  41102=>"101100000",
  41103=>"000011110",
  41104=>"010100001",
  41105=>"000000000",
  41106=>"001010001",
  41107=>"111010100",
  41108=>"111010111",
  41109=>"000111000",
  41110=>"100000100",
  41111=>"011100111",
  41112=>"111101110",
  41113=>"000010000",
  41114=>"101110101",
  41115=>"100010001",
  41116=>"111000111",
  41117=>"010110001",
  41118=>"110000010",
  41119=>"111011101",
  41120=>"110010100",
  41121=>"011100101",
  41122=>"000111011",
  41123=>"111000110",
  41124=>"111010101",
  41125=>"011110100",
  41126=>"100011000",
  41127=>"100001100",
  41128=>"001100100",
  41129=>"000011101",
  41130=>"101100101",
  41131=>"110111110",
  41132=>"011011100",
  41133=>"000011101",
  41134=>"000011000",
  41135=>"100001101",
  41136=>"000110011",
  41137=>"110100001",
  41138=>"110000110",
  41139=>"011011011",
  41140=>"010011010",
  41141=>"010011000",
  41142=>"110101001",
  41143=>"000000111",
  41144=>"100110011",
  41145=>"101011011",
  41146=>"101010101",
  41147=>"000010110",
  41148=>"111110100",
  41149=>"011110111",
  41150=>"001001111",
  41151=>"000000010",
  41152=>"000101100",
  41153=>"110001101",
  41154=>"100101111",
  41155=>"110111001",
  41156=>"011000110",
  41157=>"011101010",
  41158=>"111001010",
  41159=>"011100111",
  41160=>"010101010",
  41161=>"001110100",
  41162=>"110010110",
  41163=>"101011101",
  41164=>"111101111",
  41165=>"101000111",
  41166=>"110001101",
  41167=>"110011001",
  41168=>"111111000",
  41169=>"111010110",
  41170=>"011001110",
  41171=>"010111000",
  41172=>"111000010",
  41173=>"110001110",
  41174=>"001101101",
  41175=>"101101000",
  41176=>"101100101",
  41177=>"001010001",
  41178=>"001111100",
  41179=>"010001000",
  41180=>"110101010",
  41181=>"001010111",
  41182=>"100110011",
  41183=>"010011111",
  41184=>"001110111",
  41185=>"010011101",
  41186=>"011110110",
  41187=>"001010001",
  41188=>"101111111",
  41189=>"110111010",
  41190=>"111110101",
  41191=>"110100111",
  41192=>"011000000",
  41193=>"101011110",
  41194=>"100001110",
  41195=>"001010011",
  41196=>"111110111",
  41197=>"110101011",
  41198=>"110101101",
  41199=>"101001000",
  41200=>"010001101",
  41201=>"001100000",
  41202=>"011100010",
  41203=>"101010011",
  41204=>"010011111",
  41205=>"001100001",
  41206=>"110001010",
  41207=>"000001001",
  41208=>"100001010",
  41209=>"000101000",
  41210=>"111010010",
  41211=>"101011000",
  41212=>"100100100",
  41213=>"000100100",
  41214=>"100000100",
  41215=>"100101110",
  41216=>"010111001",
  41217=>"000101100",
  41218=>"100111011",
  41219=>"101111000",
  41220=>"100110100",
  41221=>"101001011",
  41222=>"001110000",
  41223=>"111110000",
  41224=>"100011111",
  41225=>"101101011",
  41226=>"001000001",
  41227=>"001001101",
  41228=>"000010011",
  41229=>"000111011",
  41230=>"111000000",
  41231=>"000010000",
  41232=>"000001100",
  41233=>"011001011",
  41234=>"010100010",
  41235=>"011110011",
  41236=>"100101110",
  41237=>"011001000",
  41238=>"111111000",
  41239=>"101001010",
  41240=>"011011011",
  41241=>"000011010",
  41242=>"101010100",
  41243=>"010011000",
  41244=>"000010001",
  41245=>"000001000",
  41246=>"001010011",
  41247=>"110001010",
  41248=>"101000010",
  41249=>"111011100",
  41250=>"110101100",
  41251=>"111011000",
  41252=>"011101110",
  41253=>"100101100",
  41254=>"100110100",
  41255=>"000110100",
  41256=>"000110001",
  41257=>"100000110",
  41258=>"000001100",
  41259=>"111001010",
  41260=>"111110110",
  41261=>"111110010",
  41262=>"111001111",
  41263=>"100100110",
  41264=>"101111111",
  41265=>"010111110",
  41266=>"000011110",
  41267=>"101100000",
  41268=>"011001110",
  41269=>"001100000",
  41270=>"100011001",
  41271=>"001001011",
  41272=>"111100111",
  41273=>"110010001",
  41274=>"100101110",
  41275=>"011001100",
  41276=>"110110100",
  41277=>"000101111",
  41278=>"000010000",
  41279=>"001001001",
  41280=>"011010110",
  41281=>"111100001",
  41282=>"010001101",
  41283=>"111001000",
  41284=>"110011011",
  41285=>"010000000",
  41286=>"101110000",
  41287=>"001011000",
  41288=>"011100111",
  41289=>"110110011",
  41290=>"100001111",
  41291=>"000001010",
  41292=>"000111111",
  41293=>"100111001",
  41294=>"110000011",
  41295=>"000001001",
  41296=>"100011111",
  41297=>"011110010",
  41298=>"100110111",
  41299=>"011111011",
  41300=>"111110001",
  41301=>"111010001",
  41302=>"110010010",
  41303=>"100101010",
  41304=>"010000011",
  41305=>"001010100",
  41306=>"000100110",
  41307=>"101011111",
  41308=>"011010111",
  41309=>"010010001",
  41310=>"101111101",
  41311=>"011110110",
  41312=>"110101111",
  41313=>"100100000",
  41314=>"011101111",
  41315=>"100000000",
  41316=>"110111001",
  41317=>"001101001",
  41318=>"001101010",
  41319=>"000101111",
  41320=>"111000011",
  41321=>"001100101",
  41322=>"011011000",
  41323=>"001101111",
  41324=>"110111110",
  41325=>"110100000",
  41326=>"101100100",
  41327=>"011011100",
  41328=>"010011111",
  41329=>"100011110",
  41330=>"010000001",
  41331=>"110010000",
  41332=>"011110001",
  41333=>"111111001",
  41334=>"001101101",
  41335=>"001000000",
  41336=>"010010010",
  41337=>"110101111",
  41338=>"011100001",
  41339=>"111001010",
  41340=>"100110000",
  41341=>"000100111",
  41342=>"000110100",
  41343=>"000100100",
  41344=>"111011110",
  41345=>"001110000",
  41346=>"010101011",
  41347=>"000111100",
  41348=>"001000101",
  41349=>"001111111",
  41350=>"110001011",
  41351=>"101011100",
  41352=>"111101111",
  41353=>"011000110",
  41354=>"000100001",
  41355=>"111010001",
  41356=>"010000110",
  41357=>"110100011",
  41358=>"010011010",
  41359=>"101011110",
  41360=>"101001001",
  41361=>"100000100",
  41362=>"111100101",
  41363=>"101110010",
  41364=>"100110111",
  41365=>"111101101",
  41366=>"010000101",
  41367=>"111010000",
  41368=>"011111110",
  41369=>"010000001",
  41370=>"100111010",
  41371=>"000000000",
  41372=>"000011101",
  41373=>"110100110",
  41374=>"010110001",
  41375=>"110101001",
  41376=>"001010010",
  41377=>"011001010",
  41378=>"100110010",
  41379=>"111000010",
  41380=>"011101111",
  41381=>"001010111",
  41382=>"110111000",
  41383=>"110000110",
  41384=>"000010000",
  41385=>"101011010",
  41386=>"001100000",
  41387=>"110100111",
  41388=>"101111111",
  41389=>"101001101",
  41390=>"000101110",
  41391=>"101101111",
  41392=>"110100001",
  41393=>"001000010",
  41394=>"010000000",
  41395=>"000110001",
  41396=>"010010001",
  41397=>"011110101",
  41398=>"001011111",
  41399=>"011100100",
  41400=>"001100011",
  41401=>"010001011",
  41402=>"000100100",
  41403=>"000100001",
  41404=>"101111110",
  41405=>"101001111",
  41406=>"111101010",
  41407=>"100101010",
  41408=>"011011111",
  41409=>"101010010",
  41410=>"110011101",
  41411=>"011010101",
  41412=>"010111010",
  41413=>"110010101",
  41414=>"000001111",
  41415=>"011111010",
  41416=>"100010101",
  41417=>"010011010",
  41418=>"010111111",
  41419=>"010010000",
  41420=>"000001001",
  41421=>"010010011",
  41422=>"001101000",
  41423=>"110001000",
  41424=>"010110000",
  41425=>"111001100",
  41426=>"101100000",
  41427=>"011000110",
  41428=>"101111101",
  41429=>"101111000",
  41430=>"011100010",
  41431=>"100010111",
  41432=>"001110111",
  41433=>"011100011",
  41434=>"000010110",
  41435=>"111100100",
  41436=>"101011111",
  41437=>"011111000",
  41438=>"110111111",
  41439=>"001011000",
  41440=>"100101001",
  41441=>"101011011",
  41442=>"000100110",
  41443=>"011111111",
  41444=>"101010011",
  41445=>"010110011",
  41446=>"011101000",
  41447=>"000110100",
  41448=>"101111001",
  41449=>"111101001",
  41450=>"000000110",
  41451=>"010001000",
  41452=>"000100110",
  41453=>"100001000",
  41454=>"100101111",
  41455=>"011110011",
  41456=>"000110100",
  41457=>"111100100",
  41458=>"101111000",
  41459=>"101000001",
  41460=>"101100111",
  41461=>"111001011",
  41462=>"101101111",
  41463=>"010011011",
  41464=>"010000001",
  41465=>"000110000",
  41466=>"011101010",
  41467=>"110000111",
  41468=>"001010101",
  41469=>"100010001",
  41470=>"000101110",
  41471=>"110110001",
  41472=>"011010100",
  41473=>"100001100",
  41474=>"111111000",
  41475=>"011110000",
  41476=>"110110001",
  41477=>"111000010",
  41478=>"110111011",
  41479=>"101110111",
  41480=>"010011010",
  41481=>"110000011",
  41482=>"001111111",
  41483=>"100101101",
  41484=>"111000000",
  41485=>"010000110",
  41486=>"001110110",
  41487=>"100101010",
  41488=>"010100010",
  41489=>"110010110",
  41490=>"010101110",
  41491=>"101111011",
  41492=>"000001001",
  41493=>"100001010",
  41494=>"110110111",
  41495=>"101100001",
  41496=>"100000101",
  41497=>"111100110",
  41498=>"100000000",
  41499=>"100010111",
  41500=>"101110010",
  41501=>"110010001",
  41502=>"101100110",
  41503=>"000101011",
  41504=>"100100101",
  41505=>"011000001",
  41506=>"000000101",
  41507=>"110001100",
  41508=>"010100101",
  41509=>"001110011",
  41510=>"111011111",
  41511=>"111001101",
  41512=>"010101100",
  41513=>"100001101",
  41514=>"000000100",
  41515=>"010010010",
  41516=>"001100100",
  41517=>"101011111",
  41518=>"010010101",
  41519=>"101110011",
  41520=>"010111000",
  41521=>"010011000",
  41522=>"011011001",
  41523=>"000110101",
  41524=>"111111011",
  41525=>"101000110",
  41526=>"010001101",
  41527=>"110111111",
  41528=>"011101101",
  41529=>"100010011",
  41530=>"111011110",
  41531=>"001000101",
  41532=>"100000111",
  41533=>"001010100",
  41534=>"111101100",
  41535=>"000001000",
  41536=>"010110100",
  41537=>"001110011",
  41538=>"011000100",
  41539=>"001100100",
  41540=>"000101010",
  41541=>"100001111",
  41542=>"100010011",
  41543=>"110110011",
  41544=>"101001010",
  41545=>"001010010",
  41546=>"111010000",
  41547=>"010110011",
  41548=>"100110100",
  41549=>"100010100",
  41550=>"101010011",
  41551=>"011111011",
  41552=>"001100100",
  41553=>"111011111",
  41554=>"011100001",
  41555=>"001111100",
  41556=>"010000100",
  41557=>"000100100",
  41558=>"001001100",
  41559=>"000110101",
  41560=>"010111111",
  41561=>"111010111",
  41562=>"100011101",
  41563=>"111111000",
  41564=>"010011010",
  41565=>"010010110",
  41566=>"111010111",
  41567=>"011011111",
  41568=>"101100011",
  41569=>"001010000",
  41570=>"011001000",
  41571=>"000110011",
  41572=>"110100010",
  41573=>"101110011",
  41574=>"111010011",
  41575=>"100010110",
  41576=>"010100100",
  41577=>"011101100",
  41578=>"110000110",
  41579=>"010010111",
  41580=>"010111110",
  41581=>"010101110",
  41582=>"000011101",
  41583=>"001010000",
  41584=>"111110010",
  41585=>"010011111",
  41586=>"010010110",
  41587=>"110011111",
  41588=>"011000110",
  41589=>"100001111",
  41590=>"000000000",
  41591=>"111001011",
  41592=>"100110001",
  41593=>"000101000",
  41594=>"011001000",
  41595=>"111000000",
  41596=>"111111000",
  41597=>"001010000",
  41598=>"011000011",
  41599=>"100101100",
  41600=>"011011101",
  41601=>"110011001",
  41602=>"011010111",
  41603=>"100001111",
  41604=>"110111111",
  41605=>"000100100",
  41606=>"110111010",
  41607=>"111010001",
  41608=>"011010111",
  41609=>"001110011",
  41610=>"101111010",
  41611=>"100111111",
  41612=>"110011001",
  41613=>"000001010",
  41614=>"111010011",
  41615=>"000110101",
  41616=>"000111001",
  41617=>"100000001",
  41618=>"010111000",
  41619=>"100011110",
  41620=>"010111000",
  41621=>"001001100",
  41622=>"111100011",
  41623=>"100010100",
  41624=>"100110111",
  41625=>"111101111",
  41626=>"101001100",
  41627=>"111100001",
  41628=>"111111101",
  41629=>"010100000",
  41630=>"001010011",
  41631=>"010100100",
  41632=>"001100010",
  41633=>"001101111",
  41634=>"011111110",
  41635=>"101010101",
  41636=>"101111111",
  41637=>"100110001",
  41638=>"111110011",
  41639=>"100001000",
  41640=>"110100000",
  41641=>"110101000",
  41642=>"101100110",
  41643=>"010110001",
  41644=>"100110001",
  41645=>"100001101",
  41646=>"000001000",
  41647=>"100010111",
  41648=>"111000111",
  41649=>"110010001",
  41650=>"010111111",
  41651=>"110100101",
  41652=>"010100101",
  41653=>"111111010",
  41654=>"110001101",
  41655=>"110011100",
  41656=>"110110101",
  41657=>"000001110",
  41658=>"000011000",
  41659=>"000010111",
  41660=>"100111001",
  41661=>"010011110",
  41662=>"101000110",
  41663=>"001100011",
  41664=>"111110000",
  41665=>"000110101",
  41666=>"010111011",
  41667=>"100000111",
  41668=>"000100010",
  41669=>"100010110",
  41670=>"010100000",
  41671=>"000010111",
  41672=>"100011001",
  41673=>"000010111",
  41674=>"110000100",
  41675=>"110010001",
  41676=>"010111000",
  41677=>"001101101",
  41678=>"010001111",
  41679=>"101111011",
  41680=>"111100100",
  41681=>"100000101",
  41682=>"011000101",
  41683=>"001101101",
  41684=>"111011001",
  41685=>"111101000",
  41686=>"000001001",
  41687=>"101001000",
  41688=>"010100000",
  41689=>"111101000",
  41690=>"011101111",
  41691=>"110111110",
  41692=>"101000001",
  41693=>"100001001",
  41694=>"010110010",
  41695=>"111011101",
  41696=>"101010101",
  41697=>"100110011",
  41698=>"011011011",
  41699=>"011001011",
  41700=>"001000010",
  41701=>"001111110",
  41702=>"001000100",
  41703=>"101010111",
  41704=>"000001000",
  41705=>"110110111",
  41706=>"101011000",
  41707=>"100000111",
  41708=>"011011100",
  41709=>"111010110",
  41710=>"110000001",
  41711=>"000010011",
  41712=>"110100100",
  41713=>"011011010",
  41714=>"111101010",
  41715=>"010001111",
  41716=>"100100101",
  41717=>"110110101",
  41718=>"100111010",
  41719=>"101001000",
  41720=>"111011000",
  41721=>"000111000",
  41722=>"111000111",
  41723=>"101011110",
  41724=>"101111010",
  41725=>"111110111",
  41726=>"010110000",
  41727=>"001110001",
  41728=>"000100101",
  41729=>"011101011",
  41730=>"001010001",
  41731=>"000011100",
  41732=>"110100110",
  41733=>"010000010",
  41734=>"100001110",
  41735=>"000010101",
  41736=>"001111101",
  41737=>"011001000",
  41738=>"011001111",
  41739=>"010100110",
  41740=>"010000100",
  41741=>"111111101",
  41742=>"011101001",
  41743=>"110110010",
  41744=>"011100100",
  41745=>"010000000",
  41746=>"101000100",
  41747=>"110000111",
  41748=>"110001100",
  41749=>"010100011",
  41750=>"101000111",
  41751=>"010010000",
  41752=>"011000111",
  41753=>"010011010",
  41754=>"100010100",
  41755=>"101001111",
  41756=>"100010001",
  41757=>"011010101",
  41758=>"111010111",
  41759=>"001001011",
  41760=>"100100011",
  41761=>"000001001",
  41762=>"001010110",
  41763=>"001010000",
  41764=>"011001010",
  41765=>"010001111",
  41766=>"100011010",
  41767=>"011011001",
  41768=>"000010110",
  41769=>"110111110",
  41770=>"100010000",
  41771=>"000011001",
  41772=>"011100101",
  41773=>"000001110",
  41774=>"011100011",
  41775=>"010101001",
  41776=>"010001110",
  41777=>"111011010",
  41778=>"000010001",
  41779=>"010100001",
  41780=>"110011011",
  41781=>"110111000",
  41782=>"000110010",
  41783=>"111001110",
  41784=>"111101101",
  41785=>"101000110",
  41786=>"011001010",
  41787=>"111011000",
  41788=>"100111100",
  41789=>"011010000",
  41790=>"100101010",
  41791=>"001011100",
  41792=>"101101111",
  41793=>"111000000",
  41794=>"111001111",
  41795=>"000101110",
  41796=>"011100011",
  41797=>"100100100",
  41798=>"101100000",
  41799=>"110001110",
  41800=>"000100000",
  41801=>"011111100",
  41802=>"110010010",
  41803=>"000000000",
  41804=>"111111000",
  41805=>"011000011",
  41806=>"110001000",
  41807=>"110101010",
  41808=>"101001100",
  41809=>"111111011",
  41810=>"110111110",
  41811=>"111010111",
  41812=>"110110111",
  41813=>"011101000",
  41814=>"101111111",
  41815=>"010000011",
  41816=>"100001000",
  41817=>"100000101",
  41818=>"001100101",
  41819=>"110110011",
  41820=>"001110100",
  41821=>"111111001",
  41822=>"110001100",
  41823=>"010000000",
  41824=>"100011111",
  41825=>"000001110",
  41826=>"101000010",
  41827=>"011111111",
  41828=>"110101011",
  41829=>"011101001",
  41830=>"011101010",
  41831=>"011101101",
  41832=>"000101110",
  41833=>"001000110",
  41834=>"001010001",
  41835=>"011011110",
  41836=>"000100011",
  41837=>"000011000",
  41838=>"111111001",
  41839=>"000011011",
  41840=>"010101011",
  41841=>"001111011",
  41842=>"111000110",
  41843=>"001011011",
  41844=>"011101101",
  41845=>"011100111",
  41846=>"101101011",
  41847=>"100110000",
  41848=>"101101101",
  41849=>"010001000",
  41850=>"001101000",
  41851=>"011001000",
  41852=>"000101010",
  41853=>"110001110",
  41854=>"111000111",
  41855=>"101111010",
  41856=>"011011111",
  41857=>"000100000",
  41858=>"100011110",
  41859=>"101000111",
  41860=>"001110000",
  41861=>"101010010",
  41862=>"110010110",
  41863=>"011010101",
  41864=>"010001000",
  41865=>"000100111",
  41866=>"100011001",
  41867=>"100101010",
  41868=>"101110011",
  41869=>"000101011",
  41870=>"001111001",
  41871=>"101011110",
  41872=>"110101101",
  41873=>"111111010",
  41874=>"000001010",
  41875=>"000100111",
  41876=>"000001110",
  41877=>"111101001",
  41878=>"110011111",
  41879=>"111000111",
  41880=>"100010110",
  41881=>"100101111",
  41882=>"001000110",
  41883=>"101000001",
  41884=>"001011111",
  41885=>"000011111",
  41886=>"010100010",
  41887=>"011011111",
  41888=>"000010100",
  41889=>"000011000",
  41890=>"101011000",
  41891=>"001110000",
  41892=>"110111001",
  41893=>"110001101",
  41894=>"100101101",
  41895=>"010011001",
  41896=>"101100110",
  41897=>"111111111",
  41898=>"000101100",
  41899=>"011000101",
  41900=>"010001110",
  41901=>"000000011",
  41902=>"111000101",
  41903=>"001101111",
  41904=>"100100000",
  41905=>"010001111",
  41906=>"110000001",
  41907=>"100110001",
  41908=>"100010111",
  41909=>"010111010",
  41910=>"101001110",
  41911=>"111101101",
  41912=>"111111110",
  41913=>"111100000",
  41914=>"101101011",
  41915=>"010010101",
  41916=>"111111101",
  41917=>"111100000",
  41918=>"011101001",
  41919=>"000011100",
  41920=>"011110100",
  41921=>"010110110",
  41922=>"100010111",
  41923=>"110100001",
  41924=>"001101010",
  41925=>"110110011",
  41926=>"011000101",
  41927=>"111000001",
  41928=>"100010110",
  41929=>"110001011",
  41930=>"101011011",
  41931=>"100000100",
  41932=>"011011001",
  41933=>"000110100",
  41934=>"001010000",
  41935=>"111010011",
  41936=>"110100010",
  41937=>"000010000",
  41938=>"111110011",
  41939=>"011011001",
  41940=>"000011100",
  41941=>"000100011",
  41942=>"010011000",
  41943=>"111010001",
  41944=>"101011111",
  41945=>"110101111",
  41946=>"101010110",
  41947=>"111100110",
  41948=>"011111101",
  41949=>"011001011",
  41950=>"010101100",
  41951=>"010001100",
  41952=>"110111010",
  41953=>"100111100",
  41954=>"100000000",
  41955=>"110010001",
  41956=>"011011100",
  41957=>"001001000",
  41958=>"010011010",
  41959=>"110101111",
  41960=>"001100110",
  41961=>"001110100",
  41962=>"101000000",
  41963=>"010110111",
  41964=>"101001111",
  41965=>"001000101",
  41966=>"011100010",
  41967=>"000001011",
  41968=>"001000000",
  41969=>"000011100",
  41970=>"001010001",
  41971=>"010010111",
  41972=>"110000001",
  41973=>"000000000",
  41974=>"101000100",
  41975=>"011111001",
  41976=>"111000110",
  41977=>"111011011",
  41978=>"110110011",
  41979=>"110101101",
  41980=>"010110001",
  41981=>"001010000",
  41982=>"111011001",
  41983=>"010101011",
  41984=>"001111111",
  41985=>"100100011",
  41986=>"100001100",
  41987=>"100001001",
  41988=>"111101100",
  41989=>"101101101",
  41990=>"110110111",
  41991=>"000001110",
  41992=>"110111110",
  41993=>"000010000",
  41994=>"000001011",
  41995=>"001111101",
  41996=>"110111011",
  41997=>"011010100",
  41998=>"001001111",
  41999=>"011101010",
  42000=>"111101111",
  42001=>"101010111",
  42002=>"110111011",
  42003=>"101111111",
  42004=>"101100110",
  42005=>"100000110",
  42006=>"000000001",
  42007=>"100101111",
  42008=>"100111000",
  42009=>"111101111",
  42010=>"110111111",
  42011=>"001011111",
  42012=>"000001000",
  42013=>"011001000",
  42014=>"010100010",
  42015=>"001001010",
  42016=>"011000000",
  42017=>"110011010",
  42018=>"111100100",
  42019=>"101001111",
  42020=>"010011011",
  42021=>"000110110",
  42022=>"101010011",
  42023=>"000000011",
  42024=>"010100010",
  42025=>"001001111",
  42026=>"110001110",
  42027=>"111101110",
  42028=>"101110010",
  42029=>"011100101",
  42030=>"101101111",
  42031=>"111111111",
  42032=>"010110100",
  42033=>"100110010",
  42034=>"001110000",
  42035=>"011101101",
  42036=>"011110100",
  42037=>"101010010",
  42038=>"100000011",
  42039=>"100011011",
  42040=>"111101000",
  42041=>"110110010",
  42042=>"111010001",
  42043=>"111110101",
  42044=>"010100111",
  42045=>"010000001",
  42046=>"111010011",
  42047=>"000111011",
  42048=>"010100111",
  42049=>"000111001",
  42050=>"001011011",
  42051=>"110111110",
  42052=>"100111001",
  42053=>"001111111",
  42054=>"100000110",
  42055=>"001100011",
  42056=>"011010111",
  42057=>"101001111",
  42058=>"101111110",
  42059=>"101101101",
  42060=>"111100111",
  42061=>"100110001",
  42062=>"001010000",
  42063=>"010110101",
  42064=>"010101111",
  42065=>"000100111",
  42066=>"010111010",
  42067=>"001110000",
  42068=>"101010110",
  42069=>"100110000",
  42070=>"100011010",
  42071=>"111010010",
  42072=>"101001000",
  42073=>"101001111",
  42074=>"010100110",
  42075=>"101001001",
  42076=>"111010010",
  42077=>"111011011",
  42078=>"000011111",
  42079=>"000011011",
  42080=>"011111110",
  42081=>"011101011",
  42082=>"000110000",
  42083=>"010100011",
  42084=>"000010111",
  42085=>"100001100",
  42086=>"001110101",
  42087=>"110110111",
  42088=>"010001101",
  42089=>"110001001",
  42090=>"110011001",
  42091=>"101000111",
  42092=>"101101111",
  42093=>"011101001",
  42094=>"010101110",
  42095=>"101010111",
  42096=>"000011110",
  42097=>"111010111",
  42098=>"000001011",
  42099=>"000111010",
  42100=>"010011001",
  42101=>"101011110",
  42102=>"001010111",
  42103=>"010000111",
  42104=>"110000011",
  42105=>"011001001",
  42106=>"000010101",
  42107=>"100101110",
  42108=>"100101001",
  42109=>"001110000",
  42110=>"100000011",
  42111=>"110011011",
  42112=>"111110100",
  42113=>"000000001",
  42114=>"101000100",
  42115=>"001100111",
  42116=>"000000111",
  42117=>"001010101",
  42118=>"011101001",
  42119=>"101100011",
  42120=>"110110010",
  42121=>"010000000",
  42122=>"110111111",
  42123=>"111010101",
  42124=>"111111101",
  42125=>"001000110",
  42126=>"111101011",
  42127=>"011000100",
  42128=>"000001111",
  42129=>"101011101",
  42130=>"000101100",
  42131=>"100011101",
  42132=>"000111111",
  42133=>"000100001",
  42134=>"011010101",
  42135=>"100111110",
  42136=>"011100000",
  42137=>"101001011",
  42138=>"010001011",
  42139=>"100000010",
  42140=>"100110010",
  42141=>"010001000",
  42142=>"101101111",
  42143=>"111101111",
  42144=>"000110101",
  42145=>"101101011",
  42146=>"000101111",
  42147=>"011010111",
  42148=>"101001101",
  42149=>"111111100",
  42150=>"110101001",
  42151=>"110011100",
  42152=>"010011111",
  42153=>"110101110",
  42154=>"111101001",
  42155=>"101101110",
  42156=>"001000110",
  42157=>"110111010",
  42158=>"001111010",
  42159=>"011001001",
  42160=>"111001010",
  42161=>"000100011",
  42162=>"001000010",
  42163=>"111110111",
  42164=>"110010010",
  42165=>"010010101",
  42166=>"010000101",
  42167=>"000000100",
  42168=>"111011101",
  42169=>"111010000",
  42170=>"101110001",
  42171=>"010111000",
  42172=>"001111100",
  42173=>"001001011",
  42174=>"010000110",
  42175=>"010000110",
  42176=>"011110001",
  42177=>"000100000",
  42178=>"010100100",
  42179=>"000111101",
  42180=>"111100000",
  42181=>"001111011",
  42182=>"010001001",
  42183=>"010111000",
  42184=>"100000000",
  42185=>"100111001",
  42186=>"111110111",
  42187=>"000100101",
  42188=>"011100011",
  42189=>"011101100",
  42190=>"110110101",
  42191=>"011100111",
  42192=>"100100101",
  42193=>"011101000",
  42194=>"111100100",
  42195=>"011100000",
  42196=>"000011010",
  42197=>"110100101",
  42198=>"011000001",
  42199=>"001011101",
  42200=>"100010000",
  42201=>"100010111",
  42202=>"001010110",
  42203=>"110001101",
  42204=>"110010110",
  42205=>"011110010",
  42206=>"110000000",
  42207=>"000101111",
  42208=>"001101000",
  42209=>"111111010",
  42210=>"001000010",
  42211=>"111010111",
  42212=>"010100011",
  42213=>"011011111",
  42214=>"000111111",
  42215=>"111011111",
  42216=>"110110000",
  42217=>"001001000",
  42218=>"011101111",
  42219=>"110111000",
  42220=>"111101011",
  42221=>"100001000",
  42222=>"111001000",
  42223=>"011111000",
  42224=>"010100100",
  42225=>"111000001",
  42226=>"010011110",
  42227=>"001101110",
  42228=>"111000100",
  42229=>"001000000",
  42230=>"010100000",
  42231=>"010010101",
  42232=>"010101011",
  42233=>"100000101",
  42234=>"011110010",
  42235=>"010000111",
  42236=>"101001001",
  42237=>"000100011",
  42238=>"111111111",
  42239=>"111001101",
  42240=>"100010010",
  42241=>"011111000",
  42242=>"000000100",
  42243=>"010101011",
  42244=>"000000001",
  42245=>"010001101",
  42246=>"110101110",
  42247=>"000100000",
  42248=>"110010100",
  42249=>"010111000",
  42250=>"110010010",
  42251=>"101111011",
  42252=>"011111110",
  42253=>"110110110",
  42254=>"101111100",
  42255=>"111111101",
  42256=>"111001010",
  42257=>"110100001",
  42258=>"010101111",
  42259=>"111101101",
  42260=>"111000011",
  42261=>"101101001",
  42262=>"111111111",
  42263=>"010111101",
  42264=>"011011101",
  42265=>"111011010",
  42266=>"101101001",
  42267=>"101100010",
  42268=>"010100110",
  42269=>"110001000",
  42270=>"110001000",
  42271=>"111011111",
  42272=>"111011100",
  42273=>"001001110",
  42274=>"000000001",
  42275=>"110111111",
  42276=>"001111111",
  42277=>"001001111",
  42278=>"011011010",
  42279=>"001100000",
  42280=>"110010110",
  42281=>"000111101",
  42282=>"000000001",
  42283=>"011100000",
  42284=>"001110111",
  42285=>"110010111",
  42286=>"111001001",
  42287=>"000101000",
  42288=>"010111111",
  42289=>"101010001",
  42290=>"001011000",
  42291=>"110110101",
  42292=>"000100110",
  42293=>"110001101",
  42294=>"110110011",
  42295=>"011110011",
  42296=>"111011111",
  42297=>"011000000",
  42298=>"110111011",
  42299=>"010010111",
  42300=>"000111100",
  42301=>"011000111",
  42302=>"110000110",
  42303=>"010011100",
  42304=>"111101110",
  42305=>"111111000",
  42306=>"101100000",
  42307=>"110000000",
  42308=>"110111101",
  42309=>"101011010",
  42310=>"110111111",
  42311=>"000110111",
  42312=>"111100110",
  42313=>"110001111",
  42314=>"010010000",
  42315=>"000011110",
  42316=>"001001011",
  42317=>"011110010",
  42318=>"101010000",
  42319=>"110010110",
  42320=>"110001010",
  42321=>"110010110",
  42322=>"111110111",
  42323=>"110001111",
  42324=>"000110101",
  42325=>"001001010",
  42326=>"000010101",
  42327=>"011111001",
  42328=>"111001001",
  42329=>"111011001",
  42330=>"001011110",
  42331=>"010000111",
  42332=>"110001100",
  42333=>"011001101",
  42334=>"111101001",
  42335=>"110001110",
  42336=>"011100100",
  42337=>"100110111",
  42338=>"001001111",
  42339=>"100101001",
  42340=>"000000001",
  42341=>"111010011",
  42342=>"100010000",
  42343=>"101111110",
  42344=>"001010111",
  42345=>"110011110",
  42346=>"010010111",
  42347=>"111000001",
  42348=>"000010100",
  42349=>"011101011",
  42350=>"101101111",
  42351=>"110000100",
  42352=>"000010011",
  42353=>"010001001",
  42354=>"110000111",
  42355=>"101111011",
  42356=>"100011010",
  42357=>"110111001",
  42358=>"010110100",
  42359=>"111000001",
  42360=>"111100010",
  42361=>"010101110",
  42362=>"010001100",
  42363=>"010111011",
  42364=>"110110000",
  42365=>"000101100",
  42366=>"100001111",
  42367=>"100101001",
  42368=>"110001111",
  42369=>"111111110",
  42370=>"010110100",
  42371=>"111110101",
  42372=>"000010111",
  42373=>"101111100",
  42374=>"001111000",
  42375=>"101010110",
  42376=>"000100011",
  42377=>"111111111",
  42378=>"111101011",
  42379=>"100100101",
  42380=>"011101000",
  42381=>"001101101",
  42382=>"100001000",
  42383=>"111001110",
  42384=>"100001111",
  42385=>"000111111",
  42386=>"101111101",
  42387=>"011001101",
  42388=>"001100011",
  42389=>"111001001",
  42390=>"111101011",
  42391=>"111110011",
  42392=>"010000110",
  42393=>"111111100",
  42394=>"000000000",
  42395=>"010100101",
  42396=>"100010101",
  42397=>"001110010",
  42398=>"111011001",
  42399=>"010111010",
  42400=>"000001101",
  42401=>"000101111",
  42402=>"011010011",
  42403=>"111100100",
  42404=>"000001010",
  42405=>"000101001",
  42406=>"110110000",
  42407=>"001011111",
  42408=>"101111111",
  42409=>"111100110",
  42410=>"101001110",
  42411=>"000010110",
  42412=>"111111111",
  42413=>"001000101",
  42414=>"111001001",
  42415=>"110100100",
  42416=>"101011110",
  42417=>"000000000",
  42418=>"000011111",
  42419=>"001111101",
  42420=>"010001101",
  42421=>"111000010",
  42422=>"111000111",
  42423=>"000010000",
  42424=>"111100011",
  42425=>"000111100",
  42426=>"110111100",
  42427=>"100010110",
  42428=>"001111101",
  42429=>"001111100",
  42430=>"101101011",
  42431=>"011110110",
  42432=>"111101111",
  42433=>"011100000",
  42434=>"010000000",
  42435=>"010000001",
  42436=>"010001000",
  42437=>"011100101",
  42438=>"001011100",
  42439=>"001010111",
  42440=>"001001111",
  42441=>"010011101",
  42442=>"010101000",
  42443=>"110000111",
  42444=>"011111100",
  42445=>"110010110",
  42446=>"011110000",
  42447=>"111010010",
  42448=>"110100111",
  42449=>"100010111",
  42450=>"100000100",
  42451=>"011000011",
  42452=>"010011011",
  42453=>"101110110",
  42454=>"111010111",
  42455=>"000011100",
  42456=>"101111101",
  42457=>"101101101",
  42458=>"010101101",
  42459=>"001110101",
  42460=>"110000101",
  42461=>"001101011",
  42462=>"110000001",
  42463=>"010011110",
  42464=>"101111001",
  42465=>"101000011",
  42466=>"101001110",
  42467=>"100100111",
  42468=>"010000111",
  42469=>"001000011",
  42470=>"100010011",
  42471=>"000000101",
  42472=>"011010000",
  42473=>"000100000",
  42474=>"111011100",
  42475=>"001100100",
  42476=>"100011010",
  42477=>"111101001",
  42478=>"000011001",
  42479=>"010011001",
  42480=>"100001111",
  42481=>"101111100",
  42482=>"000000100",
  42483=>"010010111",
  42484=>"000001000",
  42485=>"011101010",
  42486=>"001111100",
  42487=>"010111111",
  42488=>"100111001",
  42489=>"100011101",
  42490=>"000101100",
  42491=>"010110101",
  42492=>"111010110",
  42493=>"101011100",
  42494=>"010101111",
  42495=>"100110111",
  42496=>"001000110",
  42497=>"101011011",
  42498=>"100000100",
  42499=>"010011100",
  42500=>"011010110",
  42501=>"001111111",
  42502=>"000100001",
  42503=>"001001001",
  42504=>"000010001",
  42505=>"100010001",
  42506=>"010000000",
  42507=>"011111101",
  42508=>"100100001",
  42509=>"010001001",
  42510=>"111101101",
  42511=>"010011001",
  42512=>"000001011",
  42513=>"010111010",
  42514=>"010100001",
  42515=>"110101101",
  42516=>"110100101",
  42517=>"100110010",
  42518=>"111000111",
  42519=>"011000111",
  42520=>"111100001",
  42521=>"000100110",
  42522=>"000111111",
  42523=>"111010100",
  42524=>"011010110",
  42525=>"101011100",
  42526=>"111101100",
  42527=>"011101010",
  42528=>"000101101",
  42529=>"011110010",
  42530=>"100010101",
  42531=>"001110110",
  42532=>"000110000",
  42533=>"000101000",
  42534=>"000010000",
  42535=>"000011110",
  42536=>"010001100",
  42537=>"000001100",
  42538=>"001110101",
  42539=>"000000100",
  42540=>"101100011",
  42541=>"001110100",
  42542=>"110000101",
  42543=>"100010001",
  42544=>"000101000",
  42545=>"111101010",
  42546=>"100100011",
  42547=>"111011111",
  42548=>"100111010",
  42549=>"100001101",
  42550=>"100010010",
  42551=>"111100110",
  42552=>"111110010",
  42553=>"000110100",
  42554=>"101011101",
  42555=>"100110100",
  42556=>"111011111",
  42557=>"001001101",
  42558=>"101101101",
  42559=>"111011100",
  42560=>"011011111",
  42561=>"010000000",
  42562=>"010110100",
  42563=>"010001111",
  42564=>"100110101",
  42565=>"101111000",
  42566=>"101101010",
  42567=>"011101111",
  42568=>"100011110",
  42569=>"110000011",
  42570=>"111100111",
  42571=>"100111110",
  42572=>"011000011",
  42573=>"111111011",
  42574=>"100010000",
  42575=>"010101100",
  42576=>"100000111",
  42577=>"010101011",
  42578=>"011101101",
  42579=>"011100111",
  42580=>"101110010",
  42581=>"111111001",
  42582=>"011111111",
  42583=>"000111111",
  42584=>"101110101",
  42585=>"001100100",
  42586=>"101110111",
  42587=>"101111110",
  42588=>"011011010",
  42589=>"001011011",
  42590=>"111010110",
  42591=>"011110001",
  42592=>"000110110",
  42593=>"001111010",
  42594=>"111101101",
  42595=>"111101010",
  42596=>"001101110",
  42597=>"001001010",
  42598=>"100101001",
  42599=>"001111001",
  42600=>"111011111",
  42601=>"101101110",
  42602=>"000000101",
  42603=>"001101111",
  42604=>"111111001",
  42605=>"001011110",
  42606=>"101001000",
  42607=>"001100001",
  42608=>"110111110",
  42609=>"100101011",
  42610=>"010000011",
  42611=>"011010101",
  42612=>"001110000",
  42613=>"110010010",
  42614=>"101001000",
  42615=>"000000000",
  42616=>"110000011",
  42617=>"101110100",
  42618=>"001111000",
  42619=>"011000111",
  42620=>"000010010",
  42621=>"000110010",
  42622=>"100001101",
  42623=>"000111011",
  42624=>"110101101",
  42625=>"010000110",
  42626=>"101010011",
  42627=>"000100010",
  42628=>"001110001",
  42629=>"010111011",
  42630=>"000100010",
  42631=>"011111111",
  42632=>"110001110",
  42633=>"010001111",
  42634=>"100110100",
  42635=>"011001000",
  42636=>"011101001",
  42637=>"011111010",
  42638=>"010001010",
  42639=>"011000011",
  42640=>"011000101",
  42641=>"000110101",
  42642=>"000011000",
  42643=>"101001100",
  42644=>"101101100",
  42645=>"000011001",
  42646=>"111100001",
  42647=>"000111011",
  42648=>"111010001",
  42649=>"010101101",
  42650=>"010100010",
  42651=>"010011111",
  42652=>"001011111",
  42653=>"000000100",
  42654=>"110010101",
  42655=>"010101101",
  42656=>"010111110",
  42657=>"101001000",
  42658=>"000000000",
  42659=>"011111110",
  42660=>"000101000",
  42661=>"101101000",
  42662=>"000010100",
  42663=>"111111011",
  42664=>"011011100",
  42665=>"111100000",
  42666=>"101111000",
  42667=>"010110011",
  42668=>"001001001",
  42669=>"010100001",
  42670=>"000111000",
  42671=>"000101011",
  42672=>"100111100",
  42673=>"100111110",
  42674=>"010101111",
  42675=>"001000111",
  42676=>"001101111",
  42677=>"011011101",
  42678=>"100100111",
  42679=>"100001011",
  42680=>"001010110",
  42681=>"001101110",
  42682=>"011111000",
  42683=>"100101100",
  42684=>"011001111",
  42685=>"011001100",
  42686=>"000010111",
  42687=>"010010010",
  42688=>"101111111",
  42689=>"011101100",
  42690=>"110111110",
  42691=>"100111110",
  42692=>"111010100",
  42693=>"111001100",
  42694=>"110100000",
  42695=>"100101010",
  42696=>"010110111",
  42697=>"001110111",
  42698=>"111111100",
  42699=>"011101000",
  42700=>"000001110",
  42701=>"010000111",
  42702=>"011001001",
  42703=>"110100101",
  42704=>"000100011",
  42705=>"001101111",
  42706=>"110111100",
  42707=>"110100011",
  42708=>"111000000",
  42709=>"111111110",
  42710=>"110110000",
  42711=>"101111101",
  42712=>"010101010",
  42713=>"010111101",
  42714=>"101111111",
  42715=>"111110111",
  42716=>"101010011",
  42717=>"001100100",
  42718=>"111010100",
  42719=>"011100000",
  42720=>"010001101",
  42721=>"010011110",
  42722=>"010000011",
  42723=>"011101001",
  42724=>"101101111",
  42725=>"100000110",
  42726=>"110101000",
  42727=>"000101101",
  42728=>"001011100",
  42729=>"111011011",
  42730=>"001000100",
  42731=>"100110010",
  42732=>"110100111",
  42733=>"011001110",
  42734=>"111001111",
  42735=>"101010010",
  42736=>"000001100",
  42737=>"111111111",
  42738=>"001001101",
  42739=>"010101100",
  42740=>"111110001",
  42741=>"010101101",
  42742=>"001011001",
  42743=>"000110011",
  42744=>"110001110",
  42745=>"011010111",
  42746=>"000000011",
  42747=>"100010010",
  42748=>"000011010",
  42749=>"011000010",
  42750=>"100010111",
  42751=>"110001111",
  42752=>"000010010",
  42753=>"001110100",
  42754=>"010110010",
  42755=>"011100011",
  42756=>"001001001",
  42757=>"101001111",
  42758=>"100000100",
  42759=>"101101010",
  42760=>"111001001",
  42761=>"001110100",
  42762=>"111111110",
  42763=>"000111000",
  42764=>"111111101",
  42765=>"111000100",
  42766=>"111010011",
  42767=>"110101000",
  42768=>"010100000",
  42769=>"101010000",
  42770=>"001011010",
  42771=>"000001100",
  42772=>"111000110",
  42773=>"110001111",
  42774=>"010101101",
  42775=>"100111010",
  42776=>"011001011",
  42777=>"001111111",
  42778=>"101111110",
  42779=>"110111010",
  42780=>"110101110",
  42781=>"001101111",
  42782=>"100001110",
  42783=>"000011101",
  42784=>"111100000",
  42785=>"011100010",
  42786=>"100001010",
  42787=>"010000111",
  42788=>"110101101",
  42789=>"001101111",
  42790=>"110101000",
  42791=>"010110110",
  42792=>"000101110",
  42793=>"001001111",
  42794=>"010101000",
  42795=>"000111011",
  42796=>"001001011",
  42797=>"011011010",
  42798=>"111000111",
  42799=>"000001011",
  42800=>"111100101",
  42801=>"100100010",
  42802=>"111111101",
  42803=>"001101011",
  42804=>"101011001",
  42805=>"101000101",
  42806=>"100110010",
  42807=>"011011110",
  42808=>"100101000",
  42809=>"111111111",
  42810=>"000101100",
  42811=>"000000011",
  42812=>"000011011",
  42813=>"101011110",
  42814=>"001101110",
  42815=>"011100111",
  42816=>"111010011",
  42817=>"000111001",
  42818=>"010010010",
  42819=>"000111010",
  42820=>"011010101",
  42821=>"011101011",
  42822=>"110101011",
  42823=>"110010011",
  42824=>"111111101",
  42825=>"011101101",
  42826=>"000011101",
  42827=>"001100101",
  42828=>"010111111",
  42829=>"001001111",
  42830=>"111111010",
  42831=>"000000001",
  42832=>"101011100",
  42833=>"011001110",
  42834=>"111010111",
  42835=>"010001110",
  42836=>"001101111",
  42837=>"000100001",
  42838=>"001011001",
  42839=>"111011100",
  42840=>"011111000",
  42841=>"010101100",
  42842=>"011011110",
  42843=>"100010110",
  42844=>"111000010",
  42845=>"111011110",
  42846=>"011101111",
  42847=>"110010110",
  42848=>"110010100",
  42849=>"010101100",
  42850=>"110111111",
  42851=>"100000001",
  42852=>"101011010",
  42853=>"000000010",
  42854=>"010110001",
  42855=>"001001100",
  42856=>"000110111",
  42857=>"000110110",
  42858=>"010011011",
  42859=>"110101100",
  42860=>"110001011",
  42861=>"100101011",
  42862=>"111011000",
  42863=>"010010110",
  42864=>"001001100",
  42865=>"101111100",
  42866=>"101101010",
  42867=>"000100011",
  42868=>"011001110",
  42869=>"111111111",
  42870=>"011000111",
  42871=>"001100011",
  42872=>"010100011",
  42873=>"100001010",
  42874=>"001101000",
  42875=>"110011111",
  42876=>"010111010",
  42877=>"001000001",
  42878=>"001010111",
  42879=>"000101000",
  42880=>"010110011",
  42881=>"110111000",
  42882=>"111011110",
  42883=>"000010101",
  42884=>"111110000",
  42885=>"101000010",
  42886=>"001001101",
  42887=>"101101011",
  42888=>"101100000",
  42889=>"010100001",
  42890=>"111010010",
  42891=>"101111011",
  42892=>"000110010",
  42893=>"101010000",
  42894=>"001001000",
  42895=>"111011010",
  42896=>"100111101",
  42897=>"100001111",
  42898=>"110100111",
  42899=>"100011111",
  42900=>"011100111",
  42901=>"010100111",
  42902=>"010000100",
  42903=>"001010011",
  42904=>"000101111",
  42905=>"011111011",
  42906=>"001111101",
  42907=>"100010101",
  42908=>"100000011",
  42909=>"101101011",
  42910=>"000110101",
  42911=>"111011101",
  42912=>"011111000",
  42913=>"001001001",
  42914=>"011011101",
  42915=>"011010011",
  42916=>"011100001",
  42917=>"101101100",
  42918=>"100010000",
  42919=>"001010111",
  42920=>"011111000",
  42921=>"011110100",
  42922=>"100011111",
  42923=>"010010111",
  42924=>"110001010",
  42925=>"110111110",
  42926=>"000011110",
  42927=>"101100101",
  42928=>"100100111",
  42929=>"110111000",
  42930=>"110111111",
  42931=>"011011000",
  42932=>"000001001",
  42933=>"100000001",
  42934=>"110001001",
  42935=>"000111110",
  42936=>"100101101",
  42937=>"111001011",
  42938=>"110100010",
  42939=>"011010100",
  42940=>"010100010",
  42941=>"000100000",
  42942=>"110101111",
  42943=>"111100011",
  42944=>"110100111",
  42945=>"110011000",
  42946=>"010110010",
  42947=>"100001100",
  42948=>"111011010",
  42949=>"101101010",
  42950=>"001010000",
  42951=>"000110100",
  42952=>"110110110",
  42953=>"000010010",
  42954=>"011111110",
  42955=>"011011111",
  42956=>"101000010",
  42957=>"110100100",
  42958=>"010111111",
  42959=>"010100011",
  42960=>"100111010",
  42961=>"100001010",
  42962=>"100011110",
  42963=>"100100101",
  42964=>"101111111",
  42965=>"101111101",
  42966=>"100101011",
  42967=>"001010111",
  42968=>"001111111",
  42969=>"001100001",
  42970=>"101100001",
  42971=>"010000010",
  42972=>"101011100",
  42973=>"000110000",
  42974=>"111001000",
  42975=>"111100111",
  42976=>"011010011",
  42977=>"100011111",
  42978=>"000010010",
  42979=>"000010010",
  42980=>"011000111",
  42981=>"010000000",
  42982=>"111000111",
  42983=>"101011010",
  42984=>"011111111",
  42985=>"110001101",
  42986=>"010111011",
  42987=>"010010111",
  42988=>"001101000",
  42989=>"110000110",
  42990=>"101001001",
  42991=>"100110010",
  42992=>"011010100",
  42993=>"100110101",
  42994=>"101111111",
  42995=>"011110001",
  42996=>"010110000",
  42997=>"110001011",
  42998=>"010101011",
  42999=>"001011110",
  43000=>"111000001",
  43001=>"101111101",
  43002=>"111111011",
  43003=>"101000000",
  43004=>"100000010",
  43005=>"101111001",
  43006=>"001001000",
  43007=>"010100101",
  43008=>"010101011",
  43009=>"001010110",
  43010=>"111101111",
  43011=>"010001100",
  43012=>"011100101",
  43013=>"101111101",
  43014=>"001101101",
  43015=>"000100110",
  43016=>"111111010",
  43017=>"100100001",
  43018=>"000110001",
  43019=>"001011011",
  43020=>"100011010",
  43021=>"100101100",
  43022=>"101001011",
  43023=>"010110000",
  43024=>"110100011",
  43025=>"110110101",
  43026=>"111001110",
  43027=>"000110100",
  43028=>"100000101",
  43029=>"011000110",
  43030=>"010110000",
  43031=>"100011101",
  43032=>"111011110",
  43033=>"011100010",
  43034=>"101110011",
  43035=>"000001001",
  43036=>"100110100",
  43037=>"010100110",
  43038=>"101100100",
  43039=>"001101000",
  43040=>"111000100",
  43041=>"010100110",
  43042=>"101011110",
  43043=>"100000000",
  43044=>"101110010",
  43045=>"001101011",
  43046=>"011000010",
  43047=>"111011101",
  43048=>"100010111",
  43049=>"111100011",
  43050=>"000000101",
  43051=>"011110100",
  43052=>"111011101",
  43053=>"101001111",
  43054=>"100011001",
  43055=>"101111010",
  43056=>"100001110",
  43057=>"000000110",
  43058=>"010000111",
  43059=>"111100010",
  43060=>"010000110",
  43061=>"101101011",
  43062=>"111011110",
  43063=>"111100010",
  43064=>"011111010",
  43065=>"101100111",
  43066=>"001000100",
  43067=>"000000111",
  43068=>"111101100",
  43069=>"100101010",
  43070=>"010111111",
  43071=>"111101000",
  43072=>"011110111",
  43073=>"000000100",
  43074=>"011111101",
  43075=>"010110111",
  43076=>"101000010",
  43077=>"110110001",
  43078=>"000011001",
  43079=>"010010010",
  43080=>"010001111",
  43081=>"110110110",
  43082=>"010100101",
  43083=>"000111111",
  43084=>"001100011",
  43085=>"000010100",
  43086=>"001101010",
  43087=>"111110011",
  43088=>"100011100",
  43089=>"011000001",
  43090=>"001010010",
  43091=>"100000001",
  43092=>"011011000",
  43093=>"110100010",
  43094=>"111111011",
  43095=>"100110010",
  43096=>"100111101",
  43097=>"000010100",
  43098=>"011110010",
  43099=>"010010111",
  43100=>"011110011",
  43101=>"110001111",
  43102=>"001000110",
  43103=>"000001111",
  43104=>"011110011",
  43105=>"111011000",
  43106=>"001101000",
  43107=>"001100100",
  43108=>"000100010",
  43109=>"111001100",
  43110=>"101001100",
  43111=>"100101011",
  43112=>"100100101",
  43113=>"001110011",
  43114=>"110100011",
  43115=>"101011110",
  43116=>"100010000",
  43117=>"110111011",
  43118=>"111000010",
  43119=>"000000110",
  43120=>"001110110",
  43121=>"011000011",
  43122=>"111111101",
  43123=>"010000010",
  43124=>"111101011",
  43125=>"110110111",
  43126=>"100110000",
  43127=>"100111101",
  43128=>"000110001",
  43129=>"000010100",
  43130=>"110110011",
  43131=>"110011010",
  43132=>"111011001",
  43133=>"110100100",
  43134=>"000001000",
  43135=>"100011111",
  43136=>"101000011",
  43137=>"111011011",
  43138=>"000110110",
  43139=>"011110110",
  43140=>"100011101",
  43141=>"100001110",
  43142=>"001010001",
  43143=>"011111101",
  43144=>"101110000",
  43145=>"100000101",
  43146=>"000110110",
  43147=>"010000110",
  43148=>"111011001",
  43149=>"101100100",
  43150=>"011010010",
  43151=>"010010110",
  43152=>"110010011",
  43153=>"011111000",
  43154=>"010110001",
  43155=>"000101010",
  43156=>"010001011",
  43157=>"000100000",
  43158=>"000110011",
  43159=>"110000110",
  43160=>"001101001",
  43161=>"101010011",
  43162=>"111010101",
  43163=>"000010110",
  43164=>"000001101",
  43165=>"100100010",
  43166=>"100111010",
  43167=>"001001001",
  43168=>"000110011",
  43169=>"000100011",
  43170=>"111010100",
  43171=>"111101111",
  43172=>"000111111",
  43173=>"010000010",
  43174=>"011110000",
  43175=>"110001100",
  43176=>"010101010",
  43177=>"110100011",
  43178=>"110100110",
  43179=>"110100011",
  43180=>"101010001",
  43181=>"110101100",
  43182=>"111001001",
  43183=>"111111110",
  43184=>"001100001",
  43185=>"111011100",
  43186=>"000001110",
  43187=>"010000000",
  43188=>"101001100",
  43189=>"001010110",
  43190=>"011100111",
  43191=>"111101101",
  43192=>"010110001",
  43193=>"111100010",
  43194=>"001001111",
  43195=>"011001001",
  43196=>"011111110",
  43197=>"101011011",
  43198=>"101111001",
  43199=>"011010011",
  43200=>"101111101",
  43201=>"000010001",
  43202=>"100000001",
  43203=>"100001110",
  43204=>"110011001",
  43205=>"100110000",
  43206=>"001010100",
  43207=>"110011101",
  43208=>"001000010",
  43209=>"000101111",
  43210=>"011111101",
  43211=>"111000000",
  43212=>"010010110",
  43213=>"011001111",
  43214=>"111001000",
  43215=>"001110100",
  43216=>"111001001",
  43217=>"001110100",
  43218=>"001100001",
  43219=>"100100010",
  43220=>"111100101",
  43221=>"101010011",
  43222=>"000000000",
  43223=>"001011000",
  43224=>"010010100",
  43225=>"101100110",
  43226=>"100011010",
  43227=>"011001001",
  43228=>"111111110",
  43229=>"100000101",
  43230=>"101001001",
  43231=>"110010000",
  43232=>"001100110",
  43233=>"100010001",
  43234=>"100111000",
  43235=>"111000110",
  43236=>"110110000",
  43237=>"000010010",
  43238=>"101000000",
  43239=>"101010011",
  43240=>"010111110",
  43241=>"110110000",
  43242=>"111001001",
  43243=>"000110101",
  43244=>"011000100",
  43245=>"011100010",
  43246=>"111000101",
  43247=>"010101011",
  43248=>"111100011",
  43249=>"011011001",
  43250=>"011011011",
  43251=>"101010111",
  43252=>"001011100",
  43253=>"100010111",
  43254=>"111111110",
  43255=>"110110011",
  43256=>"101110011",
  43257=>"010010101",
  43258=>"010111110",
  43259=>"001011111",
  43260=>"101110011",
  43261=>"001001000",
  43262=>"000100000",
  43263=>"000100011",
  43264=>"110100101",
  43265=>"011101010",
  43266=>"001101111",
  43267=>"001000010",
  43268=>"101111000",
  43269=>"001011010",
  43270=>"110100100",
  43271=>"010111100",
  43272=>"011000010",
  43273=>"001000011",
  43274=>"111010111",
  43275=>"001100011",
  43276=>"101101111",
  43277=>"011100001",
  43278=>"010100111",
  43279=>"111110010",
  43280=>"111110001",
  43281=>"001011101",
  43282=>"100100011",
  43283=>"010110000",
  43284=>"100011001",
  43285=>"000110000",
  43286=>"111010100",
  43287=>"110100010",
  43288=>"001101111",
  43289=>"101010100",
  43290=>"001010011",
  43291=>"101011101",
  43292=>"101000000",
  43293=>"010100110",
  43294=>"110111111",
  43295=>"111110010",
  43296=>"011000100",
  43297=>"010111011",
  43298=>"000011000",
  43299=>"101111000",
  43300=>"111000011",
  43301=>"101100110",
  43302=>"110101111",
  43303=>"001110111",
  43304=>"011011101",
  43305=>"010010111",
  43306=>"011101110",
  43307=>"000110011",
  43308=>"111111011",
  43309=>"101011010",
  43310=>"101000110",
  43311=>"011010000",
  43312=>"010100010",
  43313=>"011011011",
  43314=>"101111000",
  43315=>"101010000",
  43316=>"010011000",
  43317=>"001010101",
  43318=>"000101000",
  43319=>"000010000",
  43320=>"110101110",
  43321=>"110111110",
  43322=>"000011010",
  43323=>"001010110",
  43324=>"001010100",
  43325=>"000010101",
  43326=>"101011011",
  43327=>"000110111",
  43328=>"110010000",
  43329=>"000010111",
  43330=>"111001011",
  43331=>"111000110",
  43332=>"010000000",
  43333=>"101111000",
  43334=>"111000101",
  43335=>"000000001",
  43336=>"111100100",
  43337=>"110111101",
  43338=>"100100001",
  43339=>"111000000",
  43340=>"001111000",
  43341=>"110110010",
  43342=>"111010011",
  43343=>"001110111",
  43344=>"000001001",
  43345=>"110000011",
  43346=>"111001001",
  43347=>"111000000",
  43348=>"010110010",
  43349=>"111001100",
  43350=>"000010100",
  43351=>"111011110",
  43352=>"100011011",
  43353=>"101100000",
  43354=>"001000101",
  43355=>"100101100",
  43356=>"100101101",
  43357=>"000000010",
  43358=>"011100100",
  43359=>"101001100",
  43360=>"001001010",
  43361=>"111010010",
  43362=>"011101000",
  43363=>"000101011",
  43364=>"101100000",
  43365=>"111010101",
  43366=>"110100101",
  43367=>"000010100",
  43368=>"000011000",
  43369=>"011011011",
  43370=>"001100110",
  43371=>"011011001",
  43372=>"001111110",
  43373=>"011001010",
  43374=>"000011100",
  43375=>"111000011",
  43376=>"010110001",
  43377=>"001000111",
  43378=>"111100100",
  43379=>"101110010",
  43380=>"000000111",
  43381=>"111110111",
  43382=>"011100010",
  43383=>"110101111",
  43384=>"001110110",
  43385=>"101111101",
  43386=>"111011101",
  43387=>"000000100",
  43388=>"010011011",
  43389=>"111010010",
  43390=>"111001100",
  43391=>"010110111",
  43392=>"010100111",
  43393=>"011001011",
  43394=>"000001000",
  43395=>"000000000",
  43396=>"100110101",
  43397=>"010011010",
  43398=>"001111010",
  43399=>"001000011",
  43400=>"101000011",
  43401=>"001011011",
  43402=>"011100100",
  43403=>"110000011",
  43404=>"101111000",
  43405=>"000000110",
  43406=>"101101000",
  43407=>"000010010",
  43408=>"100100111",
  43409=>"100011111",
  43410=>"010100110",
  43411=>"011011000",
  43412=>"000111010",
  43413=>"110100110",
  43414=>"100001011",
  43415=>"011001101",
  43416=>"101100011",
  43417=>"000001110",
  43418=>"001000011",
  43419=>"111100001",
  43420=>"101010101",
  43421=>"111101010",
  43422=>"100101100",
  43423=>"110101010",
  43424=>"000010100",
  43425=>"111110111",
  43426=>"010011100",
  43427=>"011001001",
  43428=>"101110110",
  43429=>"101101100",
  43430=>"111110000",
  43431=>"001111111",
  43432=>"100000101",
  43433=>"101111001",
  43434=>"111110010",
  43435=>"001100001",
  43436=>"001111100",
  43437=>"111010100",
  43438=>"010001011",
  43439=>"100010000",
  43440=>"111000111",
  43441=>"010111101",
  43442=>"111110111",
  43443=>"110110111",
  43444=>"110111111",
  43445=>"000001100",
  43446=>"010011000",
  43447=>"010111101",
  43448=>"110001001",
  43449=>"010011010",
  43450=>"011010111",
  43451=>"000011000",
  43452=>"001001000",
  43453=>"010101011",
  43454=>"100001100",
  43455=>"110101001",
  43456=>"111011011",
  43457=>"111011100",
  43458=>"011101011",
  43459=>"110111001",
  43460=>"111000011",
  43461=>"001001001",
  43462=>"101111101",
  43463=>"110110011",
  43464=>"100100010",
  43465=>"110110001",
  43466=>"000100001",
  43467=>"000100101",
  43468=>"110000101",
  43469=>"100111010",
  43470=>"010111011",
  43471=>"110001010",
  43472=>"100100100",
  43473=>"101111011",
  43474=>"110011110",
  43475=>"111001010",
  43476=>"110111101",
  43477=>"110000011",
  43478=>"011000001",
  43479=>"110110010",
  43480=>"110001100",
  43481=>"010111100",
  43482=>"010000100",
  43483=>"001001111",
  43484=>"101001000",
  43485=>"001010110",
  43486=>"111111101",
  43487=>"010101100",
  43488=>"010111111",
  43489=>"011101001",
  43490=>"111011110",
  43491=>"011100000",
  43492=>"110010001",
  43493=>"111101011",
  43494=>"011010010",
  43495=>"110110101",
  43496=>"110001011",
  43497=>"000011111",
  43498=>"001010001",
  43499=>"101011111",
  43500=>"111010101",
  43501=>"101101000",
  43502=>"011010011",
  43503=>"111100000",
  43504=>"110010001",
  43505=>"100111011",
  43506=>"010010100",
  43507=>"010010101",
  43508=>"001100101",
  43509=>"110000000",
  43510=>"110100110",
  43511=>"000000000",
  43512=>"001101001",
  43513=>"111101011",
  43514=>"010000100",
  43515=>"010011011",
  43516=>"101011100",
  43517=>"000011110",
  43518=>"001000110",
  43519=>"011011010",
  43520=>"011000001",
  43521=>"010011111",
  43522=>"011001110",
  43523=>"111010110",
  43524=>"111101010",
  43525=>"100101001",
  43526=>"110001001",
  43527=>"101001001",
  43528=>"110100101",
  43529=>"010010100",
  43530=>"001010110",
  43531=>"000010001",
  43532=>"100111011",
  43533=>"001110001",
  43534=>"001101000",
  43535=>"010100011",
  43536=>"011100110",
  43537=>"100010010",
  43538=>"011001101",
  43539=>"001001000",
  43540=>"000010000",
  43541=>"010010100",
  43542=>"110001010",
  43543=>"110110000",
  43544=>"000110010",
  43545=>"010000110",
  43546=>"110111111",
  43547=>"011000100",
  43548=>"101001010",
  43549=>"101101110",
  43550=>"010111010",
  43551=>"110111111",
  43552=>"001010000",
  43553=>"100011001",
  43554=>"111001000",
  43555=>"111100011",
  43556=>"001100101",
  43557=>"110011110",
  43558=>"100000111",
  43559=>"001110100",
  43560=>"111110101",
  43561=>"101110111",
  43562=>"110110111",
  43563=>"101101000",
  43564=>"001011011",
  43565=>"001100000",
  43566=>"010001001",
  43567=>"110101010",
  43568=>"110000001",
  43569=>"101101110",
  43570=>"001000110",
  43571=>"011010100",
  43572=>"000111110",
  43573=>"001011001",
  43574=>"011100001",
  43575=>"111011111",
  43576=>"101110100",
  43577=>"100100000",
  43578=>"011101011",
  43579=>"010101100",
  43580=>"100010111",
  43581=>"011110110",
  43582=>"001111000",
  43583=>"001001101",
  43584=>"010000010",
  43585=>"001000001",
  43586=>"010100010",
  43587=>"001111001",
  43588=>"010001010",
  43589=>"001001111",
  43590=>"100000001",
  43591=>"100010110",
  43592=>"101101110",
  43593=>"100000110",
  43594=>"011011110",
  43595=>"110100110",
  43596=>"110100001",
  43597=>"000100011",
  43598=>"101000010",
  43599=>"000100110",
  43600=>"011101010",
  43601=>"001010110",
  43602=>"110001111",
  43603=>"101001101",
  43604=>"101011001",
  43605=>"011011001",
  43606=>"100011001",
  43607=>"110011000",
  43608=>"001000010",
  43609=>"100011111",
  43610=>"011001001",
  43611=>"101011100",
  43612=>"001011011",
  43613=>"100010001",
  43614=>"111000110",
  43615=>"100100100",
  43616=>"100111000",
  43617=>"011100111",
  43618=>"110101000",
  43619=>"110011101",
  43620=>"001011101",
  43621=>"111000101",
  43622=>"011101010",
  43623=>"111001010",
  43624=>"100100111",
  43625=>"110101010",
  43626=>"110111001",
  43627=>"001000111",
  43628=>"010010010",
  43629=>"010010111",
  43630=>"001100110",
  43631=>"110011110",
  43632=>"101011111",
  43633=>"011010010",
  43634=>"000111101",
  43635=>"111011010",
  43636=>"000011010",
  43637=>"100100100",
  43638=>"110001101",
  43639=>"111101111",
  43640=>"101010011",
  43641=>"111101001",
  43642=>"011110100",
  43643=>"001010101",
  43644=>"001000010",
  43645=>"001100001",
  43646=>"111111101",
  43647=>"011100000",
  43648=>"110110011",
  43649=>"111010100",
  43650=>"100100010",
  43651=>"011001111",
  43652=>"110101001",
  43653=>"101100000",
  43654=>"011001010",
  43655=>"001101011",
  43656=>"101011001",
  43657=>"000101110",
  43658=>"011111000",
  43659=>"101101010",
  43660=>"011100010",
  43661=>"001011110",
  43662=>"101101100",
  43663=>"100000100",
  43664=>"000011000",
  43665=>"001010110",
  43666=>"100101000",
  43667=>"101000011",
  43668=>"100100100",
  43669=>"001010100",
  43670=>"111100101",
  43671=>"110000001",
  43672=>"000000010",
  43673=>"010100000",
  43674=>"110010111",
  43675=>"010100101",
  43676=>"010000110",
  43677=>"101001100",
  43678=>"111001011",
  43679=>"110001111",
  43680=>"001101011",
  43681=>"000110000",
  43682=>"001111101",
  43683=>"100001010",
  43684=>"001010001",
  43685=>"010010010",
  43686=>"001011100",
  43687=>"011000000",
  43688=>"110100100",
  43689=>"000100000",
  43690=>"111100110",
  43691=>"010001001",
  43692=>"100000111",
  43693=>"000001001",
  43694=>"011100101",
  43695=>"101110000",
  43696=>"100001111",
  43697=>"000010111",
  43698=>"000101110",
  43699=>"101011000",
  43700=>"010110011",
  43701=>"110111010",
  43702=>"110000111",
  43703=>"100101101",
  43704=>"011110000",
  43705=>"101011001",
  43706=>"011010011",
  43707=>"111110011",
  43708=>"101100100",
  43709=>"000000000",
  43710=>"111000000",
  43711=>"000010010",
  43712=>"010010010",
  43713=>"001000111",
  43714=>"000011011",
  43715=>"001100111",
  43716=>"101000110",
  43717=>"111010111",
  43718=>"101111000",
  43719=>"001001101",
  43720=>"000000110",
  43721=>"000000111",
  43722=>"111000001",
  43723=>"000110111",
  43724=>"010111111",
  43725=>"110110111",
  43726=>"101000111",
  43727=>"111000111",
  43728=>"101100111",
  43729=>"001101100",
  43730=>"111101001",
  43731=>"110101010",
  43732=>"010010010",
  43733=>"111011011",
  43734=>"110000111",
  43735=>"111100110",
  43736=>"000111111",
  43737=>"110101010",
  43738=>"010000010",
  43739=>"110010111",
  43740=>"001101100",
  43741=>"101111011",
  43742=>"000111010",
  43743=>"010011011",
  43744=>"101100101",
  43745=>"000100000",
  43746=>"110011101",
  43747=>"011000000",
  43748=>"010100011",
  43749=>"000111101",
  43750=>"111100001",
  43751=>"101101101",
  43752=>"001111100",
  43753=>"101001111",
  43754=>"001011110",
  43755=>"100000011",
  43756=>"111100000",
  43757=>"100010010",
  43758=>"111111010",
  43759=>"000001111",
  43760=>"110010001",
  43761=>"000110011",
  43762=>"011000001",
  43763=>"101101100",
  43764=>"001110000",
  43765=>"110010000",
  43766=>"101101101",
  43767=>"011100101",
  43768=>"000111101",
  43769=>"111000110",
  43770=>"010101111",
  43771=>"011000111",
  43772=>"110000001",
  43773=>"010110011",
  43774=>"111000101",
  43775=>"110101011",
  43776=>"011111010",
  43777=>"010000110",
  43778=>"111110010",
  43779=>"111101101",
  43780=>"000110101",
  43781=>"001000101",
  43782=>"100010101",
  43783=>"010101011",
  43784=>"010110001",
  43785=>"111111010",
  43786=>"011001011",
  43787=>"010000011",
  43788=>"001111100",
  43789=>"101101101",
  43790=>"011001101",
  43791=>"000000000",
  43792=>"101111111",
  43793=>"001011111",
  43794=>"011100011",
  43795=>"110010101",
  43796=>"000111110",
  43797=>"010111110",
  43798=>"101110111",
  43799=>"100010000",
  43800=>"100100000",
  43801=>"110110100",
  43802=>"000001010",
  43803=>"011011000",
  43804=>"110010101",
  43805=>"100001001",
  43806=>"010010001",
  43807=>"000001110",
  43808=>"101100100",
  43809=>"001100110",
  43810=>"110011101",
  43811=>"010100101",
  43812=>"111100000",
  43813=>"110001111",
  43814=>"001011110",
  43815=>"000100101",
  43816=>"000110110",
  43817=>"000010010",
  43818=>"100011101",
  43819=>"101100000",
  43820=>"011100110",
  43821=>"001000111",
  43822=>"110101011",
  43823=>"111100111",
  43824=>"000010010",
  43825=>"110001111",
  43826=>"011011011",
  43827=>"101111000",
  43828=>"010101011",
  43829=>"110110100",
  43830=>"001001010",
  43831=>"101000000",
  43832=>"100001111",
  43833=>"001010010",
  43834=>"000100101",
  43835=>"101000111",
  43836=>"000001111",
  43837=>"010000100",
  43838=>"001010101",
  43839=>"010101100",
  43840=>"101001000",
  43841=>"001101101",
  43842=>"011011010",
  43843=>"111111100",
  43844=>"000010111",
  43845=>"110011001",
  43846=>"001000100",
  43847=>"111100001",
  43848=>"101100000",
  43849=>"100011011",
  43850=>"000101100",
  43851=>"111110100",
  43852=>"101101010",
  43853=>"110111010",
  43854=>"001110011",
  43855=>"000100011",
  43856=>"000110001",
  43857=>"010100010",
  43858=>"110000000",
  43859=>"010101000",
  43860=>"001010010",
  43861=>"111101011",
  43862=>"101001101",
  43863=>"000111011",
  43864=>"011001000",
  43865=>"101000000",
  43866=>"110101111",
  43867=>"010000100",
  43868=>"111001111",
  43869=>"111011101",
  43870=>"010110100",
  43871=>"101011011",
  43872=>"010110111",
  43873=>"011111111",
  43874=>"000001000",
  43875=>"110100001",
  43876=>"011010111",
  43877=>"000000001",
  43878=>"000101100",
  43879=>"000110010",
  43880=>"111100101",
  43881=>"011100000",
  43882=>"000011111",
  43883=>"110000111",
  43884=>"100101001",
  43885=>"110111101",
  43886=>"011011111",
  43887=>"010110100",
  43888=>"110100001",
  43889=>"011101101",
  43890=>"111000001",
  43891=>"100111010",
  43892=>"010001000",
  43893=>"010110000",
  43894=>"110010100",
  43895=>"000010110",
  43896=>"111100111",
  43897=>"010110111",
  43898=>"011110001",
  43899=>"010101001",
  43900=>"110000100",
  43901=>"011100100",
  43902=>"100010001",
  43903=>"111001011",
  43904=>"110111011",
  43905=>"100100011",
  43906=>"010001110",
  43907=>"001000110",
  43908=>"011011011",
  43909=>"011000110",
  43910=>"001010000",
  43911=>"111111101",
  43912=>"010001010",
  43913=>"101100100",
  43914=>"100001010",
  43915=>"001110110",
  43916=>"111100100",
  43917=>"010010011",
  43918=>"100001010",
  43919=>"000011110",
  43920=>"011110110",
  43921=>"010110100",
  43922=>"101000000",
  43923=>"001010100",
  43924=>"011001111",
  43925=>"110000010",
  43926=>"000011010",
  43927=>"011011001",
  43928=>"011110100",
  43929=>"001110000",
  43930=>"111101010",
  43931=>"011100010",
  43932=>"110100100",
  43933=>"100110101",
  43934=>"111111011",
  43935=>"111111011",
  43936=>"100100000",
  43937=>"101011000",
  43938=>"111101000",
  43939=>"000010011",
  43940=>"111111111",
  43941=>"111111101",
  43942=>"110001001",
  43943=>"000000101",
  43944=>"110010011",
  43945=>"010111111",
  43946=>"000111011",
  43947=>"011010010",
  43948=>"000010001",
  43949=>"000000000",
  43950=>"111111110",
  43951=>"000110000",
  43952=>"000111110",
  43953=>"001000010",
  43954=>"010100010",
  43955=>"010111000",
  43956=>"000111011",
  43957=>"101100111",
  43958=>"010111011",
  43959=>"000111000",
  43960=>"101111100",
  43961=>"011111110",
  43962=>"110010111",
  43963=>"010100011",
  43964=>"011100110",
  43965=>"010101011",
  43966=>"111100101",
  43967=>"101111001",
  43968=>"111010011",
  43969=>"101110010",
  43970=>"111000010",
  43971=>"101010110",
  43972=>"010000100",
  43973=>"001010000",
  43974=>"000010100",
  43975=>"101011010",
  43976=>"101100111",
  43977=>"100010010",
  43978=>"100100101",
  43979=>"000011111",
  43980=>"100101101",
  43981=>"010011111",
  43982=>"111100000",
  43983=>"101000100",
  43984=>"101000001",
  43985=>"110110000",
  43986=>"001100010",
  43987=>"001001100",
  43988=>"000000000",
  43989=>"110001100",
  43990=>"010101010",
  43991=>"011011111",
  43992=>"010000100",
  43993=>"101100010",
  43994=>"001000110",
  43995=>"010011001",
  43996=>"100010111",
  43997=>"001000011",
  43998=>"100111011",
  43999=>"101100001",
  44000=>"101101010",
  44001=>"111010011",
  44002=>"011101101",
  44003=>"100110101",
  44004=>"011100101",
  44005=>"110111010",
  44006=>"010011010",
  44007=>"111101101",
  44008=>"110000100",
  44009=>"101101010",
  44010=>"101011011",
  44011=>"110111000",
  44012=>"011001001",
  44013=>"100000000",
  44014=>"011000100",
  44015=>"100001110",
  44016=>"110011110",
  44017=>"101010101",
  44018=>"011010011",
  44019=>"010001111",
  44020=>"001010011",
  44021=>"111011010",
  44022=>"000001011",
  44023=>"000110110",
  44024=>"010101100",
  44025=>"010100011",
  44026=>"000111011",
  44027=>"100001001",
  44028=>"110000010",
  44029=>"000111010",
  44030=>"111110111",
  44031=>"001101000",
  44032=>"110111111",
  44033=>"101101111",
  44034=>"110100000",
  44035=>"000000011",
  44036=>"010001001",
  44037=>"010100010",
  44038=>"100111110",
  44039=>"111111000",
  44040=>"110010101",
  44041=>"011111101",
  44042=>"111101101",
  44043=>"101110001",
  44044=>"000100011",
  44045=>"011100001",
  44046=>"001110110",
  44047=>"111111110",
  44048=>"101100001",
  44049=>"011010010",
  44050=>"001101011",
  44051=>"010011100",
  44052=>"100101001",
  44053=>"100101100",
  44054=>"000010111",
  44055=>"000000010",
  44056=>"000011100",
  44057=>"101100001",
  44058=>"010010101",
  44059=>"110100001",
  44060=>"100110011",
  44061=>"000011011",
  44062=>"000011001",
  44063=>"110110101",
  44064=>"110101100",
  44065=>"100111110",
  44066=>"011000011",
  44067=>"001000000",
  44068=>"110001011",
  44069=>"100010111",
  44070=>"010101000",
  44071=>"110000100",
  44072=>"110111011",
  44073=>"001101011",
  44074=>"101001100",
  44075=>"000000101",
  44076=>"101111110",
  44077=>"010011011",
  44078=>"101000101",
  44079=>"011010111",
  44080=>"111100011",
  44081=>"100001101",
  44082=>"001101110",
  44083=>"010000110",
  44084=>"111010110",
  44085=>"001000100",
  44086=>"100011010",
  44087=>"000100101",
  44088=>"100010101",
  44089=>"100000100",
  44090=>"101110011",
  44091=>"000110111",
  44092=>"000011110",
  44093=>"110010001",
  44094=>"111011010",
  44095=>"001010010",
  44096=>"100000101",
  44097=>"000001101",
  44098=>"000010010",
  44099=>"001100000",
  44100=>"011010000",
  44101=>"001100111",
  44102=>"011000000",
  44103=>"000111011",
  44104=>"100110011",
  44105=>"100010000",
  44106=>"010011110",
  44107=>"110001000",
  44108=>"111010000",
  44109=>"000111101",
  44110=>"111101110",
  44111=>"010101000",
  44112=>"111111011",
  44113=>"001010010",
  44114=>"110001000",
  44115=>"111110100",
  44116=>"111000000",
  44117=>"100001010",
  44118=>"010111001",
  44119=>"001110001",
  44120=>"111000011",
  44121=>"110001011",
  44122=>"011101111",
  44123=>"110101101",
  44124=>"000111111",
  44125=>"100000001",
  44126=>"100111101",
  44127=>"100001000",
  44128=>"000010000",
  44129=>"011111000",
  44130=>"101111011",
  44131=>"010100110",
  44132=>"110000110",
  44133=>"101001110",
  44134=>"100101110",
  44135=>"000110000",
  44136=>"000000001",
  44137=>"110001111",
  44138=>"000010100",
  44139=>"011101011",
  44140=>"111001100",
  44141=>"011111001",
  44142=>"110001111",
  44143=>"010001111",
  44144=>"110110011",
  44145=>"001111011",
  44146=>"111101110",
  44147=>"100011100",
  44148=>"000011010",
  44149=>"010011100",
  44150=>"100111100",
  44151=>"100001100",
  44152=>"001111110",
  44153=>"110101010",
  44154=>"111111011",
  44155=>"000110101",
  44156=>"000011110",
  44157=>"111111000",
  44158=>"000011100",
  44159=>"111101110",
  44160=>"111111111",
  44161=>"010101100",
  44162=>"111101001",
  44163=>"011010011",
  44164=>"100100000",
  44165=>"111010110",
  44166=>"110110001",
  44167=>"011000100",
  44168=>"011000101",
  44169=>"000110110",
  44170=>"110101010",
  44171=>"110111000",
  44172=>"000011111",
  44173=>"100101010",
  44174=>"100111111",
  44175=>"000010101",
  44176=>"010000101",
  44177=>"000001001",
  44178=>"000010010",
  44179=>"000001111",
  44180=>"001000100",
  44181=>"101010111",
  44182=>"010011001",
  44183=>"011100100",
  44184=>"000010010",
  44185=>"011110010",
  44186=>"100111010",
  44187=>"101101010",
  44188=>"101101000",
  44189=>"010111100",
  44190=>"111000001",
  44191=>"100011010",
  44192=>"101010101",
  44193=>"001101111",
  44194=>"111000110",
  44195=>"011010001",
  44196=>"010001011",
  44197=>"000001110",
  44198=>"101111100",
  44199=>"101111011",
  44200=>"011000011",
  44201=>"000010010",
  44202=>"100000101",
  44203=>"010010010",
  44204=>"100010110",
  44205=>"011010010",
  44206=>"100010100",
  44207=>"100011010",
  44208=>"101001010",
  44209=>"101111011",
  44210=>"111101110",
  44211=>"000110000",
  44212=>"000110100",
  44213=>"111001111",
  44214=>"100010100",
  44215=>"100101100",
  44216=>"001010010",
  44217=>"111000010",
  44218=>"111011100",
  44219=>"110100000",
  44220=>"111100111",
  44221=>"100011000",
  44222=>"100010100",
  44223=>"011010101",
  44224=>"011111100",
  44225=>"001101110",
  44226=>"101011111",
  44227=>"011011101",
  44228=>"101100000",
  44229=>"011010010",
  44230=>"010101101",
  44231=>"010100111",
  44232=>"100100110",
  44233=>"101101101",
  44234=>"111101111",
  44235=>"100001101",
  44236=>"001001010",
  44237=>"110000110",
  44238=>"110000111",
  44239=>"000010010",
  44240=>"111100111",
  44241=>"111000000",
  44242=>"111100111",
  44243=>"011001000",
  44244=>"101100001",
  44245=>"001101110",
  44246=>"010011100",
  44247=>"111011001",
  44248=>"101010010",
  44249=>"001110110",
  44250=>"111000111",
  44251=>"101001001",
  44252=>"110101011",
  44253=>"110001100",
  44254=>"000110000",
  44255=>"011001111",
  44256=>"011010100",
  44257=>"101101001",
  44258=>"110101110",
  44259=>"011101111",
  44260=>"011000001",
  44261=>"001011010",
  44262=>"001001101",
  44263=>"100010001",
  44264=>"000010010",
  44265=>"100100010",
  44266=>"011101011",
  44267=>"110001001",
  44268=>"010100100",
  44269=>"011110011",
  44270=>"000110010",
  44271=>"101111101",
  44272=>"110100010",
  44273=>"101001101",
  44274=>"000101111",
  44275=>"101111101",
  44276=>"101111101",
  44277=>"110000001",
  44278=>"110111000",
  44279=>"001010110",
  44280=>"000001111",
  44281=>"010111000",
  44282=>"111001111",
  44283=>"101010001",
  44284=>"000000001",
  44285=>"100010111",
  44286=>"110111111",
  44287=>"111011110",
  44288=>"110111110",
  44289=>"010110101",
  44290=>"000100110",
  44291=>"100100001",
  44292=>"111101110",
  44293=>"111011100",
  44294=>"001000100",
  44295=>"110100010",
  44296=>"011101111",
  44297=>"101010110",
  44298=>"110001111",
  44299=>"111110100",
  44300=>"101100001",
  44301=>"011010010",
  44302=>"001001110",
  44303=>"011010000",
  44304=>"101111101",
  44305=>"010111000",
  44306=>"000101110",
  44307=>"000000010",
  44308=>"011100100",
  44309=>"011111111",
  44310=>"000000111",
  44311=>"000100001",
  44312=>"111010110",
  44313=>"001111100",
  44314=>"011000100",
  44315=>"011100000",
  44316=>"111001110",
  44317=>"110110010",
  44318=>"111010101",
  44319=>"010010100",
  44320=>"111110001",
  44321=>"111010111",
  44322=>"000110010",
  44323=>"000000111",
  44324=>"100100001",
  44325=>"101101101",
  44326=>"000001111",
  44327=>"101101100",
  44328=>"111001110",
  44329=>"110011000",
  44330=>"001110000",
  44331=>"001011100",
  44332=>"111001100",
  44333=>"001011111",
  44334=>"000001000",
  44335=>"001000001",
  44336=>"111001101",
  44337=>"110110000",
  44338=>"111111100",
  44339=>"100100101",
  44340=>"001100010",
  44341=>"100101101",
  44342=>"000101010",
  44343=>"001011101",
  44344=>"001010110",
  44345=>"111110110",
  44346=>"010111110",
  44347=>"010000111",
  44348=>"111100110",
  44349=>"101010100",
  44350=>"000111000",
  44351=>"000000100",
  44352=>"101000110",
  44353=>"110011010",
  44354=>"000010111",
  44355=>"011000000",
  44356=>"101101100",
  44357=>"000011100",
  44358=>"100001010",
  44359=>"001101110",
  44360=>"010001100",
  44361=>"100000011",
  44362=>"101011101",
  44363=>"101100110",
  44364=>"101100000",
  44365=>"110010011",
  44366=>"100100001",
  44367=>"100011110",
  44368=>"001010001",
  44369=>"101000101",
  44370=>"011101000",
  44371=>"000000111",
  44372=>"100101001",
  44373=>"100111000",
  44374=>"111011000",
  44375=>"110110100",
  44376=>"000010001",
  44377=>"100100111",
  44378=>"101111011",
  44379=>"100000110",
  44380=>"001001100",
  44381=>"111100010",
  44382=>"001100011",
  44383=>"101011101",
  44384=>"001110100",
  44385=>"110101001",
  44386=>"000000100",
  44387=>"110100110",
  44388=>"011100001",
  44389=>"111101001",
  44390=>"001001111",
  44391=>"011010100",
  44392=>"000101011",
  44393=>"010011101",
  44394=>"111010100",
  44395=>"100001001",
  44396=>"000001011",
  44397=>"011101111",
  44398=>"011000011",
  44399=>"001100101",
  44400=>"110000000",
  44401=>"111010001",
  44402=>"111011001",
  44403=>"100000010",
  44404=>"010100110",
  44405=>"100111010",
  44406=>"010001111",
  44407=>"010000111",
  44408=>"001001110",
  44409=>"000110001",
  44410=>"011011101",
  44411=>"111101110",
  44412=>"110111000",
  44413=>"110010110",
  44414=>"100000110",
  44415=>"100010110",
  44416=>"101110010",
  44417=>"011100111",
  44418=>"010011011",
  44419=>"101001100",
  44420=>"010010011",
  44421=>"100011110",
  44422=>"100111011",
  44423=>"010111101",
  44424=>"100001111",
  44425=>"000100010",
  44426=>"110101001",
  44427=>"100101111",
  44428=>"101100100",
  44429=>"000010111",
  44430=>"011011001",
  44431=>"110110001",
  44432=>"000011110",
  44433=>"111000101",
  44434=>"110000010",
  44435=>"111100111",
  44436=>"101011110",
  44437=>"010001000",
  44438=>"010110110",
  44439=>"111111010",
  44440=>"000111011",
  44441=>"000000000",
  44442=>"011010111",
  44443=>"010100110",
  44444=>"101001100",
  44445=>"111110000",
  44446=>"100110110",
  44447=>"010000010",
  44448=>"001000110",
  44449=>"101010001",
  44450=>"000010010",
  44451=>"110010000",
  44452=>"110110110",
  44453=>"101100001",
  44454=>"000100000",
  44455=>"001110110",
  44456=>"001100010",
  44457=>"101001000",
  44458=>"110111000",
  44459=>"000000011",
  44460=>"100011110",
  44461=>"100010111",
  44462=>"010100111",
  44463=>"010011111",
  44464=>"111111111",
  44465=>"100111100",
  44466=>"011111000",
  44467=>"101000100",
  44468=>"010011001",
  44469=>"001010100",
  44470=>"010000010",
  44471=>"011001110",
  44472=>"111011000",
  44473=>"001010110",
  44474=>"110010000",
  44475=>"111110100",
  44476=>"100000110",
  44477=>"100001111",
  44478=>"101001100",
  44479=>"110100001",
  44480=>"010111011",
  44481=>"110111110",
  44482=>"000001000",
  44483=>"100010100",
  44484=>"000001001",
  44485=>"010010011",
  44486=>"000111110",
  44487=>"000011010",
  44488=>"110110001",
  44489=>"001011101",
  44490=>"110100010",
  44491=>"011100100",
  44492=>"000101111",
  44493=>"011011111",
  44494=>"011001111",
  44495=>"010111011",
  44496=>"000010101",
  44497=>"110000000",
  44498=>"100010010",
  44499=>"101101010",
  44500=>"011101011",
  44501=>"010011001",
  44502=>"100100111",
  44503=>"101000100",
  44504=>"001011011",
  44505=>"011100100",
  44506=>"110010110",
  44507=>"101111110",
  44508=>"101010100",
  44509=>"001000111",
  44510=>"111011101",
  44511=>"100001100",
  44512=>"001001111",
  44513=>"000001110",
  44514=>"011000110",
  44515=>"100001110",
  44516=>"111000001",
  44517=>"000010010",
  44518=>"001100101",
  44519=>"101111111",
  44520=>"100101010",
  44521=>"001100110",
  44522=>"011101100",
  44523=>"111111111",
  44524=>"011111110",
  44525=>"001100001",
  44526=>"010101011",
  44527=>"110101010",
  44528=>"000010000",
  44529=>"001111101",
  44530=>"111010100",
  44531=>"011110111",
  44532=>"011000100",
  44533=>"011000111",
  44534=>"001010010",
  44535=>"100100111",
  44536=>"011001100",
  44537=>"100100010",
  44538=>"101110001",
  44539=>"000000110",
  44540=>"001001100",
  44541=>"010000000",
  44542=>"010000101",
  44543=>"100011101",
  44544=>"110011000",
  44545=>"100000010",
  44546=>"100010111",
  44547=>"011111100",
  44548=>"111011110",
  44549=>"101110010",
  44550=>"011000011",
  44551=>"010010111",
  44552=>"001101011",
  44553=>"100110010",
  44554=>"000001110",
  44555=>"001010000",
  44556=>"111100111",
  44557=>"001100111",
  44558=>"011000010",
  44559=>"111010001",
  44560=>"111110111",
  44561=>"100110011",
  44562=>"010000111",
  44563=>"000011010",
  44564=>"100000010",
  44565=>"011111000",
  44566=>"001010111",
  44567=>"001011110",
  44568=>"001001101",
  44569=>"011100101",
  44570=>"111111100",
  44571=>"110110001",
  44572=>"010101100",
  44573=>"100010011",
  44574=>"100010001",
  44575=>"010111110",
  44576=>"101101011",
  44577=>"010011010",
  44578=>"011001001",
  44579=>"000111010",
  44580=>"011001100",
  44581=>"000110100",
  44582=>"000011101",
  44583=>"110100000",
  44584=>"011000110",
  44585=>"100011100",
  44586=>"101011101",
  44587=>"010111010",
  44588=>"001101111",
  44589=>"000000001",
  44590=>"000000010",
  44591=>"001011000",
  44592=>"101110110",
  44593=>"101111001",
  44594=>"011011100",
  44595=>"101111010",
  44596=>"100100111",
  44597=>"110111001",
  44598=>"111001111",
  44599=>"011001001",
  44600=>"111000100",
  44601=>"000100000",
  44602=>"010010101",
  44603=>"111001110",
  44604=>"000010100",
  44605=>"001000110",
  44606=>"111010100",
  44607=>"110101110",
  44608=>"010010100",
  44609=>"110001111",
  44610=>"111001111",
  44611=>"011000110",
  44612=>"101011000",
  44613=>"111011111",
  44614=>"110110000",
  44615=>"111001101",
  44616=>"001001100",
  44617=>"000110001",
  44618=>"001000001",
  44619=>"001100110",
  44620=>"010111110",
  44621=>"011010011",
  44622=>"110011111",
  44623=>"000001110",
  44624=>"010011010",
  44625=>"010001011",
  44626=>"111111101",
  44627=>"110011000",
  44628=>"100010001",
  44629=>"001000001",
  44630=>"111111000",
  44631=>"101000011",
  44632=>"111000110",
  44633=>"001010010",
  44634=>"110111111",
  44635=>"100110100",
  44636=>"101000000",
  44637=>"000110011",
  44638=>"111001011",
  44639=>"001100110",
  44640=>"110001101",
  44641=>"101111010",
  44642=>"011100110",
  44643=>"101001110",
  44644=>"000110010",
  44645=>"011001111",
  44646=>"010000110",
  44647=>"011000100",
  44648=>"001011011",
  44649=>"100000100",
  44650=>"010110000",
  44651=>"111011001",
  44652=>"101100011",
  44653=>"001101111",
  44654=>"100000010",
  44655=>"100101011",
  44656=>"111101011",
  44657=>"111111110",
  44658=>"000111111",
  44659=>"001011101",
  44660=>"111001010",
  44661=>"111111101",
  44662=>"011001010",
  44663=>"011100110",
  44664=>"010001001",
  44665=>"110110001",
  44666=>"011110010",
  44667=>"000101000",
  44668=>"010100000",
  44669=>"100001100",
  44670=>"111001000",
  44671=>"010110100",
  44672=>"010001101",
  44673=>"010111100",
  44674=>"011100011",
  44675=>"010110001",
  44676=>"011101100",
  44677=>"111100011",
  44678=>"000011101",
  44679=>"110011010",
  44680=>"110001100",
  44681=>"010100001",
  44682=>"110111010",
  44683=>"000011100",
  44684=>"010101101",
  44685=>"000000001",
  44686=>"101001000",
  44687=>"011001101",
  44688=>"011000000",
  44689=>"110010110",
  44690=>"000110001",
  44691=>"111101111",
  44692=>"000111110",
  44693=>"001010010",
  44694=>"000010110",
  44695=>"101111010",
  44696=>"011010000",
  44697=>"111011001",
  44698=>"001111001",
  44699=>"110100101",
  44700=>"000001001",
  44701=>"111101011",
  44702=>"011111001",
  44703=>"001000101",
  44704=>"001000100",
  44705=>"110010111",
  44706=>"110011101",
  44707=>"010001001",
  44708=>"100011011",
  44709=>"111111101",
  44710=>"100000001",
  44711=>"000100001",
  44712=>"011111110",
  44713=>"000100011",
  44714=>"100101101",
  44715=>"000100100",
  44716=>"110001111",
  44717=>"111001010",
  44718=>"000000001",
  44719=>"100001000",
  44720=>"010010101",
  44721=>"111100101",
  44722=>"110101101",
  44723=>"110110101",
  44724=>"101010000",
  44725=>"001010101",
  44726=>"011100010",
  44727=>"001101000",
  44728=>"000111100",
  44729=>"011010011",
  44730=>"111000111",
  44731=>"000111101",
  44732=>"011110000",
  44733=>"111111011",
  44734=>"001110011",
  44735=>"000000111",
  44736=>"000110101",
  44737=>"010010110",
  44738=>"011100100",
  44739=>"001111111",
  44740=>"100011111",
  44741=>"010010110",
  44742=>"111010010",
  44743=>"001111100",
  44744=>"100000000",
  44745=>"110111111",
  44746=>"011011111",
  44747=>"110000100",
  44748=>"110000001",
  44749=>"011101101",
  44750=>"000001111",
  44751=>"000110000",
  44752=>"000000100",
  44753=>"011101111",
  44754=>"110110100",
  44755=>"100010011",
  44756=>"110100011",
  44757=>"010011001",
  44758=>"011110101",
  44759=>"001001001",
  44760=>"011111110",
  44761=>"110000000",
  44762=>"000001001",
  44763=>"111100011",
  44764=>"011001011",
  44765=>"000101010",
  44766=>"011100101",
  44767=>"100110011",
  44768=>"001101010",
  44769=>"001000100",
  44770=>"010001100",
  44771=>"101111100",
  44772=>"111011100",
  44773=>"101100111",
  44774=>"011011010",
  44775=>"011100000",
  44776=>"101010001",
  44777=>"000000001",
  44778=>"111110001",
  44779=>"111011011",
  44780=>"110010111",
  44781=>"101111110",
  44782=>"111010111",
  44783=>"101111100",
  44784=>"001110111",
  44785=>"001101110",
  44786=>"101100001",
  44787=>"100100100",
  44788=>"110101011",
  44789=>"101100110",
  44790=>"110111100",
  44791=>"010111101",
  44792=>"001000100",
  44793=>"101011110",
  44794=>"100110001",
  44795=>"111111111",
  44796=>"111001001",
  44797=>"100111010",
  44798=>"010110100",
  44799=>"001110110",
  44800=>"011111000",
  44801=>"011110010",
  44802=>"110111110",
  44803=>"100011110",
  44804=>"001100110",
  44805=>"001011110",
  44806=>"010111011",
  44807=>"100110001",
  44808=>"010001001",
  44809=>"100010011",
  44810=>"001110111",
  44811=>"010010100",
  44812=>"111011011",
  44813=>"100000010",
  44814=>"011001000",
  44815=>"010000001",
  44816=>"010101011",
  44817=>"011111011",
  44818=>"011001101",
  44819=>"010111001",
  44820=>"010011111",
  44821=>"110110000",
  44822=>"000101010",
  44823=>"111000000",
  44824=>"001101010",
  44825=>"000100101",
  44826=>"101000000",
  44827=>"101110100",
  44828=>"001111001",
  44829=>"100010110",
  44830=>"111000101",
  44831=>"001110001",
  44832=>"110100111",
  44833=>"001001010",
  44834=>"010111110",
  44835=>"111011001",
  44836=>"000001011",
  44837=>"101100001",
  44838=>"100110010",
  44839=>"100111000",
  44840=>"001000101",
  44841=>"010100001",
  44842=>"111101011",
  44843=>"001010011",
  44844=>"001011001",
  44845=>"000000111",
  44846=>"111001100",
  44847=>"010111111",
  44848=>"000000000",
  44849=>"100011011",
  44850=>"110011111",
  44851=>"111111110",
  44852=>"101001110",
  44853=>"011001111",
  44854=>"000011011",
  44855=>"000011101",
  44856=>"110101110",
  44857=>"001011101",
  44858=>"010110010",
  44859=>"011000001",
  44860=>"000011010",
  44861=>"001110101",
  44862=>"011001100",
  44863=>"010111011",
  44864=>"111001010",
  44865=>"111101111",
  44866=>"001000111",
  44867=>"011011101",
  44868=>"000100000",
  44869=>"101010000",
  44870=>"110011010",
  44871=>"110111010",
  44872=>"010111001",
  44873=>"011111111",
  44874=>"100101011",
  44875=>"000000010",
  44876=>"011101000",
  44877=>"010110010",
  44878=>"010111010",
  44879=>"101001001",
  44880=>"111101111",
  44881=>"011101001",
  44882=>"110101011",
  44883=>"011001101",
  44884=>"101111001",
  44885=>"101001000",
  44886=>"111101101",
  44887=>"000010101",
  44888=>"000100001",
  44889=>"010110110",
  44890=>"010001001",
  44891=>"000100100",
  44892=>"111110110",
  44893=>"100001101",
  44894=>"110000001",
  44895=>"101100100",
  44896=>"000110001",
  44897=>"000111000",
  44898=>"010010111",
  44899=>"000110100",
  44900=>"010110010",
  44901=>"110000001",
  44902=>"100111100",
  44903=>"000001000",
  44904=>"100001000",
  44905=>"110000011",
  44906=>"110010011",
  44907=>"001101000",
  44908=>"010001100",
  44909=>"010111001",
  44910=>"111100010",
  44911=>"001000101",
  44912=>"010110110",
  44913=>"110111101",
  44914=>"111111100",
  44915=>"011000110",
  44916=>"110111100",
  44917=>"100001001",
  44918=>"101000011",
  44919=>"101100110",
  44920=>"111010111",
  44921=>"010010111",
  44922=>"000111011",
  44923=>"111111010",
  44924=>"001011011",
  44925=>"001101101",
  44926=>"011000011",
  44927=>"000110110",
  44928=>"001000101",
  44929=>"111101101",
  44930=>"010101011",
  44931=>"111111011",
  44932=>"010011000",
  44933=>"110011011",
  44934=>"001110001",
  44935=>"001010010",
  44936=>"010000100",
  44937=>"011011000",
  44938=>"100001011",
  44939=>"111011101",
  44940=>"111110101",
  44941=>"100010001",
  44942=>"110101101",
  44943=>"011001100",
  44944=>"100111011",
  44945=>"111001010",
  44946=>"001100101",
  44947=>"010110100",
  44948=>"001101010",
  44949=>"001101100",
  44950=>"101110000",
  44951=>"001010110",
  44952=>"001000100",
  44953=>"110100111",
  44954=>"111110011",
  44955=>"101101110",
  44956=>"111000001",
  44957=>"010100111",
  44958=>"000010111",
  44959=>"011110010",
  44960=>"000000100",
  44961=>"001101111",
  44962=>"001010101",
  44963=>"111011110",
  44964=>"100010101",
  44965=>"011001110",
  44966=>"111010110",
  44967=>"101001100",
  44968=>"111101011",
  44969=>"000010001",
  44970=>"000111011",
  44971=>"100000111",
  44972=>"110101010",
  44973=>"000000100",
  44974=>"100100100",
  44975=>"011111111",
  44976=>"111001000",
  44977=>"101011001",
  44978=>"000101111",
  44979=>"010000010",
  44980=>"001001101",
  44981=>"000000011",
  44982=>"010100010",
  44983=>"011111100",
  44984=>"100011010",
  44985=>"101011101",
  44986=>"111001111",
  44987=>"101110001",
  44988=>"001001000",
  44989=>"011000110",
  44990=>"000101100",
  44991=>"111110010",
  44992=>"000001000",
  44993=>"100001101",
  44994=>"000110000",
  44995=>"010000111",
  44996=>"111001010",
  44997=>"001001001",
  44998=>"000110101",
  44999=>"000111101",
  45000=>"110111111",
  45001=>"011100011",
  45002=>"010110110",
  45003=>"000000000",
  45004=>"111110011",
  45005=>"111001110",
  45006=>"110101010",
  45007=>"000100010",
  45008=>"101111000",
  45009=>"110011110",
  45010=>"111101011",
  45011=>"001001110",
  45012=>"000100011",
  45013=>"111100011",
  45014=>"011100000",
  45015=>"000100010",
  45016=>"011010100",
  45017=>"010110010",
  45018=>"011111111",
  45019=>"011011110",
  45020=>"101001100",
  45021=>"010000011",
  45022=>"111110101",
  45023=>"010100100",
  45024=>"000101111",
  45025=>"111010010",
  45026=>"001001001",
  45027=>"001001100",
  45028=>"001001001",
  45029=>"110000000",
  45030=>"100111110",
  45031=>"100100010",
  45032=>"001111000",
  45033=>"001000011",
  45034=>"100111000",
  45035=>"010100110",
  45036=>"100011001",
  45037=>"000110011",
  45038=>"010000000",
  45039=>"000010101",
  45040=>"001101101",
  45041=>"010001000",
  45042=>"100100100",
  45043=>"001101110",
  45044=>"011001011",
  45045=>"011000100",
  45046=>"000110001",
  45047=>"110000000",
  45048=>"000110101",
  45049=>"110100111",
  45050=>"111011111",
  45051=>"001101000",
  45052=>"011100101",
  45053=>"010111000",
  45054=>"001111000",
  45055=>"100100001",
  45056=>"111011011",
  45057=>"000001110",
  45058=>"111111000",
  45059=>"101010010",
  45060=>"101011111",
  45061=>"000110000",
  45062=>"011101001",
  45063=>"000001000",
  45064=>"101010011",
  45065=>"000100010",
  45066=>"001100010",
  45067=>"101000110",
  45068=>"011011000",
  45069=>"000000001",
  45070=>"100001001",
  45071=>"100100100",
  45072=>"000100111",
  45073=>"101010100",
  45074=>"110010101",
  45075=>"010110101",
  45076=>"110110000",
  45077=>"101111001",
  45078=>"100000101",
  45079=>"110010000",
  45080=>"111101011",
  45081=>"110100011",
  45082=>"011100010",
  45083=>"101010111",
  45084=>"101111111",
  45085=>"001110111",
  45086=>"010111110",
  45087=>"011100111",
  45088=>"111110010",
  45089=>"101111111",
  45090=>"000100111",
  45091=>"101100000",
  45092=>"111000001",
  45093=>"000110111",
  45094=>"111000100",
  45095=>"010010011",
  45096=>"010010011",
  45097=>"001110101",
  45098=>"101100011",
  45099=>"010010010",
  45100=>"001000101",
  45101=>"010000010",
  45102=>"001000010",
  45103=>"011110000",
  45104=>"101000111",
  45105=>"101011110",
  45106=>"001010000",
  45107=>"111111010",
  45108=>"100000101",
  45109=>"001001011",
  45110=>"110100010",
  45111=>"000111101",
  45112=>"111100101",
  45113=>"010010000",
  45114=>"000101001",
  45115=>"111110100",
  45116=>"111010000",
  45117=>"111010010",
  45118=>"010111000",
  45119=>"111101000",
  45120=>"011100110",
  45121=>"010011001",
  45122=>"010011000",
  45123=>"111001101",
  45124=>"010110100",
  45125=>"111111011",
  45126=>"101000100",
  45127=>"001001001",
  45128=>"101000001",
  45129=>"001001000",
  45130=>"110011110",
  45131=>"111000010",
  45132=>"000001101",
  45133=>"101111011",
  45134=>"010001111",
  45135=>"111001001",
  45136=>"000101001",
  45137=>"110010110",
  45138=>"110110000",
  45139=>"011010011",
  45140=>"001010100",
  45141=>"100000011",
  45142=>"000101101",
  45143=>"001111001",
  45144=>"111010000",
  45145=>"110101111",
  45146=>"110010100",
  45147=>"110010100",
  45148=>"000111001",
  45149=>"110100010",
  45150=>"010010110",
  45151=>"100111110",
  45152=>"010100001",
  45153=>"000000111",
  45154=>"000011111",
  45155=>"011010011",
  45156=>"000111001",
  45157=>"001001111",
  45158=>"001010010",
  45159=>"111111100",
  45160=>"111001011",
  45161=>"001010111",
  45162=>"001001011",
  45163=>"010011000",
  45164=>"101001001",
  45165=>"001000110",
  45166=>"011111100",
  45167=>"111100111",
  45168=>"111001000",
  45169=>"011001010",
  45170=>"111010000",
  45171=>"111000100",
  45172=>"011010010",
  45173=>"100111000",
  45174=>"001011001",
  45175=>"110001110",
  45176=>"000111111",
  45177=>"101010000",
  45178=>"100100011",
  45179=>"101011100",
  45180=>"001001110",
  45181=>"011010100",
  45182=>"111000010",
  45183=>"111000100",
  45184=>"110001001",
  45185=>"010111000",
  45186=>"000101001",
  45187=>"000101110",
  45188=>"111010100",
  45189=>"111001001",
  45190=>"000010000",
  45191=>"000010100",
  45192=>"000110010",
  45193=>"000101011",
  45194=>"010010000",
  45195=>"001001110",
  45196=>"101001101",
  45197=>"001101010",
  45198=>"011101101",
  45199=>"011011011",
  45200=>"001000000",
  45201=>"100011111",
  45202=>"000000001",
  45203=>"010001011",
  45204=>"000110100",
  45205=>"011001110",
  45206=>"011011100",
  45207=>"101100110",
  45208=>"000010000",
  45209=>"001111001",
  45210=>"111011000",
  45211=>"011000010",
  45212=>"101001101",
  45213=>"111100000",
  45214=>"010010000",
  45215=>"001101000",
  45216=>"000110100",
  45217=>"101100000",
  45218=>"110101111",
  45219=>"000110001",
  45220=>"100111111",
  45221=>"100001001",
  45222=>"101100101",
  45223=>"110100000",
  45224=>"111011110",
  45225=>"000110011",
  45226=>"000000100",
  45227=>"101101110",
  45228=>"110001111",
  45229=>"110001100",
  45230=>"001100000",
  45231=>"101010011",
  45232=>"100000010",
  45233=>"101000100",
  45234=>"111011010",
  45235=>"100001101",
  45236=>"110011111",
  45237=>"011001000",
  45238=>"111001000",
  45239=>"001000100",
  45240=>"000000101",
  45241=>"100101101",
  45242=>"010000001",
  45243=>"011101101",
  45244=>"001000101",
  45245=>"110001110",
  45246=>"110001111",
  45247=>"111101001",
  45248=>"001011001",
  45249=>"111100011",
  45250=>"111100110",
  45251=>"001011110",
  45252=>"010010110",
  45253=>"000010001",
  45254=>"101110111",
  45255=>"011100010",
  45256=>"000100100",
  45257=>"101110010",
  45258=>"110001110",
  45259=>"011100101",
  45260=>"101110001",
  45261=>"010100110",
  45262=>"111111100",
  45263=>"010000010",
  45264=>"101111110",
  45265=>"101010110",
  45266=>"101000111",
  45267=>"111000110",
  45268=>"011001001",
  45269=>"110001100",
  45270=>"010001001",
  45271=>"001011010",
  45272=>"101100100",
  45273=>"001110110",
  45274=>"101111010",
  45275=>"110111001",
  45276=>"010101010",
  45277=>"010000111",
  45278=>"011100000",
  45279=>"101100101",
  45280=>"010000100",
  45281=>"010100001",
  45282=>"101101110",
  45283=>"011100010",
  45284=>"111110100",
  45285=>"100101101",
  45286=>"111010101",
  45287=>"011110010",
  45288=>"000101000",
  45289=>"110111011",
  45290=>"100111001",
  45291=>"000111001",
  45292=>"110001001",
  45293=>"001100111",
  45294=>"001010110",
  45295=>"101000011",
  45296=>"001100011",
  45297=>"111001011",
  45298=>"111110001",
  45299=>"100010001",
  45300=>"111000011",
  45301=>"110101001",
  45302=>"000001110",
  45303=>"001001110",
  45304=>"010010101",
  45305=>"111100101",
  45306=>"000111011",
  45307=>"000000101",
  45308=>"000011011",
  45309=>"000100001",
  45310=>"010111010",
  45311=>"001100110",
  45312=>"111001000",
  45313=>"100001101",
  45314=>"001010110",
  45315=>"011001111",
  45316=>"101011000",
  45317=>"111111011",
  45318=>"111110100",
  45319=>"000100101",
  45320=>"001100010",
  45321=>"001111011",
  45322=>"011110110",
  45323=>"111111100",
  45324=>"001010001",
  45325=>"001100101",
  45326=>"000010111",
  45327=>"001010101",
  45328=>"111110111",
  45329=>"100000010",
  45330=>"110010000",
  45331=>"011100110",
  45332=>"011100011",
  45333=>"101110101",
  45334=>"001100100",
  45335=>"101100101",
  45336=>"100011010",
  45337=>"110111101",
  45338=>"011011111",
  45339=>"000011111",
  45340=>"000101000",
  45341=>"111010110",
  45342=>"011001000",
  45343=>"000100000",
  45344=>"100001111",
  45345=>"010000001",
  45346=>"100101000",
  45347=>"000100010",
  45348=>"111000110",
  45349=>"011100000",
  45350=>"001110010",
  45351=>"111111111",
  45352=>"110001010",
  45353=>"000111110",
  45354=>"001010001",
  45355=>"111111111",
  45356=>"101101010",
  45357=>"111011010",
  45358=>"010000000",
  45359=>"100010010",
  45360=>"110001100",
  45361=>"110000101",
  45362=>"111111111",
  45363=>"110110010",
  45364=>"101000000",
  45365=>"001010000",
  45366=>"010100001",
  45367=>"000101000",
  45368=>"110001101",
  45369=>"001111110",
  45370=>"101110101",
  45371=>"011100010",
  45372=>"101000001",
  45373=>"100110000",
  45374=>"110100110",
  45375=>"110001000",
  45376=>"001001100",
  45377=>"011110100",
  45378=>"010101110",
  45379=>"011100000",
  45380=>"111100011",
  45381=>"101010001",
  45382=>"001101001",
  45383=>"000111011",
  45384=>"010000101",
  45385=>"000000100",
  45386=>"111001011",
  45387=>"001000110",
  45388=>"111110111",
  45389=>"100000101",
  45390=>"110101000",
  45391=>"001100011",
  45392=>"011001110",
  45393=>"111001111",
  45394=>"000110010",
  45395=>"010001100",
  45396=>"011101001",
  45397=>"101000101",
  45398=>"100010100",
  45399=>"010000001",
  45400=>"100100010",
  45401=>"111110110",
  45402=>"000111000",
  45403=>"000001010",
  45404=>"010111110",
  45405=>"110100110",
  45406=>"110100000",
  45407=>"010011010",
  45408=>"001010000",
  45409=>"100010010",
  45410=>"101100011",
  45411=>"101001111",
  45412=>"101001101",
  45413=>"101111111",
  45414=>"000001000",
  45415=>"001110000",
  45416=>"101110010",
  45417=>"000010100",
  45418=>"001101101",
  45419=>"010110000",
  45420=>"001000011",
  45421=>"111110101",
  45422=>"000100000",
  45423=>"011011000",
  45424=>"010101100",
  45425=>"111001101",
  45426=>"100001111",
  45427=>"010101111",
  45428=>"010110110",
  45429=>"010011010",
  45430=>"011100111",
  45431=>"101110111",
  45432=>"101111010",
  45433=>"100101100",
  45434=>"001110000",
  45435=>"101110110",
  45436=>"000100101",
  45437=>"111100000",
  45438=>"001101111",
  45439=>"111011000",
  45440=>"110100100",
  45441=>"101110100",
  45442=>"010111101",
  45443=>"011111010",
  45444=>"000101001",
  45445=>"001110110",
  45446=>"000110001",
  45447=>"010110110",
  45448=>"000000001",
  45449=>"111100010",
  45450=>"001110000",
  45451=>"010100101",
  45452=>"111111110",
  45453=>"111000110",
  45454=>"000100110",
  45455=>"110010111",
  45456=>"001001001",
  45457=>"101101010",
  45458=>"001111000",
  45459=>"000010101",
  45460=>"001100000",
  45461=>"001010010",
  45462=>"101011010",
  45463=>"101011010",
  45464=>"001100000",
  45465=>"001100001",
  45466=>"001100001",
  45467=>"111111100",
  45468=>"011000110",
  45469=>"011010110",
  45470=>"001010101",
  45471=>"100111101",
  45472=>"001101000",
  45473=>"110110001",
  45474=>"101111100",
  45475=>"000000000",
  45476=>"100011010",
  45477=>"001000011",
  45478=>"110111000",
  45479=>"011001011",
  45480=>"100100111",
  45481=>"110000000",
  45482=>"100110111",
  45483=>"110010011",
  45484=>"100010100",
  45485=>"100000111",
  45486=>"100010111",
  45487=>"000101011",
  45488=>"000000110",
  45489=>"010011110",
  45490=>"111111000",
  45491=>"110011001",
  45492=>"100011010",
  45493=>"000100011",
  45494=>"000001111",
  45495=>"010000111",
  45496=>"000001011",
  45497=>"101100100",
  45498=>"110111100",
  45499=>"001110010",
  45500=>"000010011",
  45501=>"001001001",
  45502=>"010100111",
  45503=>"111011111",
  45504=>"001001010",
  45505=>"100110100",
  45506=>"110110010",
  45507=>"010110001",
  45508=>"000000001",
  45509=>"110110111",
  45510=>"111010011",
  45511=>"000101000",
  45512=>"110001110",
  45513=>"101011001",
  45514=>"101000001",
  45515=>"110000010",
  45516=>"001001011",
  45517=>"101000011",
  45518=>"110111010",
  45519=>"101100100",
  45520=>"000001010",
  45521=>"000100110",
  45522=>"100111111",
  45523=>"000100111",
  45524=>"111111011",
  45525=>"111001110",
  45526=>"010110001",
  45527=>"101010100",
  45528=>"111010110",
  45529=>"110010011",
  45530=>"010000110",
  45531=>"011101100",
  45532=>"000110011",
  45533=>"000000010",
  45534=>"010001011",
  45535=>"110010101",
  45536=>"111011111",
  45537=>"111000010",
  45538=>"010111010",
  45539=>"011100010",
  45540=>"001000011",
  45541=>"101000100",
  45542=>"000011101",
  45543=>"000001011",
  45544=>"101111010",
  45545=>"000111110",
  45546=>"011000101",
  45547=>"100100010",
  45548=>"011001110",
  45549=>"111100000",
  45550=>"101000100",
  45551=>"101100111",
  45552=>"011111011",
  45553=>"101100000",
  45554=>"100001100",
  45555=>"010001001",
  45556=>"101101000",
  45557=>"011111111",
  45558=>"110100010",
  45559=>"100001110",
  45560=>"110101010",
  45561=>"010001001",
  45562=>"001111101",
  45563=>"000000101",
  45564=>"010101010",
  45565=>"100110000",
  45566=>"011100010",
  45567=>"101010000",
  45568=>"110100100",
  45569=>"011000000",
  45570=>"000100001",
  45571=>"110000111",
  45572=>"010011100",
  45573=>"110000011",
  45574=>"001001110",
  45575=>"101101100",
  45576=>"111010100",
  45577=>"010000001",
  45578=>"100001011",
  45579=>"101101111",
  45580=>"110001000",
  45581=>"101101100",
  45582=>"000110111",
  45583=>"110100110",
  45584=>"001000010",
  45585=>"011010010",
  45586=>"110001100",
  45587=>"011001010",
  45588=>"001101001",
  45589=>"000100111",
  45590=>"000010001",
  45591=>"001011011",
  45592=>"110001111",
  45593=>"111010000",
  45594=>"010011001",
  45595=>"111001010",
  45596=>"110111001",
  45597=>"100111011",
  45598=>"110001000",
  45599=>"011011000",
  45600=>"010010011",
  45601=>"011000011",
  45602=>"011011011",
  45603=>"100100001",
  45604=>"111000001",
  45605=>"001100111",
  45606=>"111101111",
  45607=>"010000110",
  45608=>"110101001",
  45609=>"111010011",
  45610=>"110010110",
  45611=>"100000111",
  45612=>"001101111",
  45613=>"110011000",
  45614=>"000101001",
  45615=>"011110111",
  45616=>"000101011",
  45617=>"011101010",
  45618=>"110101111",
  45619=>"100011111",
  45620=>"010010110",
  45621=>"110110010",
  45622=>"001100011",
  45623=>"100011111",
  45624=>"111100001",
  45625=>"001001000",
  45626=>"001001010",
  45627=>"001110011",
  45628=>"111111000",
  45629=>"101110110",
  45630=>"010001010",
  45631=>"000100010",
  45632=>"010111111",
  45633=>"000100010",
  45634=>"110000101",
  45635=>"001011111",
  45636=>"000111000",
  45637=>"101101010",
  45638=>"000001011",
  45639=>"000111010",
  45640=>"110101101",
  45641=>"110101010",
  45642=>"100100111",
  45643=>"100110111",
  45644=>"011101011",
  45645=>"010011101",
  45646=>"101000100",
  45647=>"110001001",
  45648=>"101101010",
  45649=>"111001110",
  45650=>"000100110",
  45651=>"100000110",
  45652=>"001000000",
  45653=>"110100111",
  45654=>"011010110",
  45655=>"110100110",
  45656=>"010101100",
  45657=>"000101100",
  45658=>"110010010",
  45659=>"110110111",
  45660=>"101100100",
  45661=>"101010100",
  45662=>"110001111",
  45663=>"010000000",
  45664=>"011111011",
  45665=>"001100101",
  45666=>"110000111",
  45667=>"111001110",
  45668=>"110011001",
  45669=>"001110001",
  45670=>"010101011",
  45671=>"001100110",
  45672=>"011111111",
  45673=>"110110111",
  45674=>"000011001",
  45675=>"110101000",
  45676=>"100000100",
  45677=>"011100111",
  45678=>"111000101",
  45679=>"011001111",
  45680=>"011011001",
  45681=>"111010111",
  45682=>"000101101",
  45683=>"001110000",
  45684=>"001100000",
  45685=>"110000111",
  45686=>"001010100",
  45687=>"011010110",
  45688=>"011111101",
  45689=>"100011000",
  45690=>"000100101",
  45691=>"000110011",
  45692=>"101000000",
  45693=>"010001101",
  45694=>"110111101",
  45695=>"011100101",
  45696=>"010000010",
  45697=>"111000110",
  45698=>"011110010",
  45699=>"101111010",
  45700=>"001000011",
  45701=>"001110110",
  45702=>"101000011",
  45703=>"111110110",
  45704=>"100101011",
  45705=>"100010000",
  45706=>"100100111",
  45707=>"011110100",
  45708=>"100010000",
  45709=>"000100011",
  45710=>"010110101",
  45711=>"011000110",
  45712=>"010001100",
  45713=>"001110010",
  45714=>"110100111",
  45715=>"100101011",
  45716=>"011000011",
  45717=>"000011100",
  45718=>"101000011",
  45719=>"001001101",
  45720=>"010011101",
  45721=>"011010000",
  45722=>"111111011",
  45723=>"110011100",
  45724=>"001111001",
  45725=>"011100011",
  45726=>"101110100",
  45727=>"110001111",
  45728=>"100001100",
  45729=>"001100010",
  45730=>"010010000",
  45731=>"010111010",
  45732=>"110111111",
  45733=>"111000000",
  45734=>"010000111",
  45735=>"001010110",
  45736=>"111000010",
  45737=>"010100100",
  45738=>"100000100",
  45739=>"001010111",
  45740=>"011001010",
  45741=>"101101000",
  45742=>"100011110",
  45743=>"011010000",
  45744=>"100110010",
  45745=>"100110000",
  45746=>"100100110",
  45747=>"010001101",
  45748=>"101001011",
  45749=>"001011110",
  45750=>"010010111",
  45751=>"101100010",
  45752=>"000110100",
  45753=>"111110001",
  45754=>"011110101",
  45755=>"110011000",
  45756=>"100100000",
  45757=>"010000011",
  45758=>"000001100",
  45759=>"110100110",
  45760=>"001000111",
  45761=>"100110101",
  45762=>"000111110",
  45763=>"010010010",
  45764=>"101000111",
  45765=>"110001010",
  45766=>"011101110",
  45767=>"010001011",
  45768=>"101100010",
  45769=>"000000000",
  45770=>"010011100",
  45771=>"001100010",
  45772=>"100000111",
  45773=>"010111111",
  45774=>"000011001",
  45775=>"110100011",
  45776=>"111110101",
  45777=>"011001011",
  45778=>"101011011",
  45779=>"010001000",
  45780=>"010101000",
  45781=>"101000001",
  45782=>"111111011",
  45783=>"011001110",
  45784=>"110111100",
  45785=>"011011111",
  45786=>"011111100",
  45787=>"100100001",
  45788=>"011011101",
  45789=>"110010011",
  45790=>"110101101",
  45791=>"101101011",
  45792=>"111101011",
  45793=>"011010111",
  45794=>"011010001",
  45795=>"011011011",
  45796=>"100101010",
  45797=>"000000111",
  45798=>"010100001",
  45799=>"111011100",
  45800=>"111100000",
  45801=>"001101001",
  45802=>"001000111",
  45803=>"110101111",
  45804=>"111110101",
  45805=>"001010010",
  45806=>"111010000",
  45807=>"000010100",
  45808=>"110001000",
  45809=>"001001000",
  45810=>"111000101",
  45811=>"110101011",
  45812=>"000101111",
  45813=>"001101101",
  45814=>"101011100",
  45815=>"010000011",
  45816=>"111111110",
  45817=>"011111100",
  45818=>"011001011",
  45819=>"101000100",
  45820=>"111101111",
  45821=>"000111010",
  45822=>"101011100",
  45823=>"100110110",
  45824=>"001001010",
  45825=>"000010000",
  45826=>"001001101",
  45827=>"010100001",
  45828=>"101001011",
  45829=>"111101001",
  45830=>"011101001",
  45831=>"000000111",
  45832=>"000100000",
  45833=>"111010001",
  45834=>"011000000",
  45835=>"000010100",
  45836=>"011010110",
  45837=>"011110010",
  45838=>"101001010",
  45839=>"010010101",
  45840=>"001000101",
  45841=>"011111010",
  45842=>"100001111",
  45843=>"011111100",
  45844=>"101101010",
  45845=>"010010101",
  45846=>"111010010",
  45847=>"011100000",
  45848=>"101011001",
  45849=>"000000010",
  45850=>"010101010",
  45851=>"101110011",
  45852=>"001011000",
  45853=>"011011011",
  45854=>"011010100",
  45855=>"100001011",
  45856=>"100100100",
  45857=>"000000111",
  45858=>"000101000",
  45859=>"011000100",
  45860=>"001000110",
  45861=>"111101101",
  45862=>"100110001",
  45863=>"110001010",
  45864=>"110001000",
  45865=>"010011000",
  45866=>"110100010",
  45867=>"010011110",
  45868=>"010011101",
  45869=>"011110100",
  45870=>"011111100",
  45871=>"011001010",
  45872=>"011100111",
  45873=>"010001011",
  45874=>"001111000",
  45875=>"011101001",
  45876=>"111111111",
  45877=>"010011110",
  45878=>"101110100",
  45879=>"000000100",
  45880=>"111000000",
  45881=>"101010101",
  45882=>"010000100",
  45883=>"101011111",
  45884=>"000101100",
  45885=>"111100110",
  45886=>"001100000",
  45887=>"000010111",
  45888=>"010011110",
  45889=>"010111111",
  45890=>"100101111",
  45891=>"000000001",
  45892=>"001000001",
  45893=>"111101001",
  45894=>"100011011",
  45895=>"000000111",
  45896=>"101100011",
  45897=>"001010011",
  45898=>"111001100",
  45899=>"100000010",
  45900=>"100010010",
  45901=>"001001010",
  45902=>"010111101",
  45903=>"110000000",
  45904=>"111100100",
  45905=>"110101011",
  45906=>"011000000",
  45907=>"101000101",
  45908=>"011101001",
  45909=>"000101010",
  45910=>"001000001",
  45911=>"101000101",
  45912=>"001100001",
  45913=>"100110110",
  45914=>"110011101",
  45915=>"011010010",
  45916=>"011110110",
  45917=>"011010100",
  45918=>"000101111",
  45919=>"110100111",
  45920=>"010100011",
  45921=>"100100101",
  45922=>"111110111",
  45923=>"000010100",
  45924=>"101100111",
  45925=>"111001100",
  45926=>"010111110",
  45927=>"001111101",
  45928=>"101011000",
  45929=>"111000011",
  45930=>"010011111",
  45931=>"000000100",
  45932=>"000000100",
  45933=>"010010001",
  45934=>"001000010",
  45935=>"011100000",
  45936=>"000100100",
  45937=>"010110111",
  45938=>"101011101",
  45939=>"100010100",
  45940=>"000000100",
  45941=>"001111100",
  45942=>"111010011",
  45943=>"011110111",
  45944=>"101101101",
  45945=>"101011011",
  45946=>"011101100",
  45947=>"100001000",
  45948=>"010111111",
  45949=>"110100010",
  45950=>"010011000",
  45951=>"100010111",
  45952=>"011101101",
  45953=>"010100011",
  45954=>"001000101",
  45955=>"010101100",
  45956=>"000100001",
  45957=>"111110001",
  45958=>"111101001",
  45959=>"000001001",
  45960=>"010001011",
  45961=>"011100010",
  45962=>"100111111",
  45963=>"010001001",
  45964=>"101010011",
  45965=>"101011100",
  45966=>"011001001",
  45967=>"110110100",
  45968=>"111100101",
  45969=>"101011011",
  45970=>"000001111",
  45971=>"100000000",
  45972=>"111001001",
  45973=>"011011001",
  45974=>"001110111",
  45975=>"101101010",
  45976=>"000111011",
  45977=>"011101000",
  45978=>"111011000",
  45979=>"101111010",
  45980=>"100000100",
  45981=>"011000101",
  45982=>"100101000",
  45983=>"001100011",
  45984=>"101101000",
  45985=>"000110010",
  45986=>"101111111",
  45987=>"110000101",
  45988=>"100110010",
  45989=>"011100001",
  45990=>"100011100",
  45991=>"000111110",
  45992=>"111000001",
  45993=>"001101101",
  45994=>"101100011",
  45995=>"100000111",
  45996=>"011100010",
  45997=>"111011010",
  45998=>"011000110",
  45999=>"001011001",
  46000=>"011001011",
  46001=>"001011010",
  46002=>"111110111",
  46003=>"001000011",
  46004=>"000100111",
  46005=>"111000010",
  46006=>"111011100",
  46007=>"000111101",
  46008=>"000010000",
  46009=>"000010010",
  46010=>"011010100",
  46011=>"011001101",
  46012=>"100001011",
  46013=>"110000110",
  46014=>"101010000",
  46015=>"000110111",
  46016=>"000101011",
  46017=>"010011000",
  46018=>"111010010",
  46019=>"000010111",
  46020=>"100001110",
  46021=>"001100011",
  46022=>"100111111",
  46023=>"010100001",
  46024=>"011100101",
  46025=>"000100001",
  46026=>"111000101",
  46027=>"100101010",
  46028=>"000101001",
  46029=>"111001101",
  46030=>"000000011",
  46031=>"001011110",
  46032=>"011000101",
  46033=>"000010101",
  46034=>"101001011",
  46035=>"011111011",
  46036=>"001101011",
  46037=>"101010111",
  46038=>"010011000",
  46039=>"101000100",
  46040=>"101110111",
  46041=>"111000000",
  46042=>"000000001",
  46043=>"110001010",
  46044=>"010001100",
  46045=>"110101000",
  46046=>"000001110",
  46047=>"000010100",
  46048=>"011010110",
  46049=>"111111001",
  46050=>"001110111",
  46051=>"000011001",
  46052=>"000000111",
  46053=>"100011100",
  46054=>"110101110",
  46055=>"111000100",
  46056=>"000000010",
  46057=>"110101000",
  46058=>"101110001",
  46059=>"100100100",
  46060=>"010001110",
  46061=>"101101010",
  46062=>"101110111",
  46063=>"011010000",
  46064=>"010000110",
  46065=>"011001111",
  46066=>"010110110",
  46067=>"101010010",
  46068=>"111111101",
  46069=>"111100011",
  46070=>"111000100",
  46071=>"000111111",
  46072=>"011000100",
  46073=>"110111100",
  46074=>"110001111",
  46075=>"111000010",
  46076=>"000100001",
  46077=>"011011010",
  46078=>"110101111",
  46079=>"000011011",
  46080=>"000000111",
  46081=>"001010110",
  46082=>"001110101",
  46083=>"001011000",
  46084=>"101000111",
  46085=>"000110000",
  46086=>"100011000",
  46087=>"011101010",
  46088=>"111010110",
  46089=>"001111101",
  46090=>"111011000",
  46091=>"011101010",
  46092=>"110110001",
  46093=>"000001001",
  46094=>"110001110",
  46095=>"001000000",
  46096=>"011000000",
  46097=>"011011011",
  46098=>"001000000",
  46099=>"101110111",
  46100=>"001000011",
  46101=>"110111001",
  46102=>"101110111",
  46103=>"000111101",
  46104=>"100110001",
  46105=>"011001101",
  46106=>"010010001",
  46107=>"111011110",
  46108=>"111011011",
  46109=>"110110010",
  46110=>"011001100",
  46111=>"111001011",
  46112=>"110110101",
  46113=>"000010110",
  46114=>"011100100",
  46115=>"001110111",
  46116=>"001100010",
  46117=>"110111011",
  46118=>"100010100",
  46119=>"111110001",
  46120=>"110111101",
  46121=>"101110001",
  46122=>"110011000",
  46123=>"001001000",
  46124=>"001011100",
  46125=>"110111000",
  46126=>"000111110",
  46127=>"000110010",
  46128=>"111000100",
  46129=>"110011000",
  46130=>"111110011",
  46131=>"100010111",
  46132=>"100001000",
  46133=>"111010100",
  46134=>"101100001",
  46135=>"111011011",
  46136=>"101100001",
  46137=>"101000010",
  46138=>"010001101",
  46139=>"000010011",
  46140=>"101101001",
  46141=>"001011111",
  46142=>"110110100",
  46143=>"000000100",
  46144=>"111011001",
  46145=>"101000111",
  46146=>"100111111",
  46147=>"010111001",
  46148=>"000110010",
  46149=>"001000011",
  46150=>"011000111",
  46151=>"001111100",
  46152=>"010111011",
  46153=>"001101101",
  46154=>"111100011",
  46155=>"010101011",
  46156=>"110001101",
  46157=>"100000110",
  46158=>"000100000",
  46159=>"101011111",
  46160=>"010001111",
  46161=>"011111110",
  46162=>"100101110",
  46163=>"101110111",
  46164=>"011001111",
  46165=>"101101101",
  46166=>"010010000",
  46167=>"100111011",
  46168=>"010101011",
  46169=>"110111111",
  46170=>"000110101",
  46171=>"011100011",
  46172=>"000001010",
  46173=>"011111100",
  46174=>"011001101",
  46175=>"011111000",
  46176=>"001111011",
  46177=>"111011011",
  46178=>"010101111",
  46179=>"001110100",
  46180=>"010110110",
  46181=>"101101101",
  46182=>"011010101",
  46183=>"001011100",
  46184=>"000010011",
  46185=>"101111010",
  46186=>"111010001",
  46187=>"110110010",
  46188=>"011110110",
  46189=>"001111100",
  46190=>"110000000",
  46191=>"000010101",
  46192=>"001001001",
  46193=>"110001000",
  46194=>"101101001",
  46195=>"010000101",
  46196=>"101100101",
  46197=>"111100000",
  46198=>"000010110",
  46199=>"111100000",
  46200=>"100111000",
  46201=>"000111101",
  46202=>"000110011",
  46203=>"001101110",
  46204=>"111100010",
  46205=>"111110100",
  46206=>"111010100",
  46207=>"101111001",
  46208=>"101111011",
  46209=>"111101110",
  46210=>"111101111",
  46211=>"001101111",
  46212=>"001110111",
  46213=>"001000100",
  46214=>"111110110",
  46215=>"010010111",
  46216=>"100000101",
  46217=>"101110110",
  46218=>"001000011",
  46219=>"101010001",
  46220=>"110000100",
  46221=>"011010100",
  46222=>"001000001",
  46223=>"011111011",
  46224=>"110011100",
  46225=>"100001001",
  46226=>"010011010",
  46227=>"101011011",
  46228=>"111110010",
  46229=>"011000100",
  46230=>"001100111",
  46231=>"001111110",
  46232=>"100010100",
  46233=>"010001010",
  46234=>"100011011",
  46235=>"001001001",
  46236=>"101111111",
  46237=>"000110100",
  46238=>"001010100",
  46239=>"111001010",
  46240=>"101000011",
  46241=>"111100101",
  46242=>"111100111",
  46243=>"010001010",
  46244=>"011101101",
  46245=>"101111110",
  46246=>"100001110",
  46247=>"000010111",
  46248=>"000100100",
  46249=>"001110001",
  46250=>"100011100",
  46251=>"011010110",
  46252=>"011000000",
  46253=>"001001110",
  46254=>"111010000",
  46255=>"010010000",
  46256=>"110101001",
  46257=>"101010110",
  46258=>"010100111",
  46259=>"000110100",
  46260=>"001001101",
  46261=>"101101111",
  46262=>"110110001",
  46263=>"000100001",
  46264=>"010100100",
  46265=>"100101101",
  46266=>"000010100",
  46267=>"010110111",
  46268=>"101000010",
  46269=>"010011000",
  46270=>"001101001",
  46271=>"100001010",
  46272=>"001100110",
  46273=>"110000101",
  46274=>"001110001",
  46275=>"000000100",
  46276=>"100111010",
  46277=>"010011011",
  46278=>"001100101",
  46279=>"111010000",
  46280=>"011000100",
  46281=>"100111111",
  46282=>"101010010",
  46283=>"100100111",
  46284=>"011111101",
  46285=>"111101111",
  46286=>"001011010",
  46287=>"101101010",
  46288=>"010100010",
  46289=>"000101001",
  46290=>"010101001",
  46291=>"111110010",
  46292=>"000100101",
  46293=>"110000110",
  46294=>"011110000",
  46295=>"011001011",
  46296=>"110010110",
  46297=>"111011111",
  46298=>"001010101",
  46299=>"101101110",
  46300=>"100011000",
  46301=>"111000001",
  46302=>"001110000",
  46303=>"010000010",
  46304=>"010010010",
  46305=>"011101101",
  46306=>"111010001",
  46307=>"110000001",
  46308=>"011111011",
  46309=>"010101011",
  46310=>"100010010",
  46311=>"101110000",
  46312=>"001000001",
  46313=>"010101001",
  46314=>"011011100",
  46315=>"111010111",
  46316=>"001100001",
  46317=>"100000111",
  46318=>"111001101",
  46319=>"101111001",
  46320=>"111100101",
  46321=>"100111111",
  46322=>"010111000",
  46323=>"100001010",
  46324=>"101001001",
  46325=>"111111000",
  46326=>"000000111",
  46327=>"100111011",
  46328=>"000010010",
  46329=>"101100001",
  46330=>"110010110",
  46331=>"001001011",
  46332=>"011100001",
  46333=>"111101101",
  46334=>"110010111",
  46335=>"100111110",
  46336=>"011110111",
  46337=>"001101100",
  46338=>"101111101",
  46339=>"110110011",
  46340=>"101000101",
  46341=>"000010000",
  46342=>"010101101",
  46343=>"100110011",
  46344=>"110100100",
  46345=>"010010001",
  46346=>"001100010",
  46347=>"100111111",
  46348=>"110111000",
  46349=>"100011011",
  46350=>"111110101",
  46351=>"100010011",
  46352=>"000011100",
  46353=>"100110011",
  46354=>"010000000",
  46355=>"111011111",
  46356=>"111101011",
  46357=>"001110010",
  46358=>"000010001",
  46359=>"101000001",
  46360=>"001010111",
  46361=>"011011101",
  46362=>"101000010",
  46363=>"001000100",
  46364=>"100000100",
  46365=>"101000011",
  46366=>"011111111",
  46367=>"010010110",
  46368=>"011000010",
  46369=>"001000100",
  46370=>"111011111",
  46371=>"111011111",
  46372=>"111001100",
  46373=>"110101111",
  46374=>"001010000",
  46375=>"111110011",
  46376=>"111001000",
  46377=>"111111011",
  46378=>"001101011",
  46379=>"101000001",
  46380=>"000001000",
  46381=>"010111110",
  46382=>"101100010",
  46383=>"101100010",
  46384=>"110011111",
  46385=>"010011000",
  46386=>"110010111",
  46387=>"110010000",
  46388=>"010100011",
  46389=>"000011011",
  46390=>"000010111",
  46391=>"011111110",
  46392=>"111111110",
  46393=>"101010110",
  46394=>"110101110",
  46395=>"011000101",
  46396=>"000010000",
  46397=>"010111101",
  46398=>"000010011",
  46399=>"011011111",
  46400=>"111111110",
  46401=>"100101010",
  46402=>"010100101",
  46403=>"111000110",
  46404=>"011101110",
  46405=>"010010110",
  46406=>"101100001",
  46407=>"100101001",
  46408=>"010100110",
  46409=>"101000010",
  46410=>"111001010",
  46411=>"110111001",
  46412=>"010001001",
  46413=>"111111111",
  46414=>"101110010",
  46415=>"011101010",
  46416=>"010000100",
  46417=>"111111011",
  46418=>"111011111",
  46419=>"100100011",
  46420=>"111101101",
  46421=>"111110011",
  46422=>"110101100",
  46423=>"010100000",
  46424=>"101111000",
  46425=>"011010100",
  46426=>"000001010",
  46427=>"010000010",
  46428=>"001000011",
  46429=>"110100110",
  46430=>"011110101",
  46431=>"011111000",
  46432=>"111000011",
  46433=>"010001011",
  46434=>"111000110",
  46435=>"111101101",
  46436=>"010100111",
  46437=>"110100010",
  46438=>"001000111",
  46439=>"001011011",
  46440=>"101000111",
  46441=>"010000100",
  46442=>"100101111",
  46443=>"001110000",
  46444=>"100100010",
  46445=>"000010011",
  46446=>"000100000",
  46447=>"011101000",
  46448=>"011010101",
  46449=>"001011111",
  46450=>"000111010",
  46451=>"010111000",
  46452=>"010100000",
  46453=>"110001110",
  46454=>"000011101",
  46455=>"111001111",
  46456=>"110011100",
  46457=>"001101110",
  46458=>"111000010",
  46459=>"010010011",
  46460=>"010000101",
  46461=>"111010111",
  46462=>"100001001",
  46463=>"001010111",
  46464=>"111101100",
  46465=>"110010011",
  46466=>"110101010",
  46467=>"010111111",
  46468=>"010010011",
  46469=>"100010101",
  46470=>"110111010",
  46471=>"100101010",
  46472=>"000110101",
  46473=>"010110010",
  46474=>"011010011",
  46475=>"011111110",
  46476=>"000000001",
  46477=>"000100111",
  46478=>"100111001",
  46479=>"101100001",
  46480=>"010000101",
  46481=>"111011000",
  46482=>"011101110",
  46483=>"011000011",
  46484=>"101111001",
  46485=>"010010010",
  46486=>"001001101",
  46487=>"000101011",
  46488=>"011011100",
  46489=>"110010111",
  46490=>"111110011",
  46491=>"100000010",
  46492=>"111000001",
  46493=>"001000111",
  46494=>"011111010",
  46495=>"101110001",
  46496=>"101000000",
  46497=>"011000110",
  46498=>"001010000",
  46499=>"000101001",
  46500=>"100111100",
  46501=>"010000011",
  46502=>"011110110",
  46503=>"101100101",
  46504=>"111111000",
  46505=>"011110000",
  46506=>"101100111",
  46507=>"011001001",
  46508=>"001010100",
  46509=>"111111110",
  46510=>"110001011",
  46511=>"010100111",
  46512=>"100111101",
  46513=>"110101110",
  46514=>"010001010",
  46515=>"000001011",
  46516=>"000111100",
  46517=>"111001001",
  46518=>"100011101",
  46519=>"111110001",
  46520=>"001011111",
  46521=>"010110010",
  46522=>"001010101",
  46523=>"100110110",
  46524=>"010001101",
  46525=>"111110011",
  46526=>"000001111",
  46527=>"001110111",
  46528=>"100001010",
  46529=>"000101000",
  46530=>"011100111",
  46531=>"001001110",
  46532=>"010110111",
  46533=>"101100101",
  46534=>"110001010",
  46535=>"011000010",
  46536=>"110110101",
  46537=>"011101010",
  46538=>"010010100",
  46539=>"010011010",
  46540=>"111111001",
  46541=>"010010100",
  46542=>"110011001",
  46543=>"111110111",
  46544=>"000110110",
  46545=>"110001011",
  46546=>"000011110",
  46547=>"000001000",
  46548=>"110111110",
  46549=>"111110101",
  46550=>"000100111",
  46551=>"110110100",
  46552=>"100110000",
  46553=>"111011000",
  46554=>"101100000",
  46555=>"000000100",
  46556=>"110000101",
  46557=>"101101010",
  46558=>"110101111",
  46559=>"011010101",
  46560=>"101110010",
  46561=>"010000000",
  46562=>"111001001",
  46563=>"001101010",
  46564=>"101000011",
  46565=>"001101100",
  46566=>"110001101",
  46567=>"100001000",
  46568=>"011000010",
  46569=>"111110110",
  46570=>"000100100",
  46571=>"000000000",
  46572=>"001000110",
  46573=>"000000001",
  46574=>"100101011",
  46575=>"000010001",
  46576=>"101000001",
  46577=>"100100101",
  46578=>"100110100",
  46579=>"010001111",
  46580=>"111000010",
  46581=>"111010001",
  46582=>"101011110",
  46583=>"100010011",
  46584=>"000000100",
  46585=>"111000011",
  46586=>"101110000",
  46587=>"011000000",
  46588=>"100010101",
  46589=>"010110010",
  46590=>"101010011",
  46591=>"001100101",
  46592=>"100100101",
  46593=>"011011100",
  46594=>"000110111",
  46595=>"001000101",
  46596=>"011101100",
  46597=>"000100111",
  46598=>"001110001",
  46599=>"101011011",
  46600=>"111000011",
  46601=>"111111001",
  46602=>"000011101",
  46603=>"101111111",
  46604=>"001100010",
  46605=>"001111110",
  46606=>"010100100",
  46607=>"000101001",
  46608=>"001000101",
  46609=>"101111001",
  46610=>"110000001",
  46611=>"101111000",
  46612=>"000010011",
  46613=>"111111110",
  46614=>"100010110",
  46615=>"100010011",
  46616=>"000010001",
  46617=>"001011101",
  46618=>"100101000",
  46619=>"100010100",
  46620=>"000010110",
  46621=>"000001000",
  46622=>"000000000",
  46623=>"000111001",
  46624=>"101011110",
  46625=>"100101111",
  46626=>"000111001",
  46627=>"011101010",
  46628=>"100011010",
  46629=>"010111110",
  46630=>"011111000",
  46631=>"011101011",
  46632=>"010001101",
  46633=>"000110101",
  46634=>"110101010",
  46635=>"101001110",
  46636=>"110001110",
  46637=>"110100001",
  46638=>"111011000",
  46639=>"111001011",
  46640=>"101000101",
  46641=>"000000111",
  46642=>"111111110",
  46643=>"010011100",
  46644=>"000001010",
  46645=>"001010000",
  46646=>"111001001",
  46647=>"101100011",
  46648=>"010001000",
  46649=>"101100000",
  46650=>"001011110",
  46651=>"011110101",
  46652=>"001110000",
  46653=>"110001000",
  46654=>"101001111",
  46655=>"111100000",
  46656=>"110101011",
  46657=>"111111111",
  46658=>"001011011",
  46659=>"001110101",
  46660=>"101010010",
  46661=>"000101100",
  46662=>"010111100",
  46663=>"000101000",
  46664=>"110011111",
  46665=>"110011011",
  46666=>"100101001",
  46667=>"100001101",
  46668=>"101111011",
  46669=>"000110111",
  46670=>"111010110",
  46671=>"101110110",
  46672=>"111010001",
  46673=>"111101110",
  46674=>"100110010",
  46675=>"101001010",
  46676=>"000100111",
  46677=>"000100010",
  46678=>"001000000",
  46679=>"100000000",
  46680=>"110111111",
  46681=>"000101111",
  46682=>"111010000",
  46683=>"010110011",
  46684=>"110010110",
  46685=>"000000101",
  46686=>"010100001",
  46687=>"100111111",
  46688=>"111010011",
  46689=>"110110010",
  46690=>"010111010",
  46691=>"000101100",
  46692=>"000110000",
  46693=>"001111111",
  46694=>"011110111",
  46695=>"000000101",
  46696=>"100010110",
  46697=>"011011100",
  46698=>"100111010",
  46699=>"010001000",
  46700=>"100111111",
  46701=>"010110110",
  46702=>"000001110",
  46703=>"110101000",
  46704=>"111001111",
  46705=>"101111000",
  46706=>"111101010",
  46707=>"110000011",
  46708=>"101000000",
  46709=>"100111100",
  46710=>"111110111",
  46711=>"110011101",
  46712=>"001000000",
  46713=>"111000111",
  46714=>"000100000",
  46715=>"100100100",
  46716=>"101100000",
  46717=>"110011101",
  46718=>"010000100",
  46719=>"111010110",
  46720=>"111000010",
  46721=>"011010011",
  46722=>"001010100",
  46723=>"111011010",
  46724=>"011010011",
  46725=>"001111111",
  46726=>"111100000",
  46727=>"110101011",
  46728=>"110101011",
  46729=>"100010110",
  46730=>"001010010",
  46731=>"111011101",
  46732=>"111011111",
  46733=>"110110100",
  46734=>"100001000",
  46735=>"111100011",
  46736=>"001111011",
  46737=>"111111011",
  46738=>"011001000",
  46739=>"111001001",
  46740=>"011101100",
  46741=>"001100111",
  46742=>"111100111",
  46743=>"000101011",
  46744=>"011010011",
  46745=>"111111001",
  46746=>"110011101",
  46747=>"011110100",
  46748=>"011101011",
  46749=>"100011100",
  46750=>"010100001",
  46751=>"001100101",
  46752=>"001000010",
  46753=>"000011111",
  46754=>"101111001",
  46755=>"101010010",
  46756=>"001001111",
  46757=>"000100010",
  46758=>"101111100",
  46759=>"100010011",
  46760=>"111111001",
  46761=>"000101000",
  46762=>"011110001",
  46763=>"101100011",
  46764=>"101100001",
  46765=>"011101000",
  46766=>"010000100",
  46767=>"000100101",
  46768=>"011010101",
  46769=>"100011100",
  46770=>"101001110",
  46771=>"010001000",
  46772=>"001010110",
  46773=>"000100001",
  46774=>"100100010",
  46775=>"111101111",
  46776=>"110100000",
  46777=>"101000100",
  46778=>"101011111",
  46779=>"000110110",
  46780=>"011101001",
  46781=>"010110011",
  46782=>"001101111",
  46783=>"000110010",
  46784=>"011000001",
  46785=>"011010000",
  46786=>"100101010",
  46787=>"000100101",
  46788=>"111110001",
  46789=>"101100111",
  46790=>"101011001",
  46791=>"010111101",
  46792=>"011001001",
  46793=>"101010111",
  46794=>"000011111",
  46795=>"001110011",
  46796=>"001011010",
  46797=>"000010011",
  46798=>"100010011",
  46799=>"011001011",
  46800=>"110000001",
  46801=>"101100111",
  46802=>"010010111",
  46803=>"100011000",
  46804=>"010000011",
  46805=>"010110000",
  46806=>"010010001",
  46807=>"000011100",
  46808=>"000111001",
  46809=>"111101101",
  46810=>"101101111",
  46811=>"100001000",
  46812=>"111011011",
  46813=>"111010111",
  46814=>"110101011",
  46815=>"111001001",
  46816=>"000000111",
  46817=>"100001101",
  46818=>"101000000",
  46819=>"011111001",
  46820=>"110010111",
  46821=>"001000000",
  46822=>"010001001",
  46823=>"101111000",
  46824=>"111100101",
  46825=>"110110010",
  46826=>"110101000",
  46827=>"110100000",
  46828=>"111000100",
  46829=>"100100011",
  46830=>"001100011",
  46831=>"000101010",
  46832=>"011000100",
  46833=>"110011011",
  46834=>"110101110",
  46835=>"110101110",
  46836=>"101100010",
  46837=>"101111001",
  46838=>"001111101",
  46839=>"110111110",
  46840=>"110010110",
  46841=>"011101010",
  46842=>"111001100",
  46843=>"111010010",
  46844=>"010100011",
  46845=>"010111100",
  46846=>"000000001",
  46847=>"101100011",
  46848=>"000111001",
  46849=>"011001011",
  46850=>"111110001",
  46851=>"000111010",
  46852=>"111010001",
  46853=>"000110101",
  46854=>"100010110",
  46855=>"011111011",
  46856=>"001100010",
  46857=>"001000011",
  46858=>"111111111",
  46859=>"100011010",
  46860=>"111100001",
  46861=>"010001011",
  46862=>"000111101",
  46863=>"111110010",
  46864=>"111101011",
  46865=>"010110000",
  46866=>"000111001",
  46867=>"110000001",
  46868=>"100001000",
  46869=>"101100001",
  46870=>"010011111",
  46871=>"101110101",
  46872=>"000100000",
  46873=>"000000110",
  46874=>"100101111",
  46875=>"101000111",
  46876=>"001010101",
  46877=>"011001000",
  46878=>"001000001",
  46879=>"110000001",
  46880=>"001001110",
  46881=>"101110101",
  46882=>"100001110",
  46883=>"110101010",
  46884=>"010100100",
  46885=>"000100010",
  46886=>"001001111",
  46887=>"101100110",
  46888=>"011010011",
  46889=>"111100100",
  46890=>"010000100",
  46891=>"110000110",
  46892=>"110101000",
  46893=>"000010111",
  46894=>"100000100",
  46895=>"110110101",
  46896=>"110000011",
  46897=>"001110001",
  46898=>"011111011",
  46899=>"010111111",
  46900=>"110100110",
  46901=>"110000100",
  46902=>"001100110",
  46903=>"101001100",
  46904=>"011001111",
  46905=>"000010000",
  46906=>"111101110",
  46907=>"100111100",
  46908=>"010101110",
  46909=>"101100101",
  46910=>"100111110",
  46911=>"101111001",
  46912=>"110010001",
  46913=>"111011100",
  46914=>"010100000",
  46915=>"000100110",
  46916=>"010100111",
  46917=>"001111000",
  46918=>"000101011",
  46919=>"110110011",
  46920=>"001011111",
  46921=>"110001111",
  46922=>"100111110",
  46923=>"001111000",
  46924=>"000111011",
  46925=>"100100010",
  46926=>"111110110",
  46927=>"100000000",
  46928=>"110000111",
  46929=>"001111111",
  46930=>"000010101",
  46931=>"101000000",
  46932=>"100010110",
  46933=>"011111001",
  46934=>"010110110",
  46935=>"011101100",
  46936=>"000000100",
  46937=>"101110100",
  46938=>"001001010",
  46939=>"010111111",
  46940=>"000000111",
  46941=>"010110100",
  46942=>"001000111",
  46943=>"000000101",
  46944=>"111111110",
  46945=>"110100101",
  46946=>"001101111",
  46947=>"000011110",
  46948=>"011000001",
  46949=>"100000001",
  46950=>"000010010",
  46951=>"111110101",
  46952=>"011101101",
  46953=>"000111010",
  46954=>"011000100",
  46955=>"100000000",
  46956=>"111101100",
  46957=>"011111011",
  46958=>"000100010",
  46959=>"011100001",
  46960=>"100100110",
  46961=>"001010111",
  46962=>"100110001",
  46963=>"101100101",
  46964=>"000101111",
  46965=>"101000110",
  46966=>"100011001",
  46967=>"000100010",
  46968=>"100011001",
  46969=>"101101011",
  46970=>"101100100",
  46971=>"010000110",
  46972=>"000011100",
  46973=>"111000011",
  46974=>"011110101",
  46975=>"011001100",
  46976=>"101111110",
  46977=>"111000011",
  46978=>"011011101",
  46979=>"110000000",
  46980=>"111011111",
  46981=>"110000110",
  46982=>"110001100",
  46983=>"011001010",
  46984=>"000100001",
  46985=>"100111111",
  46986=>"100001110",
  46987=>"001100100",
  46988=>"011100100",
  46989=>"011111010",
  46990=>"010111101",
  46991=>"100000111",
  46992=>"100100001",
  46993=>"111111001",
  46994=>"000110111",
  46995=>"010111110",
  46996=>"110000100",
  46997=>"101111110",
  46998=>"011100001",
  46999=>"100110010",
  47000=>"001000101",
  47001=>"010001111",
  47002=>"111111001",
  47003=>"000110000",
  47004=>"000010110",
  47005=>"001001100",
  47006=>"100001000",
  47007=>"010010010",
  47008=>"001111010",
  47009=>"111001000",
  47010=>"010011100",
  47011=>"000011010",
  47012=>"101101000",
  47013=>"111111011",
  47014=>"111010011",
  47015=>"111000000",
  47016=>"100011010",
  47017=>"101111101",
  47018=>"110111110",
  47019=>"110100100",
  47020=>"100010110",
  47021=>"000111001",
  47022=>"111000011",
  47023=>"111111011",
  47024=>"000110110",
  47025=>"110110111",
  47026=>"011110000",
  47027=>"001000100",
  47028=>"111101101",
  47029=>"110000111",
  47030=>"000001011",
  47031=>"010111111",
  47032=>"011111001",
  47033=>"110001011",
  47034=>"111101111",
  47035=>"001011010",
  47036=>"111000100",
  47037=>"100001101",
  47038=>"110001010",
  47039=>"111011101",
  47040=>"100000011",
  47041=>"010101000",
  47042=>"100001010",
  47043=>"101101110",
  47044=>"101111101",
  47045=>"000101100",
  47046=>"101000111",
  47047=>"010001001",
  47048=>"100100001",
  47049=>"001001000",
  47050=>"000111000",
  47051=>"111000101",
  47052=>"111011001",
  47053=>"110001000",
  47054=>"000111011",
  47055=>"000101001",
  47056=>"100001100",
  47057=>"001010101",
  47058=>"001010010",
  47059=>"011100011",
  47060=>"001100011",
  47061=>"000000100",
  47062=>"000011011",
  47063=>"010110001",
  47064=>"101111110",
  47065=>"010011000",
  47066=>"000111101",
  47067=>"001100010",
  47068=>"001000110",
  47069=>"000000010",
  47070=>"010110111",
  47071=>"100001110",
  47072=>"001010111",
  47073=>"011000111",
  47074=>"001101001",
  47075=>"100111100",
  47076=>"011101011",
  47077=>"001000000",
  47078=>"101110111",
  47079=>"001111100",
  47080=>"100000001",
  47081=>"011001011",
  47082=>"000011010",
  47083=>"000111101",
  47084=>"000001010",
  47085=>"101110100",
  47086=>"001111111",
  47087=>"101110111",
  47088=>"110010100",
  47089=>"100111000",
  47090=>"001010101",
  47091=>"001001100",
  47092=>"001110111",
  47093=>"000111111",
  47094=>"110010001",
  47095=>"100000010",
  47096=>"110111100",
  47097=>"010111111",
  47098=>"001001100",
  47099=>"100010001",
  47100=>"110011010",
  47101=>"110011000",
  47102=>"001100101",
  47103=>"111110110",
  47104=>"010111000",
  47105=>"111000110",
  47106=>"100101011",
  47107=>"110000000",
  47108=>"100010110",
  47109=>"111000010",
  47110=>"100011010",
  47111=>"000111011",
  47112=>"101100111",
  47113=>"101111011",
  47114=>"101110001",
  47115=>"110100010",
  47116=>"111110000",
  47117=>"011001100",
  47118=>"001100010",
  47119=>"100111100",
  47120=>"101010110",
  47121=>"010111011",
  47122=>"011111100",
  47123=>"110001111",
  47124=>"110001100",
  47125=>"000010100",
  47126=>"000100001",
  47127=>"000110000",
  47128=>"010101010",
  47129=>"011110011",
  47130=>"011011011",
  47131=>"111001100",
  47132=>"000100100",
  47133=>"010101101",
  47134=>"010001010",
  47135=>"000010011",
  47136=>"110001011",
  47137=>"110001000",
  47138=>"000000111",
  47139=>"000010000",
  47140=>"010101101",
  47141=>"111110100",
  47142=>"010110110",
  47143=>"101000001",
  47144=>"001110100",
  47145=>"010101011",
  47146=>"001100010",
  47147=>"000100101",
  47148=>"101001001",
  47149=>"010000010",
  47150=>"010100000",
  47151=>"111010010",
  47152=>"000011110",
  47153=>"110000010",
  47154=>"000110001",
  47155=>"110101000",
  47156=>"110000010",
  47157=>"010100001",
  47158=>"000000000",
  47159=>"110011010",
  47160=>"011000001",
  47161=>"110101110",
  47162=>"011010011",
  47163=>"001100011",
  47164=>"110101110",
  47165=>"111111000",
  47166=>"111111100",
  47167=>"100001100",
  47168=>"000011011",
  47169=>"000100111",
  47170=>"011100000",
  47171=>"111000000",
  47172=>"011100101",
  47173=>"111101001",
  47174=>"100000000",
  47175=>"010001100",
  47176=>"000011010",
  47177=>"100011101",
  47178=>"110111010",
  47179=>"010000010",
  47180=>"010000110",
  47181=>"010001001",
  47182=>"001001101",
  47183=>"001100110",
  47184=>"101011010",
  47185=>"000000100",
  47186=>"011010111",
  47187=>"000001000",
  47188=>"110110000",
  47189=>"011100000",
  47190=>"010110000",
  47191=>"000000000",
  47192=>"100110101",
  47193=>"100110010",
  47194=>"110110101",
  47195=>"101100011",
  47196=>"001100110",
  47197=>"001011111",
  47198=>"001111110",
  47199=>"100001010",
  47200=>"111011001",
  47201=>"111111111",
  47202=>"001101010",
  47203=>"100101000",
  47204=>"000000100",
  47205=>"111100010",
  47206=>"110010001",
  47207=>"110100110",
  47208=>"110100110",
  47209=>"101001000",
  47210=>"001101110",
  47211=>"100001100",
  47212=>"010011011",
  47213=>"001110010",
  47214=>"100000001",
  47215=>"101011011",
  47216=>"101101010",
  47217=>"111110110",
  47218=>"111010011",
  47219=>"000110001",
  47220=>"010111100",
  47221=>"000010011",
  47222=>"011111110",
  47223=>"000011100",
  47224=>"001000111",
  47225=>"111011011",
  47226=>"100011010",
  47227=>"111110101",
  47228=>"110011001",
  47229=>"101111111",
  47230=>"001100000",
  47231=>"100010001",
  47232=>"100010100",
  47233=>"111101100",
  47234=>"111101011",
  47235=>"101111101",
  47236=>"101011110",
  47237=>"100110111",
  47238=>"000001010",
  47239=>"111000010",
  47240=>"011000111",
  47241=>"101000010",
  47242=>"010011100",
  47243=>"011111001",
  47244=>"000100111",
  47245=>"110111000",
  47246=>"000100111",
  47247=>"000001111",
  47248=>"101011011",
  47249=>"110000100",
  47250=>"101111111",
  47251=>"000010010",
  47252=>"101010011",
  47253=>"001110111",
  47254=>"100011001",
  47255=>"101011110",
  47256=>"000111101",
  47257=>"100111011",
  47258=>"101111011",
  47259=>"010010110",
  47260=>"111111100",
  47261=>"100000010",
  47262=>"100101011",
  47263=>"001110001",
  47264=>"001101100",
  47265=>"001100011",
  47266=>"010010101",
  47267=>"110100111",
  47268=>"011000100",
  47269=>"010100101",
  47270=>"111111101",
  47271=>"001110000",
  47272=>"111010010",
  47273=>"001100001",
  47274=>"001000011",
  47275=>"111010010",
  47276=>"111011100",
  47277=>"001111100",
  47278=>"000100001",
  47279=>"100101101",
  47280=>"111110010",
  47281=>"011111011",
  47282=>"000101011",
  47283=>"000110110",
  47284=>"111001101",
  47285=>"111111111",
  47286=>"100101111",
  47287=>"001000001",
  47288=>"110000100",
  47289=>"000110010",
  47290=>"001010010",
  47291=>"101110100",
  47292=>"011001001",
  47293=>"000111010",
  47294=>"110010100",
  47295=>"111111101",
  47296=>"111010011",
  47297=>"101001010",
  47298=>"100111001",
  47299=>"101110010",
  47300=>"001111001",
  47301=>"010001010",
  47302=>"011010100",
  47303=>"100000101",
  47304=>"110110101",
  47305=>"110000001",
  47306=>"110111111",
  47307=>"101110110",
  47308=>"010100011",
  47309=>"010000011",
  47310=>"000000010",
  47311=>"111110011",
  47312=>"010000000",
  47313=>"110001111",
  47314=>"011100100",
  47315=>"001111011",
  47316=>"100111000",
  47317=>"111011101",
  47318=>"011010011",
  47319=>"101011011",
  47320=>"011000010",
  47321=>"111110110",
  47322=>"111100011",
  47323=>"000100111",
  47324=>"000011111",
  47325=>"001110000",
  47326=>"110000011",
  47327=>"000000010",
  47328=>"110110011",
  47329=>"110001011",
  47330=>"111000001",
  47331=>"110010011",
  47332=>"000010010",
  47333=>"001001111",
  47334=>"001110010",
  47335=>"100010111",
  47336=>"111101100",
  47337=>"001000101",
  47338=>"011010000",
  47339=>"100101011",
  47340=>"010000000",
  47341=>"011000001",
  47342=>"010111101",
  47343=>"011110111",
  47344=>"111101001",
  47345=>"110110101",
  47346=>"110101001",
  47347=>"000101111",
  47348=>"010100110",
  47349=>"110110101",
  47350=>"111100111",
  47351=>"000010000",
  47352=>"111111000",
  47353=>"000001001",
  47354=>"111000111",
  47355=>"111011010",
  47356=>"110101010",
  47357=>"000110111",
  47358=>"110111110",
  47359=>"101011000",
  47360=>"000010111",
  47361=>"001100110",
  47362=>"000110000",
  47363=>"001110111",
  47364=>"011011001",
  47365=>"101110101",
  47366=>"001010001",
  47367=>"001110010",
  47368=>"010001100",
  47369=>"001000011",
  47370=>"010000010",
  47371=>"001101010",
  47372=>"010111000",
  47373=>"000000010",
  47374=>"010001000",
  47375=>"110000111",
  47376=>"001110000",
  47377=>"010110011",
  47378=>"110110010",
  47379=>"011011010",
  47380=>"011100110",
  47381=>"010110011",
  47382=>"000101011",
  47383=>"111000111",
  47384=>"010110111",
  47385=>"010000111",
  47386=>"111000010",
  47387=>"110010111",
  47388=>"000111100",
  47389=>"111111000",
  47390=>"110101111",
  47391=>"110110111",
  47392=>"111101101",
  47393=>"000101011",
  47394=>"110111111",
  47395=>"011000011",
  47396=>"111100100",
  47397=>"100000111",
  47398=>"110101001",
  47399=>"001100011",
  47400=>"011101100",
  47401=>"111101111",
  47402=>"111000010",
  47403=>"101000000",
  47404=>"110111100",
  47405=>"101011000",
  47406=>"011001010",
  47407=>"110110011",
  47408=>"110100100",
  47409=>"001011000",
  47410=>"110110010",
  47411=>"111111111",
  47412=>"000111101",
  47413=>"001110110",
  47414=>"011001000",
  47415=>"001111001",
  47416=>"000110001",
  47417=>"110000010",
  47418=>"101011110",
  47419=>"110011111",
  47420=>"111111111",
  47421=>"011000001",
  47422=>"001110100",
  47423=>"000011010",
  47424=>"111010001",
  47425=>"010011000",
  47426=>"111101101",
  47427=>"000010001",
  47428=>"100011111",
  47429=>"001111101",
  47430=>"000000110",
  47431=>"111110011",
  47432=>"011101101",
  47433=>"010000011",
  47434=>"101001111",
  47435=>"001001110",
  47436=>"110110100",
  47437=>"100100000",
  47438=>"101101101",
  47439=>"011000100",
  47440=>"010111101",
  47441=>"101000101",
  47442=>"010001111",
  47443=>"110110111",
  47444=>"000111100",
  47445=>"111110110",
  47446=>"110110010",
  47447=>"000010000",
  47448=>"011010100",
  47449=>"101010110",
  47450=>"011001110",
  47451=>"000010000",
  47452=>"111110001",
  47453=>"101101111",
  47454=>"100101000",
  47455=>"010100010",
  47456=>"000010111",
  47457=>"000010000",
  47458=>"101011101",
  47459=>"101010001",
  47460=>"101111110",
  47461=>"111101111",
  47462=>"101100000",
  47463=>"011011100",
  47464=>"110001100",
  47465=>"000000111",
  47466=>"101111111",
  47467=>"010001010",
  47468=>"101101010",
  47469=>"100010001",
  47470=>"111110000",
  47471=>"001100000",
  47472=>"010100100",
  47473=>"101111011",
  47474=>"011101110",
  47475=>"111011101",
  47476=>"111011001",
  47477=>"101010000",
  47478=>"110111000",
  47479=>"111101010",
  47480=>"001100011",
  47481=>"111010000",
  47482=>"000100101",
  47483=>"000110111",
  47484=>"010111110",
  47485=>"011111111",
  47486=>"001110011",
  47487=>"010100000",
  47488=>"110010110",
  47489=>"101000101",
  47490=>"100111111",
  47491=>"010101011",
  47492=>"100111110",
  47493=>"010011101",
  47494=>"000001011",
  47495=>"001111010",
  47496=>"111111010",
  47497=>"000110110",
  47498=>"011011111",
  47499=>"111011110",
  47500=>"100101110",
  47501=>"101001100",
  47502=>"100100000",
  47503=>"111000100",
  47504=>"000100011",
  47505=>"000100000",
  47506=>"001101100",
  47507=>"000101100",
  47508=>"000000000",
  47509=>"001110000",
  47510=>"010000100",
  47511=>"000111010",
  47512=>"101010001",
  47513=>"000000011",
  47514=>"100111000",
  47515=>"110000100",
  47516=>"110110101",
  47517=>"001111111",
  47518=>"011100110",
  47519=>"011000001",
  47520=>"100100000",
  47521=>"111100000",
  47522=>"100001110",
  47523=>"100101110",
  47524=>"100111110",
  47525=>"101011000",
  47526=>"111000100",
  47527=>"011110111",
  47528=>"101111110",
  47529=>"000100101",
  47530=>"100111101",
  47531=>"010011000",
  47532=>"100001101",
  47533=>"000110110",
  47534=>"100000111",
  47535=>"010110001",
  47536=>"000000100",
  47537=>"001000011",
  47538=>"110110111",
  47539=>"000000001",
  47540=>"000100010",
  47541=>"011100010",
  47542=>"011010111",
  47543=>"101110100",
  47544=>"101011010",
  47545=>"010111000",
  47546=>"101111111",
  47547=>"111111011",
  47548=>"111000110",
  47549=>"100111110",
  47550=>"101010111",
  47551=>"010010101",
  47552=>"000010000",
  47553=>"101000101",
  47554=>"001001000",
  47555=>"001111111",
  47556=>"100000000",
  47557=>"001010100",
  47558=>"100010100",
  47559=>"001000000",
  47560=>"110111010",
  47561=>"110110011",
  47562=>"000010011",
  47563=>"000011111",
  47564=>"000110111",
  47565=>"010110100",
  47566=>"000010001",
  47567=>"000100000",
  47568=>"111111010",
  47569=>"111101100",
  47570=>"000100101",
  47571=>"011101111",
  47572=>"011100000",
  47573=>"101011100",
  47574=>"000111100",
  47575=>"111111010",
  47576=>"111010001",
  47577=>"110111010",
  47578=>"110100110",
  47579=>"101010000",
  47580=>"011010010",
  47581=>"111111010",
  47582=>"000100000",
  47583=>"110010101",
  47584=>"001000000",
  47585=>"001000010",
  47586=>"001100100",
  47587=>"001000110",
  47588=>"000001101",
  47589=>"011110000",
  47590=>"101011110",
  47591=>"100000001",
  47592=>"001011001",
  47593=>"000001000",
  47594=>"000001010",
  47595=>"100011111",
  47596=>"011100010",
  47597=>"010001101",
  47598=>"010010000",
  47599=>"110010100",
  47600=>"100000000",
  47601=>"110000110",
  47602=>"111101011",
  47603=>"000101111",
  47604=>"111111000",
  47605=>"000111110",
  47606=>"100000011",
  47607=>"000010011",
  47608=>"011111100",
  47609=>"100011100",
  47610=>"110111100",
  47611=>"110110111",
  47612=>"001100001",
  47613=>"111111000",
  47614=>"101011101",
  47615=>"110001001",
  47616=>"000010010",
  47617=>"100010000",
  47618=>"111010011",
  47619=>"011001101",
  47620=>"101101001",
  47621=>"101011100",
  47622=>"011111011",
  47623=>"000100010",
  47624=>"000101001",
  47625=>"010001011",
  47626=>"110101101",
  47627=>"011000110",
  47628=>"100100110",
  47629=>"110010110",
  47630=>"000001100",
  47631=>"101000111",
  47632=>"011100100",
  47633=>"111111010",
  47634=>"011010011",
  47635=>"100000000",
  47636=>"111110001",
  47637=>"011011010",
  47638=>"111100001",
  47639=>"101110111",
  47640=>"110100100",
  47641=>"001001000",
  47642=>"000101011",
  47643=>"110010000",
  47644=>"101010101",
  47645=>"101010110",
  47646=>"101010100",
  47647=>"111011110",
  47648=>"111001111",
  47649=>"110000011",
  47650=>"000101000",
  47651=>"000111010",
  47652=>"000101000",
  47653=>"011000010",
  47654=>"000101100",
  47655=>"111110111",
  47656=>"100101110",
  47657=>"000100001",
  47658=>"110011001",
  47659=>"111001100",
  47660=>"011001110",
  47661=>"110011101",
  47662=>"001101111",
  47663=>"001001110",
  47664=>"110110100",
  47665=>"110101000",
  47666=>"011111100",
  47667=>"101110010",
  47668=>"110000000",
  47669=>"010110100",
  47670=>"000000010",
  47671=>"100101000",
  47672=>"111111000",
  47673=>"011000010",
  47674=>"000010110",
  47675=>"111000101",
  47676=>"101101110",
  47677=>"001000011",
  47678=>"010100000",
  47679=>"001011110",
  47680=>"000110111",
  47681=>"101010110",
  47682=>"011100000",
  47683=>"001010110",
  47684=>"000100010",
  47685=>"001100000",
  47686=>"001011001",
  47687=>"010110100",
  47688=>"011010100",
  47689=>"001111011",
  47690=>"101011010",
  47691=>"111111100",
  47692=>"010101010",
  47693=>"010110011",
  47694=>"101110101",
  47695=>"111111001",
  47696=>"111010011",
  47697=>"000011100",
  47698=>"010001010",
  47699=>"010011111",
  47700=>"010101000",
  47701=>"000000101",
  47702=>"110010101",
  47703=>"010010110",
  47704=>"001101010",
  47705=>"100000100",
  47706=>"110101001",
  47707=>"000000000",
  47708=>"110101111",
  47709=>"000100111",
  47710=>"101101010",
  47711=>"011010010",
  47712=>"100111111",
  47713=>"101001000",
  47714=>"000110110",
  47715=>"110011000",
  47716=>"110110100",
  47717=>"100110011",
  47718=>"001100111",
  47719=>"000000111",
  47720=>"111000001",
  47721=>"111111000",
  47722=>"011011011",
  47723=>"001000001",
  47724=>"010100010",
  47725=>"011001111",
  47726=>"110000010",
  47727=>"110010011",
  47728=>"101000011",
  47729=>"010100011",
  47730=>"110100101",
  47731=>"111001100",
  47732=>"110001010",
  47733=>"101001010",
  47734=>"001000011",
  47735=>"011011111",
  47736=>"000011011",
  47737=>"001110010",
  47738=>"001101110",
  47739=>"000010100",
  47740=>"010010101",
  47741=>"111010110",
  47742=>"001110001",
  47743=>"111100100",
  47744=>"001010000",
  47745=>"001000000",
  47746=>"000010100",
  47747=>"111111010",
  47748=>"011001000",
  47749=>"110100000",
  47750=>"000111001",
  47751=>"001111001",
  47752=>"001011111",
  47753=>"110101010",
  47754=>"110011001",
  47755=>"111110101",
  47756=>"011000000",
  47757=>"110001000",
  47758=>"011110000",
  47759=>"100010111",
  47760=>"000111010",
  47761=>"000011111",
  47762=>"010000111",
  47763=>"110011000",
  47764=>"010011111",
  47765=>"011101000",
  47766=>"011001110",
  47767=>"011101100",
  47768=>"111000100",
  47769=>"101111110",
  47770=>"001001111",
  47771=>"110000000",
  47772=>"000101000",
  47773=>"000011111",
  47774=>"111000101",
  47775=>"100000010",
  47776=>"000100000",
  47777=>"101111110",
  47778=>"100001001",
  47779=>"100011111",
  47780=>"001111111",
  47781=>"011011111",
  47782=>"010111010",
  47783=>"100110011",
  47784=>"011100001",
  47785=>"101100001",
  47786=>"000100100",
  47787=>"011111111",
  47788=>"100010011",
  47789=>"011100001",
  47790=>"100100000",
  47791=>"111111101",
  47792=>"101010010",
  47793=>"000011101",
  47794=>"110110100",
  47795=>"100101001",
  47796=>"000110001",
  47797=>"000110011",
  47798=>"010011111",
  47799=>"010001001",
  47800=>"101101101",
  47801=>"001011001",
  47802=>"010100110",
  47803=>"100011000",
  47804=>"000001001",
  47805=>"111110111",
  47806=>"011111010",
  47807=>"111001100",
  47808=>"110010101",
  47809=>"010011110",
  47810=>"111100000",
  47811=>"011000111",
  47812=>"101111101",
  47813=>"100111111",
  47814=>"001111000",
  47815=>"101010010",
  47816=>"111111111",
  47817=>"010101110",
  47818=>"001111000",
  47819=>"001101011",
  47820=>"010100000",
  47821=>"111110101",
  47822=>"001100100",
  47823=>"010010111",
  47824=>"111010110",
  47825=>"110111110",
  47826=>"110010011",
  47827=>"000100101",
  47828=>"001000110",
  47829=>"000101000",
  47830=>"010001000",
  47831=>"100000011",
  47832=>"101111100",
  47833=>"010100001",
  47834=>"010000010",
  47835=>"111000111",
  47836=>"111000100",
  47837=>"010011000",
  47838=>"101001111",
  47839=>"110110011",
  47840=>"110011111",
  47841=>"101110111",
  47842=>"010111000",
  47843=>"001010001",
  47844=>"010010010",
  47845=>"000101000",
  47846=>"101010010",
  47847=>"000000101",
  47848=>"001011010",
  47849=>"001001000",
  47850=>"001011111",
  47851=>"101100011",
  47852=>"001100010",
  47853=>"110101001",
  47854=>"110111100",
  47855=>"010010010",
  47856=>"011001001",
  47857=>"010110001",
  47858=>"011001111",
  47859=>"000010000",
  47860=>"001100001",
  47861=>"111010001",
  47862=>"110001110",
  47863=>"111111110",
  47864=>"100101100",
  47865=>"100000101",
  47866=>"110100001",
  47867=>"111111000",
  47868=>"101110010",
  47869=>"101010111",
  47870=>"011001000",
  47871=>"000001010",
  47872=>"000110000",
  47873=>"101001010",
  47874=>"101000110",
  47875=>"000001000",
  47876=>"100101101",
  47877=>"011111111",
  47878=>"111001110",
  47879=>"010001101",
  47880=>"100100000",
  47881=>"011010110",
  47882=>"101011000",
  47883=>"001011110",
  47884=>"101101000",
  47885=>"100111110",
  47886=>"100011101",
  47887=>"111011000",
  47888=>"100001101",
  47889=>"010001001",
  47890=>"110100011",
  47891=>"100010001",
  47892=>"111110100",
  47893=>"101100111",
  47894=>"110010010",
  47895=>"100001010",
  47896=>"010110001",
  47897=>"000000100",
  47898=>"110011011",
  47899=>"001110111",
  47900=>"001011000",
  47901=>"110011010",
  47902=>"100100110",
  47903=>"111100111",
  47904=>"000101100",
  47905=>"110000000",
  47906=>"110011110",
  47907=>"101110100",
  47908=>"101110111",
  47909=>"001100100",
  47910=>"000000111",
  47911=>"010010111",
  47912=>"011110100",
  47913=>"010010111",
  47914=>"100100011",
  47915=>"010001101",
  47916=>"011011100",
  47917=>"111010111",
  47918=>"010011001",
  47919=>"011101101",
  47920=>"010011001",
  47921=>"010000000",
  47922=>"110110110",
  47923=>"000110101",
  47924=>"111111101",
  47925=>"000001000",
  47926=>"010001101",
  47927=>"011010000",
  47928=>"001001001",
  47929=>"111000110",
  47930=>"001010100",
  47931=>"001111100",
  47932=>"100101000",
  47933=>"100000100",
  47934=>"000001010",
  47935=>"111111011",
  47936=>"010100111",
  47937=>"111111110",
  47938=>"000000010",
  47939=>"001111000",
  47940=>"111100001",
  47941=>"001111101",
  47942=>"000001000",
  47943=>"111011101",
  47944=>"001100011",
  47945=>"011110001",
  47946=>"100101000",
  47947=>"000001000",
  47948=>"101000000",
  47949=>"010010011",
  47950=>"011011110",
  47951=>"000011000",
  47952=>"000010110",
  47953=>"000101100",
  47954=>"100110010",
  47955=>"010111000",
  47956=>"100010011",
  47957=>"000100001",
  47958=>"000010000",
  47959=>"101000111",
  47960=>"100011001",
  47961=>"111000010",
  47962=>"001110110",
  47963=>"110110011",
  47964=>"101111111",
  47965=>"010000000",
  47966=>"001001000",
  47967=>"010100100",
  47968=>"010111011",
  47969=>"000110110",
  47970=>"010101000",
  47971=>"010101011",
  47972=>"110111000",
  47973=>"110110010",
  47974=>"110100010",
  47975=>"101100001",
  47976=>"101111110",
  47977=>"110111101",
  47978=>"001101010",
  47979=>"110011000",
  47980=>"110011001",
  47981=>"001101110",
  47982=>"111001110",
  47983=>"011011111",
  47984=>"001101001",
  47985=>"001111101",
  47986=>"000110000",
  47987=>"110100101",
  47988=>"001011011",
  47989=>"100001100",
  47990=>"010010000",
  47991=>"100001001",
  47992=>"111111110",
  47993=>"010001111",
  47994=>"000111101",
  47995=>"101000111",
  47996=>"000000100",
  47997=>"111101111",
  47998=>"111011110",
  47999=>"101010100",
  48000=>"001010001",
  48001=>"001110111",
  48002=>"100101101",
  48003=>"100100010",
  48004=>"100001000",
  48005=>"010101100",
  48006=>"111111111",
  48007=>"100111000",
  48008=>"010111000",
  48009=>"100011101",
  48010=>"110010100",
  48011=>"111100111",
  48012=>"111001011",
  48013=>"011000011",
  48014=>"111101101",
  48015=>"100000001",
  48016=>"010100111",
  48017=>"110001001",
  48018=>"011000010",
  48019=>"100010011",
  48020=>"100111010",
  48021=>"101111110",
  48022=>"110101010",
  48023=>"111001001",
  48024=>"001111000",
  48025=>"100011000",
  48026=>"110100100",
  48027=>"010001111",
  48028=>"000100101",
  48029=>"100001011",
  48030=>"000111011",
  48031=>"111111000",
  48032=>"000001011",
  48033=>"001111101",
  48034=>"111001111",
  48035=>"100110001",
  48036=>"100000001",
  48037=>"010100011",
  48038=>"011101001",
  48039=>"001100011",
  48040=>"011011000",
  48041=>"111111100",
  48042=>"000001101",
  48043=>"010100111",
  48044=>"000101101",
  48045=>"000110101",
  48046=>"010010110",
  48047=>"110000100",
  48048=>"011000010",
  48049=>"111100100",
  48050=>"110001011",
  48051=>"101001000",
  48052=>"000101111",
  48053=>"000001000",
  48054=>"010111111",
  48055=>"111100100",
  48056=>"011000010",
  48057=>"101000011",
  48058=>"010100111",
  48059=>"011001001",
  48060=>"000000100",
  48061=>"000110110",
  48062=>"100001011",
  48063=>"101110010",
  48064=>"111010111",
  48065=>"111111111",
  48066=>"100000010",
  48067=>"101110100",
  48068=>"111001100",
  48069=>"100110000",
  48070=>"010101111",
  48071=>"111010101",
  48072=>"001010111",
  48073=>"110001001",
  48074=>"011111010",
  48075=>"000010000",
  48076=>"011011011",
  48077=>"001100111",
  48078=>"101110010",
  48079=>"111010100",
  48080=>"101000101",
  48081=>"011001100",
  48082=>"010101001",
  48083=>"001010010",
  48084=>"000000001",
  48085=>"101010011",
  48086=>"000100100",
  48087=>"100001101",
  48088=>"000100101",
  48089=>"011101000",
  48090=>"010111101",
  48091=>"101000100",
  48092=>"000000000",
  48093=>"101010100",
  48094=>"010100001",
  48095=>"100000100",
  48096=>"001101010",
  48097=>"111001100",
  48098=>"000000011",
  48099=>"100010111",
  48100=>"111010010",
  48101=>"010101000",
  48102=>"101110111",
  48103=>"000001101",
  48104=>"100010111",
  48105=>"100110001",
  48106=>"001000010",
  48107=>"001100011",
  48108=>"101111111",
  48109=>"011000111",
  48110=>"100001000",
  48111=>"010010100",
  48112=>"010011010",
  48113=>"010110101",
  48114=>"100101001",
  48115=>"101011010",
  48116=>"011100111",
  48117=>"111010000",
  48118=>"011100101",
  48119=>"001111011",
  48120=>"111001010",
  48121=>"011100101",
  48122=>"111100110",
  48123=>"000111011",
  48124=>"110000100",
  48125=>"001110111",
  48126=>"101011000",
  48127=>"001101100",
  48128=>"000000100",
  48129=>"010011110",
  48130=>"001001001",
  48131=>"100100010",
  48132=>"101111110",
  48133=>"000110001",
  48134=>"101101011",
  48135=>"010101100",
  48136=>"010001010",
  48137=>"111011011",
  48138=>"011101010",
  48139=>"000101011",
  48140=>"001111010",
  48141=>"110011100",
  48142=>"000001000",
  48143=>"101001001",
  48144=>"100011011",
  48145=>"010010100",
  48146=>"111110100",
  48147=>"100111111",
  48148=>"101100100",
  48149=>"000100011",
  48150=>"011101011",
  48151=>"011111101",
  48152=>"000011001",
  48153=>"100010001",
  48154=>"011011111",
  48155=>"000011110",
  48156=>"010101111",
  48157=>"011101101",
  48158=>"011000011",
  48159=>"001010101",
  48160=>"010110110",
  48161=>"000110011",
  48162=>"100000101",
  48163=>"001001100",
  48164=>"100101000",
  48165=>"101010110",
  48166=>"001110111",
  48167=>"000100010",
  48168=>"101001011",
  48169=>"010011000",
  48170=>"001100100",
  48171=>"110011011",
  48172=>"010110101",
  48173=>"000010011",
  48174=>"000101011",
  48175=>"111010110",
  48176=>"101110101",
  48177=>"011001000",
  48178=>"001101001",
  48179=>"111111111",
  48180=>"111010011",
  48181=>"101010001",
  48182=>"111101000",
  48183=>"100111111",
  48184=>"010101110",
  48185=>"111111010",
  48186=>"000101101",
  48187=>"000101000",
  48188=>"000101111",
  48189=>"000100111",
  48190=>"101000000",
  48191=>"000101110",
  48192=>"111000100",
  48193=>"110001010",
  48194=>"001110100",
  48195=>"000110000",
  48196=>"000100011",
  48197=>"000001000",
  48198=>"110001010",
  48199=>"101111011",
  48200=>"010001011",
  48201=>"000001100",
  48202=>"010101000",
  48203=>"000100010",
  48204=>"001110000",
  48205=>"010000100",
  48206=>"010111011",
  48207=>"010101010",
  48208=>"011111101",
  48209=>"100000111",
  48210=>"000110100",
  48211=>"110010100",
  48212=>"100101101",
  48213=>"010010101",
  48214=>"101110000",
  48215=>"110000100",
  48216=>"011111110",
  48217=>"000000100",
  48218=>"000000111",
  48219=>"000101001",
  48220=>"001000010",
  48221=>"100001000",
  48222=>"111110100",
  48223=>"100000000",
  48224=>"000101001",
  48225=>"011010110",
  48226=>"101000100",
  48227=>"000010010",
  48228=>"100100001",
  48229=>"101100111",
  48230=>"100111010",
  48231=>"110011001",
  48232=>"010001111",
  48233=>"000001000",
  48234=>"101001001",
  48235=>"100111111",
  48236=>"011010110",
  48237=>"110101111",
  48238=>"011010001",
  48239=>"100101001",
  48240=>"100110010",
  48241=>"011101101",
  48242=>"100101000",
  48243=>"010111100",
  48244=>"110011011",
  48245=>"000001000",
  48246=>"000000110",
  48247=>"111111001",
  48248=>"110111011",
  48249=>"101111010",
  48250=>"000001011",
  48251=>"011111010",
  48252=>"110011010",
  48253=>"010011111",
  48254=>"001001000",
  48255=>"110000011",
  48256=>"010011101",
  48257=>"110100010",
  48258=>"011000101",
  48259=>"100101111",
  48260=>"000001010",
  48261=>"001101100",
  48262=>"011111101",
  48263=>"111101101",
  48264=>"011011010",
  48265=>"100100001",
  48266=>"011111000",
  48267=>"001000100",
  48268=>"110101001",
  48269=>"000110101",
  48270=>"000100001",
  48271=>"110011011",
  48272=>"011010011",
  48273=>"000010000",
  48274=>"111110000",
  48275=>"011111011",
  48276=>"001110000",
  48277=>"001101110",
  48278=>"001000000",
  48279=>"101111111",
  48280=>"011001010",
  48281=>"111110111",
  48282=>"111100001",
  48283=>"000110111",
  48284=>"010010011",
  48285=>"101011010",
  48286=>"000011000",
  48287=>"111011110",
  48288=>"101011001",
  48289=>"001100001",
  48290=>"010111100",
  48291=>"110000101",
  48292=>"110100111",
  48293=>"001001101",
  48294=>"001100111",
  48295=>"111110100",
  48296=>"110000000",
  48297=>"011100111",
  48298=>"010101000",
  48299=>"000100000",
  48300=>"111111110",
  48301=>"110011110",
  48302=>"101111011",
  48303=>"011111011",
  48304=>"001100110",
  48305=>"001010101",
  48306=>"000101110",
  48307=>"100011001",
  48308=>"010001010",
  48309=>"001000001",
  48310=>"001110101",
  48311=>"000001010",
  48312=>"000111110",
  48313=>"100100011",
  48314=>"001010000",
  48315=>"000001100",
  48316=>"010001110",
  48317=>"101101111",
  48318=>"111010101",
  48319=>"001010101",
  48320=>"111110111",
  48321=>"000101110",
  48322=>"100000000",
  48323=>"100111101",
  48324=>"110111110",
  48325=>"010011111",
  48326=>"110011000",
  48327=>"011001000",
  48328=>"001011111",
  48329=>"001011000",
  48330=>"011000001",
  48331=>"111011110",
  48332=>"111000000",
  48333=>"010010110",
  48334=>"110011101",
  48335=>"001010001",
  48336=>"101100010",
  48337=>"000100110",
  48338=>"000010100",
  48339=>"010110001",
  48340=>"110101110",
  48341=>"010101010",
  48342=>"111111100",
  48343=>"001111001",
  48344=>"001110001",
  48345=>"011000011",
  48346=>"100011111",
  48347=>"011100011",
  48348=>"100001011",
  48349=>"100001100",
  48350=>"001101101",
  48351=>"100000010",
  48352=>"001011101",
  48353=>"011101101",
  48354=>"010011001",
  48355=>"110000100",
  48356=>"110100100",
  48357=>"110101001",
  48358=>"001100010",
  48359=>"000110011",
  48360=>"010010110",
  48361=>"100001101",
  48362=>"111111011",
  48363=>"110010111",
  48364=>"000010101",
  48365=>"000001100",
  48366=>"001001001",
  48367=>"001000100",
  48368=>"100010011",
  48369=>"111001001",
  48370=>"110001001",
  48371=>"010001100",
  48372=>"110111100",
  48373=>"100100100",
  48374=>"010001011",
  48375=>"011111100",
  48376=>"111111000",
  48377=>"001010111",
  48378=>"000011100",
  48379=>"000111011",
  48380=>"011011100",
  48381=>"010111010",
  48382=>"111010000",
  48383=>"001110110",
  48384=>"111010011",
  48385=>"101011011",
  48386=>"011000000",
  48387=>"111001110",
  48388=>"111111000",
  48389=>"101011001",
  48390=>"101001100",
  48391=>"011111100",
  48392=>"011011100",
  48393=>"101111111",
  48394=>"001011100",
  48395=>"001101000",
  48396=>"011111000",
  48397=>"010111111",
  48398=>"010100100",
  48399=>"001010101",
  48400=>"011011010",
  48401=>"001111110",
  48402=>"001101000",
  48403=>"010001011",
  48404=>"010101001",
  48405=>"000100010",
  48406=>"100001110",
  48407=>"111001000",
  48408=>"010100010",
  48409=>"110110111",
  48410=>"101011011",
  48411=>"100001001",
  48412=>"011101101",
  48413=>"011001111",
  48414=>"010010011",
  48415=>"010101000",
  48416=>"100001010",
  48417=>"010111100",
  48418=>"010010010",
  48419=>"000000011",
  48420=>"011110101",
  48421=>"000110110",
  48422=>"111010000",
  48423=>"000100001",
  48424=>"010000111",
  48425=>"100100101",
  48426=>"001100011",
  48427=>"011011101",
  48428=>"111110011",
  48429=>"000010000",
  48430=>"100000010",
  48431=>"000000100",
  48432=>"001110000",
  48433=>"001100110",
  48434=>"001100010",
  48435=>"101101000",
  48436=>"001000000",
  48437=>"001011000",
  48438=>"011101111",
  48439=>"110000101",
  48440=>"100100001",
  48441=>"000001101",
  48442=>"001011010",
  48443=>"110000001",
  48444=>"110001110",
  48445=>"000010111",
  48446=>"001111101",
  48447=>"110110000",
  48448=>"111000000",
  48449=>"000000010",
  48450=>"100100111",
  48451=>"000001000",
  48452=>"001110100",
  48453=>"100000111",
  48454=>"111101101",
  48455=>"111011111",
  48456=>"011111110",
  48457=>"001101001",
  48458=>"100000100",
  48459=>"100001101",
  48460=>"110101110",
  48461=>"101111001",
  48462=>"001001110",
  48463=>"100001001",
  48464=>"001011101",
  48465=>"011110110",
  48466=>"000001001",
  48467=>"010010111",
  48468=>"000010010",
  48469=>"111111111",
  48470=>"110101100",
  48471=>"100111000",
  48472=>"011100000",
  48473=>"110010010",
  48474=>"100000010",
  48475=>"101010000",
  48476=>"111110101",
  48477=>"111001001",
  48478=>"111011100",
  48479=>"101010111",
  48480=>"101100001",
  48481=>"000111100",
  48482=>"011111010",
  48483=>"111000011",
  48484=>"100000000",
  48485=>"010101001",
  48486=>"100010000",
  48487=>"101011110",
  48488=>"100000010",
  48489=>"010011000",
  48490=>"011010001",
  48491=>"111101011",
  48492=>"011111000",
  48493=>"001111111",
  48494=>"100111011",
  48495=>"100100011",
  48496=>"110111010",
  48497=>"101101001",
  48498=>"011111111",
  48499=>"111110001",
  48500=>"100000110",
  48501=>"001001110",
  48502=>"011011111",
  48503=>"000101111",
  48504=>"001111011",
  48505=>"001010010",
  48506=>"011010010",
  48507=>"101001111",
  48508=>"100011000",
  48509=>"000110011",
  48510=>"000111000",
  48511=>"000011010",
  48512=>"010001001",
  48513=>"101111001",
  48514=>"101011011",
  48515=>"000000001",
  48516=>"001000111",
  48517=>"010010000",
  48518=>"010110010",
  48519=>"001010100",
  48520=>"111101000",
  48521=>"111110101",
  48522=>"011100010",
  48523=>"010001000",
  48524=>"100010010",
  48525=>"011000101",
  48526=>"110111100",
  48527=>"100100000",
  48528=>"100110100",
  48529=>"011110110",
  48530=>"110111110",
  48531=>"010110110",
  48532=>"001001110",
  48533=>"010001010",
  48534=>"010010001",
  48535=>"110011101",
  48536=>"001101111",
  48537=>"101001111",
  48538=>"010000110",
  48539=>"000000111",
  48540=>"010110010",
  48541=>"000110001",
  48542=>"011101100",
  48543=>"000001110",
  48544=>"101010101",
  48545=>"001000011",
  48546=>"001011001",
  48547=>"100001100",
  48548=>"001000100",
  48549=>"011000001",
  48550=>"000001101",
  48551=>"100011111",
  48552=>"011100101",
  48553=>"101010101",
  48554=>"110110110",
  48555=>"011010110",
  48556=>"101001001",
  48557=>"011011000",
  48558=>"110001101",
  48559=>"010111000",
  48560=>"010110100",
  48561=>"100010010",
  48562=>"001001001",
  48563=>"001100101",
  48564=>"111110010",
  48565=>"010110100",
  48566=>"000011100",
  48567=>"010100001",
  48568=>"001110110",
  48569=>"010001100",
  48570=>"000001000",
  48571=>"111000001",
  48572=>"100011000",
  48573=>"001110001",
  48574=>"000000010",
  48575=>"001101101",
  48576=>"111011111",
  48577=>"111110000",
  48578=>"000110110",
  48579=>"101000101",
  48580=>"000000010",
  48581=>"111100101",
  48582=>"000001111",
  48583=>"010110100",
  48584=>"111001010",
  48585=>"000010000",
  48586=>"001001011",
  48587=>"001100110",
  48588=>"011111100",
  48589=>"010100101",
  48590=>"001110000",
  48591=>"010011001",
  48592=>"101010101",
  48593=>"011110010",
  48594=>"100001011",
  48595=>"000101000",
  48596=>"001111110",
  48597=>"100110001",
  48598=>"011111001",
  48599=>"010010010",
  48600=>"001111101",
  48601=>"111010111",
  48602=>"000000010",
  48603=>"011001001",
  48604=>"010110101",
  48605=>"011001011",
  48606=>"111100001",
  48607=>"001011111",
  48608=>"111011010",
  48609=>"001011011",
  48610=>"010111110",
  48611=>"011000111",
  48612=>"111010100",
  48613=>"001011001",
  48614=>"010101000",
  48615=>"101001000",
  48616=>"110000110",
  48617=>"000000111",
  48618=>"101100110",
  48619=>"100100111",
  48620=>"000010001",
  48621=>"001010010",
  48622=>"000111011",
  48623=>"110010100",
  48624=>"111100100",
  48625=>"111010010",
  48626=>"011101000",
  48627=>"001100010",
  48628=>"101100100",
  48629=>"111010111",
  48630=>"110110100",
  48631=>"100001101",
  48632=>"110111111",
  48633=>"010100010",
  48634=>"000101100",
  48635=>"010110000",
  48636=>"101101001",
  48637=>"101100100",
  48638=>"111001000",
  48639=>"101100110",
  48640=>"111111000",
  48641=>"100000100",
  48642=>"011111001",
  48643=>"000100001",
  48644=>"001010100",
  48645=>"001110000",
  48646=>"100111111",
  48647=>"000100110",
  48648=>"000010111",
  48649=>"100001011",
  48650=>"110010011",
  48651=>"010011101",
  48652=>"010000011",
  48653=>"100011111",
  48654=>"010111100",
  48655=>"111110111",
  48656=>"000010000",
  48657=>"011101011",
  48658=>"110000100",
  48659=>"110110110",
  48660=>"000010110",
  48661=>"010001010",
  48662=>"111101101",
  48663=>"001010011",
  48664=>"100001000",
  48665=>"010101000",
  48666=>"001001000",
  48667=>"011011010",
  48668=>"010000110",
  48669=>"111001001",
  48670=>"010110001",
  48671=>"000100010",
  48672=>"011101000",
  48673=>"100100000",
  48674=>"000100111",
  48675=>"001011101",
  48676=>"110111000",
  48677=>"100101101",
  48678=>"000000001",
  48679=>"000100011",
  48680=>"100101010",
  48681=>"100110011",
  48682=>"110111101",
  48683=>"100111111",
  48684=>"011010011",
  48685=>"101111100",
  48686=>"000100110",
  48687=>"101000010",
  48688=>"001101010",
  48689=>"011010001",
  48690=>"100011011",
  48691=>"100110111",
  48692=>"100001000",
  48693=>"111011011",
  48694=>"010111011",
  48695=>"000001000",
  48696=>"011100001",
  48697=>"011101000",
  48698=>"000110011",
  48699=>"001010111",
  48700=>"110100100",
  48701=>"001101111",
  48702=>"010111011",
  48703=>"101101101",
  48704=>"100010101",
  48705=>"100101010",
  48706=>"000000011",
  48707=>"010011000",
  48708=>"101100100",
  48709=>"010111011",
  48710=>"000100110",
  48711=>"001111110",
  48712=>"001010110",
  48713=>"010010111",
  48714=>"111001101",
  48715=>"010111110",
  48716=>"000101101",
  48717=>"100111001",
  48718=>"011001101",
  48719=>"111010110",
  48720=>"011110011",
  48721=>"111001010",
  48722=>"101001111",
  48723=>"111101101",
  48724=>"100100000",
  48725=>"110110101",
  48726=>"011111101",
  48727=>"001010010",
  48728=>"001101101",
  48729=>"011011111",
  48730=>"111000101",
  48731=>"000010001",
  48732=>"100011010",
  48733=>"010110010",
  48734=>"101010100",
  48735=>"001101100",
  48736=>"101100100",
  48737=>"010001011",
  48738=>"111011111",
  48739=>"000101000",
  48740=>"100100101",
  48741=>"000000000",
  48742=>"101111010",
  48743=>"010000000",
  48744=>"001111100",
  48745=>"000100100",
  48746=>"001011110",
  48747=>"110001000",
  48748=>"011100101",
  48749=>"001000011",
  48750=>"100100011",
  48751=>"001101111",
  48752=>"100110101",
  48753=>"101000111",
  48754=>"100000011",
  48755=>"101100001",
  48756=>"000000010",
  48757=>"111101111",
  48758=>"011110100",
  48759=>"101110001",
  48760=>"100000010",
  48761=>"011101100",
  48762=>"110000000",
  48763=>"000100011",
  48764=>"011010010",
  48765=>"100100000",
  48766=>"001001101",
  48767=>"100111111",
  48768=>"010110010",
  48769=>"010011000",
  48770=>"010011001",
  48771=>"001001101",
  48772=>"100000111",
  48773=>"111101100",
  48774=>"001011010",
  48775=>"110010111",
  48776=>"101111001",
  48777=>"001000010",
  48778=>"010011110",
  48779=>"001101111",
  48780=>"001101110",
  48781=>"001001110",
  48782=>"001100000",
  48783=>"111011010",
  48784=>"110110101",
  48785=>"010100010",
  48786=>"010110110",
  48787=>"011110111",
  48788=>"010101111",
  48789=>"001010101",
  48790=>"111111101",
  48791=>"010101111",
  48792=>"100011000",
  48793=>"111011010",
  48794=>"010110100",
  48795=>"110001111",
  48796=>"111011010",
  48797=>"100001111",
  48798=>"110001001",
  48799=>"101111101",
  48800=>"001101000",
  48801=>"001110100",
  48802=>"011011111",
  48803=>"011011000",
  48804=>"101100000",
  48805=>"111000100",
  48806=>"110010100",
  48807=>"101000101",
  48808=>"011101011",
  48809=>"100111101",
  48810=>"001010110",
  48811=>"000110101",
  48812=>"110000000",
  48813=>"001001011",
  48814=>"011110110",
  48815=>"101001100",
  48816=>"010001000",
  48817=>"100101111",
  48818=>"011010001",
  48819=>"101111010",
  48820=>"010011001",
  48821=>"001001110",
  48822=>"011011011",
  48823=>"010011001",
  48824=>"100100001",
  48825=>"000100011",
  48826=>"010110100",
  48827=>"110111101",
  48828=>"010100011",
  48829=>"001010110",
  48830=>"100000011",
  48831=>"010110000",
  48832=>"001110011",
  48833=>"001101000",
  48834=>"101101000",
  48835=>"000001001",
  48836=>"001111100",
  48837=>"010110111",
  48838=>"011001100",
  48839=>"110111100",
  48840=>"101111000",
  48841=>"110011101",
  48842=>"110001111",
  48843=>"111001101",
  48844=>"001111100",
  48845=>"101100101",
  48846=>"110100100",
  48847=>"100010110",
  48848=>"010100010",
  48849=>"111000011",
  48850=>"110011010",
  48851=>"011001001",
  48852=>"111000000",
  48853=>"000110101",
  48854=>"001101100",
  48855=>"010011110",
  48856=>"000110010",
  48857=>"000011000",
  48858=>"001000111",
  48859=>"000111100",
  48860=>"110100111",
  48861=>"110110001",
  48862=>"111001111",
  48863=>"010110101",
  48864=>"100011101",
  48865=>"100111111",
  48866=>"111101001",
  48867=>"011101010",
  48868=>"001001011",
  48869=>"111100100",
  48870=>"000110111",
  48871=>"011111101",
  48872=>"101010011",
  48873=>"101000101",
  48874=>"011100000",
  48875=>"010001101",
  48876=>"101010001",
  48877=>"000000101",
  48878=>"111111100",
  48879=>"001111111",
  48880=>"111000100",
  48881=>"100010010",
  48882=>"000101011",
  48883=>"011110110",
  48884=>"111010011",
  48885=>"101110000",
  48886=>"110010101",
  48887=>"001010011",
  48888=>"011000111",
  48889=>"101011100",
  48890=>"101101001",
  48891=>"111110101",
  48892=>"100101111",
  48893=>"101011111",
  48894=>"100000010",
  48895=>"000000011",
  48896=>"110010110",
  48897=>"011101011",
  48898=>"001100111",
  48899=>"000100101",
  48900=>"011000110",
  48901=>"101100110",
  48902=>"111000111",
  48903=>"011001101",
  48904=>"001010010",
  48905=>"001100010",
  48906=>"100010000",
  48907=>"000001111",
  48908=>"110001101",
  48909=>"001110111",
  48910=>"000000001",
  48911=>"100001011",
  48912=>"000000100",
  48913=>"100100010",
  48914=>"111011011",
  48915=>"100100000",
  48916=>"100100101",
  48917=>"000010101",
  48918=>"100000000",
  48919=>"101010110",
  48920=>"111110100",
  48921=>"101011110",
  48922=>"100000000",
  48923=>"110001011",
  48924=>"011100111",
  48925=>"101111000",
  48926=>"010110111",
  48927=>"111000011",
  48928=>"010100000",
  48929=>"000010011",
  48930=>"000010000",
  48931=>"101010001",
  48932=>"110101110",
  48933=>"111100110",
  48934=>"010011010",
  48935=>"101101111",
  48936=>"011110001",
  48937=>"010100111",
  48938=>"000101101",
  48939=>"101100011",
  48940=>"001011001",
  48941=>"110111111",
  48942=>"000011100",
  48943=>"000100110",
  48944=>"010011101",
  48945=>"101100001",
  48946=>"000011101",
  48947=>"111111010",
  48948=>"011111010",
  48949=>"111010000",
  48950=>"110011010",
  48951=>"000101001",
  48952=>"001110001",
  48953=>"000101010",
  48954=>"000001011",
  48955=>"011101011",
  48956=>"101000010",
  48957=>"110110110",
  48958=>"111010010",
  48959=>"000011101",
  48960=>"110000010",
  48961=>"110000000",
  48962=>"100000001",
  48963=>"000101011",
  48964=>"101000000",
  48965=>"011111100",
  48966=>"110101110",
  48967=>"011101011",
  48968=>"110111111",
  48969=>"000010100",
  48970=>"110101011",
  48971=>"010100101",
  48972=>"110010110",
  48973=>"111100001",
  48974=>"110011000",
  48975=>"101100100",
  48976=>"110101110",
  48977=>"110001000",
  48978=>"010001010",
  48979=>"110110000",
  48980=>"000000001",
  48981=>"011001110",
  48982=>"100111011",
  48983=>"100100101",
  48984=>"010100010",
  48985=>"010101100",
  48986=>"000000000",
  48987=>"001111111",
  48988=>"001000010",
  48989=>"101000001",
  48990=>"101010110",
  48991=>"100110101",
  48992=>"111000011",
  48993=>"010101100",
  48994=>"000101011",
  48995=>"001010101",
  48996=>"001111000",
  48997=>"001101000",
  48998=>"001100100",
  48999=>"010001100",
  49000=>"100011110",
  49001=>"101101101",
  49002=>"101001010",
  49003=>"110001101",
  49004=>"011101000",
  49005=>"010010101",
  49006=>"100101000",
  49007=>"101110000",
  49008=>"010010100",
  49009=>"010001100",
  49010=>"001001000",
  49011=>"100110000",
  49012=>"010101000",
  49013=>"001010001",
  49014=>"101000101",
  49015=>"101100000",
  49016=>"010110011",
  49017=>"001110011",
  49018=>"111101001",
  49019=>"111011000",
  49020=>"000110111",
  49021=>"001110111",
  49022=>"100011010",
  49023=>"100111111",
  49024=>"101100001",
  49025=>"001111110",
  49026=>"110111100",
  49027=>"010011010",
  49028=>"001101000",
  49029=>"101011000",
  49030=>"110000101",
  49031=>"110111000",
  49032=>"011110110",
  49033=>"001000110",
  49034=>"001000010",
  49035=>"000110100",
  49036=>"110100111",
  49037=>"000000011",
  49038=>"010010010",
  49039=>"100110111",
  49040=>"100001111",
  49041=>"010000110",
  49042=>"111011010",
  49043=>"101000010",
  49044=>"000010101",
  49045=>"111101101",
  49046=>"000101101",
  49047=>"100100110",
  49048=>"010011111",
  49049=>"000011011",
  49050=>"110111001",
  49051=>"101110110",
  49052=>"111001111",
  49053=>"111111011",
  49054=>"011000011",
  49055=>"001111111",
  49056=>"001110100",
  49057=>"001000111",
  49058=>"011001101",
  49059=>"000010000",
  49060=>"100011111",
  49061=>"111011110",
  49062=>"110100010",
  49063=>"011010011",
  49064=>"111100010",
  49065=>"110010001",
  49066=>"100110110",
  49067=>"001001110",
  49068=>"011100101",
  49069=>"001101110",
  49070=>"010001001",
  49071=>"101100110",
  49072=>"111010000",
  49073=>"000000110",
  49074=>"010001101",
  49075=>"101001001",
  49076=>"111100001",
  49077=>"110101000",
  49078=>"111111101",
  49079=>"010101110",
  49080=>"101000111",
  49081=>"011111011",
  49082=>"110111001",
  49083=>"011111000",
  49084=>"100011001",
  49085=>"110011010",
  49086=>"001100011",
  49087=>"011000000",
  49088=>"011001010",
  49089=>"100010100",
  49090=>"010111110",
  49091=>"010101110",
  49092=>"010010100",
  49093=>"111010011",
  49094=>"011101111",
  49095=>"000110100",
  49096=>"000011101",
  49097=>"000000110",
  49098=>"111000110",
  49099=>"011001011",
  49100=>"111110111",
  49101=>"100001001",
  49102=>"101100000",
  49103=>"000101010",
  49104=>"100001001",
  49105=>"000000011",
  49106=>"001100010",
  49107=>"101000001",
  49108=>"000100110",
  49109=>"110000101",
  49110=>"000011000",
  49111=>"101111010",
  49112=>"111000011",
  49113=>"011110000",
  49114=>"000001111",
  49115=>"100110101",
  49116=>"010011000",
  49117=>"011010100",
  49118=>"010101000",
  49119=>"000000010",
  49120=>"001001111",
  49121=>"101011010",
  49122=>"110101001",
  49123=>"110110011",
  49124=>"010011111",
  49125=>"011010011",
  49126=>"001110001",
  49127=>"100110011",
  49128=>"110010000",
  49129=>"101010001",
  49130=>"111000111",
  49131=>"101010100",
  49132=>"011011000",
  49133=>"000101110",
  49134=>"100110101",
  49135=>"100010010",
  49136=>"010001000",
  49137=>"111111100",
  49138=>"010110011",
  49139=>"000011111",
  49140=>"001101000",
  49141=>"000100101",
  49142=>"001011000",
  49143=>"011101100",
  49144=>"111110011",
  49145=>"111111001",
  49146=>"001001110",
  49147=>"001110110",
  49148=>"100101011",
  49149=>"101110101",
  49150=>"010101111",
  49151=>"001001110",
  49152=>"001010111",
  49153=>"011111000",
  49154=>"001111101",
  49155=>"010000001",
  49156=>"000001101",
  49157=>"110111110",
  49158=>"010110000",
  49159=>"011000100",
  49160=>"100101111",
  49161=>"110011011",
  49162=>"100000010",
  49163=>"001010100",
  49164=>"110000101",
  49165=>"110111011",
  49166=>"001101111",
  49167=>"011100011",
  49168=>"010110000",
  49169=>"000000101",
  49170=>"000000000",
  49171=>"100101100",
  49172=>"111010111",
  49173=>"001001110",
  49174=>"111011001",
  49175=>"000110001",
  49176=>"001011111",
  49177=>"100010110",
  49178=>"000011001",
  49179=>"100110001",
  49180=>"000101010",
  49181=>"100111010",
  49182=>"001111100",
  49183=>"101000100",
  49184=>"110100111",
  49185=>"001001011",
  49186=>"011000010",
  49187=>"110010010",
  49188=>"101100010",
  49189=>"010111100",
  49190=>"010001101",
  49191=>"110100101",
  49192=>"100011010",
  49193=>"011010010",
  49194=>"101101110",
  49195=>"010111100",
  49196=>"111110101",
  49197=>"110111101",
  49198=>"011010000",
  49199=>"000111111",
  49200=>"101010011",
  49201=>"010111101",
  49202=>"100111000",
  49203=>"010101100",
  49204=>"010000001",
  49205=>"010000000",
  49206=>"000101100",
  49207=>"111001001",
  49208=>"101101100",
  49209=>"010011110",
  49210=>"100100100",
  49211=>"110001011",
  49212=>"100010101",
  49213=>"001011110",
  49214=>"100101001",
  49215=>"110111011",
  49216=>"001011111",
  49217=>"000000101",
  49218=>"010001000",
  49219=>"000101100",
  49220=>"111110110",
  49221=>"111101101",
  49222=>"101011110",
  49223=>"111110111",
  49224=>"111000000",
  49225=>"000000010",
  49226=>"001000101",
  49227=>"101110001",
  49228=>"100110101",
  49229=>"101100110",
  49230=>"001001011",
  49231=>"100010010",
  49232=>"100010011",
  49233=>"000111001",
  49234=>"001111110",
  49235=>"000010101",
  49236=>"010011010",
  49237=>"000101000",
  49238=>"010110100",
  49239=>"100101101",
  49240=>"101101011",
  49241=>"001110101",
  49242=>"011010111",
  49243=>"011001100",
  49244=>"011010111",
  49245=>"111111111",
  49246=>"101001010",
  49247=>"001010010",
  49248=>"010111101",
  49249=>"001010010",
  49250=>"110011111",
  49251=>"100000001",
  49252=>"000100111",
  49253=>"111111110",
  49254=>"000100001",
  49255=>"000011110",
  49256=>"101110010",
  49257=>"101000100",
  49258=>"101010100",
  49259=>"011110001",
  49260=>"100001110",
  49261=>"000001001",
  49262=>"110100111",
  49263=>"100101000",
  49264=>"110001111",
  49265=>"001010110",
  49266=>"110111101",
  49267=>"110101110",
  49268=>"000111110",
  49269=>"010111000",
  49270=>"111100011",
  49271=>"101111100",
  49272=>"000011010",
  49273=>"010010110",
  49274=>"010011010",
  49275=>"011110000",
  49276=>"001111011",
  49277=>"010110100",
  49278=>"011100110",
  49279=>"000000011",
  49280=>"011101011",
  49281=>"111001101",
  49282=>"111111101",
  49283=>"001010100",
  49284=>"110010011",
  49285=>"110100011",
  49286=>"101000011",
  49287=>"010100111",
  49288=>"011101101",
  49289=>"000011000",
  49290=>"001010010",
  49291=>"101110010",
  49292=>"100100010",
  49293=>"011110010",
  49294=>"101010001",
  49295=>"110011000",
  49296=>"111011100",
  49297=>"011010010",
  49298=>"011010111",
  49299=>"001111010",
  49300=>"011010001",
  49301=>"001111010",
  49302=>"000110100",
  49303=>"110010110",
  49304=>"000000000",
  49305=>"001110100",
  49306=>"011000111",
  49307=>"000000100",
  49308=>"001111010",
  49309=>"010111000",
  49310=>"011001110",
  49311=>"000111001",
  49312=>"001111100",
  49313=>"111110010",
  49314=>"010001110",
  49315=>"111011001",
  49316=>"000111010",
  49317=>"000101011",
  49318=>"111001110",
  49319=>"100101111",
  49320=>"000110111",
  49321=>"110101111",
  49322=>"001001111",
  49323=>"101011101",
  49324=>"001100000",
  49325=>"011010100",
  49326=>"000011111",
  49327=>"101100000",
  49328=>"100000010",
  49329=>"010001111",
  49330=>"001100100",
  49331=>"101000100",
  49332=>"010011111",
  49333=>"000110001",
  49334=>"101110101",
  49335=>"000011011",
  49336=>"111111000",
  49337=>"110110011",
  49338=>"100001100",
  49339=>"010101001",
  49340=>"000010001",
  49341=>"010000010",
  49342=>"001101100",
  49343=>"010100000",
  49344=>"001110111",
  49345=>"100000111",
  49346=>"101011101",
  49347=>"110111100",
  49348=>"000110010",
  49349=>"110100010",
  49350=>"111101000",
  49351=>"111111111",
  49352=>"110101111",
  49353=>"001000110",
  49354=>"010011101",
  49355=>"100110001",
  49356=>"000101001",
  49357=>"000110101",
  49358=>"100000000",
  49359=>"011010100",
  49360=>"011101011",
  49361=>"111111100",
  49362=>"010101101",
  49363=>"111001110",
  49364=>"100010001",
  49365=>"100001001",
  49366=>"010110110",
  49367=>"111101110",
  49368=>"111101011",
  49369=>"100111001",
  49370=>"010100010",
  49371=>"111011100",
  49372=>"000000000",
  49373=>"111110010",
  49374=>"011110110",
  49375=>"000010101",
  49376=>"000000110",
  49377=>"000010010",
  49378=>"111100010",
  49379=>"001000000",
  49380=>"110011101",
  49381=>"100000110",
  49382=>"001010011",
  49383=>"000111111",
  49384=>"010011111",
  49385=>"101111101",
  49386=>"000000000",
  49387=>"010101000",
  49388=>"111110111",
  49389=>"000110011",
  49390=>"101000001",
  49391=>"001001010",
  49392=>"001000011",
  49393=>"111010000",
  49394=>"101100110",
  49395=>"011100011",
  49396=>"000000011",
  49397=>"011110011",
  49398=>"000000001",
  49399=>"001111100",
  49400=>"101101110",
  49401=>"100110111",
  49402=>"101100000",
  49403=>"010010100",
  49404=>"001000001",
  49405=>"001101110",
  49406=>"000000111",
  49407=>"000111111",
  49408=>"110101001",
  49409=>"111011001",
  49410=>"100111100",
  49411=>"111001011",
  49412=>"111011011",
  49413=>"101111100",
  49414=>"001010111",
  49415=>"110100010",
  49416=>"001110101",
  49417=>"111001111",
  49418=>"111010100",
  49419=>"101100100",
  49420=>"000100101",
  49421=>"110011000",
  49422=>"011110010",
  49423=>"001000100",
  49424=>"000110100",
  49425=>"000101000",
  49426=>"101110000",
  49427=>"101101011",
  49428=>"111110000",
  49429=>"111001110",
  49430=>"101001011",
  49431=>"101000000",
  49432=>"000000101",
  49433=>"101110000",
  49434=>"100101011",
  49435=>"100110001",
  49436=>"111100001",
  49437=>"000111110",
  49438=>"010010000",
  49439=>"100000111",
  49440=>"000011011",
  49441=>"000100101",
  49442=>"010001010",
  49443=>"000000010",
  49444=>"001111101",
  49445=>"111010000",
  49446=>"001000001",
  49447=>"110001111",
  49448=>"011101110",
  49449=>"000011011",
  49450=>"010111011",
  49451=>"011100001",
  49452=>"010101001",
  49453=>"011110110",
  49454=>"101000001",
  49455=>"001100000",
  49456=>"110101001",
  49457=>"100011100",
  49458=>"110101110",
  49459=>"000000010",
  49460=>"001101000",
  49461=>"101111000",
  49462=>"110111001",
  49463=>"010100011",
  49464=>"110010111",
  49465=>"100000010",
  49466=>"010001001",
  49467=>"100101100",
  49468=>"011010000",
  49469=>"111111010",
  49470=>"010101101",
  49471=>"010111011",
  49472=>"011100000",
  49473=>"001100011",
  49474=>"101110100",
  49475=>"010001111",
  49476=>"011011001",
  49477=>"011111101",
  49478=>"110001010",
  49479=>"111110101",
  49480=>"100110000",
  49481=>"011111010",
  49482=>"001011011",
  49483=>"001000100",
  49484=>"101011010",
  49485=>"110010000",
  49486=>"101001010",
  49487=>"000101000",
  49488=>"010111111",
  49489=>"011011010",
  49490=>"011000000",
  49491=>"000111101",
  49492=>"101111010",
  49493=>"100100010",
  49494=>"010100111",
  49495=>"110111100",
  49496=>"000010101",
  49497=>"110000100",
  49498=>"100101100",
  49499=>"000000000",
  49500=>"111001000",
  49501=>"000111110",
  49502=>"010101000",
  49503=>"101100100",
  49504=>"111111001",
  49505=>"100111011",
  49506=>"111010001",
  49507=>"000111101",
  49508=>"000100101",
  49509=>"000000001",
  49510=>"000100110",
  49511=>"100001000",
  49512=>"100111101",
  49513=>"110111111",
  49514=>"011111101",
  49515=>"101100011",
  49516=>"110111001",
  49517=>"111111000",
  49518=>"100011010",
  49519=>"000111111",
  49520=>"111010101",
  49521=>"001001001",
  49522=>"011001001",
  49523=>"000100111",
  49524=>"011101111",
  49525=>"111110000",
  49526=>"111011110",
  49527=>"110110000",
  49528=>"000011100",
  49529=>"101010000",
  49530=>"101001010",
  49531=>"000101010",
  49532=>"101011111",
  49533=>"011010000",
  49534=>"111000101",
  49535=>"100111001",
  49536=>"101101110",
  49537=>"011110001",
  49538=>"011101101",
  49539=>"010110000",
  49540=>"111010100",
  49541=>"110000111",
  49542=>"110111100",
  49543=>"100101000",
  49544=>"010111101",
  49545=>"001101010",
  49546=>"110100000",
  49547=>"011111101",
  49548=>"101110010",
  49549=>"011000011",
  49550=>"111011101",
  49551=>"110111000",
  49552=>"001011010",
  49553=>"111100010",
  49554=>"101101100",
  49555=>"010101010",
  49556=>"011011100",
  49557=>"000001011",
  49558=>"111110000",
  49559=>"111011000",
  49560=>"110101001",
  49561=>"011100010",
  49562=>"010100000",
  49563=>"010000100",
  49564=>"000000100",
  49565=>"110011000",
  49566=>"111110000",
  49567=>"010101001",
  49568=>"011110110",
  49569=>"111110011",
  49570=>"010111101",
  49571=>"001001010",
  49572=>"111101011",
  49573=>"011000011",
  49574=>"110101101",
  49575=>"010001001",
  49576=>"001000100",
  49577=>"101101001",
  49578=>"110001100",
  49579=>"000010000",
  49580=>"011100011",
  49581=>"011111100",
  49582=>"001110001",
  49583=>"110011001",
  49584=>"101001010",
  49585=>"001101101",
  49586=>"100101110",
  49587=>"110010100",
  49588=>"001110110",
  49589=>"100001111",
  49590=>"011111100",
  49591=>"101011101",
  49592=>"010000011",
  49593=>"000111111",
  49594=>"010100011",
  49595=>"010110111",
  49596=>"110001111",
  49597=>"111100100",
  49598=>"101110001",
  49599=>"001110011",
  49600=>"111011001",
  49601=>"011010001",
  49602=>"010011110",
  49603=>"110010010",
  49604=>"111101111",
  49605=>"100101011",
  49606=>"111100000",
  49607=>"000101110",
  49608=>"000100111",
  49609=>"111110011",
  49610=>"111110010",
  49611=>"110110111",
  49612=>"000100011",
  49613=>"100011011",
  49614=>"101101011",
  49615=>"010001010",
  49616=>"100110101",
  49617=>"110001101",
  49618=>"101011011",
  49619=>"001011001",
  49620=>"001010101",
  49621=>"110010010",
  49622=>"000110010",
  49623=>"000000011",
  49624=>"111101100",
  49625=>"010111011",
  49626=>"000010011",
  49627=>"101011110",
  49628=>"000111110",
  49629=>"011101101",
  49630=>"011011001",
  49631=>"110110110",
  49632=>"001000100",
  49633=>"101000100",
  49634=>"000101111",
  49635=>"010010101",
  49636=>"001111001",
  49637=>"010011011",
  49638=>"000101111",
  49639=>"111111111",
  49640=>"111100010",
  49641=>"101100101",
  49642=>"110011001",
  49643=>"000100000",
  49644=>"000100010",
  49645=>"111010100",
  49646=>"000100001",
  49647=>"000010011",
  49648=>"101011100",
  49649=>"010011110",
  49650=>"001001011",
  49651=>"110101011",
  49652=>"111000000",
  49653=>"100111111",
  49654=>"011010001",
  49655=>"011111011",
  49656=>"100011010",
  49657=>"111111010",
  49658=>"111100000",
  49659=>"001100000",
  49660=>"110111111",
  49661=>"101000000",
  49662=>"001010000",
  49663=>"101010001",
  49664=>"000101001",
  49665=>"001010101",
  49666=>"110001101",
  49667=>"010110010",
  49668=>"101110011",
  49669=>"100010000",
  49670=>"011001001",
  49671=>"100000110",
  49672=>"100111101",
  49673=>"011001001",
  49674=>"111110010",
  49675=>"100100011",
  49676=>"011111100",
  49677=>"010011110",
  49678=>"011101001",
  49679=>"101100000",
  49680=>"111000101",
  49681=>"101100011",
  49682=>"111100010",
  49683=>"111110000",
  49684=>"011001101",
  49685=>"011001110",
  49686=>"100011101",
  49687=>"011011000",
  49688=>"100000001",
  49689=>"001001110",
  49690=>"001000010",
  49691=>"111100011",
  49692=>"111010011",
  49693=>"111001100",
  49694=>"011100101",
  49695=>"001001001",
  49696=>"000101110",
  49697=>"101100101",
  49698=>"100100111",
  49699=>"010001011",
  49700=>"111111110",
  49701=>"010110011",
  49702=>"100010110",
  49703=>"001001001",
  49704=>"010010010",
  49705=>"111000111",
  49706=>"001101001",
  49707=>"000100010",
  49708=>"101010011",
  49709=>"000010110",
  49710=>"100010110",
  49711=>"001011001",
  49712=>"000001000",
  49713=>"101000111",
  49714=>"110010100",
  49715=>"100010011",
  49716=>"110000101",
  49717=>"100011101",
  49718=>"011100001",
  49719=>"111010111",
  49720=>"101011101",
  49721=>"100110100",
  49722=>"101100000",
  49723=>"111010000",
  49724=>"001011011",
  49725=>"001110111",
  49726=>"000101110",
  49727=>"111000111",
  49728=>"110011010",
  49729=>"101000001",
  49730=>"010010110",
  49731=>"101100000",
  49732=>"101011100",
  49733=>"010111111",
  49734=>"000011111",
  49735=>"101010111",
  49736=>"111111000",
  49737=>"000111101",
  49738=>"110000000",
  49739=>"110001001",
  49740=>"100001010",
  49741=>"010101011",
  49742=>"101110000",
  49743=>"100000101",
  49744=>"010010110",
  49745=>"010011100",
  49746=>"110001000",
  49747=>"111000110",
  49748=>"101001000",
  49749=>"011000100",
  49750=>"101010101",
  49751=>"000010000",
  49752=>"010010101",
  49753=>"100000100",
  49754=>"001011100",
  49755=>"101100111",
  49756=>"100000100",
  49757=>"000101010",
  49758=>"100001101",
  49759=>"110101011",
  49760=>"000111111",
  49761=>"011010100",
  49762=>"110011010",
  49763=>"111100100",
  49764=>"111011000",
  49765=>"011001111",
  49766=>"110110000",
  49767=>"000011011",
  49768=>"111011101",
  49769=>"110111011",
  49770=>"001101010",
  49771=>"110100110",
  49772=>"100110011",
  49773=>"011011010",
  49774=>"011010001",
  49775=>"110101001",
  49776=>"000001111",
  49777=>"000001000",
  49778=>"100110000",
  49779=>"000110100",
  49780=>"111000010",
  49781=>"001101010",
  49782=>"001100000",
  49783=>"100100111",
  49784=>"101110100",
  49785=>"011111000",
  49786=>"111001110",
  49787=>"000100100",
  49788=>"100101111",
  49789=>"101100000",
  49790=>"101100111",
  49791=>"011101001",
  49792=>"001100110",
  49793=>"101111111",
  49794=>"111110101",
  49795=>"000011011",
  49796=>"001111111",
  49797=>"010110110",
  49798=>"001000010",
  49799=>"001011001",
  49800=>"110110111",
  49801=>"010100001",
  49802=>"111100100",
  49803=>"111001001",
  49804=>"011000000",
  49805=>"011001101",
  49806=>"011001000",
  49807=>"100000100",
  49808=>"111100000",
  49809=>"000101111",
  49810=>"101000000",
  49811=>"111011100",
  49812=>"100000111",
  49813=>"001000011",
  49814=>"001101110",
  49815=>"110111110",
  49816=>"001110110",
  49817=>"001110011",
  49818=>"101110010",
  49819=>"010111010",
  49820=>"000010000",
  49821=>"111001101",
  49822=>"010011000",
  49823=>"111100001",
  49824=>"010000001",
  49825=>"000101100",
  49826=>"111001101",
  49827=>"000111111",
  49828=>"110010010",
  49829=>"111101100",
  49830=>"000101001",
  49831=>"010000111",
  49832=>"011111100",
  49833=>"010000110",
  49834=>"111111001",
  49835=>"101111010",
  49836=>"001011001",
  49837=>"111010110",
  49838=>"001010101",
  49839=>"100000001",
  49840=>"111101011",
  49841=>"111010100",
  49842=>"100111111",
  49843=>"010010011",
  49844=>"110111001",
  49845=>"101100011",
  49846=>"111010110",
  49847=>"111110010",
  49848=>"110111111",
  49849=>"111110001",
  49850=>"101001111",
  49851=>"110010110",
  49852=>"001001010",
  49853=>"001011100",
  49854=>"011000010",
  49855=>"000001001",
  49856=>"010101011",
  49857=>"011101001",
  49858=>"110101011",
  49859=>"100100010",
  49860=>"100011101",
  49861=>"111011111",
  49862=>"010000000",
  49863=>"000101010",
  49864=>"110011000",
  49865=>"100101100",
  49866=>"010101101",
  49867=>"000011001",
  49868=>"010110100",
  49869=>"010010000",
  49870=>"001001101",
  49871=>"011111100",
  49872=>"110000110",
  49873=>"101001111",
  49874=>"010101111",
  49875=>"010011010",
  49876=>"111111010",
  49877=>"111011111",
  49878=>"001101110",
  49879=>"100111000",
  49880=>"010100001",
  49881=>"111001111",
  49882=>"010000100",
  49883=>"111001111",
  49884=>"110101011",
  49885=>"111100011",
  49886=>"111010000",
  49887=>"110110010",
  49888=>"000000101",
  49889=>"000100010",
  49890=>"111011000",
  49891=>"000110010",
  49892=>"111011010",
  49893=>"111011110",
  49894=>"001101101",
  49895=>"000100000",
  49896=>"110100100",
  49897=>"101001111",
  49898=>"111101101",
  49899=>"011110111",
  49900=>"000000101",
  49901=>"000110100",
  49902=>"101101001",
  49903=>"011010000",
  49904=>"111001001",
  49905=>"100000101",
  49906=>"100110110",
  49907=>"010000100",
  49908=>"100001010",
  49909=>"110001000",
  49910=>"111001000",
  49911=>"101010100",
  49912=>"011010001",
  49913=>"011011011",
  49914=>"100011111",
  49915=>"110001110",
  49916=>"101100001",
  49917=>"100100000",
  49918=>"011101000",
  49919=>"100010000",
  49920=>"111010101",
  49921=>"100011111",
  49922=>"110010010",
  49923=>"100110111",
  49924=>"101100110",
  49925=>"001000001",
  49926=>"111101000",
  49927=>"110010101",
  49928=>"101000100",
  49929=>"111101101",
  49930=>"111101010",
  49931=>"001011110",
  49932=>"011001011",
  49933=>"111100101",
  49934=>"000110100",
  49935=>"000110111",
  49936=>"000100111",
  49937=>"001010010",
  49938=>"101011110",
  49939=>"100110100",
  49940=>"000111110",
  49941=>"100100000",
  49942=>"011100111",
  49943=>"010111000",
  49944=>"110010010",
  49945=>"001100101",
  49946=>"101100000",
  49947=>"111001010",
  49948=>"101001000",
  49949=>"111011000",
  49950=>"001110001",
  49951=>"100101011",
  49952=>"011000100",
  49953=>"111111101",
  49954=>"001110101",
  49955=>"100001010",
  49956=>"011100001",
  49957=>"010010110",
  49958=>"011101000",
  49959=>"001010001",
  49960=>"111101101",
  49961=>"101110011",
  49962=>"000011111",
  49963=>"011001110",
  49964=>"100000011",
  49965=>"010001000",
  49966=>"101010001",
  49967=>"001000111",
  49968=>"010000110",
  49969=>"010111000",
  49970=>"101110010",
  49971=>"010010100",
  49972=>"111011100",
  49973=>"010101000",
  49974=>"010101111",
  49975=>"001011011",
  49976=>"101110011",
  49977=>"101010000",
  49978=>"001111110",
  49979=>"011111010",
  49980=>"010100011",
  49981=>"010111010",
  49982=>"101000010",
  49983=>"011001000",
  49984=>"111101011",
  49985=>"100100111",
  49986=>"010010001",
  49987=>"011100100",
  49988=>"110011001",
  49989=>"111000001",
  49990=>"001000000",
  49991=>"010100000",
  49992=>"011111000",
  49993=>"000010101",
  49994=>"100110011",
  49995=>"110001001",
  49996=>"101010101",
  49997=>"110000101",
  49998=>"110100100",
  49999=>"100001001",
  50000=>"011010011",
  50001=>"000001011",
  50002=>"110100010",
  50003=>"110000001",
  50004=>"010001101",
  50005=>"111000001",
  50006=>"000100111",
  50007=>"101101100",
  50008=>"001011111",
  50009=>"000111010",
  50010=>"001110101",
  50011=>"110000001",
  50012=>"101110100",
  50013=>"111100001",
  50014=>"101011001",
  50015=>"100101110",
  50016=>"110000100",
  50017=>"011111010",
  50018=>"001100111",
  50019=>"110110011",
  50020=>"100000101",
  50021=>"111010010",
  50022=>"010001111",
  50023=>"100111110",
  50024=>"110100111",
  50025=>"010000000",
  50026=>"011111101",
  50027=>"000001010",
  50028=>"100111010",
  50029=>"001101010",
  50030=>"001101111",
  50031=>"100011010",
  50032=>"010000100",
  50033=>"010110101",
  50034=>"010010100",
  50035=>"001101111",
  50036=>"011111100",
  50037=>"100000011",
  50038=>"111110010",
  50039=>"110010001",
  50040=>"100111001",
  50041=>"010001111",
  50042=>"010111101",
  50043=>"010010000",
  50044=>"000111111",
  50045=>"100000100",
  50046=>"110010000",
  50047=>"100101001",
  50048=>"111111000",
  50049=>"011011100",
  50050=>"110011010",
  50051=>"110110011",
  50052=>"010110001",
  50053=>"111010100",
  50054=>"110100110",
  50055=>"100110110",
  50056=>"110110011",
  50057=>"011000100",
  50058=>"100101110",
  50059=>"111100100",
  50060=>"000111111",
  50061=>"010100000",
  50062=>"100001110",
  50063=>"011011010",
  50064=>"000000101",
  50065=>"100101100",
  50066=>"001101000",
  50067=>"100001000",
  50068=>"110101101",
  50069=>"001010010",
  50070=>"010111111",
  50071=>"011111000",
  50072=>"110000011",
  50073=>"000100010",
  50074=>"100000010",
  50075=>"010001010",
  50076=>"101001000",
  50077=>"101010100",
  50078=>"010011100",
  50079=>"000110011",
  50080=>"011000010",
  50081=>"011110000",
  50082=>"110100110",
  50083=>"011100111",
  50084=>"001001101",
  50085=>"101011001",
  50086=>"010111111",
  50087=>"010011110",
  50088=>"010110100",
  50089=>"000110010",
  50090=>"110111010",
  50091=>"001010011",
  50092=>"011000100",
  50093=>"000001110",
  50094=>"101000110",
  50095=>"011101111",
  50096=>"001001111",
  50097=>"111111110",
  50098=>"011010011",
  50099=>"100010001",
  50100=>"100110011",
  50101=>"001011111",
  50102=>"110011010",
  50103=>"010110101",
  50104=>"101001010",
  50105=>"010001100",
  50106=>"001001100",
  50107=>"011010111",
  50108=>"100011000",
  50109=>"100000011",
  50110=>"111011100",
  50111=>"010100111",
  50112=>"111111111",
  50113=>"010110101",
  50114=>"000101110",
  50115=>"011011001",
  50116=>"101111101",
  50117=>"010001011",
  50118=>"111010011",
  50119=>"111111010",
  50120=>"111011100",
  50121=>"001100100",
  50122=>"101101110",
  50123=>"101011011",
  50124=>"001000000",
  50125=>"110101100",
  50126=>"010110100",
  50127=>"011000101",
  50128=>"111001000",
  50129=>"000010000",
  50130=>"111100100",
  50131=>"101000001",
  50132=>"001011101",
  50133=>"111110111",
  50134=>"001101111",
  50135=>"101000010",
  50136=>"000101101",
  50137=>"010101001",
  50138=>"010011001",
  50139=>"000001101",
  50140=>"110000111",
  50141=>"001010001",
  50142=>"101110011",
  50143=>"111100100",
  50144=>"010101001",
  50145=>"111100100",
  50146=>"101110011",
  50147=>"111111110",
  50148=>"100011000",
  50149=>"111111100",
  50150=>"000001010",
  50151=>"110101001",
  50152=>"111001100",
  50153=>"010111010",
  50154=>"001011010",
  50155=>"111110100",
  50156=>"110010100",
  50157=>"000100110",
  50158=>"011111001",
  50159=>"001101101",
  50160=>"110100011",
  50161=>"010011001",
  50162=>"011100100",
  50163=>"101000111",
  50164=>"111100111",
  50165=>"100000000",
  50166=>"101110000",
  50167=>"010111110",
  50168=>"101111010",
  50169=>"010100000",
  50170=>"100100101",
  50171=>"110100000",
  50172=>"100110001",
  50173=>"110010001",
  50174=>"101111110",
  50175=>"110001100",
  50176=>"001001000",
  50177=>"011101011",
  50178=>"000010100",
  50179=>"011111100",
  50180=>"110001010",
  50181=>"101101011",
  50182=>"001010110",
  50183=>"101100000",
  50184=>"011011100",
  50185=>"100100110",
  50186=>"111000101",
  50187=>"010111110",
  50188=>"111000000",
  50189=>"000001000",
  50190=>"101000111",
  50191=>"111011111",
  50192=>"111000111",
  50193=>"000110100",
  50194=>"110101000",
  50195=>"010111111",
  50196=>"100011110",
  50197=>"110000101",
  50198=>"110001010",
  50199=>"000100010",
  50200=>"110000001",
  50201=>"111001101",
  50202=>"011100100",
  50203=>"011010111",
  50204=>"101010001",
  50205=>"000100111",
  50206=>"111110100",
  50207=>"011110001",
  50208=>"011110010",
  50209=>"000001111",
  50210=>"111011010",
  50211=>"011110110",
  50212=>"010111111",
  50213=>"100001011",
  50214=>"000000011",
  50215=>"100101011",
  50216=>"011000010",
  50217=>"000000111",
  50218=>"010100101",
  50219=>"101010001",
  50220=>"011001000",
  50221=>"101011000",
  50222=>"000011101",
  50223=>"001000100",
  50224=>"110101100",
  50225=>"010101000",
  50226=>"000100000",
  50227=>"100011010",
  50228=>"011000010",
  50229=>"101101010",
  50230=>"101001101",
  50231=>"010111010",
  50232=>"100000100",
  50233=>"100001111",
  50234=>"100011101",
  50235=>"110101101",
  50236=>"001100010",
  50237=>"110100100",
  50238=>"111011000",
  50239=>"001001010",
  50240=>"011010001",
  50241=>"000110101",
  50242=>"011111100",
  50243=>"001011010",
  50244=>"101101101",
  50245=>"010100110",
  50246=>"100101100",
  50247=>"100101111",
  50248=>"101010110",
  50249=>"110100101",
  50250=>"001100111",
  50251=>"001100011",
  50252=>"100001010",
  50253=>"111001010",
  50254=>"111111111",
  50255=>"100100000",
  50256=>"010110010",
  50257=>"100011111",
  50258=>"100001001",
  50259=>"101011000",
  50260=>"110111000",
  50261=>"111010010",
  50262=>"010011110",
  50263=>"100011111",
  50264=>"011001000",
  50265=>"010100101",
  50266=>"101011100",
  50267=>"010000010",
  50268=>"100011101",
  50269=>"001000100",
  50270=>"000110110",
  50271=>"100011000",
  50272=>"111101101",
  50273=>"111111101",
  50274=>"011111001",
  50275=>"001100000",
  50276=>"011010001",
  50277=>"101101101",
  50278=>"101010011",
  50279=>"001111111",
  50280=>"001101100",
  50281=>"111001010",
  50282=>"110000011",
  50283=>"010111011",
  50284=>"011101011",
  50285=>"011110100",
  50286=>"110110110",
  50287=>"011000111",
  50288=>"000000011",
  50289=>"000101000",
  50290=>"011001011",
  50291=>"111100110",
  50292=>"000011010",
  50293=>"110011001",
  50294=>"100100110",
  50295=>"011100010",
  50296=>"011010000",
  50297=>"110101000",
  50298=>"000100100",
  50299=>"101001111",
  50300=>"011000011",
  50301=>"001010001",
  50302=>"011110111",
  50303=>"010110110",
  50304=>"111001100",
  50305=>"110101111",
  50306=>"000111010",
  50307=>"001001011",
  50308=>"000001000",
  50309=>"100010010",
  50310=>"111010001",
  50311=>"011110000",
  50312=>"000000001",
  50313=>"100001101",
  50314=>"011100100",
  50315=>"101010000",
  50316=>"110001101",
  50317=>"101000001",
  50318=>"101110100",
  50319=>"101110100",
  50320=>"011111101",
  50321=>"101100111",
  50322=>"101010111",
  50323=>"111011110",
  50324=>"000001111",
  50325=>"011010000",
  50326=>"011010011",
  50327=>"100001101",
  50328=>"000000100",
  50329=>"101011110",
  50330=>"111111011",
  50331=>"011000101",
  50332=>"001100001",
  50333=>"010010011",
  50334=>"101000111",
  50335=>"111011010",
  50336=>"001100010",
  50337=>"110110101",
  50338=>"111000100",
  50339=>"100010101",
  50340=>"010001011",
  50341=>"100101000",
  50342=>"100101111",
  50343=>"001100100",
  50344=>"110001111",
  50345=>"100101001",
  50346=>"111111011",
  50347=>"001100011",
  50348=>"011111110",
  50349=>"010010000",
  50350=>"101110100",
  50351=>"010011110",
  50352=>"110011000",
  50353=>"000011010",
  50354=>"001000010",
  50355=>"011100100",
  50356=>"110100010",
  50357=>"101010100",
  50358=>"010010011",
  50359=>"000000000",
  50360=>"000001010",
  50361=>"000001001",
  50362=>"000100010",
  50363=>"001111110",
  50364=>"111110000",
  50365=>"010010010",
  50366=>"100100111",
  50367=>"011100000",
  50368=>"110110101",
  50369=>"111001001",
  50370=>"001111000",
  50371=>"101110010",
  50372=>"010001111",
  50373=>"001000010",
  50374=>"010000100",
  50375=>"001010111",
  50376=>"011011000",
  50377=>"100010001",
  50378=>"001000010",
  50379=>"101010010",
  50380=>"010001010",
  50381=>"110010000",
  50382=>"000010001",
  50383=>"111101010",
  50384=>"111101111",
  50385=>"011001001",
  50386=>"100101000",
  50387=>"001111001",
  50388=>"100000110",
  50389=>"101100110",
  50390=>"110110100",
  50391=>"010011010",
  50392=>"110001101",
  50393=>"101011011",
  50394=>"000101001",
  50395=>"010000111",
  50396=>"011111011",
  50397=>"101000010",
  50398=>"000100011",
  50399=>"010110111",
  50400=>"101011101",
  50401=>"101111110",
  50402=>"001100000",
  50403=>"001000100",
  50404=>"101110010",
  50405=>"011001100",
  50406=>"001011010",
  50407=>"111001111",
  50408=>"100100000",
  50409=>"001101001",
  50410=>"100001101",
  50411=>"101011011",
  50412=>"000111000",
  50413=>"010101110",
  50414=>"101111011",
  50415=>"000011100",
  50416=>"001010101",
  50417=>"110110110",
  50418=>"011001000",
  50419=>"010011010",
  50420=>"010100100",
  50421=>"010000011",
  50422=>"101001110",
  50423=>"111011111",
  50424=>"000011111",
  50425=>"010110011",
  50426=>"110110111",
  50427=>"010011000",
  50428=>"010000111",
  50429=>"101110110",
  50430=>"001111010",
  50431=>"000100000",
  50432=>"010010100",
  50433=>"001011010",
  50434=>"110100101",
  50435=>"100001101",
  50436=>"000101000",
  50437=>"101001101",
  50438=>"101000110",
  50439=>"111001101",
  50440=>"000101001",
  50441=>"011110111",
  50442=>"100010101",
  50443=>"011000010",
  50444=>"101001101",
  50445=>"000110000",
  50446=>"110000000",
  50447=>"000111101",
  50448=>"100000101",
  50449=>"000011110",
  50450=>"000111111",
  50451=>"000111001",
  50452=>"011010000",
  50453=>"011000001",
  50454=>"100001101",
  50455=>"010100110",
  50456=>"100000010",
  50457=>"001100010",
  50458=>"001001110",
  50459=>"001000010",
  50460=>"010111011",
  50461=>"101001111",
  50462=>"111110111",
  50463=>"100010100",
  50464=>"001000100",
  50465=>"001111010",
  50466=>"000010001",
  50467=>"110101101",
  50468=>"100111110",
  50469=>"000111110",
  50470=>"101000001",
  50471=>"010010001",
  50472=>"100111100",
  50473=>"111010101",
  50474=>"010010011",
  50475=>"000100010",
  50476=>"000001010",
  50477=>"011000000",
  50478=>"001000011",
  50479=>"100101110",
  50480=>"101001101",
  50481=>"010011000",
  50482=>"000000111",
  50483=>"010110101",
  50484=>"000001001",
  50485=>"011100000",
  50486=>"011001100",
  50487=>"111001001",
  50488=>"000101001",
  50489=>"100111100",
  50490=>"000110010",
  50491=>"100010011",
  50492=>"000101011",
  50493=>"111011111",
  50494=>"111000111",
  50495=>"110101101",
  50496=>"000100000",
  50497=>"011001111",
  50498=>"100100111",
  50499=>"111011111",
  50500=>"000011011",
  50501=>"111111001",
  50502=>"101010110",
  50503=>"111111101",
  50504=>"100000101",
  50505=>"101011010",
  50506=>"110110001",
  50507=>"010101011",
  50508=>"011000001",
  50509=>"101011101",
  50510=>"111110111",
  50511=>"101111100",
  50512=>"000000000",
  50513=>"001100110",
  50514=>"111110101",
  50515=>"000000111",
  50516=>"000100000",
  50517=>"000000111",
  50518=>"001110101",
  50519=>"001101011",
  50520=>"000101001",
  50521=>"000100110",
  50522=>"010100001",
  50523=>"100000001",
  50524=>"010100010",
  50525=>"010111101",
  50526=>"010100001",
  50527=>"010101001",
  50528=>"001111000",
  50529=>"001000001",
  50530=>"101001101",
  50531=>"001000001",
  50532=>"100000010",
  50533=>"111000001",
  50534=>"101111101",
  50535=>"100001110",
  50536=>"111100000",
  50537=>"000101101",
  50538=>"011100010",
  50539=>"100101010",
  50540=>"101000101",
  50541=>"111001011",
  50542=>"110011011",
  50543=>"111011101",
  50544=>"110000110",
  50545=>"101110011",
  50546=>"110110010",
  50547=>"100100111",
  50548=>"101100111",
  50549=>"010010000",
  50550=>"100010111",
  50551=>"100010011",
  50552=>"000010110",
  50553=>"010111111",
  50554=>"000100010",
  50555=>"101000001",
  50556=>"010111110",
  50557=>"000010011",
  50558=>"010110111",
  50559=>"000111001",
  50560=>"111001101",
  50561=>"100010110",
  50562=>"001100000",
  50563=>"011010110",
  50564=>"000011000",
  50565=>"000100001",
  50566=>"111110111",
  50567=>"111101001",
  50568=>"110000100",
  50569=>"101000111",
  50570=>"001110000",
  50571=>"100000011",
  50572=>"101001011",
  50573=>"110011000",
  50574=>"011110000",
  50575=>"010001110",
  50576=>"001011110",
  50577=>"010000010",
  50578=>"110101101",
  50579=>"100100101",
  50580=>"010010000",
  50581=>"110101010",
  50582=>"011010101",
  50583=>"100000110",
  50584=>"001110111",
  50585=>"010111000",
  50586=>"010000011",
  50587=>"111111000",
  50588=>"111011101",
  50589=>"111111010",
  50590=>"000011100",
  50591=>"011001000",
  50592=>"010101110",
  50593=>"000000000",
  50594=>"010111000",
  50595=>"000000000",
  50596=>"011101110",
  50597=>"000010010",
  50598=>"011011010",
  50599=>"000000100",
  50600=>"011111110",
  50601=>"010011010",
  50602=>"000011101",
  50603=>"101011011",
  50604=>"010101011",
  50605=>"011101111",
  50606=>"101001000",
  50607=>"010100000",
  50608=>"111011111",
  50609=>"011000110",
  50610=>"001100101",
  50611=>"001000011",
  50612=>"001010011",
  50613=>"111011100",
  50614=>"000111100",
  50615=>"011010011",
  50616=>"001010011",
  50617=>"110111010",
  50618=>"010001101",
  50619=>"011011111",
  50620=>"110110101",
  50621=>"101101010",
  50622=>"001100011",
  50623=>"001110000",
  50624=>"001011110",
  50625=>"100101001",
  50626=>"111110011",
  50627=>"010111010",
  50628=>"010011110",
  50629=>"110010000",
  50630=>"011010100",
  50631=>"000101011",
  50632=>"000001010",
  50633=>"101110011",
  50634=>"110100111",
  50635=>"100011111",
  50636=>"000110001",
  50637=>"001001101",
  50638=>"101001110",
  50639=>"100010010",
  50640=>"100111110",
  50641=>"100010101",
  50642=>"000111000",
  50643=>"011000100",
  50644=>"000100010",
  50645=>"000010010",
  50646=>"110011000",
  50647=>"010000100",
  50648=>"111110011",
  50649=>"000010000",
  50650=>"000000100",
  50651=>"110111101",
  50652=>"100011000",
  50653=>"101101110",
  50654=>"110010110",
  50655=>"001100010",
  50656=>"111001110",
  50657=>"111100111",
  50658=>"011111010",
  50659=>"000010110",
  50660=>"110101110",
  50661=>"111101111",
  50662=>"101111010",
  50663=>"110011100",
  50664=>"000000000",
  50665=>"010110011",
  50666=>"111010001",
  50667=>"010101110",
  50668=>"100000011",
  50669=>"000010000",
  50670=>"000010000",
  50671=>"001100100",
  50672=>"000010000",
  50673=>"100111001",
  50674=>"100100111",
  50675=>"110010010",
  50676=>"001100101",
  50677=>"100000001",
  50678=>"110011011",
  50679=>"100111000",
  50680=>"000001000",
  50681=>"110000110",
  50682=>"000000111",
  50683=>"110000101",
  50684=>"011100101",
  50685=>"001010000",
  50686=>"010010010",
  50687=>"101110101",
  50688=>"101100001",
  50689=>"011101101",
  50690=>"110011110",
  50691=>"001000111",
  50692=>"110111010",
  50693=>"000101011",
  50694=>"100011001",
  50695=>"011100010",
  50696=>"011000011",
  50697=>"000110001",
  50698=>"101100101",
  50699=>"000000010",
  50700=>"110000110",
  50701=>"100001010",
  50702=>"110100101",
  50703=>"011001101",
  50704=>"101011101",
  50705=>"001000101",
  50706=>"001001011",
  50707=>"001101001",
  50708=>"111011000",
  50709=>"111010010",
  50710=>"110110001",
  50711=>"101011111",
  50712=>"111000100",
  50713=>"011110111",
  50714=>"011001001",
  50715=>"110111010",
  50716=>"101101101",
  50717=>"001000101",
  50718=>"111111100",
  50719=>"010000001",
  50720=>"110001001",
  50721=>"110111001",
  50722=>"011101110",
  50723=>"000110001",
  50724=>"001001111",
  50725=>"001001110",
  50726=>"110101000",
  50727=>"101001001",
  50728=>"011100000",
  50729=>"100111101",
  50730=>"000110011",
  50731=>"010010010",
  50732=>"000101100",
  50733=>"001010001",
  50734=>"000011000",
  50735=>"000010000",
  50736=>"001110111",
  50737=>"100111111",
  50738=>"011100110",
  50739=>"001100111",
  50740=>"101101100",
  50741=>"101011000",
  50742=>"110110100",
  50743=>"110000011",
  50744=>"011000011",
  50745=>"001111111",
  50746=>"101100011",
  50747=>"001000011",
  50748=>"001000110",
  50749=>"101011110",
  50750=>"011100000",
  50751=>"000010110",
  50752=>"010000101",
  50753=>"000101010",
  50754=>"111010011",
  50755=>"001100111",
  50756=>"100000010",
  50757=>"000101100",
  50758=>"001000001",
  50759=>"111001001",
  50760=>"111010100",
  50761=>"010101111",
  50762=>"010101110",
  50763=>"000000111",
  50764=>"000110010",
  50765=>"001101001",
  50766=>"111000101",
  50767=>"100111000",
  50768=>"100100001",
  50769=>"000101010",
  50770=>"101001110",
  50771=>"001100000",
  50772=>"000011001",
  50773=>"000111001",
  50774=>"110101000",
  50775=>"000110010",
  50776=>"101110000",
  50777=>"000000110",
  50778=>"010101010",
  50779=>"110101100",
  50780=>"111011010",
  50781=>"001111101",
  50782=>"001111110",
  50783=>"000000001",
  50784=>"111010111",
  50785=>"000001001",
  50786=>"110110001",
  50787=>"101100000",
  50788=>"010010001",
  50789=>"101000110",
  50790=>"010000110",
  50791=>"111110100",
  50792=>"100110110",
  50793=>"111101000",
  50794=>"100111101",
  50795=>"000011000",
  50796=>"011110011",
  50797=>"011011011",
  50798=>"101001001",
  50799=>"010010011",
  50800=>"111001000",
  50801=>"000100001",
  50802=>"011100100",
  50803=>"101101011",
  50804=>"110001000",
  50805=>"011100101",
  50806=>"001010111",
  50807=>"000010010",
  50808=>"110011110",
  50809=>"011111111",
  50810=>"011001000",
  50811=>"110011111",
  50812=>"000110010",
  50813=>"011001010",
  50814=>"000100101",
  50815=>"111100010",
  50816=>"000011101",
  50817=>"011011100",
  50818=>"100000010",
  50819=>"100111101",
  50820=>"100110001",
  50821=>"010010001",
  50822=>"111101011",
  50823=>"101001011",
  50824=>"001000001",
  50825=>"100001000",
  50826=>"011111111",
  50827=>"011111100",
  50828=>"101101010",
  50829=>"001000010",
  50830=>"100011111",
  50831=>"101100001",
  50832=>"100101000",
  50833=>"110100100",
  50834=>"101010010",
  50835=>"010111000",
  50836=>"000100001",
  50837=>"100110100",
  50838=>"101001111",
  50839=>"101110100",
  50840=>"011101100",
  50841=>"010010001",
  50842=>"011001010",
  50843=>"011111001",
  50844=>"101101001",
  50845=>"111010101",
  50846=>"111011011",
  50847=>"110011010",
  50848=>"110011011",
  50849=>"110100011",
  50850=>"110101000",
  50851=>"101001010",
  50852=>"000000101",
  50853=>"100101010",
  50854=>"010110110",
  50855=>"000101110",
  50856=>"000110100",
  50857=>"111100100",
  50858=>"111000101",
  50859=>"100101110",
  50860=>"011110001",
  50861=>"010011010",
  50862=>"111001111",
  50863=>"001100111",
  50864=>"010100111",
  50865=>"101010110",
  50866=>"001001110",
  50867=>"100100100",
  50868=>"000111100",
  50869=>"111110100",
  50870=>"111111000",
  50871=>"001111111",
  50872=>"011010010",
  50873=>"000110011",
  50874=>"010011100",
  50875=>"001000110",
  50876=>"001001110",
  50877=>"010001111",
  50878=>"001111011",
  50879=>"110011110",
  50880=>"111111111",
  50881=>"000110010",
  50882=>"000110101",
  50883=>"110101100",
  50884=>"010011101",
  50885=>"011111110",
  50886=>"110100011",
  50887=>"000111110",
  50888=>"101000110",
  50889=>"111000100",
  50890=>"010011010",
  50891=>"001001010",
  50892=>"001000001",
  50893=>"110001101",
  50894=>"000000110",
  50895=>"111110101",
  50896=>"011100000",
  50897=>"001001110",
  50898=>"001100000",
  50899=>"010010110",
  50900=>"100001011",
  50901=>"100101110",
  50902=>"000110010",
  50903=>"010010010",
  50904=>"110110011",
  50905=>"100001010",
  50906=>"110100001",
  50907=>"011001100",
  50908=>"001100101",
  50909=>"000110010",
  50910=>"010001110",
  50911=>"010111101",
  50912=>"110010110",
  50913=>"001111100",
  50914=>"111100001",
  50915=>"110100111",
  50916=>"001010011",
  50917=>"101111110",
  50918=>"110111000",
  50919=>"011010111",
  50920=>"110111111",
  50921=>"100100011",
  50922=>"001000000",
  50923=>"110000110",
  50924=>"001011111",
  50925=>"111001100",
  50926=>"010100100",
  50927=>"000011110",
  50928=>"100110100",
  50929=>"111100110",
  50930=>"100000111",
  50931=>"101001001",
  50932=>"111001101",
  50933=>"111011001",
  50934=>"001110010",
  50935=>"011100001",
  50936=>"111011101",
  50937=>"001110101",
  50938=>"101000100",
  50939=>"101001000",
  50940=>"101011000",
  50941=>"010111110",
  50942=>"110101011",
  50943=>"100011001",
  50944=>"000011111",
  50945=>"001111000",
  50946=>"010110000",
  50947=>"001100111",
  50948=>"100000100",
  50949=>"101000100",
  50950=>"001111000",
  50951=>"101010101",
  50952=>"011011100",
  50953=>"010101011",
  50954=>"001101111",
  50955=>"101100010",
  50956=>"010010110",
  50957=>"100010001",
  50958=>"111100011",
  50959=>"100001101",
  50960=>"101010000",
  50961=>"100100000",
  50962=>"010010101",
  50963=>"011011111",
  50964=>"101100011",
  50965=>"100110100",
  50966=>"010100001",
  50967=>"001110100",
  50968=>"101000010",
  50969=>"110010000",
  50970=>"010101101",
  50971=>"010011001",
  50972=>"101110000",
  50973=>"010100011",
  50974=>"101110110",
  50975=>"010010000",
  50976=>"010101010",
  50977=>"111010111",
  50978=>"000011000",
  50979=>"100111110",
  50980=>"110100100",
  50981=>"100001001",
  50982=>"010111101",
  50983=>"100011010",
  50984=>"000001111",
  50985=>"100110010",
  50986=>"010111011",
  50987=>"000111010",
  50988=>"110110000",
  50989=>"000110010",
  50990=>"110010111",
  50991=>"111110011",
  50992=>"000110001",
  50993=>"000001101",
  50994=>"100111110",
  50995=>"011000000",
  50996=>"000010000",
  50997=>"111111011",
  50998=>"111101010",
  50999=>"110100001",
  51000=>"110110001",
  51001=>"011101111",
  51002=>"000000100",
  51003=>"110101000",
  51004=>"000101100",
  51005=>"011100010",
  51006=>"111000000",
  51007=>"000101101",
  51008=>"011011011",
  51009=>"000111001",
  51010=>"000000111",
  51011=>"111111011",
  51012=>"011101001",
  51013=>"101110111",
  51014=>"000101110",
  51015=>"000011110",
  51016=>"110010110",
  51017=>"110011111",
  51018=>"001110011",
  51019=>"111100100",
  51020=>"101000011",
  51021=>"000101110",
  51022=>"110111010",
  51023=>"010111001",
  51024=>"010010111",
  51025=>"111101001",
  51026=>"000010111",
  51027=>"010001101",
  51028=>"111110011",
  51029=>"011111001",
  51030=>"010000001",
  51031=>"011111100",
  51032=>"111011111",
  51033=>"110000100",
  51034=>"110110111",
  51035=>"100110101",
  51036=>"011111111",
  51037=>"000011101",
  51038=>"010001100",
  51039=>"101101100",
  51040=>"010001000",
  51041=>"011110001",
  51042=>"000001000",
  51043=>"110000010",
  51044=>"010101011",
  51045=>"000100001",
  51046=>"011110110",
  51047=>"000010100",
  51048=>"000010000",
  51049=>"001011100",
  51050=>"001100011",
  51051=>"000011001",
  51052=>"101111111",
  51053=>"010011010",
  51054=>"110101000",
  51055=>"011101001",
  51056=>"011000010",
  51057=>"000100110",
  51058=>"000100010",
  51059=>"000100101",
  51060=>"111010100",
  51061=>"010100000",
  51062=>"000110001",
  51063=>"110011111",
  51064=>"000010000",
  51065=>"110101010",
  51066=>"111000000",
  51067=>"011110011",
  51068=>"000010110",
  51069=>"111000101",
  51070=>"110111110",
  51071=>"111110001",
  51072=>"000111110",
  51073=>"000101001",
  51074=>"100100100",
  51075=>"110101110",
  51076=>"110111010",
  51077=>"011101001",
  51078=>"101100011",
  51079=>"010110011",
  51080=>"010011110",
  51081=>"100011010",
  51082=>"000111001",
  51083=>"000100011",
  51084=>"111011101",
  51085=>"011011010",
  51086=>"011110000",
  51087=>"010010011",
  51088=>"100110001",
  51089=>"000110010",
  51090=>"101000111",
  51091=>"111110101",
  51092=>"101100010",
  51093=>"100110111",
  51094=>"001000110",
  51095=>"111111010",
  51096=>"001111111",
  51097=>"111110110",
  51098=>"000100010",
  51099=>"101100111",
  51100=>"011100000",
  51101=>"011100000",
  51102=>"101101100",
  51103=>"111100000",
  51104=>"100100001",
  51105=>"101110000",
  51106=>"001000001",
  51107=>"001000001",
  51108=>"000010000",
  51109=>"011000111",
  51110=>"011100110",
  51111=>"100011111",
  51112=>"000010110",
  51113=>"111111111",
  51114=>"110110101",
  51115=>"101100010",
  51116=>"001001000",
  51117=>"100010101",
  51118=>"101101100",
  51119=>"000000011",
  51120=>"110010110",
  51121=>"110001100",
  51122=>"000101111",
  51123=>"100000001",
  51124=>"111111111",
  51125=>"010001011",
  51126=>"100101001",
  51127=>"100110111",
  51128=>"100100000",
  51129=>"010010110",
  51130=>"101111111",
  51131=>"001001111",
  51132=>"010111111",
  51133=>"110000110",
  51134=>"111111110",
  51135=>"011111000",
  51136=>"110110011",
  51137=>"110111001",
  51138=>"110110000",
  51139=>"111001110",
  51140=>"000111111",
  51141=>"101010110",
  51142=>"001110010",
  51143=>"000010110",
  51144=>"011111111",
  51145=>"010001000",
  51146=>"010111001",
  51147=>"011100011",
  51148=>"111011110",
  51149=>"010100000",
  51150=>"100000110",
  51151=>"001000001",
  51152=>"100100111",
  51153=>"011110001",
  51154=>"000110111",
  51155=>"010100000",
  51156=>"000010010",
  51157=>"110101100",
  51158=>"101011010",
  51159=>"010100010",
  51160=>"001010111",
  51161=>"001010000",
  51162=>"111000001",
  51163=>"100010100",
  51164=>"001001011",
  51165=>"100101001",
  51166=>"110010011",
  51167=>"110010101",
  51168=>"001011000",
  51169=>"011000010",
  51170=>"010011000",
  51171=>"111000010",
  51172=>"001000100",
  51173=>"000010000",
  51174=>"011101010",
  51175=>"111111000",
  51176=>"011100111",
  51177=>"010111110",
  51178=>"011001111",
  51179=>"101001101",
  51180=>"111110110",
  51181=>"101101110",
  51182=>"010000111",
  51183=>"000001011",
  51184=>"111000000",
  51185=>"110001001",
  51186=>"101111101",
  51187=>"001000101",
  51188=>"100000000",
  51189=>"110110100",
  51190=>"010001001",
  51191=>"000101011",
  51192=>"110010111",
  51193=>"101101011",
  51194=>"110100101",
  51195=>"101001000",
  51196=>"011000111",
  51197=>"110100110",
  51198=>"110011010",
  51199=>"100010011",
  51200=>"000011100",
  51201=>"011011100",
  51202=>"101101000",
  51203=>"001010101",
  51204=>"101001010",
  51205=>"100111111",
  51206=>"011000010",
  51207=>"111111110",
  51208=>"001000100",
  51209=>"101001001",
  51210=>"111110010",
  51211=>"010010101",
  51212=>"001011011",
  51213=>"110110100",
  51214=>"001010010",
  51215=>"111111000",
  51216=>"000010001",
  51217=>"110101010",
  51218=>"001010110",
  51219=>"110011110",
  51220=>"001101011",
  51221=>"110100110",
  51222=>"010100110",
  51223=>"000100101",
  51224=>"001001011",
  51225=>"100011000",
  51226=>"101110101",
  51227=>"000111111",
  51228=>"001100001",
  51229=>"000010011",
  51230=>"000111110",
  51231=>"010010110",
  51232=>"001001001",
  51233=>"100111001",
  51234=>"100101111",
  51235=>"001111010",
  51236=>"000001110",
  51237=>"111011000",
  51238=>"001000100",
  51239=>"111110001",
  51240=>"010111010",
  51241=>"001001100",
  51242=>"001010011",
  51243=>"111011000",
  51244=>"010110111",
  51245=>"010111001",
  51246=>"000111110",
  51247=>"101000111",
  51248=>"110111101",
  51249=>"001000000",
  51250=>"001110000",
  51251=>"000100010",
  51252=>"000000010",
  51253=>"001111111",
  51254=>"111010010",
  51255=>"110110111",
  51256=>"001000111",
  51257=>"000000000",
  51258=>"100001111",
  51259=>"110000110",
  51260=>"111101111",
  51261=>"000100111",
  51262=>"010000110",
  51263=>"110011111",
  51264=>"101101101",
  51265=>"000100001",
  51266=>"011110101",
  51267=>"111010111",
  51268=>"001010111",
  51269=>"000010111",
  51270=>"101101010",
  51271=>"000110000",
  51272=>"101011010",
  51273=>"101101010",
  51274=>"010110110",
  51275=>"000011000",
  51276=>"001110101",
  51277=>"010110110",
  51278=>"011011101",
  51279=>"100100101",
  51280=>"010111011",
  51281=>"010011011",
  51282=>"010100001",
  51283=>"001000000",
  51284=>"000111100",
  51285=>"100101000",
  51286=>"100111000",
  51287=>"000001010",
  51288=>"010011000",
  51289=>"010011101",
  51290=>"110110100",
  51291=>"110010101",
  51292=>"001111010",
  51293=>"110000010",
  51294=>"000000010",
  51295=>"000001110",
  51296=>"010010100",
  51297=>"000000111",
  51298=>"101100110",
  51299=>"010000011",
  51300=>"111010110",
  51301=>"100000101",
  51302=>"111110011",
  51303=>"010001011",
  51304=>"100111001",
  51305=>"111010110",
  51306=>"010101001",
  51307=>"100011110",
  51308=>"111000010",
  51309=>"100100100",
  51310=>"101000101",
  51311=>"101010101",
  51312=>"001010111",
  51313=>"011101011",
  51314=>"010011111",
  51315=>"001100110",
  51316=>"001110001",
  51317=>"000111010",
  51318=>"111001100",
  51319=>"100101101",
  51320=>"011000011",
  51321=>"011010001",
  51322=>"011001100",
  51323=>"000101100",
  51324=>"010110011",
  51325=>"000111010",
  51326=>"000010111",
  51327=>"110100010",
  51328=>"011010011",
  51329=>"101100010",
  51330=>"001010011",
  51331=>"100110110",
  51332=>"001111011",
  51333=>"101111010",
  51334=>"101000000",
  51335=>"110110010",
  51336=>"101111011",
  51337=>"000010000",
  51338=>"010100110",
  51339=>"111111111",
  51340=>"100000010",
  51341=>"110001101",
  51342=>"111011111",
  51343=>"101101100",
  51344=>"001010111",
  51345=>"101101000",
  51346=>"100111001",
  51347=>"101111000",
  51348=>"010101111",
  51349=>"010110101",
  51350=>"000110110",
  51351=>"010111000",
  51352=>"111100101",
  51353=>"111100100",
  51354=>"000111110",
  51355=>"111110001",
  51356=>"000010101",
  51357=>"101110101",
  51358=>"010010100",
  51359=>"011101011",
  51360=>"100010110",
  51361=>"100110111",
  51362=>"110001001",
  51363=>"001111001",
  51364=>"010011100",
  51365=>"101100110",
  51366=>"000001000",
  51367=>"001110000",
  51368=>"010011010",
  51369=>"101101010",
  51370=>"111011011",
  51371=>"110000111",
  51372=>"101100100",
  51373=>"001101001",
  51374=>"011010011",
  51375=>"011000100",
  51376=>"110001100",
  51377=>"110011110",
  51378=>"001000101",
  51379=>"101010111",
  51380=>"111100000",
  51381=>"110100101",
  51382=>"001111001",
  51383=>"011011000",
  51384=>"000100110",
  51385=>"011111001",
  51386=>"001011110",
  51387=>"011100101",
  51388=>"001101110",
  51389=>"101110011",
  51390=>"010000011",
  51391=>"110100010",
  51392=>"110000001",
  51393=>"010000110",
  51394=>"000010000",
  51395=>"110111101",
  51396=>"001100000",
  51397=>"100110011",
  51398=>"000110111",
  51399=>"110110011",
  51400=>"100011010",
  51401=>"010101011",
  51402=>"110101111",
  51403=>"011100001",
  51404=>"100010010",
  51405=>"110000101",
  51406=>"000011011",
  51407=>"110011100",
  51408=>"010011101",
  51409=>"111110001",
  51410=>"000010100",
  51411=>"001100111",
  51412=>"101010110",
  51413=>"101111111",
  51414=>"001011010",
  51415=>"001101101",
  51416=>"110000110",
  51417=>"011000111",
  51418=>"100010010",
  51419=>"001001100",
  51420=>"000011011",
  51421=>"010010111",
  51422=>"111110110",
  51423=>"111100111",
  51424=>"111111001",
  51425=>"011010110",
  51426=>"110010000",
  51427=>"011000110",
  51428=>"110000100",
  51429=>"101101011",
  51430=>"011111110",
  51431=>"110000010",
  51432=>"111101111",
  51433=>"010101111",
  51434=>"111110001",
  51435=>"000001101",
  51436=>"101100001",
  51437=>"011100011",
  51438=>"111101001",
  51439=>"011001110",
  51440=>"000101111",
  51441=>"101111011",
  51442=>"010001101",
  51443=>"111111010",
  51444=>"001100100",
  51445=>"101011011",
  51446=>"111101101",
  51447=>"000101110",
  51448=>"100111110",
  51449=>"010111110",
  51450=>"000010101",
  51451=>"100010001",
  51452=>"000000000",
  51453=>"011011001",
  51454=>"100100000",
  51455=>"000011000",
  51456=>"100111111",
  51457=>"100110111",
  51458=>"111101100",
  51459=>"000001110",
  51460=>"101011001",
  51461=>"111010010",
  51462=>"101101010",
  51463=>"111011100",
  51464=>"111100010",
  51465=>"100011011",
  51466=>"011110010",
  51467=>"010111010",
  51468=>"000110111",
  51469=>"101010100",
  51470=>"110111011",
  51471=>"000000010",
  51472=>"001000111",
  51473=>"000111111",
  51474=>"011100010",
  51475=>"100111110",
  51476=>"111110101",
  51477=>"110111011",
  51478=>"101011110",
  51479=>"000001011",
  51480=>"011011101",
  51481=>"110011100",
  51482=>"110000111",
  51483=>"101011000",
  51484=>"111001111",
  51485=>"001111101",
  51486=>"011011101",
  51487=>"000010101",
  51488=>"111101001",
  51489=>"101000000",
  51490=>"101001111",
  51491=>"011001111",
  51492=>"010010000",
  51493=>"100000111",
  51494=>"011010010",
  51495=>"101111101",
  51496=>"001010110",
  51497=>"000111111",
  51498=>"101101101",
  51499=>"101001001",
  51500=>"100001001",
  51501=>"101010100",
  51502=>"100010100",
  51503=>"011110011",
  51504=>"011010000",
  51505=>"000010010",
  51506=>"100100101",
  51507=>"010000110",
  51508=>"010110110",
  51509=>"001110111",
  51510=>"010110011",
  51511=>"010001000",
  51512=>"011001101",
  51513=>"100001101",
  51514=>"001111101",
  51515=>"011011011",
  51516=>"010111010",
  51517=>"011110100",
  51518=>"000011001",
  51519=>"011111000",
  51520=>"000101000",
  51521=>"101101111",
  51522=>"101000000",
  51523=>"110011000",
  51524=>"111011111",
  51525=>"101101100",
  51526=>"111000010",
  51527=>"101100000",
  51528=>"111101101",
  51529=>"010100010",
  51530=>"000011111",
  51531=>"001011010",
  51532=>"000010001",
  51533=>"101111111",
  51534=>"110000010",
  51535=>"000000101",
  51536=>"101111000",
  51537=>"010100110",
  51538=>"000100111",
  51539=>"011100000",
  51540=>"010110001",
  51541=>"011110100",
  51542=>"010011101",
  51543=>"010000000",
  51544=>"101001110",
  51545=>"110000100",
  51546=>"011001000",
  51547=>"010000111",
  51548=>"101100110",
  51549=>"111101101",
  51550=>"000001110",
  51551=>"111011010",
  51552=>"011100111",
  51553=>"001000111",
  51554=>"000011001",
  51555=>"100000100",
  51556=>"100111101",
  51557=>"000011000",
  51558=>"001100000",
  51559=>"101101111",
  51560=>"000001011",
  51561=>"110010010",
  51562=>"101111111",
  51563=>"000111000",
  51564=>"001101111",
  51565=>"000101110",
  51566=>"101001001",
  51567=>"011010010",
  51568=>"111110010",
  51569=>"100101110",
  51570=>"110000001",
  51571=>"010111101",
  51572=>"110101101",
  51573=>"011101111",
  51574=>"110101110",
  51575=>"000011001",
  51576=>"100101010",
  51577=>"111011101",
  51578=>"001111001",
  51579=>"000001000",
  51580=>"101011101",
  51581=>"111110010",
  51582=>"010111000",
  51583=>"100100100",
  51584=>"011100111",
  51585=>"111010010",
  51586=>"010011001",
  51587=>"111101010",
  51588=>"111111011",
  51589=>"100100111",
  51590=>"011111111",
  51591=>"010100011",
  51592=>"010101010",
  51593=>"001111010",
  51594=>"001110001",
  51595=>"111100001",
  51596=>"000101101",
  51597=>"010011001",
  51598=>"110000100",
  51599=>"011111100",
  51600=>"111010100",
  51601=>"110000100",
  51602=>"000101001",
  51603=>"010100010",
  51604=>"110111001",
  51605=>"001010101",
  51606=>"000010010",
  51607=>"100010011",
  51608=>"001100101",
  51609=>"011000100",
  51610=>"011100011",
  51611=>"001111101",
  51612=>"010100111",
  51613=>"011011001",
  51614=>"011011011",
  51615=>"100101000",
  51616=>"011110000",
  51617=>"010010100",
  51618=>"101000010",
  51619=>"111101111",
  51620=>"001000100",
  51621=>"000001011",
  51622=>"101001001",
  51623=>"110011100",
  51624=>"101010001",
  51625=>"010001001",
  51626=>"101101011",
  51627=>"001100111",
  51628=>"011000000",
  51629=>"111000010",
  51630=>"101001010",
  51631=>"010010000",
  51632=>"011100011",
  51633=>"001101000",
  51634=>"011001000",
  51635=>"001010001",
  51636=>"111111001",
  51637=>"110010110",
  51638=>"000011001",
  51639=>"100010100",
  51640=>"101100101",
  51641=>"110000110",
  51642=>"010000000",
  51643=>"100001011",
  51644=>"011111010",
  51645=>"111101010",
  51646=>"100110001",
  51647=>"101100111",
  51648=>"001000111",
  51649=>"010100101",
  51650=>"111011100",
  51651=>"010100111",
  51652=>"011110111",
  51653=>"000100101",
  51654=>"101101100",
  51655=>"011010111",
  51656=>"010000000",
  51657=>"101011011",
  51658=>"011010110",
  51659=>"101100001",
  51660=>"001110010",
  51661=>"101000101",
  51662=>"001101010",
  51663=>"001010001",
  51664=>"000011000",
  51665=>"010000110",
  51666=>"100001000",
  51667=>"000110000",
  51668=>"000011111",
  51669=>"011001110",
  51670=>"101110110",
  51671=>"000100011",
  51672=>"111001100",
  51673=>"100000000",
  51674=>"000001110",
  51675=>"101111000",
  51676=>"001011000",
  51677=>"100110101",
  51678=>"010110100",
  51679=>"101001100",
  51680=>"011000001",
  51681=>"000011111",
  51682=>"000010010",
  51683=>"111110011",
  51684=>"001010011",
  51685=>"010010110",
  51686=>"110011100",
  51687=>"000110111",
  51688=>"101100010",
  51689=>"001101000",
  51690=>"100001001",
  51691=>"110011111",
  51692=>"010001011",
  51693=>"110110010",
  51694=>"000110011",
  51695=>"111110010",
  51696=>"111101100",
  51697=>"110011110",
  51698=>"110111001",
  51699=>"011011110",
  51700=>"101000010",
  51701=>"101000000",
  51702=>"011001110",
  51703=>"011100000",
  51704=>"011001100",
  51705=>"010001001",
  51706=>"111000010",
  51707=>"101110011",
  51708=>"010001011",
  51709=>"100101110",
  51710=>"110010101",
  51711=>"111011101",
  51712=>"111010000",
  51713=>"011100110",
  51714=>"001000110",
  51715=>"110111001",
  51716=>"111101101",
  51717=>"001001000",
  51718=>"111110000",
  51719=>"000000011",
  51720=>"110100001",
  51721=>"110001010",
  51722=>"111110010",
  51723=>"010101000",
  51724=>"100000100",
  51725=>"110111011",
  51726=>"000011110",
  51727=>"111111000",
  51728=>"100011001",
  51729=>"000011001",
  51730=>"001111100",
  51731=>"111111010",
  51732=>"101010011",
  51733=>"100100010",
  51734=>"110010111",
  51735=>"111010000",
  51736=>"000001101",
  51737=>"111101001",
  51738=>"100101000",
  51739=>"111101000",
  51740=>"100000011",
  51741=>"100001000",
  51742=>"101011111",
  51743=>"110100110",
  51744=>"000011100",
  51745=>"100100100",
  51746=>"001111000",
  51747=>"000111010",
  51748=>"111001010",
  51749=>"011011011",
  51750=>"011000001",
  51751=>"100001100",
  51752=>"101011101",
  51753=>"010110111",
  51754=>"111100011",
  51755=>"111110111",
  51756=>"111011001",
  51757=>"101000011",
  51758=>"010110101",
  51759=>"011001000",
  51760=>"011110010",
  51761=>"100111011",
  51762=>"100100000",
  51763=>"011001010",
  51764=>"000011100",
  51765=>"111000011",
  51766=>"000101111",
  51767=>"001111011",
  51768=>"101010101",
  51769=>"000101100",
  51770=>"100110110",
  51771=>"101000001",
  51772=>"001000101",
  51773=>"000100010",
  51774=>"110000101",
  51775=>"101111111",
  51776=>"111101100",
  51777=>"010101101",
  51778=>"000001000",
  51779=>"011111001",
  51780=>"001000001",
  51781=>"010011000",
  51782=>"000100001",
  51783=>"001011110",
  51784=>"100100100",
  51785=>"111101010",
  51786=>"010011110",
  51787=>"010101000",
  51788=>"001011100",
  51789=>"000010010",
  51790=>"011111010",
  51791=>"110010110",
  51792=>"101110011",
  51793=>"111101000",
  51794=>"101001000",
  51795=>"101111011",
  51796=>"111100111",
  51797=>"000001000",
  51798=>"000001000",
  51799=>"011001110",
  51800=>"011101010",
  51801=>"010001000",
  51802=>"100011011",
  51803=>"111100111",
  51804=>"101010101",
  51805=>"000000101",
  51806=>"001000001",
  51807=>"111101111",
  51808=>"010001101",
  51809=>"110110001",
  51810=>"100111010",
  51811=>"000011110",
  51812=>"100000001",
  51813=>"110110100",
  51814=>"101101010",
  51815=>"101000111",
  51816=>"011100000",
  51817=>"011000101",
  51818=>"100100100",
  51819=>"000101001",
  51820=>"101010011",
  51821=>"010110011",
  51822=>"001111101",
  51823=>"100010111",
  51824=>"011101110",
  51825=>"000100001",
  51826=>"111010011",
  51827=>"101101101",
  51828=>"100001000",
  51829=>"010001111",
  51830=>"100111010",
  51831=>"100010111",
  51832=>"000101111",
  51833=>"000000100",
  51834=>"000010111",
  51835=>"000111101",
  51836=>"011000101",
  51837=>"011101110",
  51838=>"110110000",
  51839=>"100110010",
  51840=>"011110011",
  51841=>"101010001",
  51842=>"111001111",
  51843=>"110000111",
  51844=>"011011010",
  51845=>"000101001",
  51846=>"011110010",
  51847=>"110110110",
  51848=>"101010101",
  51849=>"111100001",
  51850=>"111110111",
  51851=>"011011011",
  51852=>"011101000",
  51853=>"110011000",
  51854=>"000100001",
  51855=>"010000100",
  51856=>"111100110",
  51857=>"110011110",
  51858=>"101011111",
  51859=>"010111001",
  51860=>"100101100",
  51861=>"100110100",
  51862=>"010010001",
  51863=>"101011100",
  51864=>"001111111",
  51865=>"001100101",
  51866=>"110010101",
  51867=>"111110001",
  51868=>"000100111",
  51869=>"000001001",
  51870=>"111010010",
  51871=>"111111111",
  51872=>"111110110",
  51873=>"100010000",
  51874=>"111010011",
  51875=>"100001110",
  51876=>"110101010",
  51877=>"001011010",
  51878=>"000010111",
  51879=>"011100001",
  51880=>"101001011",
  51881=>"011001100",
  51882=>"000110011",
  51883=>"000001010",
  51884=>"001111101",
  51885=>"011110000",
  51886=>"000010010",
  51887=>"111010010",
  51888=>"100000011",
  51889=>"111011111",
  51890=>"000100000",
  51891=>"101000110",
  51892=>"101101001",
  51893=>"001101110",
  51894=>"011011111",
  51895=>"011111000",
  51896=>"111011101",
  51897=>"000000100",
  51898=>"010001000",
  51899=>"011000000",
  51900=>"111000010",
  51901=>"100100000",
  51902=>"101000010",
  51903=>"000111010",
  51904=>"001110111",
  51905=>"010111001",
  51906=>"101110101",
  51907=>"111100100",
  51908=>"000100011",
  51909=>"111111000",
  51910=>"011011111",
  51911=>"101110100",
  51912=>"110000001",
  51913=>"100010011",
  51914=>"100000011",
  51915=>"000111000",
  51916=>"001001010",
  51917=>"110000000",
  51918=>"111101100",
  51919=>"100001101",
  51920=>"000101101",
  51921=>"010001111",
  51922=>"111111110",
  51923=>"010101011",
  51924=>"010111000",
  51925=>"110100101",
  51926=>"101000100",
  51927=>"000010010",
  51928=>"010110101",
  51929=>"101101001",
  51930=>"011110101",
  51931=>"100111000",
  51932=>"011000110",
  51933=>"000010111",
  51934=>"101110111",
  51935=>"100111101",
  51936=>"100100001",
  51937=>"101001010",
  51938=>"110110100",
  51939=>"100000001",
  51940=>"110110001",
  51941=>"111001100",
  51942=>"111010010",
  51943=>"010001001",
  51944=>"101101000",
  51945=>"000001000",
  51946=>"011000001",
  51947=>"010110111",
  51948=>"000001110",
  51949=>"010100010",
  51950=>"101101101",
  51951=>"010100011",
  51952=>"101011101",
  51953=>"111001010",
  51954=>"110011111",
  51955=>"110111010",
  51956=>"110011010",
  51957=>"110111111",
  51958=>"100100011",
  51959=>"111010100",
  51960=>"001011110",
  51961=>"110001001",
  51962=>"000000101",
  51963=>"011000011",
  51964=>"000110100",
  51965=>"000011010",
  51966=>"111000001",
  51967=>"011010100",
  51968=>"100011110",
  51969=>"010111000",
  51970=>"110100011",
  51971=>"100100111",
  51972=>"100100011",
  51973=>"000010011",
  51974=>"111111111",
  51975=>"101100100",
  51976=>"001000010",
  51977=>"101001111",
  51978=>"010001111",
  51979=>"111110111",
  51980=>"110110101",
  51981=>"010001100",
  51982=>"011010000",
  51983=>"001101111",
  51984=>"010100010",
  51985=>"001001110",
  51986=>"001010110",
  51987=>"010111001",
  51988=>"000110111",
  51989=>"011011000",
  51990=>"011010101",
  51991=>"000010011",
  51992=>"101000010",
  51993=>"000000000",
  51994=>"000000100",
  51995=>"011010010",
  51996=>"100100001",
  51997=>"111101011",
  51998=>"000010011",
  51999=>"000100101",
  52000=>"000111110",
  52001=>"010001010",
  52002=>"100001101",
  52003=>"101000000",
  52004=>"011100101",
  52005=>"111001011",
  52006=>"111100110",
  52007=>"010111010",
  52008=>"110100101",
  52009=>"111111111",
  52010=>"101010010",
  52011=>"011010110",
  52012=>"011101100",
  52013=>"000010010",
  52014=>"101101000",
  52015=>"100110000",
  52016=>"001001011",
  52017=>"101001000",
  52018=>"001101100",
  52019=>"101011000",
  52020=>"011010101",
  52021=>"111110000",
  52022=>"000010000",
  52023=>"011000111",
  52024=>"010101000",
  52025=>"001110001",
  52026=>"000101011",
  52027=>"111001000",
  52028=>"110100110",
  52029=>"000111111",
  52030=>"110110111",
  52031=>"000111110",
  52032=>"011010100",
  52033=>"101010100",
  52034=>"100101101",
  52035=>"100111100",
  52036=>"010000110",
  52037=>"001000011",
  52038=>"011110010",
  52039=>"110111010",
  52040=>"111000100",
  52041=>"110110001",
  52042=>"101100010",
  52043=>"000011010",
  52044=>"011011100",
  52045=>"111111101",
  52046=>"101100011",
  52047=>"001011101",
  52048=>"010110010",
  52049=>"011010010",
  52050=>"010000001",
  52051=>"011101000",
  52052=>"011101000",
  52053=>"110000110",
  52054=>"110001000",
  52055=>"100001101",
  52056=>"111000111",
  52057=>"110010000",
  52058=>"010111110",
  52059=>"110011110",
  52060=>"001101100",
  52061=>"111000110",
  52062=>"010001010",
  52063=>"000001110",
  52064=>"000000101",
  52065=>"011000000",
  52066=>"000110010",
  52067=>"100101010",
  52068=>"111100001",
  52069=>"101001000",
  52070=>"100001100",
  52071=>"011101101",
  52072=>"100100001",
  52073=>"110111111",
  52074=>"001111000",
  52075=>"000001011",
  52076=>"101110101",
  52077=>"110001011",
  52078=>"101100010",
  52079=>"110011101",
  52080=>"010011100",
  52081=>"111001000",
  52082=>"001111100",
  52083=>"010000010",
  52084=>"010011100",
  52085=>"100010000",
  52086=>"100001100",
  52087=>"011001011",
  52088=>"011100011",
  52089=>"010011011",
  52090=>"000111111",
  52091=>"110111100",
  52092=>"101111000",
  52093=>"100111010",
  52094=>"011101101",
  52095=>"110101101",
  52096=>"101011010",
  52097=>"011101011",
  52098=>"010001100",
  52099=>"000110010",
  52100=>"000110111",
  52101=>"001110100",
  52102=>"111111011",
  52103=>"111011010",
  52104=>"000000000",
  52105=>"000011111",
  52106=>"011101001",
  52107=>"110000010",
  52108=>"101111011",
  52109=>"100000000",
  52110=>"000101000",
  52111=>"001010110",
  52112=>"000010001",
  52113=>"011110111",
  52114=>"111100000",
  52115=>"110010110",
  52116=>"110100101",
  52117=>"001100110",
  52118=>"110000011",
  52119=>"100100110",
  52120=>"011010110",
  52121=>"100101001",
  52122=>"000010100",
  52123=>"100001101",
  52124=>"110000001",
  52125=>"101100010",
  52126=>"011101001",
  52127=>"110111010",
  52128=>"001000111",
  52129=>"010001110",
  52130=>"010111011",
  52131=>"011001001",
  52132=>"011100001",
  52133=>"011011011",
  52134=>"011010100",
  52135=>"111111011",
  52136=>"111000000",
  52137=>"000111011",
  52138=>"010101010",
  52139=>"000100110",
  52140=>"000000111",
  52141=>"001100001",
  52142=>"111011001",
  52143=>"110111001",
  52144=>"001010111",
  52145=>"001101011",
  52146=>"111000011",
  52147=>"011110011",
  52148=>"010010010",
  52149=>"011110001",
  52150=>"111110100",
  52151=>"110111011",
  52152=>"011100110",
  52153=>"010101010",
  52154=>"111101101",
  52155=>"110110011",
  52156=>"100100000",
  52157=>"100011110",
  52158=>"111000110",
  52159=>"011110010",
  52160=>"010111010",
  52161=>"011000100",
  52162=>"000000001",
  52163=>"001110100",
  52164=>"001100110",
  52165=>"110100101",
  52166=>"101100011",
  52167=>"101110111",
  52168=>"001001011",
  52169=>"010111000",
  52170=>"011011000",
  52171=>"100011011",
  52172=>"011000011",
  52173=>"100101110",
  52174=>"000110100",
  52175=>"110110011",
  52176=>"100001111",
  52177=>"011100110",
  52178=>"010100001",
  52179=>"001100000",
  52180=>"000111001",
  52181=>"101001100",
  52182=>"100011001",
  52183=>"010010011",
  52184=>"010000101",
  52185=>"101100011",
  52186=>"100101100",
  52187=>"010011001",
  52188=>"100010011",
  52189=>"010011001",
  52190=>"100000001",
  52191=>"010110111",
  52192=>"111010010",
  52193=>"110001110",
  52194=>"101111100",
  52195=>"100111110",
  52196=>"010001000",
  52197=>"111101010",
  52198=>"010010110",
  52199=>"000100101",
  52200=>"101100110",
  52201=>"000000111",
  52202=>"001111101",
  52203=>"000000001",
  52204=>"000110001",
  52205=>"000001000",
  52206=>"101111000",
  52207=>"101110111",
  52208=>"001010000",
  52209=>"101101100",
  52210=>"000101011",
  52211=>"010000101",
  52212=>"111100100",
  52213=>"100010100",
  52214=>"000011011",
  52215=>"110010101",
  52216=>"101010110",
  52217=>"111000101",
  52218=>"001110000",
  52219=>"111001110",
  52220=>"000000100",
  52221=>"010111110",
  52222=>"011101010",
  52223=>"101011100",
  52224=>"101000000",
  52225=>"110001000",
  52226=>"011101010",
  52227=>"001001100",
  52228=>"110010000",
  52229=>"011010001",
  52230=>"101110010",
  52231=>"001000000",
  52232=>"100101111",
  52233=>"100111010",
  52234=>"000100011",
  52235=>"101100000",
  52236=>"010110000",
  52237=>"011111101",
  52238=>"010101101",
  52239=>"100001101",
  52240=>"010011001",
  52241=>"010011110",
  52242=>"001000011",
  52243=>"010111100",
  52244=>"101101010",
  52245=>"000101110",
  52246=>"110110011",
  52247=>"100010000",
  52248=>"111000001",
  52249=>"010110110",
  52250=>"101101010",
  52251=>"011010011",
  52252=>"101010111",
  52253=>"110101000",
  52254=>"000110101",
  52255=>"101000111",
  52256=>"000011110",
  52257=>"001100101",
  52258=>"101000010",
  52259=>"010010100",
  52260=>"111101100",
  52261=>"100000010",
  52262=>"100011001",
  52263=>"010000001",
  52264=>"011110000",
  52265=>"000111100",
  52266=>"100110010",
  52267=>"001101010",
  52268=>"110001111",
  52269=>"011110101",
  52270=>"111011000",
  52271=>"101011101",
  52272=>"111001010",
  52273=>"111111011",
  52274=>"110010110",
  52275=>"110110101",
  52276=>"100000010",
  52277=>"100001010",
  52278=>"110100001",
  52279=>"111000110",
  52280=>"011010100",
  52281=>"111000001",
  52282=>"001000011",
  52283=>"001110100",
  52284=>"001111010",
  52285=>"110110010",
  52286=>"111100111",
  52287=>"000110110",
  52288=>"000010101",
  52289=>"001100101",
  52290=>"110101110",
  52291=>"000000100",
  52292=>"110101001",
  52293=>"110010000",
  52294=>"111010011",
  52295=>"101101110",
  52296=>"000010011",
  52297=>"100111110",
  52298=>"101011000",
  52299=>"011000101",
  52300=>"111111001",
  52301=>"111011100",
  52302=>"111111101",
  52303=>"100101000",
  52304=>"000100100",
  52305=>"010110110",
  52306=>"001111000",
  52307=>"110010110",
  52308=>"001001100",
  52309=>"111101000",
  52310=>"001001011",
  52311=>"000101000",
  52312=>"010000101",
  52313=>"100001001",
  52314=>"110100100",
  52315=>"001010101",
  52316=>"001110001",
  52317=>"100101101",
  52318=>"111010001",
  52319=>"101111011",
  52320=>"111000010",
  52321=>"101100110",
  52322=>"100001000",
  52323=>"011101100",
  52324=>"001000110",
  52325=>"001000110",
  52326=>"011000100",
  52327=>"111100101",
  52328=>"000101111",
  52329=>"100010110",
  52330=>"110010000",
  52331=>"010100001",
  52332=>"100001000",
  52333=>"010011101",
  52334=>"101101001",
  52335=>"101100001",
  52336=>"101110100",
  52337=>"101000111",
  52338=>"111001001",
  52339=>"100000010",
  52340=>"110111111",
  52341=>"111011010",
  52342=>"100101101",
  52343=>"011110100",
  52344=>"011011110",
  52345=>"100100111",
  52346=>"011000110",
  52347=>"000010011",
  52348=>"111001101",
  52349=>"101011011",
  52350=>"100100000",
  52351=>"110011110",
  52352=>"101101011",
  52353=>"000101000",
  52354=>"001010000",
  52355=>"011110100",
  52356=>"000100101",
  52357=>"100011101",
  52358=>"011001010",
  52359=>"001110000",
  52360=>"100010110",
  52361=>"111101011",
  52362=>"101010001",
  52363=>"011100100",
  52364=>"001011001",
  52365=>"001010010",
  52366=>"111000001",
  52367=>"000000011",
  52368=>"000100101",
  52369=>"011011101",
  52370=>"111101110",
  52371=>"001000000",
  52372=>"001001010",
  52373=>"100111011",
  52374=>"100100111",
  52375=>"010100100",
  52376=>"001100000",
  52377=>"110101000",
  52378=>"111101111",
  52379=>"101010111",
  52380=>"001111101",
  52381=>"010100110",
  52382=>"001100100",
  52383=>"000101101",
  52384=>"101000110",
  52385=>"001100100",
  52386=>"000000101",
  52387=>"000110100",
  52388=>"010101010",
  52389=>"001100111",
  52390=>"000111110",
  52391=>"111010100",
  52392=>"110101111",
  52393=>"100011010",
  52394=>"000101011",
  52395=>"101010000",
  52396=>"111011110",
  52397=>"001111100",
  52398=>"001010101",
  52399=>"100001010",
  52400=>"101111010",
  52401=>"000101101",
  52402=>"111010000",
  52403=>"001110110",
  52404=>"101100110",
  52405=>"011100100",
  52406=>"100111101",
  52407=>"000000101",
  52408=>"101110010",
  52409=>"001010001",
  52410=>"101001100",
  52411=>"001100011",
  52412=>"110001100",
  52413=>"101100011",
  52414=>"010100010",
  52415=>"001000001",
  52416=>"100100111",
  52417=>"101000001",
  52418=>"001101101",
  52419=>"010010000",
  52420=>"011100010",
  52421=>"101110010",
  52422=>"000101000",
  52423=>"001111110",
  52424=>"101011111",
  52425=>"011110010",
  52426=>"111000100",
  52427=>"011001001",
  52428=>"011100110",
  52429=>"101011000",
  52430=>"100111000",
  52431=>"010110011",
  52432=>"111111010",
  52433=>"001110101",
  52434=>"100011111",
  52435=>"110001110",
  52436=>"010100011",
  52437=>"110111100",
  52438=>"011000010",
  52439=>"011111100",
  52440=>"010000010",
  52441=>"110111110",
  52442=>"111010101",
  52443=>"101010011",
  52444=>"010101101",
  52445=>"111110111",
  52446=>"100001000",
  52447=>"111000111",
  52448=>"001110011",
  52449=>"100001110",
  52450=>"011100010",
  52451=>"100101101",
  52452=>"010001111",
  52453=>"000111000",
  52454=>"110110101",
  52455=>"010010100",
  52456=>"011100001",
  52457=>"010111110",
  52458=>"000111001",
  52459=>"000001000",
  52460=>"110111100",
  52461=>"010111110",
  52462=>"111101110",
  52463=>"100111010",
  52464=>"100010101",
  52465=>"011101001",
  52466=>"011011001",
  52467=>"000001000",
  52468=>"101110001",
  52469=>"011010111",
  52470=>"100000110",
  52471=>"111001110",
  52472=>"011111111",
  52473=>"110001110",
  52474=>"111001101",
  52475=>"101001101",
  52476=>"010101011",
  52477=>"000111110",
  52478=>"010100111",
  52479=>"010000010",
  52480=>"000110011",
  52481=>"101011110",
  52482=>"000011011",
  52483=>"001101101",
  52484=>"100101100",
  52485=>"011110100",
  52486=>"000010000",
  52487=>"001110010",
  52488=>"101010000",
  52489=>"000011000",
  52490=>"111011011",
  52491=>"000011100",
  52492=>"001001110",
  52493=>"101110000",
  52494=>"100010110",
  52495=>"010010001",
  52496=>"011111001",
  52497=>"111000011",
  52498=>"110101001",
  52499=>"101101010",
  52500=>"001101110",
  52501=>"111010000",
  52502=>"111011001",
  52503=>"011000110",
  52504=>"101101100",
  52505=>"010001011",
  52506=>"111110100",
  52507=>"100011111",
  52508=>"100000010",
  52509=>"010010000",
  52510=>"000111001",
  52511=>"100100010",
  52512=>"011101011",
  52513=>"000111001",
  52514=>"101000100",
  52515=>"010011011",
  52516=>"011101000",
  52517=>"100011100",
  52518=>"011100111",
  52519=>"101111000",
  52520=>"110000110",
  52521=>"000110011",
  52522=>"111101010",
  52523=>"100101100",
  52524=>"001010100",
  52525=>"011010101",
  52526=>"001101110",
  52527=>"111101111",
  52528=>"100000001",
  52529=>"101010110",
  52530=>"110110110",
  52531=>"101000100",
  52532=>"101111110",
  52533=>"000101110",
  52534=>"111011100",
  52535=>"010101100",
  52536=>"010001111",
  52537=>"010111011",
  52538=>"111100111",
  52539=>"001100110",
  52540=>"000111001",
  52541=>"110000010",
  52542=>"010100011",
  52543=>"111110011",
  52544=>"010111000",
  52545=>"110110010",
  52546=>"100111011",
  52547=>"111001010",
  52548=>"001010110",
  52549=>"101011001",
  52550=>"000110011",
  52551=>"100101111",
  52552=>"100100100",
  52553=>"001101000",
  52554=>"100000010",
  52555=>"000000000",
  52556=>"111100101",
  52557=>"111001001",
  52558=>"100000001",
  52559=>"101011110",
  52560=>"010101110",
  52561=>"001111001",
  52562=>"010000010",
  52563=>"111000000",
  52564=>"001111001",
  52565=>"100110111",
  52566=>"011010001",
  52567=>"101111000",
  52568=>"010011111",
  52569=>"011111100",
  52570=>"001000101",
  52571=>"000100111",
  52572=>"111010110",
  52573=>"000110011",
  52574=>"101110101",
  52575=>"101111001",
  52576=>"000111110",
  52577=>"000110100",
  52578=>"010010110",
  52579=>"000011100",
  52580=>"010100100",
  52581=>"010000000",
  52582=>"100010101",
  52583=>"111001111",
  52584=>"111011111",
  52585=>"110010011",
  52586=>"000101001",
  52587=>"011111110",
  52588=>"111011010",
  52589=>"101010001",
  52590=>"001000100",
  52591=>"100011110",
  52592=>"000110101",
  52593=>"010101001",
  52594=>"110010011",
  52595=>"011110101",
  52596=>"010001111",
  52597=>"100110101",
  52598=>"011110101",
  52599=>"101111111",
  52600=>"100100100",
  52601=>"111000001",
  52602=>"011111101",
  52603=>"010100011",
  52604=>"100001111",
  52605=>"111110010",
  52606=>"100000010",
  52607=>"100111010",
  52608=>"101001111",
  52609=>"100101001",
  52610=>"011111110",
  52611=>"100100111",
  52612=>"011111101",
  52613=>"011011100",
  52614=>"010010010",
  52615=>"101001010",
  52616=>"110001000",
  52617=>"000000010",
  52618=>"100101111",
  52619=>"001011010",
  52620=>"101101011",
  52621=>"000001000",
  52622=>"101110010",
  52623=>"101111000",
  52624=>"111101010",
  52625=>"000000010",
  52626=>"000010001",
  52627=>"010000000",
  52628=>"111111000",
  52629=>"110001010",
  52630=>"011010001",
  52631=>"100011001",
  52632=>"110101101",
  52633=>"000110001",
  52634=>"111011111",
  52635=>"010101100",
  52636=>"101000110",
  52637=>"100100111",
  52638=>"100101100",
  52639=>"101111000",
  52640=>"011011110",
  52641=>"100000110",
  52642=>"110001111",
  52643=>"001000000",
  52644=>"110110101",
  52645=>"101000101",
  52646=>"000110100",
  52647=>"010110101",
  52648=>"000101001",
  52649=>"101010011",
  52650=>"000000111",
  52651=>"111110010",
  52652=>"100011010",
  52653=>"111010101",
  52654=>"110111101",
  52655=>"000110001",
  52656=>"101000000",
  52657=>"000100011",
  52658=>"101011111",
  52659=>"110111111",
  52660=>"010110111",
  52661=>"100001011",
  52662=>"010010011",
  52663=>"000110001",
  52664=>"100001110",
  52665=>"111011111",
  52666=>"101000101",
  52667=>"100110101",
  52668=>"110101111",
  52669=>"001111100",
  52670=>"010110100",
  52671=>"000010011",
  52672=>"001000011",
  52673=>"010000011",
  52674=>"110101000",
  52675=>"111110100",
  52676=>"100101101",
  52677=>"110110110",
  52678=>"010101111",
  52679=>"101000111",
  52680=>"001111010",
  52681=>"001011111",
  52682=>"110001011",
  52683=>"010101010",
  52684=>"000001000",
  52685=>"101000011",
  52686=>"010000110",
  52687=>"101101100",
  52688=>"001011000",
  52689=>"111000001",
  52690=>"000110110",
  52691=>"001101011",
  52692=>"100011101",
  52693=>"101000011",
  52694=>"101111000",
  52695=>"010010010",
  52696=>"010101100",
  52697=>"011010010",
  52698=>"111000001",
  52699=>"101111111",
  52700=>"101010100",
  52701=>"010010100",
  52702=>"000111100",
  52703=>"011111111",
  52704=>"001111111",
  52705=>"011010101",
  52706=>"000101100",
  52707=>"010001000",
  52708=>"000001101",
  52709=>"101110011",
  52710=>"101011100",
  52711=>"010100010",
  52712=>"101001011",
  52713=>"000111101",
  52714=>"110111110",
  52715=>"111011011",
  52716=>"001111001",
  52717=>"101010000",
  52718=>"101101101",
  52719=>"000010001",
  52720=>"110101010",
  52721=>"111111111",
  52722=>"100111110",
  52723=>"011111100",
  52724=>"011100000",
  52725=>"101110001",
  52726=>"101011101",
  52727=>"001110101",
  52728=>"101001111",
  52729=>"011110011",
  52730=>"000000000",
  52731=>"010110110",
  52732=>"000110101",
  52733=>"110101010",
  52734=>"110100111",
  52735=>"010010110",
  52736=>"101001101",
  52737=>"101111101",
  52738=>"101100110",
  52739=>"001000010",
  52740=>"000000110",
  52741=>"111011100",
  52742=>"110001110",
  52743=>"011101001",
  52744=>"100011100",
  52745=>"111010001",
  52746=>"110101110",
  52747=>"010101000",
  52748=>"000110110",
  52749=>"000110110",
  52750=>"100011110",
  52751=>"001111001",
  52752=>"110110000",
  52753=>"111011010",
  52754=>"101001100",
  52755=>"001110010",
  52756=>"101010011",
  52757=>"000010001",
  52758=>"011000100",
  52759=>"000000000",
  52760=>"000110000",
  52761=>"100001011",
  52762=>"011110100",
  52763=>"001011011",
  52764=>"011000011",
  52765=>"000011001",
  52766=>"101000100",
  52767=>"101010000",
  52768=>"010010101",
  52769=>"010000000",
  52770=>"001010001",
  52771=>"001100000",
  52772=>"011000000",
  52773=>"101111001",
  52774=>"101010011",
  52775=>"010001101",
  52776=>"000011110",
  52777=>"001010000",
  52778=>"101111101",
  52779=>"010001000",
  52780=>"100010010",
  52781=>"111111100",
  52782=>"000010010",
  52783=>"001101110",
  52784=>"110110101",
  52785=>"001110101",
  52786=>"011000110",
  52787=>"111001001",
  52788=>"011011111",
  52789=>"110111110",
  52790=>"111110111",
  52791=>"011100000",
  52792=>"111010001",
  52793=>"001111010",
  52794=>"101011001",
  52795=>"111101111",
  52796=>"111101010",
  52797=>"011001110",
  52798=>"010000100",
  52799=>"111011111",
  52800=>"101000001",
  52801=>"001011110",
  52802=>"000000000",
  52803=>"101111001",
  52804=>"100101100",
  52805=>"001000110",
  52806=>"011011101",
  52807=>"100001111",
  52808=>"000011001",
  52809=>"001100000",
  52810=>"110001111",
  52811=>"111011101",
  52812=>"001001111",
  52813=>"000000111",
  52814=>"000001111",
  52815=>"111001100",
  52816=>"010000100",
  52817=>"111001101",
  52818=>"011011111",
  52819=>"111101110",
  52820=>"000100111",
  52821=>"001111100",
  52822=>"010111101",
  52823=>"101100000",
  52824=>"110010100",
  52825=>"110100101",
  52826=>"010111010",
  52827=>"101001001",
  52828=>"000111010",
  52829=>"000000111",
  52830=>"101011111",
  52831=>"010110100",
  52832=>"101110110",
  52833=>"101111010",
  52834=>"010010001",
  52835=>"111111001",
  52836=>"101111011",
  52837=>"001100110",
  52838=>"000110011",
  52839=>"100000010",
  52840=>"001001110",
  52841=>"010011111",
  52842=>"100000011",
  52843=>"101101100",
  52844=>"000111011",
  52845=>"100011101",
  52846=>"011100111",
  52847=>"101110101",
  52848=>"110000111",
  52849=>"110111100",
  52850=>"110000101",
  52851=>"011110100",
  52852=>"010001010",
  52853=>"100010000",
  52854=>"101110001",
  52855=>"001101000",
  52856=>"100100001",
  52857=>"011101011",
  52858=>"011011110",
  52859=>"110110101",
  52860=>"000111001",
  52861=>"101110110",
  52862=>"111101110",
  52863=>"011011010",
  52864=>"011010101",
  52865=>"001011101",
  52866=>"111100101",
  52867=>"001010000",
  52868=>"001001100",
  52869=>"000010110",
  52870=>"111111011",
  52871=>"111101010",
  52872=>"010111111",
  52873=>"000001111",
  52874=>"101111111",
  52875=>"000000100",
  52876=>"101010010",
  52877=>"010000111",
  52878=>"000110100",
  52879=>"000010011",
  52880=>"000111110",
  52881=>"111010001",
  52882=>"100111110",
  52883=>"010001110",
  52884=>"001100100",
  52885=>"111101010",
  52886=>"110101000",
  52887=>"111100110",
  52888=>"001000100",
  52889=>"000010010",
  52890=>"010101100",
  52891=>"101000100",
  52892=>"010000110",
  52893=>"101110100",
  52894=>"100111100",
  52895=>"101001111",
  52896=>"000011100",
  52897=>"001001111",
  52898=>"011100010",
  52899=>"101101000",
  52900=>"111100010",
  52901=>"000111100",
  52902=>"111111110",
  52903=>"011101110",
  52904=>"101100100",
  52905=>"001011010",
  52906=>"000111101",
  52907=>"101010000",
  52908=>"100110101",
  52909=>"011011000",
  52910=>"001011001",
  52911=>"010001001",
  52912=>"010001111",
  52913=>"000111101",
  52914=>"101010011",
  52915=>"000110100",
  52916=>"110111001",
  52917=>"101000011",
  52918=>"101000101",
  52919=>"101011110",
  52920=>"011111110",
  52921=>"110010011",
  52922=>"000101111",
  52923=>"000100101",
  52924=>"001111100",
  52925=>"001100001",
  52926=>"100011110",
  52927=>"101111110",
  52928=>"111111100",
  52929=>"101101111",
  52930=>"000101101",
  52931=>"001110100",
  52932=>"111110100",
  52933=>"001010100",
  52934=>"101001000",
  52935=>"011101101",
  52936=>"010000000",
  52937=>"101011000",
  52938=>"100010100",
  52939=>"110000001",
  52940=>"111110100",
  52941=>"000001101",
  52942=>"100000001",
  52943=>"111010100",
  52944=>"000001011",
  52945=>"000110010",
  52946=>"001001000",
  52947=>"101100101",
  52948=>"010110110",
  52949=>"000111101",
  52950=>"111001100",
  52951=>"010011011",
  52952=>"100001010",
  52953=>"011000101",
  52954=>"110101010",
  52955=>"000101001",
  52956=>"111100101",
  52957=>"000110010",
  52958=>"110000010",
  52959=>"111111101",
  52960=>"011001001",
  52961=>"101011011",
  52962=>"111111100",
  52963=>"001001101",
  52964=>"111111011",
  52965=>"011100000",
  52966=>"100000111",
  52967=>"101000001",
  52968=>"101000101",
  52969=>"011001110",
  52970=>"110111001",
  52971=>"111101001",
  52972=>"110011110",
  52973=>"111001110",
  52974=>"000011001",
  52975=>"001010000",
  52976=>"000001000",
  52977=>"111110011",
  52978=>"110101111",
  52979=>"001001111",
  52980=>"010011011",
  52981=>"011011000",
  52982=>"010110000",
  52983=>"111001010",
  52984=>"000011011",
  52985=>"001101001",
  52986=>"001111101",
  52987=>"010001110",
  52988=>"010000111",
  52989=>"101110101",
  52990=>"010000111",
  52991=>"000010010",
  52992=>"111001011",
  52993=>"001001110",
  52994=>"100101100",
  52995=>"100001000",
  52996=>"011110011",
  52997=>"000001111",
  52998=>"110001011",
  52999=>"011010000",
  53000=>"011000111",
  53001=>"000101110",
  53002=>"011111101",
  53003=>"001001001",
  53004=>"111010110",
  53005=>"101111111",
  53006=>"111011110",
  53007=>"010010000",
  53008=>"011000100",
  53009=>"000011111",
  53010=>"110000111",
  53011=>"001111101",
  53012=>"010000100",
  53013=>"001000101",
  53014=>"100101010",
  53015=>"100110001",
  53016=>"110110010",
  53017=>"101101110",
  53018=>"110111010",
  53019=>"111000011",
  53020=>"101000110",
  53021=>"111101111",
  53022=>"000100010",
  53023=>"000000111",
  53024=>"101001111",
  53025=>"100011110",
  53026=>"101111011",
  53027=>"100001001",
  53028=>"100101011",
  53029=>"001000111",
  53030=>"100000011",
  53031=>"101000110",
  53032=>"101000010",
  53033=>"010110101",
  53034=>"001111101",
  53035=>"001111100",
  53036=>"100001010",
  53037=>"001110011",
  53038=>"010110101",
  53039=>"011010110",
  53040=>"100001111",
  53041=>"100101011",
  53042=>"000010011",
  53043=>"001011011",
  53044=>"111001101",
  53045=>"101000010",
  53046=>"011011100",
  53047=>"100010001",
  53048=>"011101110",
  53049=>"111101001",
  53050=>"000101110",
  53051=>"001000111",
  53052=>"100010011",
  53053=>"000100100",
  53054=>"110000100",
  53055=>"000110000",
  53056=>"000100101",
  53057=>"011111110",
  53058=>"001101101",
  53059=>"001000101",
  53060=>"101111100",
  53061=>"001110000",
  53062=>"011111100",
  53063=>"010111000",
  53064=>"000011010",
  53065=>"111000100",
  53066=>"100101111",
  53067=>"000100011",
  53068=>"000110001",
  53069=>"111110110",
  53070=>"110000001",
  53071=>"110010100",
  53072=>"010100111",
  53073=>"100110111",
  53074=>"001110000",
  53075=>"001100101",
  53076=>"010101000",
  53077=>"001011001",
  53078=>"101111000",
  53079=>"100000011",
  53080=>"010111111",
  53081=>"010100000",
  53082=>"111101010",
  53083=>"110010000",
  53084=>"101111001",
  53085=>"111110111",
  53086=>"110101100",
  53087=>"110010011",
  53088=>"110101111",
  53089=>"010100000",
  53090=>"100010100",
  53091=>"111011000",
  53092=>"011111010",
  53093=>"000010110",
  53094=>"001110101",
  53095=>"111011001",
  53096=>"000010010",
  53097=>"110011101",
  53098=>"111100011",
  53099=>"100000101",
  53100=>"011000100",
  53101=>"011110001",
  53102=>"010001011",
  53103=>"110111001",
  53104=>"110110011",
  53105=>"110001111",
  53106=>"101000001",
  53107=>"111101101",
  53108=>"101111010",
  53109=>"100000101",
  53110=>"111111111",
  53111=>"001100100",
  53112=>"101101001",
  53113=>"100000001",
  53114=>"110001000",
  53115=>"011011111",
  53116=>"000000100",
  53117=>"111111001",
  53118=>"001001100",
  53119=>"111110001",
  53120=>"010110011",
  53121=>"100101100",
  53122=>"000100011",
  53123=>"001101110",
  53124=>"000000010",
  53125=>"111010010",
  53126=>"100000001",
  53127=>"101000100",
  53128=>"110001011",
  53129=>"000001110",
  53130=>"010110010",
  53131=>"001100111",
  53132=>"110001101",
  53133=>"110110111",
  53134=>"111000000",
  53135=>"011000110",
  53136=>"000010001",
  53137=>"010010101",
  53138=>"001101010",
  53139=>"011110011",
  53140=>"000011111",
  53141=>"111111010",
  53142=>"110101001",
  53143=>"100101110",
  53144=>"000010100",
  53145=>"100000001",
  53146=>"001011100",
  53147=>"011100000",
  53148=>"000110111",
  53149=>"010100110",
  53150=>"100010010",
  53151=>"011010100",
  53152=>"111011011",
  53153=>"110000010",
  53154=>"111011100",
  53155=>"111001101",
  53156=>"010110011",
  53157=>"100010110",
  53158=>"110000101",
  53159=>"111010111",
  53160=>"001111000",
  53161=>"001111101",
  53162=>"100010010",
  53163=>"111010110",
  53164=>"010100110",
  53165=>"010010001",
  53166=>"001111101",
  53167=>"110100100",
  53168=>"010010001",
  53169=>"100011000",
  53170=>"011110101",
  53171=>"101010010",
  53172=>"100011000",
  53173=>"011101110",
  53174=>"001100011",
  53175=>"001110111",
  53176=>"000110000",
  53177=>"011101111",
  53178=>"111101100",
  53179=>"110100000",
  53180=>"010110110",
  53181=>"001011110",
  53182=>"110101101",
  53183=>"001010010",
  53184=>"001111111",
  53185=>"000111000",
  53186=>"101101111",
  53187=>"111000010",
  53188=>"000110000",
  53189=>"011001111",
  53190=>"000100110",
  53191=>"111110111",
  53192=>"101100011",
  53193=>"010100011",
  53194=>"010001001",
  53195=>"000101101",
  53196=>"011110011",
  53197=>"101000000",
  53198=>"010000101",
  53199=>"011001001",
  53200=>"110000111",
  53201=>"000011010",
  53202=>"110111000",
  53203=>"000011110",
  53204=>"010110100",
  53205=>"111001011",
  53206=>"011011110",
  53207=>"000110101",
  53208=>"000000100",
  53209=>"000001101",
  53210=>"100001010",
  53211=>"111111110",
  53212=>"011101100",
  53213=>"101110101",
  53214=>"010101011",
  53215=>"010110000",
  53216=>"000011101",
  53217=>"101011111",
  53218=>"111011100",
  53219=>"101111100",
  53220=>"010110110",
  53221=>"101110111",
  53222=>"001000000",
  53223=>"110010001",
  53224=>"001010011",
  53225=>"001110100",
  53226=>"001010100",
  53227=>"111111111",
  53228=>"100111001",
  53229=>"101001001",
  53230=>"011010010",
  53231=>"101011111",
  53232=>"000001101",
  53233=>"000110101",
  53234=>"010000000",
  53235=>"101011111",
  53236=>"000011011",
  53237=>"000001111",
  53238=>"111001110",
  53239=>"110111010",
  53240=>"001100011",
  53241=>"100110101",
  53242=>"111110010",
  53243=>"110100101",
  53244=>"000111001",
  53245=>"101011111",
  53246=>"010110110",
  53247=>"100110000",
  53248=>"111000110",
  53249=>"010110001",
  53250=>"010010100",
  53251=>"011100001",
  53252=>"000101101",
  53253=>"100110110",
  53254=>"010010000",
  53255=>"010000000",
  53256=>"010011000",
  53257=>"110100011",
  53258=>"010100001",
  53259=>"111101000",
  53260=>"111011101",
  53261=>"001011100",
  53262=>"010010110",
  53263=>"111010111",
  53264=>"100110000",
  53265=>"001011110",
  53266=>"101000100",
  53267=>"100110010",
  53268=>"110000101",
  53269=>"000011101",
  53270=>"011010110",
  53271=>"100100000",
  53272=>"111111111",
  53273=>"011101101",
  53274=>"110110010",
  53275=>"110001011",
  53276=>"101110100",
  53277=>"001111100",
  53278=>"011010111",
  53279=>"011010001",
  53280=>"100010010",
  53281=>"111011000",
  53282=>"010000011",
  53283=>"010001111",
  53284=>"010110100",
  53285=>"000110101",
  53286=>"110110001",
  53287=>"000101011",
  53288=>"101101010",
  53289=>"111100110",
  53290=>"111011111",
  53291=>"001111010",
  53292=>"100111011",
  53293=>"111000110",
  53294=>"000010000",
  53295=>"111011000",
  53296=>"100100001",
  53297=>"001111111",
  53298=>"010011011",
  53299=>"001110111",
  53300=>"000000011",
  53301=>"011111000",
  53302=>"000101001",
  53303=>"110111111",
  53304=>"110000000",
  53305=>"000100010",
  53306=>"101001011",
  53307=>"110100110",
  53308=>"100101000",
  53309=>"001101101",
  53310=>"011110011",
  53311=>"000100001",
  53312=>"100101100",
  53313=>"000010011",
  53314=>"000110100",
  53315=>"000100100",
  53316=>"010100101",
  53317=>"100111100",
  53318=>"101010111",
  53319=>"001111110",
  53320=>"100101111",
  53321=>"110011001",
  53322=>"010001111",
  53323=>"100110001",
  53324=>"001101000",
  53325=>"101011111",
  53326=>"010111101",
  53327=>"110111101",
  53328=>"001100111",
  53329=>"101111010",
  53330=>"101001010",
  53331=>"010101010",
  53332=>"010010000",
  53333=>"110001000",
  53334=>"101101011",
  53335=>"101101110",
  53336=>"111111110",
  53337=>"011000101",
  53338=>"101001010",
  53339=>"100110011",
  53340=>"111101101",
  53341=>"000100111",
  53342=>"110000110",
  53343=>"011000001",
  53344=>"010111110",
  53345=>"101010011",
  53346=>"101111111",
  53347=>"110110010",
  53348=>"011010100",
  53349=>"110000110",
  53350=>"001100110",
  53351=>"000001000",
  53352=>"111110100",
  53353=>"010111001",
  53354=>"111111000",
  53355=>"010100001",
  53356=>"000101011",
  53357=>"110101100",
  53358=>"100101100",
  53359=>"100100111",
  53360=>"011011100",
  53361=>"010000100",
  53362=>"100001011",
  53363=>"111001110",
  53364=>"001101111",
  53365=>"010010110",
  53366=>"010101011",
  53367=>"010000111",
  53368=>"001010000",
  53369=>"011101100",
  53370=>"111011111",
  53371=>"110110110",
  53372=>"000000001",
  53373=>"110111111",
  53374=>"100001101",
  53375=>"000101010",
  53376=>"110010111",
  53377=>"111010000",
  53378=>"000100001",
  53379=>"101110101",
  53380=>"000001101",
  53381=>"110011000",
  53382=>"111101111",
  53383=>"111110011",
  53384=>"011100010",
  53385=>"110111000",
  53386=>"111001100",
  53387=>"010100101",
  53388=>"011000010",
  53389=>"100100001",
  53390=>"000101000",
  53391=>"000101010",
  53392=>"101111010",
  53393=>"101101010",
  53394=>"111111110",
  53395=>"111111101",
  53396=>"110010001",
  53397=>"011001001",
  53398=>"010000010",
  53399=>"011110000",
  53400=>"111000100",
  53401=>"101000110",
  53402=>"011111111",
  53403=>"000011110",
  53404=>"110111010",
  53405=>"010110110",
  53406=>"111111101",
  53407=>"100000110",
  53408=>"111000000",
  53409=>"000001011",
  53410=>"111011011",
  53411=>"110100000",
  53412=>"111111110",
  53413=>"011011100",
  53414=>"110000011",
  53415=>"001010100",
  53416=>"100100100",
  53417=>"011000110",
  53418=>"000110110",
  53419=>"001000000",
  53420=>"110100001",
  53421=>"110000000",
  53422=>"011100001",
  53423=>"101111011",
  53424=>"001010010",
  53425=>"110000110",
  53426=>"001011101",
  53427=>"000010010",
  53428=>"101111011",
  53429=>"011001001",
  53430=>"101100111",
  53431=>"000011110",
  53432=>"011001111",
  53433=>"110010000",
  53434=>"010100001",
  53435=>"001111001",
  53436=>"100111100",
  53437=>"000000000",
  53438=>"010010100",
  53439=>"011101011",
  53440=>"001010111",
  53441=>"001101101",
  53442=>"001100001",
  53443=>"011011001",
  53444=>"000101101",
  53445=>"110001000",
  53446=>"111010101",
  53447=>"000100000",
  53448=>"101111111",
  53449=>"010101011",
  53450=>"001011010",
  53451=>"111111101",
  53452=>"011011000",
  53453=>"111000110",
  53454=>"100110111",
  53455=>"001001100",
  53456=>"100100100",
  53457=>"001101100",
  53458=>"110110001",
  53459=>"111100010",
  53460=>"001110000",
  53461=>"001100110",
  53462=>"010110000",
  53463=>"000111000",
  53464=>"101011101",
  53465=>"111110111",
  53466=>"111000001",
  53467=>"011000001",
  53468=>"110111001",
  53469=>"100001100",
  53470=>"000111101",
  53471=>"100100001",
  53472=>"001111110",
  53473=>"110100101",
  53474=>"010011011",
  53475=>"011100110",
  53476=>"110111000",
  53477=>"000001001",
  53478=>"111100101",
  53479=>"111110100",
  53480=>"100110011",
  53481=>"000110011",
  53482=>"101101010",
  53483=>"111110011",
  53484=>"111111111",
  53485=>"000101111",
  53486=>"000010010",
  53487=>"110010101",
  53488=>"111001100",
  53489=>"011101011",
  53490=>"100010011",
  53491=>"011001110",
  53492=>"100011101",
  53493=>"110100111",
  53494=>"011100101",
  53495=>"110101000",
  53496=>"000001111",
  53497=>"110011010",
  53498=>"111110000",
  53499=>"100101101",
  53500=>"011100110",
  53501=>"101001110",
  53502=>"111001101",
  53503=>"010000101",
  53504=>"100001001",
  53505=>"110101000",
  53506=>"001100011",
  53507=>"001100000",
  53508=>"100101001",
  53509=>"010110000",
  53510=>"110001011",
  53511=>"000011010",
  53512=>"010111101",
  53513=>"010100010",
  53514=>"111011101",
  53515=>"111110110",
  53516=>"111111111",
  53517=>"111100110",
  53518=>"110101011",
  53519=>"111110100",
  53520=>"001011010",
  53521=>"011001011",
  53522=>"001111111",
  53523=>"111101101",
  53524=>"001010001",
  53525=>"111111111",
  53526=>"000111111",
  53527=>"101111001",
  53528=>"100011100",
  53529=>"111101101",
  53530=>"100111010",
  53531=>"111010010",
  53532=>"011111000",
  53533=>"011111010",
  53534=>"110000111",
  53535=>"011010000",
  53536=>"010000100",
  53537=>"001100111",
  53538=>"101010100",
  53539=>"111110011",
  53540=>"101000100",
  53541=>"111100110",
  53542=>"110001000",
  53543=>"011100001",
  53544=>"001100111",
  53545=>"011001110",
  53546=>"000101110",
  53547=>"011101011",
  53548=>"101100011",
  53549=>"101110011",
  53550=>"011011001",
  53551=>"110101110",
  53552=>"101110110",
  53553=>"110101001",
  53554=>"010111011",
  53555=>"001001111",
  53556=>"101110101",
  53557=>"110011010",
  53558=>"101101101",
  53559=>"111001100",
  53560=>"000010000",
  53561=>"010001000",
  53562=>"001111010",
  53563=>"000000100",
  53564=>"010100011",
  53565=>"110110011",
  53566=>"000001110",
  53567=>"010111010",
  53568=>"010100001",
  53569=>"011101010",
  53570=>"001011001",
  53571=>"010010110",
  53572=>"011011111",
  53573=>"101000111",
  53574=>"000001011",
  53575=>"010100110",
  53576=>"000001000",
  53577=>"101111110",
  53578=>"110100100",
  53579=>"001110110",
  53580=>"100101010",
  53581=>"001011100",
  53582=>"100111100",
  53583=>"101110000",
  53584=>"111111101",
  53585=>"110111000",
  53586=>"101111111",
  53587=>"110110111",
  53588=>"001011010",
  53589=>"110001100",
  53590=>"011001100",
  53591=>"111101101",
  53592=>"010011110",
  53593=>"000101010",
  53594=>"111110001",
  53595=>"001001010",
  53596=>"010001110",
  53597=>"100111111",
  53598=>"000001010",
  53599=>"000001100",
  53600=>"001010001",
  53601=>"101101111",
  53602=>"101101111",
  53603=>"000000011",
  53604=>"000010000",
  53605=>"010100011",
  53606=>"100011101",
  53607=>"010000001",
  53608=>"110011100",
  53609=>"111100010",
  53610=>"010100000",
  53611=>"111010001",
  53612=>"011011000",
  53613=>"100111110",
  53614=>"011110000",
  53615=>"001000110",
  53616=>"111000001",
  53617=>"010011101",
  53618=>"011111100",
  53619=>"001011111",
  53620=>"001100100",
  53621=>"101000010",
  53622=>"000001010",
  53623=>"010110001",
  53624=>"110001111",
  53625=>"010011100",
  53626=>"000011000",
  53627=>"011111011",
  53628=>"011010110",
  53629=>"010101101",
  53630=>"010111111",
  53631=>"010001110",
  53632=>"101110011",
  53633=>"000110110",
  53634=>"111001101",
  53635=>"111011111",
  53636=>"110011111",
  53637=>"011101011",
  53638=>"000010101",
  53639=>"110100010",
  53640=>"000110101",
  53641=>"001001001",
  53642=>"001001110",
  53643=>"011110111",
  53644=>"011000101",
  53645=>"101110100",
  53646=>"111111100",
  53647=>"010100000",
  53648=>"110011001",
  53649=>"000101111",
  53650=>"000000000",
  53651=>"001001000",
  53652=>"100111100",
  53653=>"111100101",
  53654=>"011100010",
  53655=>"111110011",
  53656=>"011101111",
  53657=>"100111100",
  53658=>"101001011",
  53659=>"000101110",
  53660=>"111111100",
  53661=>"100101111",
  53662=>"011110011",
  53663=>"111100101",
  53664=>"011000101",
  53665=>"110001011",
  53666=>"001100101",
  53667=>"010100001",
  53668=>"110001110",
  53669=>"001010100",
  53670=>"110010110",
  53671=>"001011100",
  53672=>"111110111",
  53673=>"101100011",
  53674=>"110000100",
  53675=>"001011000",
  53676=>"110011011",
  53677=>"111011111",
  53678=>"010000010",
  53679=>"000100100",
  53680=>"011011110",
  53681=>"000001011",
  53682=>"100111000",
  53683=>"111101111",
  53684=>"001010000",
  53685=>"010011001",
  53686=>"011111010",
  53687=>"101111011",
  53688=>"101010100",
  53689=>"011000100",
  53690=>"111100000",
  53691=>"001010010",
  53692=>"101111110",
  53693=>"110010010",
  53694=>"010111111",
  53695=>"111000100",
  53696=>"100001101",
  53697=>"110010001",
  53698=>"010000011",
  53699=>"011100111",
  53700=>"110101011",
  53701=>"000001011",
  53702=>"110111100",
  53703=>"111001000",
  53704=>"000100111",
  53705=>"110001111",
  53706=>"100000110",
  53707=>"101000001",
  53708=>"110010011",
  53709=>"010101001",
  53710=>"000100001",
  53711=>"111000110",
  53712=>"011001111",
  53713=>"001100110",
  53714=>"010100011",
  53715=>"100110100",
  53716=>"010110110",
  53717=>"111111110",
  53718=>"101010010",
  53719=>"111110110",
  53720=>"101001001",
  53721=>"110100110",
  53722=>"000111100",
  53723=>"010011000",
  53724=>"110000001",
  53725=>"100000011",
  53726=>"011111100",
  53727=>"001110011",
  53728=>"000001001",
  53729=>"000000000",
  53730=>"110011101",
  53731=>"000011010",
  53732=>"101110001",
  53733=>"101100001",
  53734=>"100001000",
  53735=>"010100011",
  53736=>"001010100",
  53737=>"011001001",
  53738=>"110011010",
  53739=>"010001100",
  53740=>"110001100",
  53741=>"011011010",
  53742=>"011111011",
  53743=>"011011010",
  53744=>"010010111",
  53745=>"000101011",
  53746=>"111001000",
  53747=>"000001111",
  53748=>"101010100",
  53749=>"110000111",
  53750=>"011111101",
  53751=>"110111101",
  53752=>"111000010",
  53753=>"010101011",
  53754=>"011010100",
  53755=>"000110110",
  53756=>"000101101",
  53757=>"111010010",
  53758=>"101111010",
  53759=>"000000111",
  53760=>"110101011",
  53761=>"001011111",
  53762=>"010110111",
  53763=>"011100100",
  53764=>"110000101",
  53765=>"101110110",
  53766=>"100111010",
  53767=>"001100100",
  53768=>"001010101",
  53769=>"100011000",
  53770=>"111010100",
  53771=>"001001001",
  53772=>"110010010",
  53773=>"000011001",
  53774=>"010110000",
  53775=>"011011000",
  53776=>"000000110",
  53777=>"110101111",
  53778=>"111110110",
  53779=>"000001010",
  53780=>"111111111",
  53781=>"100000001",
  53782=>"001111100",
  53783=>"100101110",
  53784=>"010011101",
  53785=>"101110000",
  53786=>"100111111",
  53787=>"001110000",
  53788=>"110110000",
  53789=>"100001000",
  53790=>"010101000",
  53791=>"111101111",
  53792=>"001010100",
  53793=>"000100001",
  53794=>"110011111",
  53795=>"000111101",
  53796=>"110111010",
  53797=>"111000110",
  53798=>"011000101",
  53799=>"010101001",
  53800=>"000100111",
  53801=>"001010111",
  53802=>"001000001",
  53803=>"010111011",
  53804=>"100101110",
  53805=>"000010011",
  53806=>"101100100",
  53807=>"111000100",
  53808=>"111010000",
  53809=>"010010001",
  53810=>"101010001",
  53811=>"001111111",
  53812=>"011100111",
  53813=>"010110110",
  53814=>"110010010",
  53815=>"101101110",
  53816=>"111111110",
  53817=>"001000110",
  53818=>"111100101",
  53819=>"010111001",
  53820=>"100110111",
  53821=>"000111110",
  53822=>"100010100",
  53823=>"101000001",
  53824=>"110000010",
  53825=>"001010101",
  53826=>"001001000",
  53827=>"110011111",
  53828=>"101001111",
  53829=>"001111001",
  53830=>"010001010",
  53831=>"000000101",
  53832=>"100000000",
  53833=>"010111001",
  53834=>"111000000",
  53835=>"101000111",
  53836=>"101110010",
  53837=>"110100110",
  53838=>"101110101",
  53839=>"110110011",
  53840=>"010001100",
  53841=>"101001111",
  53842=>"011010011",
  53843=>"100000010",
  53844=>"001000000",
  53845=>"000001110",
  53846=>"010010111",
  53847=>"110111001",
  53848=>"000110011",
  53849=>"110010100",
  53850=>"001100010",
  53851=>"100001111",
  53852=>"001110000",
  53853=>"100100110",
  53854=>"000110111",
  53855=>"100000000",
  53856=>"111011101",
  53857=>"101111101",
  53858=>"010110001",
  53859=>"101000100",
  53860=>"101011011",
  53861=>"010100111",
  53862=>"000111111",
  53863=>"010100010",
  53864=>"000101001",
  53865=>"101001101",
  53866=>"001110001",
  53867=>"111111000",
  53868=>"100100111",
  53869=>"000100101",
  53870=>"111100011",
  53871=>"011010000",
  53872=>"111100101",
  53873=>"110001001",
  53874=>"000000010",
  53875=>"000110101",
  53876=>"001111100",
  53877=>"110001000",
  53878=>"101111011",
  53879=>"100100100",
  53880=>"011000000",
  53881=>"011011111",
  53882=>"110111110",
  53883=>"000010101",
  53884=>"010011001",
  53885=>"110110110",
  53886=>"101000111",
  53887=>"010101011",
  53888=>"011111100",
  53889=>"000011010",
  53890=>"000111101",
  53891=>"001101000",
  53892=>"001001010",
  53893=>"010001110",
  53894=>"001000001",
  53895=>"111010111",
  53896=>"000100110",
  53897=>"010010110",
  53898=>"001100101",
  53899=>"111100111",
  53900=>"000011100",
  53901=>"100000110",
  53902=>"111111101",
  53903=>"011110001",
  53904=>"010111111",
  53905=>"101000011",
  53906=>"101011011",
  53907=>"000001010",
  53908=>"110010000",
  53909=>"001110000",
  53910=>"011101000",
  53911=>"010010000",
  53912=>"101001001",
  53913=>"010001000",
  53914=>"000000111",
  53915=>"001000001",
  53916=>"101111100",
  53917=>"110111001",
  53918=>"101001001",
  53919=>"100000111",
  53920=>"100101001",
  53921=>"110000111",
  53922=>"101001000",
  53923=>"111100100",
  53924=>"111100111",
  53925=>"011111110",
  53926=>"101100010",
  53927=>"010010101",
  53928=>"000101000",
  53929=>"110101001",
  53930=>"111011010",
  53931=>"111011110",
  53932=>"110011010",
  53933=>"100101011",
  53934=>"001100001",
  53935=>"000000000",
  53936=>"000111101",
  53937=>"110011101",
  53938=>"110101001",
  53939=>"111100001",
  53940=>"001010110",
  53941=>"010110110",
  53942=>"010110110",
  53943=>"011100101",
  53944=>"011011100",
  53945=>"001101001",
  53946=>"110111111",
  53947=>"100101011",
  53948=>"100000111",
  53949=>"101011000",
  53950=>"000101110",
  53951=>"011010010",
  53952=>"110110101",
  53953=>"011101000",
  53954=>"111101111",
  53955=>"010110101",
  53956=>"111101011",
  53957=>"000011010",
  53958=>"111111101",
  53959=>"111011011",
  53960=>"001101111",
  53961=>"100000111",
  53962=>"100000011",
  53963=>"100100111",
  53964=>"111011111",
  53965=>"010101011",
  53966=>"000101001",
  53967=>"111101010",
  53968=>"011111010",
  53969=>"111100101",
  53970=>"101000011",
  53971=>"101101100",
  53972=>"000000110",
  53973=>"110001111",
  53974=>"011001100",
  53975=>"010001100",
  53976=>"101001110",
  53977=>"001011001",
  53978=>"100001001",
  53979=>"010011001",
  53980=>"110001111",
  53981=>"110110110",
  53982=>"000000011",
  53983=>"010111010",
  53984=>"011100110",
  53985=>"001011010",
  53986=>"000001101",
  53987=>"101110001",
  53988=>"101111100",
  53989=>"010100110",
  53990=>"111111001",
  53991=>"100000010",
  53992=>"001101110",
  53993=>"011010101",
  53994=>"110110101",
  53995=>"011100010",
  53996=>"101111110",
  53997=>"101100011",
  53998=>"000010100",
  53999=>"101000100",
  54000=>"001100111",
  54001=>"100101110",
  54002=>"100111110",
  54003=>"010100100",
  54004=>"010100001",
  54005=>"011010110",
  54006=>"111110010",
  54007=>"101100001",
  54008=>"111110001",
  54009=>"100111011",
  54010=>"110001100",
  54011=>"101011101",
  54012=>"111101011",
  54013=>"100011100",
  54014=>"110000011",
  54015=>"110001101",
  54016=>"111000010",
  54017=>"110001011",
  54018=>"101110111",
  54019=>"010001111",
  54020=>"101110111",
  54021=>"101011110",
  54022=>"000001010",
  54023=>"111110001",
  54024=>"101101001",
  54025=>"000001000",
  54026=>"000001000",
  54027=>"001001110",
  54028=>"101101100",
  54029=>"110100001",
  54030=>"111001100",
  54031=>"101111000",
  54032=>"001011110",
  54033=>"110001111",
  54034=>"100110111",
  54035=>"110100001",
  54036=>"110000010",
  54037=>"010000000",
  54038=>"111101101",
  54039=>"100101000",
  54040=>"010001000",
  54041=>"100010000",
  54042=>"000001001",
  54043=>"010100110",
  54044=>"100101001",
  54045=>"000110011",
  54046=>"001100011",
  54047=>"011001001",
  54048=>"111100001",
  54049=>"101111001",
  54050=>"101011010",
  54051=>"110110100",
  54052=>"101111000",
  54053=>"100100111",
  54054=>"111110001",
  54055=>"000000110",
  54056=>"101100111",
  54057=>"010100001",
  54058=>"001100010",
  54059=>"110100101",
  54060=>"010001111",
  54061=>"000000101",
  54062=>"000011110",
  54063=>"111001100",
  54064=>"110100100",
  54065=>"100001110",
  54066=>"111111110",
  54067=>"011000000",
  54068=>"110111100",
  54069=>"110001100",
  54070=>"111111101",
  54071=>"100110011",
  54072=>"110111100",
  54073=>"010110011",
  54074=>"010000101",
  54075=>"001001010",
  54076=>"011011100",
  54077=>"111101110",
  54078=>"010111101",
  54079=>"011110001",
  54080=>"011001100",
  54081=>"011000111",
  54082=>"110100110",
  54083=>"100111110",
  54084=>"000010000",
  54085=>"000111001",
  54086=>"011010100",
  54087=>"010011100",
  54088=>"101001000",
  54089=>"111011000",
  54090=>"011110000",
  54091=>"100110001",
  54092=>"011010000",
  54093=>"000001001",
  54094=>"100110110",
  54095=>"000001010",
  54096=>"101101111",
  54097=>"100110100",
  54098=>"001000001",
  54099=>"100011101",
  54100=>"001000011",
  54101=>"100100111",
  54102=>"110011100",
  54103=>"011001001",
  54104=>"011000101",
  54105=>"010010001",
  54106=>"101011000",
  54107=>"001001111",
  54108=>"110110111",
  54109=>"000100100",
  54110=>"100101000",
  54111=>"001010010",
  54112=>"001000000",
  54113=>"101111011",
  54114=>"001001011",
  54115=>"010101101",
  54116=>"110100010",
  54117=>"010011000",
  54118=>"001111001",
  54119=>"110111001",
  54120=>"010110100",
  54121=>"000011011",
  54122=>"011111110",
  54123=>"011100010",
  54124=>"111010111",
  54125=>"010110110",
  54126=>"110011011",
  54127=>"101110010",
  54128=>"001011111",
  54129=>"010101111",
  54130=>"110101001",
  54131=>"110101100",
  54132=>"000101000",
  54133=>"011111000",
  54134=>"110001010",
  54135=>"011011110",
  54136=>"000000011",
  54137=>"101110000",
  54138=>"000001111",
  54139=>"001111101",
  54140=>"101111011",
  54141=>"111000101",
  54142=>"011000111",
  54143=>"011011101",
  54144=>"110000111",
  54145=>"001111011",
  54146=>"011101100",
  54147=>"100110011",
  54148=>"010110100",
  54149=>"001011001",
  54150=>"111101011",
  54151=>"010100100",
  54152=>"010000001",
  54153=>"101010010",
  54154=>"001001100",
  54155=>"100000110",
  54156=>"110111001",
  54157=>"000010001",
  54158=>"001001000",
  54159=>"101110000",
  54160=>"100101011",
  54161=>"111100101",
  54162=>"110100011",
  54163=>"000011111",
  54164=>"010110011",
  54165=>"101010111",
  54166=>"110110110",
  54167=>"000010101",
  54168=>"111001111",
  54169=>"000111000",
  54170=>"100001010",
  54171=>"011100101",
  54172=>"100000100",
  54173=>"001101000",
  54174=>"010101011",
  54175=>"011001110",
  54176=>"100011110",
  54177=>"111111101",
  54178=>"100011010",
  54179=>"100000100",
  54180=>"010101010",
  54181=>"011101100",
  54182=>"100100100",
  54183=>"001111001",
  54184=>"101010001",
  54185=>"001110111",
  54186=>"010000001",
  54187=>"101000001",
  54188=>"110011001",
  54189=>"010010000",
  54190=>"011001011",
  54191=>"011010110",
  54192=>"000001111",
  54193=>"011101001",
  54194=>"001111110",
  54195=>"001001010",
  54196=>"110001010",
  54197=>"100001100",
  54198=>"000011000",
  54199=>"110101000",
  54200=>"010000111",
  54201=>"111001111",
  54202=>"101110101",
  54203=>"110110110",
  54204=>"010001111",
  54205=>"011101100",
  54206=>"001110001",
  54207=>"001100101",
  54208=>"101111011",
  54209=>"101001001",
  54210=>"000011101",
  54211=>"010111001",
  54212=>"000000111",
  54213=>"001001101",
  54214=>"101101000",
  54215=>"000001100",
  54216=>"001111011",
  54217=>"001100001",
  54218=>"100011101",
  54219=>"010000011",
  54220=>"111000011",
  54221=>"011010011",
  54222=>"010110100",
  54223=>"101011001",
  54224=>"001110110",
  54225=>"000001110",
  54226=>"010011001",
  54227=>"101111001",
  54228=>"101111001",
  54229=>"101000001",
  54230=>"010000000",
  54231=>"101011110",
  54232=>"010100001",
  54233=>"100101110",
  54234=>"010011111",
  54235=>"111110011",
  54236=>"000100110",
  54237=>"010011100",
  54238=>"100010111",
  54239=>"101000010",
  54240=>"111010000",
  54241=>"100011010",
  54242=>"000000011",
  54243=>"100001100",
  54244=>"101000101",
  54245=>"011000111",
  54246=>"100011101",
  54247=>"010010010",
  54248=>"001001111",
  54249=>"000101000",
  54250=>"000110010",
  54251=>"101100100",
  54252=>"000000101",
  54253=>"010110001",
  54254=>"100110111",
  54255=>"010001100",
  54256=>"100001001",
  54257=>"011011011",
  54258=>"101100010",
  54259=>"100100011",
  54260=>"000010001",
  54261=>"000101110",
  54262=>"010011111",
  54263=>"011000011",
  54264=>"000001011",
  54265=>"111110100",
  54266=>"110101011",
  54267=>"001011101",
  54268=>"101010110",
  54269=>"010100111",
  54270=>"100110001",
  54271=>"001001111",
  54272=>"010010111",
  54273=>"010111000",
  54274=>"011010111",
  54275=>"111000111",
  54276=>"101010111",
  54277=>"010011000",
  54278=>"100111010",
  54279=>"001010110",
  54280=>"000101110",
  54281=>"111001010",
  54282=>"000010011",
  54283=>"111110010",
  54284=>"110110100",
  54285=>"110011000",
  54286=>"101110100",
  54287=>"000001000",
  54288=>"011001101",
  54289=>"111110000",
  54290=>"110001010",
  54291=>"110001010",
  54292=>"000101100",
  54293=>"011001100",
  54294=>"011000011",
  54295=>"010010011",
  54296=>"011110011",
  54297=>"000010111",
  54298=>"100100110",
  54299=>"011010101",
  54300=>"011011010",
  54301=>"000000101",
  54302=>"110000100",
  54303=>"000100100",
  54304=>"110101001",
  54305=>"000001001",
  54306=>"110000110",
  54307=>"011000010",
  54308=>"101111111",
  54309=>"100100100",
  54310=>"110011001",
  54311=>"100000000",
  54312=>"001001000",
  54313=>"010011001",
  54314=>"101000111",
  54315=>"010010011",
  54316=>"011001001",
  54317=>"011110110",
  54318=>"111101110",
  54319=>"010110000",
  54320=>"001110011",
  54321=>"001001011",
  54322=>"000110110",
  54323=>"000111010",
  54324=>"100001001",
  54325=>"111101110",
  54326=>"011000010",
  54327=>"111111010",
  54328=>"000100100",
  54329=>"000001011",
  54330=>"010110001",
  54331=>"111011011",
  54332=>"000111100",
  54333=>"010010111",
  54334=>"100100000",
  54335=>"101001110",
  54336=>"100000111",
  54337=>"001010100",
  54338=>"000001010",
  54339=>"100011111",
  54340=>"100111000",
  54341=>"111100000",
  54342=>"111000100",
  54343=>"110000011",
  54344=>"001001101",
  54345=>"000001010",
  54346=>"101100100",
  54347=>"110001101",
  54348=>"101100110",
  54349=>"001010011",
  54350=>"011011011",
  54351=>"010111111",
  54352=>"101111111",
  54353=>"000100100",
  54354=>"010010111",
  54355=>"000100001",
  54356=>"011001101",
  54357=>"110111101",
  54358=>"010111011",
  54359=>"101001110",
  54360=>"100111111",
  54361=>"011011110",
  54362=>"010000111",
  54363=>"100100110",
  54364=>"000001001",
  54365=>"100000011",
  54366=>"000101000",
  54367=>"001000010",
  54368=>"011111010",
  54369=>"101001101",
  54370=>"110000101",
  54371=>"100000010",
  54372=>"011001010",
  54373=>"111100111",
  54374=>"100000010",
  54375=>"001001010",
  54376=>"000001010",
  54377=>"010111000",
  54378=>"000010100",
  54379=>"100100010",
  54380=>"000001111",
  54381=>"001110010",
  54382=>"010101100",
  54383=>"100110101",
  54384=>"101011011",
  54385=>"100110011",
  54386=>"000001111",
  54387=>"011110011",
  54388=>"000011111",
  54389=>"110101111",
  54390=>"101101100",
  54391=>"000010000",
  54392=>"011011001",
  54393=>"010100111",
  54394=>"001110110",
  54395=>"010000001",
  54396=>"010111010",
  54397=>"001011000",
  54398=>"110001000",
  54399=>"000101101",
  54400=>"111101001",
  54401=>"011111111",
  54402=>"100101010",
  54403=>"110101000",
  54404=>"111001010",
  54405=>"010001001",
  54406=>"011011100",
  54407=>"000000011",
  54408=>"101010001",
  54409=>"010010101",
  54410=>"011000100",
  54411=>"000101000",
  54412=>"111111110",
  54413=>"000010000",
  54414=>"001111000",
  54415=>"110011110",
  54416=>"011110010",
  54417=>"010011111",
  54418=>"100100011",
  54419=>"111110101",
  54420=>"110111001",
  54421=>"100100110",
  54422=>"111110010",
  54423=>"101100101",
  54424=>"100110000",
  54425=>"000100110",
  54426=>"001011101",
  54427=>"000000010",
  54428=>"111000010",
  54429=>"110110000",
  54430=>"001001001",
  54431=>"000100100",
  54432=>"011010110",
  54433=>"000001101",
  54434=>"111000000",
  54435=>"101000111",
  54436=>"001101011",
  54437=>"101100111",
  54438=>"111001100",
  54439=>"011011101",
  54440=>"001000110",
  54441=>"100001000",
  54442=>"001010110",
  54443=>"110010100",
  54444=>"110010000",
  54445=>"011010001",
  54446=>"001011001",
  54447=>"010010001",
  54448=>"111010101",
  54449=>"111110011",
  54450=>"111101100",
  54451=>"110101000",
  54452=>"100001010",
  54453=>"001110111",
  54454=>"111010111",
  54455=>"100101010",
  54456=>"010000010",
  54457=>"001001010",
  54458=>"100110111",
  54459=>"100100110",
  54460=>"010000001",
  54461=>"010000000",
  54462=>"101001110",
  54463=>"111010011",
  54464=>"100010101",
  54465=>"000100000",
  54466=>"000010001",
  54467=>"101101111",
  54468=>"101100000",
  54469=>"101011001",
  54470=>"001000000",
  54471=>"111111100",
  54472=>"110111010",
  54473=>"001110001",
  54474=>"000001111",
  54475=>"101111000",
  54476=>"111010101",
  54477=>"011010010",
  54478=>"001101100",
  54479=>"101101000",
  54480=>"001011000",
  54481=>"010111010",
  54482=>"010110000",
  54483=>"010101010",
  54484=>"011100001",
  54485=>"111110000",
  54486=>"111000011",
  54487=>"000001000",
  54488=>"000000011",
  54489=>"010100010",
  54490=>"001001010",
  54491=>"011001101",
  54492=>"001111000",
  54493=>"011101000",
  54494=>"001000001",
  54495=>"110111110",
  54496=>"000100010",
  54497=>"010000010",
  54498=>"111000101",
  54499=>"000001101",
  54500=>"111000110",
  54501=>"100001111",
  54502=>"001111010",
  54503=>"010111011",
  54504=>"101001101",
  54505=>"111011010",
  54506=>"010011111",
  54507=>"110101110",
  54508=>"001000010",
  54509=>"010111101",
  54510=>"100111110",
  54511=>"001100000",
  54512=>"111000010",
  54513=>"011110100",
  54514=>"000110100",
  54515=>"011000010",
  54516=>"010100001",
  54517=>"100000011",
  54518=>"011111000",
  54519=>"001101011",
  54520=>"001111101",
  54521=>"000111101",
  54522=>"101000101",
  54523=>"001001001",
  54524=>"101000111",
  54525=>"001101000",
  54526=>"111101000",
  54527=>"110100010",
  54528=>"100001111",
  54529=>"100100101",
  54530=>"000101110",
  54531=>"101010101",
  54532=>"010011010",
  54533=>"000100110",
  54534=>"111110111",
  54535=>"010010101",
  54536=>"101111110",
  54537=>"001100111",
  54538=>"111110100",
  54539=>"100110110",
  54540=>"101110010",
  54541=>"100111001",
  54542=>"111000001",
  54543=>"000001100",
  54544=>"111111001",
  54545=>"111111110",
  54546=>"101001110",
  54547=>"100101101",
  54548=>"101001110",
  54549=>"100011101",
  54550=>"010000101",
  54551=>"111000000",
  54552=>"101011110",
  54553=>"001010001",
  54554=>"111100111",
  54555=>"110000110",
  54556=>"100010010",
  54557=>"100001010",
  54558=>"001100000",
  54559=>"100000010",
  54560=>"110000110",
  54561=>"010001000",
  54562=>"110110100",
  54563=>"100000001",
  54564=>"111011101",
  54565=>"010000001",
  54566=>"001110110",
  54567=>"000111111",
  54568=>"001101011",
  54569=>"011010010",
  54570=>"100100001",
  54571=>"011111111",
  54572=>"101111000",
  54573=>"101110111",
  54574=>"011011111",
  54575=>"100010100",
  54576=>"010101101",
  54577=>"110011110",
  54578=>"111010111",
  54579=>"111100011",
  54580=>"001111011",
  54581=>"011101110",
  54582=>"111100000",
  54583=>"011011101",
  54584=>"111011010",
  54585=>"100111100",
  54586=>"000101001",
  54587=>"101111000",
  54588=>"100000011",
  54589=>"010110110",
  54590=>"100000001",
  54591=>"111000110",
  54592=>"100100010",
  54593=>"011000010",
  54594=>"000011011",
  54595=>"010100000",
  54596=>"111111110",
  54597=>"100000010",
  54598=>"110001101",
  54599=>"111101010",
  54600=>"101000000",
  54601=>"000001000",
  54602=>"010100100",
  54603=>"010000010",
  54604=>"010101111",
  54605=>"100111111",
  54606=>"100010101",
  54607=>"101100011",
  54608=>"010000101",
  54609=>"100011100",
  54610=>"011100100",
  54611=>"000101111",
  54612=>"000110000",
  54613=>"100100001",
  54614=>"011010001",
  54615=>"000100110",
  54616=>"011001000",
  54617=>"110011001",
  54618=>"000010000",
  54619=>"100011110",
  54620=>"111000100",
  54621=>"110011001",
  54622=>"100100101",
  54623=>"111001011",
  54624=>"100101001",
  54625=>"011000010",
  54626=>"010001010",
  54627=>"100000101",
  54628=>"110001000",
  54629=>"010111100",
  54630=>"101101110",
  54631=>"011000000",
  54632=>"001000011",
  54633=>"000000001",
  54634=>"100101001",
  54635=>"000101110",
  54636=>"111001010",
  54637=>"000001110",
  54638=>"111000111",
  54639=>"001010001",
  54640=>"110001000",
  54641=>"110111000",
  54642=>"011000100",
  54643=>"110010011",
  54644=>"011000000",
  54645=>"000011001",
  54646=>"010011100",
  54647=>"010110101",
  54648=>"001011011",
  54649=>"001011000",
  54650=>"001101111",
  54651=>"111110111",
  54652=>"011111111",
  54653=>"001011110",
  54654=>"110101000",
  54655=>"010011100",
  54656=>"010010000",
  54657=>"001000011",
  54658=>"001000110",
  54659=>"011101101",
  54660=>"101010011",
  54661=>"000001010",
  54662=>"101100010",
  54663=>"000101000",
  54664=>"100110011",
  54665=>"100111110",
  54666=>"101100010",
  54667=>"000101111",
  54668=>"010011110",
  54669=>"000100010",
  54670=>"100101001",
  54671=>"001111010",
  54672=>"000110101",
  54673=>"010100001",
  54674=>"110111000",
  54675=>"110001001",
  54676=>"101001110",
  54677=>"010010000",
  54678=>"011111111",
  54679=>"111011000",
  54680=>"101111010",
  54681=>"101100101",
  54682=>"010110101",
  54683=>"100100101",
  54684=>"011101101",
  54685=>"111111111",
  54686=>"111100110",
  54687=>"001101001",
  54688=>"111110010",
  54689=>"111100101",
  54690=>"110100010",
  54691=>"100001000",
  54692=>"100001110",
  54693=>"110001001",
  54694=>"001100111",
  54695=>"011110110",
  54696=>"100110110",
  54697=>"101110101",
  54698=>"100001000",
  54699=>"110001111",
  54700=>"000001111",
  54701=>"010110101",
  54702=>"101011100",
  54703=>"011100101",
  54704=>"100000101",
  54705=>"000110100",
  54706=>"110111111",
  54707=>"110101111",
  54708=>"111011111",
  54709=>"101011011",
  54710=>"000001011",
  54711=>"110111011",
  54712=>"010101101",
  54713=>"010010000",
  54714=>"100000000",
  54715=>"011110011",
  54716=>"101111111",
  54717=>"101110110",
  54718=>"000011011",
  54719=>"000111101",
  54720=>"000001000",
  54721=>"010100111",
  54722=>"110100010",
  54723=>"110001110",
  54724=>"000010010",
  54725=>"111001111",
  54726=>"010010101",
  54727=>"101111110",
  54728=>"100001010",
  54729=>"100010001",
  54730=>"010100011",
  54731=>"100001011",
  54732=>"011110111",
  54733=>"010000000",
  54734=>"101000001",
  54735=>"010001110",
  54736=>"100110100",
  54737=>"111000000",
  54738=>"011001000",
  54739=>"001010111",
  54740=>"010111111",
  54741=>"110000000",
  54742=>"011001001",
  54743=>"100100111",
  54744=>"101101011",
  54745=>"010111011",
  54746=>"101011110",
  54747=>"110001110",
  54748=>"100000110",
  54749=>"101011001",
  54750=>"000011000",
  54751=>"101010000",
  54752=>"100100100",
  54753=>"011011001",
  54754=>"010011010",
  54755=>"011000000",
  54756=>"111100100",
  54757=>"111010001",
  54758=>"000100010",
  54759=>"101110111",
  54760=>"000010000",
  54761=>"010011001",
  54762=>"111111110",
  54763=>"100101010",
  54764=>"010100001",
  54765=>"110000111",
  54766=>"001101110",
  54767=>"101011100",
  54768=>"110110000",
  54769=>"010001111",
  54770=>"010110100",
  54771=>"011111010",
  54772=>"010110000",
  54773=>"011101111",
  54774=>"101111000",
  54775=>"010011110",
  54776=>"111000000",
  54777=>"000101110",
  54778=>"001101101",
  54779=>"100011100",
  54780=>"010111001",
  54781=>"101011000",
  54782=>"111101000",
  54783=>"101100000",
  54784=>"000001110",
  54785=>"101010101",
  54786=>"111010101",
  54787=>"000011111",
  54788=>"101111101",
  54789=>"001111010",
  54790=>"111001100",
  54791=>"000011110",
  54792=>"001000111",
  54793=>"101000010",
  54794=>"101011011",
  54795=>"111101101",
  54796=>"001000100",
  54797=>"001100101",
  54798=>"000100000",
  54799=>"111111011",
  54800=>"110011001",
  54801=>"010011011",
  54802=>"010101110",
  54803=>"100001100",
  54804=>"001010000",
  54805=>"101010110",
  54806=>"000110100",
  54807=>"111001101",
  54808=>"010000111",
  54809=>"000001110",
  54810=>"111001001",
  54811=>"100011110",
  54812=>"111100010",
  54813=>"001001000",
  54814=>"111100111",
  54815=>"101111111",
  54816=>"111011111",
  54817=>"001101001",
  54818=>"101000011",
  54819=>"011010110",
  54820=>"100111110",
  54821=>"011001101",
  54822=>"110110001",
  54823=>"100010011",
  54824=>"000000011",
  54825=>"100001101",
  54826=>"101110001",
  54827=>"010111000",
  54828=>"001001011",
  54829=>"001110100",
  54830=>"000001100",
  54831=>"101111111",
  54832=>"100100011",
  54833=>"110100011",
  54834=>"111000101",
  54835=>"001001000",
  54836=>"010000001",
  54837=>"101100001",
  54838=>"111000001",
  54839=>"011001000",
  54840=>"111111001",
  54841=>"110111010",
  54842=>"101000001",
  54843=>"101101011",
  54844=>"010110111",
  54845=>"100001111",
  54846=>"001100100",
  54847=>"101101100",
  54848=>"100000101",
  54849=>"001010000",
  54850=>"110100110",
  54851=>"011001001",
  54852=>"100111111",
  54853=>"110111001",
  54854=>"010111000",
  54855=>"001001010",
  54856=>"110110010",
  54857=>"110000100",
  54858=>"111111011",
  54859=>"010110111",
  54860=>"010111000",
  54861=>"010001010",
  54862=>"111001111",
  54863=>"100110111",
  54864=>"101100011",
  54865=>"100010110",
  54866=>"000101101",
  54867=>"010111100",
  54868=>"011010010",
  54869=>"101000101",
  54870=>"001001001",
  54871=>"010011010",
  54872=>"001011000",
  54873=>"101111110",
  54874=>"000000001",
  54875=>"000100110",
  54876=>"100001111",
  54877=>"100101001",
  54878=>"110010111",
  54879=>"001000100",
  54880=>"001101000",
  54881=>"100101010",
  54882=>"101111100",
  54883=>"111000001",
  54884=>"001110110",
  54885=>"011010100",
  54886=>"100110101",
  54887=>"001101011",
  54888=>"101110101",
  54889=>"010110110",
  54890=>"000011101",
  54891=>"111100001",
  54892=>"001001010",
  54893=>"010001100",
  54894=>"001001000",
  54895=>"001011010",
  54896=>"011111110",
  54897=>"000011010",
  54898=>"110000110",
  54899=>"011011110",
  54900=>"001000111",
  54901=>"101101100",
  54902=>"001110000",
  54903=>"011011001",
  54904=>"010011001",
  54905=>"100000110",
  54906=>"000101001",
  54907=>"000111010",
  54908=>"111010010",
  54909=>"111111010",
  54910=>"000111100",
  54911=>"100010000",
  54912=>"010011111",
  54913=>"010000101",
  54914=>"010111001",
  54915=>"111101101",
  54916=>"010000110",
  54917=>"100110010",
  54918=>"101011011",
  54919=>"010101010",
  54920=>"011110000",
  54921=>"000101111",
  54922=>"000011011",
  54923=>"011001010",
  54924=>"101110011",
  54925=>"100010010",
  54926=>"010110101",
  54927=>"000011110",
  54928=>"010010111",
  54929=>"100000101",
  54930=>"111000000",
  54931=>"101001000",
  54932=>"100100010",
  54933=>"000110100",
  54934=>"111010011",
  54935=>"101001001",
  54936=>"011111000",
  54937=>"000101010",
  54938=>"100000011",
  54939=>"010010101",
  54940=>"100111010",
  54941=>"001010101",
  54942=>"111011111",
  54943=>"100001011",
  54944=>"100010100",
  54945=>"000100000",
  54946=>"100010001",
  54947=>"001000001",
  54948=>"101101000",
  54949=>"111100011",
  54950=>"001000000",
  54951=>"000000000",
  54952=>"111011011",
  54953=>"000100110",
  54954=>"010001011",
  54955=>"110010011",
  54956=>"011000010",
  54957=>"110011000",
  54958=>"001100111",
  54959=>"111000010",
  54960=>"000110110",
  54961=>"100001110",
  54962=>"001101000",
  54963=>"001111111",
  54964=>"111101011",
  54965=>"010011010",
  54966=>"000111101",
  54967=>"011010111",
  54968=>"011100000",
  54969=>"011001110",
  54970=>"110000100",
  54971=>"001100100",
  54972=>"110111111",
  54973=>"011110101",
  54974=>"000011110",
  54975=>"000001011",
  54976=>"011010110",
  54977=>"100111011",
  54978=>"010101101",
  54979=>"000010111",
  54980=>"100001011",
  54981=>"011100011",
  54982=>"111000010",
  54983=>"000101011",
  54984=>"011111000",
  54985=>"100000010",
  54986=>"111110111",
  54987=>"000001101",
  54988=>"100111000",
  54989=>"010010110",
  54990=>"010100000",
  54991=>"001111011",
  54992=>"000101111",
  54993=>"001001100",
  54994=>"100011111",
  54995=>"111101110",
  54996=>"101010000",
  54997=>"100100001",
  54998=>"011101001",
  54999=>"010001011",
  55000=>"011110011",
  55001=>"010011000",
  55002=>"010011000",
  55003=>"001101010",
  55004=>"010110000",
  55005=>"111111111",
  55006=>"101100101",
  55007=>"110101001",
  55008=>"001110010",
  55009=>"000000001",
  55010=>"001110010",
  55011=>"010101100",
  55012=>"010011011",
  55013=>"110000010",
  55014=>"001101011",
  55015=>"100010011",
  55016=>"100110000",
  55017=>"100110001",
  55018=>"100101100",
  55019=>"100100100",
  55020=>"000110111",
  55021=>"111010000",
  55022=>"010101110",
  55023=>"110011001",
  55024=>"111000001",
  55025=>"111011101",
  55026=>"111111010",
  55027=>"101110100",
  55028=>"011100100",
  55029=>"000000000",
  55030=>"100001010",
  55031=>"010000111",
  55032=>"010100011",
  55033=>"111010001",
  55034=>"101111000",
  55035=>"101010111",
  55036=>"100110110",
  55037=>"110110001",
  55038=>"100011101",
  55039=>"010110010",
  55040=>"101101111",
  55041=>"110110011",
  55042=>"100111101",
  55043=>"000010000",
  55044=>"101001000",
  55045=>"001010001",
  55046=>"100001011",
  55047=>"010101111",
  55048=>"101110100",
  55049=>"110101000",
  55050=>"011110011",
  55051=>"101110111",
  55052=>"110111010",
  55053=>"000001010",
  55054=>"100000010",
  55055=>"001101001",
  55056=>"011001011",
  55057=>"011101110",
  55058=>"111110110",
  55059=>"001000101",
  55060=>"000000101",
  55061=>"101100100",
  55062=>"000000111",
  55063=>"001101000",
  55064=>"101111011",
  55065=>"100010101",
  55066=>"010000001",
  55067=>"011011100",
  55068=>"110111010",
  55069=>"111011111",
  55070=>"110011100",
  55071=>"011110111",
  55072=>"111001111",
  55073=>"000001011",
  55074=>"011001110",
  55075=>"011101001",
  55076=>"110001000",
  55077=>"000111101",
  55078=>"011000010",
  55079=>"100100010",
  55080=>"000001000",
  55081=>"001000110",
  55082=>"110011101",
  55083=>"100010000",
  55084=>"001111010",
  55085=>"101011111",
  55086=>"111001001",
  55087=>"011000101",
  55088=>"101101000",
  55089=>"010001110",
  55090=>"101010011",
  55091=>"010010000",
  55092=>"111001110",
  55093=>"000010100",
  55094=>"100110111",
  55095=>"101011101",
  55096=>"100101111",
  55097=>"001010101",
  55098=>"011000010",
  55099=>"100111011",
  55100=>"111011001",
  55101=>"110011011",
  55102=>"010000000",
  55103=>"011110010",
  55104=>"011101000",
  55105=>"010001101",
  55106=>"100000000",
  55107=>"000010110",
  55108=>"111010001",
  55109=>"010110000",
  55110=>"000101010",
  55111=>"110101101",
  55112=>"001111101",
  55113=>"101011101",
  55114=>"100011110",
  55115=>"100001000",
  55116=>"001100001",
  55117=>"000111001",
  55118=>"111011010",
  55119=>"011111001",
  55120=>"000010110",
  55121=>"000110011",
  55122=>"000100001",
  55123=>"011111010",
  55124=>"101111011",
  55125=>"010000110",
  55126=>"101100000",
  55127=>"000011011",
  55128=>"110000000",
  55129=>"010110110",
  55130=>"100001001",
  55131=>"001000100",
  55132=>"101011001",
  55133=>"010110011",
  55134=>"011101111",
  55135=>"001100101",
  55136=>"000110001",
  55137=>"111000010",
  55138=>"111010010",
  55139=>"000011111",
  55140=>"110010010",
  55141=>"101011011",
  55142=>"011001110",
  55143=>"111001000",
  55144=>"101111011",
  55145=>"011000000",
  55146=>"001111100",
  55147=>"010001100",
  55148=>"000110110",
  55149=>"001100100",
  55150=>"100100001",
  55151=>"011010111",
  55152=>"000111010",
  55153=>"011100000",
  55154=>"010010000",
  55155=>"001000110",
  55156=>"001111010",
  55157=>"001010011",
  55158=>"010100011",
  55159=>"100101111",
  55160=>"001101100",
  55161=>"110101110",
  55162=>"001110011",
  55163=>"101101001",
  55164=>"100101101",
  55165=>"111101011",
  55166=>"100100010",
  55167=>"111110100",
  55168=>"000010111",
  55169=>"110111111",
  55170=>"101011110",
  55171=>"001011111",
  55172=>"010111110",
  55173=>"010000000",
  55174=>"101100011",
  55175=>"100000011",
  55176=>"010000011",
  55177=>"011110000",
  55178=>"010100011",
  55179=>"111011101",
  55180=>"100001000",
  55181=>"001000001",
  55182=>"011100100",
  55183=>"110111110",
  55184=>"110010000",
  55185=>"100100000",
  55186=>"110000001",
  55187=>"011011011",
  55188=>"101101000",
  55189=>"110100010",
  55190=>"001000101",
  55191=>"011110110",
  55192=>"101100101",
  55193=>"110100110",
  55194=>"001011111",
  55195=>"000110100",
  55196=>"000000111",
  55197=>"101000010",
  55198=>"100010100",
  55199=>"011001100",
  55200=>"001110101",
  55201=>"100001110",
  55202=>"001001101",
  55203=>"100001110",
  55204=>"000101000",
  55205=>"101001100",
  55206=>"001001101",
  55207=>"001000101",
  55208=>"000010100",
  55209=>"100000000",
  55210=>"011011100",
  55211=>"000011010",
  55212=>"111110010",
  55213=>"000100110",
  55214=>"111111111",
  55215=>"100011111",
  55216=>"000000011",
  55217=>"011100001",
  55218=>"001101101",
  55219=>"110000010",
  55220=>"100101011",
  55221=>"000000000",
  55222=>"101011101",
  55223=>"001101110",
  55224=>"101110011",
  55225=>"111011101",
  55226=>"011000111",
  55227=>"010001010",
  55228=>"000000001",
  55229=>"100011000",
  55230=>"010111000",
  55231=>"110011010",
  55232=>"010010100",
  55233=>"111110110",
  55234=>"010110111",
  55235=>"101011000",
  55236=>"111000111",
  55237=>"010000111",
  55238=>"111101100",
  55239=>"010101010",
  55240=>"110101111",
  55241=>"100010111",
  55242=>"100111110",
  55243=>"101100001",
  55244=>"100010001",
  55245=>"000000101",
  55246=>"101110100",
  55247=>"010101000",
  55248=>"101101110",
  55249=>"000011011",
  55250=>"000011111",
  55251=>"011111100",
  55252=>"000001011",
  55253=>"100001001",
  55254=>"000110001",
  55255=>"110101110",
  55256=>"110000000",
  55257=>"111110001",
  55258=>"000000100",
  55259=>"111100011",
  55260=>"000101110",
  55261=>"000101010",
  55262=>"010110111",
  55263=>"010100011",
  55264=>"111110011",
  55265=>"001100101",
  55266=>"110010110",
  55267=>"110100000",
  55268=>"000110000",
  55269=>"101100111",
  55270=>"001110111",
  55271=>"101011010",
  55272=>"010100110",
  55273=>"111110000",
  55274=>"100000001",
  55275=>"100000111",
  55276=>"100000010",
  55277=>"001111101",
  55278=>"100000010",
  55279=>"111011111",
  55280=>"111000110",
  55281=>"110101100",
  55282=>"010001111",
  55283=>"010011010",
  55284=>"010001111",
  55285=>"111110110",
  55286=>"111001010",
  55287=>"010100110",
  55288=>"100011001",
  55289=>"001100001",
  55290=>"110010101",
  55291=>"100001000",
  55292=>"011010100",
  55293=>"011110000",
  55294=>"111101110",
  55295=>"101100100",
  55296=>"001001101",
  55297=>"011010001",
  55298=>"000010011",
  55299=>"110111101",
  55300=>"010010111",
  55301=>"100110100",
  55302=>"011001010",
  55303=>"110000000",
  55304=>"010010000",
  55305=>"101110110",
  55306=>"010010100",
  55307=>"001011010",
  55308=>"111011000",
  55309=>"101110011",
  55310=>"010111000",
  55311=>"011111010",
  55312=>"110101000",
  55313=>"100111101",
  55314=>"111110000",
  55315=>"101010111",
  55316=>"001100111",
  55317=>"110001011",
  55318=>"001000101",
  55319=>"011100110",
  55320=>"001011001",
  55321=>"100011001",
  55322=>"011000101",
  55323=>"010001100",
  55324=>"111000100",
  55325=>"010110110",
  55326=>"010110100",
  55327=>"011000100",
  55328=>"001010000",
  55329=>"110000000",
  55330=>"010100000",
  55331=>"001000100",
  55332=>"010011000",
  55333=>"010001001",
  55334=>"111101100",
  55335=>"100101110",
  55336=>"111101110",
  55337=>"100000010",
  55338=>"011011101",
  55339=>"100110101",
  55340=>"000111101",
  55341=>"100010000",
  55342=>"011101001",
  55343=>"011100010",
  55344=>"000001101",
  55345=>"100001111",
  55346=>"101111111",
  55347=>"111100001",
  55348=>"001110110",
  55349=>"110110001",
  55350=>"010001101",
  55351=>"100000100",
  55352=>"001011100",
  55353=>"111011000",
  55354=>"010011110",
  55355=>"110100110",
  55356=>"101101110",
  55357=>"100001111",
  55358=>"001010011",
  55359=>"111101010",
  55360=>"101111000",
  55361=>"011101001",
  55362=>"001011110",
  55363=>"000000010",
  55364=>"100100110",
  55365=>"100110110",
  55366=>"011111010",
  55367=>"110110111",
  55368=>"110001100",
  55369=>"011000010",
  55370=>"101111011",
  55371=>"111110011",
  55372=>"110011101",
  55373=>"100001011",
  55374=>"000110101",
  55375=>"111101101",
  55376=>"100111001",
  55377=>"101001110",
  55378=>"101100000",
  55379=>"001110100",
  55380=>"000100110",
  55381=>"110011000",
  55382=>"001101110",
  55383=>"101001001",
  55384=>"001111111",
  55385=>"111000100",
  55386=>"001101001",
  55387=>"101110001",
  55388=>"011111111",
  55389=>"000110010",
  55390=>"010101100",
  55391=>"100110101",
  55392=>"011000000",
  55393=>"011101000",
  55394=>"011011110",
  55395=>"111111111",
  55396=>"000011011",
  55397=>"110010000",
  55398=>"011100000",
  55399=>"100110100",
  55400=>"111101111",
  55401=>"111101110",
  55402=>"011011101",
  55403=>"100011000",
  55404=>"111110101",
  55405=>"111111100",
  55406=>"110000110",
  55407=>"010110111",
  55408=>"000111001",
  55409=>"001001110",
  55410=>"111001010",
  55411=>"010011110",
  55412=>"111101101",
  55413=>"110011111",
  55414=>"101010000",
  55415=>"101011001",
  55416=>"111011111",
  55417=>"001001001",
  55418=>"111101110",
  55419=>"010001010",
  55420=>"111100010",
  55421=>"001011010",
  55422=>"001100011",
  55423=>"110110100",
  55424=>"011101001",
  55425=>"110000100",
  55426=>"001001010",
  55427=>"010110000",
  55428=>"001000000",
  55429=>"111100100",
  55430=>"000100110",
  55431=>"100010010",
  55432=>"010101101",
  55433=>"011010011",
  55434=>"100111000",
  55435=>"000111111",
  55436=>"100000010",
  55437=>"101001111",
  55438=>"010100110",
  55439=>"110010101",
  55440=>"101010100",
  55441=>"100100100",
  55442=>"010011101",
  55443=>"110110010",
  55444=>"111111101",
  55445=>"111110001",
  55446=>"000110111",
  55447=>"110101011",
  55448=>"110000100",
  55449=>"010010000",
  55450=>"101001011",
  55451=>"001111011",
  55452=>"010001000",
  55453=>"111101001",
  55454=>"111001000",
  55455=>"100010100",
  55456=>"111011111",
  55457=>"100111100",
  55458=>"000100010",
  55459=>"110111101",
  55460=>"001000010",
  55461=>"011011010",
  55462=>"110101000",
  55463=>"101110111",
  55464=>"110101000",
  55465=>"101011000",
  55466=>"001101000",
  55467=>"100000110",
  55468=>"111110101",
  55469=>"000111001",
  55470=>"010011100",
  55471=>"100011011",
  55472=>"001010001",
  55473=>"001000000",
  55474=>"000010011",
  55475=>"011101100",
  55476=>"111111110",
  55477=>"000001101",
  55478=>"000010100",
  55479=>"010110000",
  55480=>"100100011",
  55481=>"011100001",
  55482=>"000110010",
  55483=>"011011011",
  55484=>"111100000",
  55485=>"100111100",
  55486=>"010011101",
  55487=>"010111000",
  55488=>"000101001",
  55489=>"100000001",
  55490=>"101000000",
  55491=>"000000110",
  55492=>"101100101",
  55493=>"110100110",
  55494=>"101100110",
  55495=>"110110100",
  55496=>"100001011",
  55497=>"010001110",
  55498=>"110010011",
  55499=>"110110110",
  55500=>"100010111",
  55501=>"000100110",
  55502=>"111101110",
  55503=>"010100111",
  55504=>"011101011",
  55505=>"100100111",
  55506=>"000010001",
  55507=>"101100111",
  55508=>"101110110",
  55509=>"010101000",
  55510=>"011001010",
  55511=>"010001010",
  55512=>"011110011",
  55513=>"110000110",
  55514=>"111000011",
  55515=>"101100100",
  55516=>"011000111",
  55517=>"011111010",
  55518=>"110010010",
  55519=>"001110001",
  55520=>"100111110",
  55521=>"000011111",
  55522=>"000011011",
  55523=>"011010100",
  55524=>"011110111",
  55525=>"110111110",
  55526=>"111101111",
  55527=>"011000000",
  55528=>"100011100",
  55529=>"001101100",
  55530=>"000100011",
  55531=>"000001011",
  55532=>"101100100",
  55533=>"111100011",
  55534=>"100100011",
  55535=>"010111110",
  55536=>"010000010",
  55537=>"000011110",
  55538=>"011001101",
  55539=>"100101001",
  55540=>"011011011",
  55541=>"101011010",
  55542=>"110111111",
  55543=>"110101011",
  55544=>"110111000",
  55545=>"100101011",
  55546=>"110000010",
  55547=>"110010101",
  55548=>"000100110",
  55549=>"101010111",
  55550=>"101000100",
  55551=>"010001011",
  55552=>"111111100",
  55553=>"010111001",
  55554=>"010000110",
  55555=>"001011111",
  55556=>"011111000",
  55557=>"111110000",
  55558=>"110100100",
  55559=>"100001000",
  55560=>"101000100",
  55561=>"100010000",
  55562=>"111000011",
  55563=>"100001110",
  55564=>"010000110",
  55565=>"101111101",
  55566=>"101000101",
  55567=>"101100101",
  55568=>"000001011",
  55569=>"001011111",
  55570=>"011001101",
  55571=>"010100000",
  55572=>"100010000",
  55573=>"000001110",
  55574=>"000110010",
  55575=>"111011000",
  55576=>"011101100",
  55577=>"011110010",
  55578=>"101111010",
  55579=>"001101001",
  55580=>"010000001",
  55581=>"001011011",
  55582=>"111111110",
  55583=>"110001001",
  55584=>"001010000",
  55585=>"000111010",
  55586=>"111111101",
  55587=>"110000010",
  55588=>"100101001",
  55589=>"000101001",
  55590=>"001011001",
  55591=>"111001111",
  55592=>"000100111",
  55593=>"100110010",
  55594=>"100110011",
  55595=>"010011001",
  55596=>"101010001",
  55597=>"101101101",
  55598=>"110111110",
  55599=>"101010010",
  55600=>"000101000",
  55601=>"010100011",
  55602=>"011101010",
  55603=>"101001100",
  55604=>"110001110",
  55605=>"100101110",
  55606=>"100010000",
  55607=>"011011011",
  55608=>"001001010",
  55609=>"000100000",
  55610=>"110010000",
  55611=>"011000110",
  55612=>"100101000",
  55613=>"000101101",
  55614=>"010000110",
  55615=>"011111100",
  55616=>"111111011",
  55617=>"100101110",
  55618=>"111011001",
  55619=>"100011111",
  55620=>"111111111",
  55621=>"100001010",
  55622=>"111110110",
  55623=>"101111010",
  55624=>"111000010",
  55625=>"001000010",
  55626=>"111110000",
  55627=>"101000101",
  55628=>"100011001",
  55629=>"111100111",
  55630=>"010010010",
  55631=>"011110001",
  55632=>"101100111",
  55633=>"000100011",
  55634=>"011111010",
  55635=>"000010110",
  55636=>"011110100",
  55637=>"110101111",
  55638=>"001111101",
  55639=>"100001000",
  55640=>"110111111",
  55641=>"011000001",
  55642=>"010100011",
  55643=>"111001101",
  55644=>"011100100",
  55645=>"111110101",
  55646=>"101101001",
  55647=>"001111000",
  55648=>"000110101",
  55649=>"000001100",
  55650=>"000001011",
  55651=>"001001110",
  55652=>"101101101",
  55653=>"101011111",
  55654=>"101001110",
  55655=>"101001110",
  55656=>"110110011",
  55657=>"011101111",
  55658=>"000000101",
  55659=>"111100000",
  55660=>"000111111",
  55661=>"110001000",
  55662=>"101101000",
  55663=>"100011010",
  55664=>"111111001",
  55665=>"100001010",
  55666=>"100010110",
  55667=>"011111100",
  55668=>"000000010",
  55669=>"000010000",
  55670=>"111001111",
  55671=>"100001010",
  55672=>"110110000",
  55673=>"000100110",
  55674=>"011011000",
  55675=>"010000000",
  55676=>"000111000",
  55677=>"011101101",
  55678=>"001000011",
  55679=>"111110011",
  55680=>"101100100",
  55681=>"111010010",
  55682=>"100010001",
  55683=>"001001000",
  55684=>"110000110",
  55685=>"111011101",
  55686=>"001000010",
  55687=>"100010110",
  55688=>"000100111",
  55689=>"111001100",
  55690=>"100000100",
  55691=>"000111111",
  55692=>"101110011",
  55693=>"011000101",
  55694=>"000000010",
  55695=>"101101011",
  55696=>"101101001",
  55697=>"000011000",
  55698=>"111111000",
  55699=>"000010101",
  55700=>"111011111",
  55701=>"000011101",
  55702=>"100001011",
  55703=>"001000000",
  55704=>"101111111",
  55705=>"001000001",
  55706=>"011000001",
  55707=>"101101000",
  55708=>"010001101",
  55709=>"011010100",
  55710=>"011110000",
  55711=>"010100000",
  55712=>"001111111",
  55713=>"100001100",
  55714=>"111010100",
  55715=>"110100111",
  55716=>"100100001",
  55717=>"101110111",
  55718=>"111001001",
  55719=>"111001001",
  55720=>"111010010",
  55721=>"010010111",
  55722=>"001000001",
  55723=>"010001001",
  55724=>"010010111",
  55725=>"101010110",
  55726=>"000011011",
  55727=>"100101110",
  55728=>"101010110",
  55729=>"111100000",
  55730=>"001001110",
  55731=>"001011010",
  55732=>"110111111",
  55733=>"110100101",
  55734=>"110011100",
  55735=>"010101101",
  55736=>"011111011",
  55737=>"101101101",
  55738=>"011000111",
  55739=>"000001100",
  55740=>"111100111",
  55741=>"011110010",
  55742=>"000110010",
  55743=>"111010001",
  55744=>"011110010",
  55745=>"101001101",
  55746=>"000110000",
  55747=>"000101001",
  55748=>"100110011",
  55749=>"110100010",
  55750=>"000110111",
  55751=>"111000111",
  55752=>"111111001",
  55753=>"000011000",
  55754=>"101111111",
  55755=>"011000001",
  55756=>"101110111",
  55757=>"000001000",
  55758=>"010000100",
  55759=>"110010011",
  55760=>"011000010",
  55761=>"011001111",
  55762=>"100011000",
  55763=>"100110011",
  55764=>"101100111",
  55765=>"010010100",
  55766=>"000100000",
  55767=>"111010111",
  55768=>"000111011",
  55769=>"111101100",
  55770=>"010011101",
  55771=>"000111111",
  55772=>"011101010",
  55773=>"110010010",
  55774=>"011100100",
  55775=>"111101111",
  55776=>"011110110",
  55777=>"100000110",
  55778=>"011010111",
  55779=>"000011001",
  55780=>"101110000",
  55781=>"000000111",
  55782=>"010000001",
  55783=>"000011111",
  55784=>"111011100",
  55785=>"100111111",
  55786=>"110110110",
  55787=>"011101010",
  55788=>"001100111",
  55789=>"001000000",
  55790=>"110111111",
  55791=>"000100101",
  55792=>"010101110",
  55793=>"110100100",
  55794=>"100011001",
  55795=>"101001001",
  55796=>"100000010",
  55797=>"010101010",
  55798=>"011101100",
  55799=>"010001001",
  55800=>"011100011",
  55801=>"000011101",
  55802=>"110110111",
  55803=>"000001101",
  55804=>"001110001",
  55805=>"111110100",
  55806=>"010100001",
  55807=>"010101110",
  55808=>"100010011",
  55809=>"100010011",
  55810=>"111111011",
  55811=>"001001100",
  55812=>"000011000",
  55813=>"000100001",
  55814=>"010111001",
  55815=>"100000100",
  55816=>"000101011",
  55817=>"000000001",
  55818=>"100100010",
  55819=>"111011011",
  55820=>"010011010",
  55821=>"000001011",
  55822=>"000110110",
  55823=>"001110011",
  55824=>"000011101",
  55825=>"001111110",
  55826=>"100100101",
  55827=>"000011001",
  55828=>"111110011",
  55829=>"101001000",
  55830=>"111100111",
  55831=>"011010000",
  55832=>"000001101",
  55833=>"111000110",
  55834=>"010100001",
  55835=>"010101101",
  55836=>"000001100",
  55837=>"000111101",
  55838=>"000000010",
  55839=>"111101100",
  55840=>"111000011",
  55841=>"000010111",
  55842=>"100100010",
  55843=>"011001011",
  55844=>"100001001",
  55845=>"110000101",
  55846=>"011000001",
  55847=>"000010101",
  55848=>"111001110",
  55849=>"011011000",
  55850=>"100111001",
  55851=>"111011010",
  55852=>"111011000",
  55853=>"110101011",
  55854=>"111001010",
  55855=>"100011000",
  55856=>"101110010",
  55857=>"100000001",
  55858=>"111010011",
  55859=>"111001001",
  55860=>"001100000",
  55861=>"111000100",
  55862=>"111011000",
  55863=>"000001001",
  55864=>"000011101",
  55865=>"000011001",
  55866=>"101001110",
  55867=>"000111010",
  55868=>"111111110",
  55869=>"000100011",
  55870=>"000001000",
  55871=>"000001110",
  55872=>"001011110",
  55873=>"000000011",
  55874=>"000000011",
  55875=>"000010001",
  55876=>"010010111",
  55877=>"100101111",
  55878=>"001111110",
  55879=>"000000110",
  55880=>"001000111",
  55881=>"011011100",
  55882=>"000110010",
  55883=>"100110110",
  55884=>"110111010",
  55885=>"101011010",
  55886=>"001010001",
  55887=>"011010101",
  55888=>"001000001",
  55889=>"001001000",
  55890=>"101101010",
  55891=>"001011001",
  55892=>"000011111",
  55893=>"101011010",
  55894=>"101000111",
  55895=>"100001110",
  55896=>"000000100",
  55897=>"100101111",
  55898=>"010101010",
  55899=>"111000000",
  55900=>"101100111",
  55901=>"100111011",
  55902=>"111010111",
  55903=>"000111101",
  55904=>"100101001",
  55905=>"100101100",
  55906=>"000101000",
  55907=>"011010001",
  55908=>"001100110",
  55909=>"001000000",
  55910=>"001110101",
  55911=>"000110011",
  55912=>"101100101",
  55913=>"010011111",
  55914=>"001100001",
  55915=>"111101100",
  55916=>"110111001",
  55917=>"101100000",
  55918=>"000001110",
  55919=>"100101000",
  55920=>"001000111",
  55921=>"100000111",
  55922=>"111100100",
  55923=>"101100101",
  55924=>"001011010",
  55925=>"000001110",
  55926=>"111000011",
  55927=>"110101100",
  55928=>"000111000",
  55929=>"111010100",
  55930=>"110100110",
  55931=>"000111010",
  55932=>"011011110",
  55933=>"000000100",
  55934=>"010001101",
  55935=>"001101100",
  55936=>"001000011",
  55937=>"011111100",
  55938=>"110000101",
  55939=>"001011000",
  55940=>"111010000",
  55941=>"100110000",
  55942=>"001100010",
  55943=>"011000010",
  55944=>"010111110",
  55945=>"010000111",
  55946=>"000010000",
  55947=>"001111000",
  55948=>"100101000",
  55949=>"011010000",
  55950=>"110001101",
  55951=>"001110110",
  55952=>"100010100",
  55953=>"010010110",
  55954=>"011111111",
  55955=>"111101010",
  55956=>"011111010",
  55957=>"011110010",
  55958=>"101110010",
  55959=>"000010100",
  55960=>"001110100",
  55961=>"001001011",
  55962=>"111000001",
  55963=>"110101111",
  55964=>"001010110",
  55965=>"100111111",
  55966=>"101110110",
  55967=>"111111111",
  55968=>"110101100",
  55969=>"110000001",
  55970=>"110111100",
  55971=>"111010110",
  55972=>"010100011",
  55973=>"110011010",
  55974=>"110101110",
  55975=>"001000100",
  55976=>"000011010",
  55977=>"000111010",
  55978=>"110101100",
  55979=>"000101000",
  55980=>"011000110",
  55981=>"010100000",
  55982=>"111011100",
  55983=>"011110101",
  55984=>"010000111",
  55985=>"100101100",
  55986=>"001110001",
  55987=>"101001111",
  55988=>"011111001",
  55989=>"010100001",
  55990=>"111101111",
  55991=>"001001100",
  55992=>"111111010",
  55993=>"010001011",
  55994=>"110001001",
  55995=>"101011010",
  55996=>"110110111",
  55997=>"101101100",
  55998=>"001101111",
  55999=>"010110101",
  56000=>"101000110",
  56001=>"101110010",
  56002=>"000110000",
  56003=>"110000010",
  56004=>"010111001",
  56005=>"010101001",
  56006=>"010111111",
  56007=>"001100110",
  56008=>"111011001",
  56009=>"001111101",
  56010=>"011001011",
  56011=>"111111111",
  56012=>"000111000",
  56013=>"000000110",
  56014=>"000011110",
  56015=>"000001001",
  56016=>"010000000",
  56017=>"110110000",
  56018=>"010101110",
  56019=>"000010100",
  56020=>"110001101",
  56021=>"001110001",
  56022=>"101011000",
  56023=>"110111110",
  56024=>"001010111",
  56025=>"010011110",
  56026=>"011010101",
  56027=>"111000100",
  56028=>"011101001",
  56029=>"000100011",
  56030=>"111101101",
  56031=>"001001001",
  56032=>"001011110",
  56033=>"001100100",
  56034=>"011111101",
  56035=>"000010100",
  56036=>"000100011",
  56037=>"001111011",
  56038=>"001010010",
  56039=>"010101101",
  56040=>"000100111",
  56041=>"011110100",
  56042=>"000111110",
  56043=>"011110010",
  56044=>"000011101",
  56045=>"100111011",
  56046=>"111010100",
  56047=>"111111011",
  56048=>"111011111",
  56049=>"100101111",
  56050=>"100100101",
  56051=>"001010001",
  56052=>"010011101",
  56053=>"110011111",
  56054=>"100110110",
  56055=>"100000111",
  56056=>"011000011",
  56057=>"010010000",
  56058=>"110000101",
  56059=>"011100000",
  56060=>"111011110",
  56061=>"011000011",
  56062=>"011101101",
  56063=>"001011110",
  56064=>"010011000",
  56065=>"010010010",
  56066=>"100100100",
  56067=>"010001010",
  56068=>"010000100",
  56069=>"000000010",
  56070=>"100110110",
  56071=>"000011100",
  56072=>"001001101",
  56073=>"011100100",
  56074=>"000011010",
  56075=>"011011100",
  56076=>"110110100",
  56077=>"101001010",
  56078=>"000111011",
  56079=>"011010100",
  56080=>"110001010",
  56081=>"100000101",
  56082=>"101011100",
  56083=>"001001111",
  56084=>"100000011",
  56085=>"001011010",
  56086=>"011001001",
  56087=>"100001101",
  56088=>"001001101",
  56089=>"011011000",
  56090=>"001010000",
  56091=>"001111011",
  56092=>"000011111",
  56093=>"000100010",
  56094=>"111011010",
  56095=>"101100100",
  56096=>"101010101",
  56097=>"111101001",
  56098=>"000101010",
  56099=>"111001010",
  56100=>"010111110",
  56101=>"100001100",
  56102=>"110111110",
  56103=>"011100010",
  56104=>"011011110",
  56105=>"111111110",
  56106=>"001111001",
  56107=>"110010111",
  56108=>"110000111",
  56109=>"000100101",
  56110=>"000000110",
  56111=>"101000110",
  56112=>"001100101",
  56113=>"111000011",
  56114=>"100001100",
  56115=>"001000110",
  56116=>"111000011",
  56117=>"000101101",
  56118=>"100101011",
  56119=>"000110001",
  56120=>"011011001",
  56121=>"101011000",
  56122=>"100101010",
  56123=>"111000100",
  56124=>"110010001",
  56125=>"100111101",
  56126=>"000100100",
  56127=>"010001000",
  56128=>"111100001",
  56129=>"110001011",
  56130=>"110110110",
  56131=>"001100101",
  56132=>"101111101",
  56133=>"010000100",
  56134=>"111100101",
  56135=>"110011001",
  56136=>"101010111",
  56137=>"011000001",
  56138=>"111000011",
  56139=>"000110000",
  56140=>"100101101",
  56141=>"001101000",
  56142=>"100100001",
  56143=>"100000010",
  56144=>"101101001",
  56145=>"000001000",
  56146=>"000001011",
  56147=>"011010011",
  56148=>"100100000",
  56149=>"000101000",
  56150=>"011100110",
  56151=>"111011111",
  56152=>"110010100",
  56153=>"011011010",
  56154=>"101111101",
  56155=>"010010101",
  56156=>"110001011",
  56157=>"100111110",
  56158=>"100111001",
  56159=>"011011001",
  56160=>"101001110",
  56161=>"111101001",
  56162=>"001111100",
  56163=>"010001101",
  56164=>"011110111",
  56165=>"110010111",
  56166=>"000011111",
  56167=>"001011110",
  56168=>"011000010",
  56169=>"101100111",
  56170=>"010101110",
  56171=>"011111000",
  56172=>"000110111",
  56173=>"001100000",
  56174=>"010101011",
  56175=>"101010010",
  56176=>"111001101",
  56177=>"000101100",
  56178=>"110000000",
  56179=>"010000110",
  56180=>"100101100",
  56181=>"001111111",
  56182=>"111010010",
  56183=>"001010101",
  56184=>"011001101",
  56185=>"011110010",
  56186=>"000111101",
  56187=>"111011100",
  56188=>"010001111",
  56189=>"101011000",
  56190=>"000000100",
  56191=>"111011111",
  56192=>"000111000",
  56193=>"101011111",
  56194=>"001100101",
  56195=>"000100000",
  56196=>"110011111",
  56197=>"110010101",
  56198=>"101100101",
  56199=>"101100001",
  56200=>"111100010",
  56201=>"100000010",
  56202=>"001101100",
  56203=>"110110101",
  56204=>"010110000",
  56205=>"000100001",
  56206=>"111010000",
  56207=>"100110010",
  56208=>"000110100",
  56209=>"001101100",
  56210=>"011011110",
  56211=>"011011010",
  56212=>"100010010",
  56213=>"100110110",
  56214=>"011000110",
  56215=>"111100010",
  56216=>"011111000",
  56217=>"000111011",
  56218=>"110101100",
  56219=>"010011110",
  56220=>"101000111",
  56221=>"001000101",
  56222=>"100001001",
  56223=>"101001001",
  56224=>"111000010",
  56225=>"111111111",
  56226=>"110011101",
  56227=>"100110101",
  56228=>"110000100",
  56229=>"000011000",
  56230=>"000111111",
  56231=>"100111111",
  56232=>"110110110",
  56233=>"000100000",
  56234=>"101100101",
  56235=>"111011011",
  56236=>"101111000",
  56237=>"101101101",
  56238=>"100011110",
  56239=>"100111010",
  56240=>"011001000",
  56241=>"010111110",
  56242=>"110110110",
  56243=>"111101011",
  56244=>"011001010",
  56245=>"100110010",
  56246=>"001111111",
  56247=>"010000010",
  56248=>"110000000",
  56249=>"101110000",
  56250=>"110010100",
  56251=>"001111111",
  56252=>"000110101",
  56253=>"000101111",
  56254=>"111011001",
  56255=>"111111101",
  56256=>"000011001",
  56257=>"010111110",
  56258=>"010011111",
  56259=>"101001000",
  56260=>"010110111",
  56261=>"011101010",
  56262=>"011101100",
  56263=>"111010110",
  56264=>"100101010",
  56265=>"011100100",
  56266=>"001110001",
  56267=>"111111000",
  56268=>"010010110",
  56269=>"101011001",
  56270=>"100011110",
  56271=>"110111111",
  56272=>"110000011",
  56273=>"110100110",
  56274=>"010110100",
  56275=>"100001100",
  56276=>"001000000",
  56277=>"001011000",
  56278=>"101000010",
  56279=>"111000101",
  56280=>"010010000",
  56281=>"010101010",
  56282=>"110111100",
  56283=>"111101010",
  56284=>"111110101",
  56285=>"110100100",
  56286=>"110110110",
  56287=>"001001110",
  56288=>"010111010",
  56289=>"000110001",
  56290=>"010101001",
  56291=>"101101110",
  56292=>"001001101",
  56293=>"101111101",
  56294=>"100100011",
  56295=>"000000010",
  56296=>"010011000",
  56297=>"000111101",
  56298=>"010110001",
  56299=>"111111100",
  56300=>"110111011",
  56301=>"101111100",
  56302=>"100101011",
  56303=>"000101000",
  56304=>"011100010",
  56305=>"010100100",
  56306=>"101100110",
  56307=>"101101110",
  56308=>"000011101",
  56309=>"001100110",
  56310=>"001110010",
  56311=>"011110001",
  56312=>"110111011",
  56313=>"001010010",
  56314=>"000110000",
  56315=>"111111110",
  56316=>"010100000",
  56317=>"111100110",
  56318=>"101010101",
  56319=>"011110111",
  56320=>"011011011",
  56321=>"100100001",
  56322=>"110001010",
  56323=>"110110101",
  56324=>"000100111",
  56325=>"001001011",
  56326=>"011101101",
  56327=>"111000010",
  56328=>"011110100",
  56329=>"001000110",
  56330=>"110000111",
  56331=>"100110110",
  56332=>"000111011",
  56333=>"111100001",
  56334=>"000110011",
  56335=>"010101100",
  56336=>"010001100",
  56337=>"100010010",
  56338=>"000110000",
  56339=>"011110110",
  56340=>"010001111",
  56341=>"010110011",
  56342=>"000001110",
  56343=>"000111111",
  56344=>"111000110",
  56345=>"010000101",
  56346=>"000101111",
  56347=>"011011111",
  56348=>"011111101",
  56349=>"010110001",
  56350=>"111110111",
  56351=>"011111111",
  56352=>"001100001",
  56353=>"111001101",
  56354=>"110010011",
  56355=>"100000101",
  56356=>"101111111",
  56357=>"011001110",
  56358=>"111010110",
  56359=>"111011100",
  56360=>"010100101",
  56361=>"010101001",
  56362=>"110110000",
  56363=>"000000100",
  56364=>"101011000",
  56365=>"010101100",
  56366=>"010011010",
  56367=>"101110101",
  56368=>"111010011",
  56369=>"101100000",
  56370=>"011001001",
  56371=>"111010111",
  56372=>"011100000",
  56373=>"111110011",
  56374=>"101111000",
  56375=>"101111111",
  56376=>"100011100",
  56377=>"010111101",
  56378=>"111011110",
  56379=>"110110110",
  56380=>"000000001",
  56381=>"000101011",
  56382=>"111100101",
  56383=>"011101010",
  56384=>"100100101",
  56385=>"000000010",
  56386=>"110100010",
  56387=>"001010100",
  56388=>"010100010",
  56389=>"011001111",
  56390=>"000001110",
  56391=>"000100001",
  56392=>"001001010",
  56393=>"111100000",
  56394=>"111000001",
  56395=>"100010001",
  56396=>"111110101",
  56397=>"100001100",
  56398=>"010111100",
  56399=>"000000001",
  56400=>"001000101",
  56401=>"010001110",
  56402=>"010001001",
  56403=>"001011001",
  56404=>"111001011",
  56405=>"001010101",
  56406=>"001000110",
  56407=>"100110001",
  56408=>"010011100",
  56409=>"000111011",
  56410=>"100001110",
  56411=>"101010001",
  56412=>"000010100",
  56413=>"011010010",
  56414=>"110000110",
  56415=>"100000100",
  56416=>"110010001",
  56417=>"011000000",
  56418=>"110000100",
  56419=>"010010010",
  56420=>"111000011",
  56421=>"001101001",
  56422=>"011001001",
  56423=>"100100011",
  56424=>"110100100",
  56425=>"101001001",
  56426=>"011110101",
  56427=>"011111111",
  56428=>"110110111",
  56429=>"001101100",
  56430=>"011110010",
  56431=>"010000000",
  56432=>"110110111",
  56433=>"110011101",
  56434=>"001000100",
  56435=>"110011011",
  56436=>"001100000",
  56437=>"101101010",
  56438=>"000111111",
  56439=>"101100101",
  56440=>"001001010",
  56441=>"000011100",
  56442=>"100101100",
  56443=>"110011001",
  56444=>"001011101",
  56445=>"001110110",
  56446=>"000010000",
  56447=>"101110010",
  56448=>"000101100",
  56449=>"100010100",
  56450=>"110001010",
  56451=>"000101000",
  56452=>"100010011",
  56453=>"110111101",
  56454=>"111110001",
  56455=>"111011011",
  56456=>"111001011",
  56457=>"100011110",
  56458=>"011110011",
  56459=>"110100011",
  56460=>"010001111",
  56461=>"000010101",
  56462=>"011111000",
  56463=>"001010111",
  56464=>"101011110",
  56465=>"011011110",
  56466=>"110101000",
  56467=>"110101010",
  56468=>"010111101",
  56469=>"010000010",
  56470=>"101001100",
  56471=>"010001011",
  56472=>"011011010",
  56473=>"110010100",
  56474=>"010101110",
  56475=>"101100001",
  56476=>"110010010",
  56477=>"010100100",
  56478=>"110111101",
  56479=>"010010111",
  56480=>"011010000",
  56481=>"111111100",
  56482=>"100001110",
  56483=>"001000101",
  56484=>"001110000",
  56485=>"001011100",
  56486=>"011110010",
  56487=>"111111101",
  56488=>"001110011",
  56489=>"011001000",
  56490=>"010011100",
  56491=>"110001011",
  56492=>"000111100",
  56493=>"010010011",
  56494=>"011101101",
  56495=>"011111011",
  56496=>"111111001",
  56497=>"011100111",
  56498=>"101010000",
  56499=>"001100000",
  56500=>"000010100",
  56501=>"111111110",
  56502=>"000011000",
  56503=>"000101011",
  56504=>"100101001",
  56505=>"000111001",
  56506=>"000000110",
  56507=>"111101100",
  56508=>"000011001",
  56509=>"101100010",
  56510=>"101101010",
  56511=>"000011101",
  56512=>"011010111",
  56513=>"111000000",
  56514=>"111010110",
  56515=>"001110010",
  56516=>"111100001",
  56517=>"010000011",
  56518=>"101101011",
  56519=>"000101110",
  56520=>"001110001",
  56521=>"000010111",
  56522=>"111011100",
  56523=>"110110011",
  56524=>"110001111",
  56525=>"000110001",
  56526=>"011001011",
  56527=>"101110101",
  56528=>"011110011",
  56529=>"010101100",
  56530=>"110010001",
  56531=>"110001101",
  56532=>"000000000",
  56533=>"011000000",
  56534=>"011001001",
  56535=>"001101001",
  56536=>"111111100",
  56537=>"000111000",
  56538=>"110000000",
  56539=>"101110101",
  56540=>"101100010",
  56541=>"101111001",
  56542=>"001100001",
  56543=>"111110001",
  56544=>"100000100",
  56545=>"101001000",
  56546=>"010100111",
  56547=>"010010111",
  56548=>"110101000",
  56549=>"110011110",
  56550=>"111011111",
  56551=>"100001110",
  56552=>"011110010",
  56553=>"101000110",
  56554=>"100101111",
  56555=>"100000100",
  56556=>"000001001",
  56557=>"110101010",
  56558=>"111011111",
  56559=>"011101011",
  56560=>"110111111",
  56561=>"111101111",
  56562=>"010100101",
  56563=>"100111100",
  56564=>"101101110",
  56565=>"010010110",
  56566=>"010100110",
  56567=>"110000001",
  56568=>"100000000",
  56569=>"001111101",
  56570=>"001001101",
  56571=>"000011110",
  56572=>"110001010",
  56573=>"111101101",
  56574=>"000011010",
  56575=>"110110010",
  56576=>"110101000",
  56577=>"001101000",
  56578=>"111001000",
  56579=>"100001010",
  56580=>"000001100",
  56581=>"001010101",
  56582=>"111111101",
  56583=>"111100000",
  56584=>"100010110",
  56585=>"001110110",
  56586=>"101111111",
  56587=>"111110011",
  56588=>"111000100",
  56589=>"111110000",
  56590=>"111001001",
  56591=>"000000000",
  56592=>"000110001",
  56593=>"000011001",
  56594=>"000111010",
  56595=>"001111001",
  56596=>"011001001",
  56597=>"011011010",
  56598=>"100000001",
  56599=>"010101111",
  56600=>"000000010",
  56601=>"011100101",
  56602=>"100110110",
  56603=>"100110001",
  56604=>"000101111",
  56605=>"111111000",
  56606=>"010010001",
  56607=>"101000000",
  56608=>"111001100",
  56609=>"000100111",
  56610=>"001100101",
  56611=>"111011111",
  56612=>"000100001",
  56613=>"100001011",
  56614=>"010110101",
  56615=>"010010011",
  56616=>"011001110",
  56617=>"010001111",
  56618=>"000010110",
  56619=>"011101101",
  56620=>"100110100",
  56621=>"100011110",
  56622=>"100100000",
  56623=>"101111100",
  56624=>"101010011",
  56625=>"001100010",
  56626=>"111110101",
  56627=>"010110110",
  56628=>"101110001",
  56629=>"000001000",
  56630=>"010010010",
  56631=>"100110101",
  56632=>"010000111",
  56633=>"101100000",
  56634=>"010101100",
  56635=>"110110111",
  56636=>"000000011",
  56637=>"000111010",
  56638=>"000000110",
  56639=>"011101101",
  56640=>"001010011",
  56641=>"010001100",
  56642=>"001001101",
  56643=>"110000000",
  56644=>"110110100",
  56645=>"100111110",
  56646=>"000000000",
  56647=>"101100000",
  56648=>"001001111",
  56649=>"010100101",
  56650=>"001000000",
  56651=>"000001011",
  56652=>"101010100",
  56653=>"100101110",
  56654=>"100000010",
  56655=>"101111001",
  56656=>"001010000",
  56657=>"000010001",
  56658=>"011101111",
  56659=>"100000100",
  56660=>"101101101",
  56661=>"010111110",
  56662=>"000010011",
  56663=>"011011101",
  56664=>"011010000",
  56665=>"001000110",
  56666=>"000011111",
  56667=>"001000011",
  56668=>"101101101",
  56669=>"111111010",
  56670=>"010101010",
  56671=>"011001100",
  56672=>"011011110",
  56673=>"010111100",
  56674=>"111101110",
  56675=>"111110000",
  56676=>"010100111",
  56677=>"110100000",
  56678=>"001000100",
  56679=>"110110010",
  56680=>"001000011",
  56681=>"000010111",
  56682=>"011101101",
  56683=>"110010111",
  56684=>"100011110",
  56685=>"000011011",
  56686=>"111100001",
  56687=>"100010100",
  56688=>"010101111",
  56689=>"010101111",
  56690=>"000101010",
  56691=>"100011000",
  56692=>"100110111",
  56693=>"011011010",
  56694=>"111110111",
  56695=>"111110000",
  56696=>"011001100",
  56697=>"101110110",
  56698=>"111001000",
  56699=>"001000010",
  56700=>"100101101",
  56701=>"111111111",
  56702=>"011100000",
  56703=>"101110111",
  56704=>"111101111",
  56705=>"100111110",
  56706=>"011111101",
  56707=>"101000001",
  56708=>"101011010",
  56709=>"101001101",
  56710=>"110110001",
  56711=>"110000001",
  56712=>"011111010",
  56713=>"011100010",
  56714=>"100011010",
  56715=>"111110111",
  56716=>"110011111",
  56717=>"011011110",
  56718=>"000011101",
  56719=>"101100100",
  56720=>"000000111",
  56721=>"101101111",
  56722=>"111000010",
  56723=>"111010111",
  56724=>"110000001",
  56725=>"010011100",
  56726=>"000000010",
  56727=>"000111111",
  56728=>"110001101",
  56729=>"011110111",
  56730=>"100000000",
  56731=>"110101100",
  56732=>"111001010",
  56733=>"001001000",
  56734=>"010110111",
  56735=>"100100100",
  56736=>"001000000",
  56737=>"000111110",
  56738=>"001110011",
  56739=>"011000010",
  56740=>"001110000",
  56741=>"101000001",
  56742=>"000000110",
  56743=>"110000011",
  56744=>"001101000",
  56745=>"010100000",
  56746=>"011101110",
  56747=>"110100110",
  56748=>"111110110",
  56749=>"100001000",
  56750=>"110010000",
  56751=>"010000000",
  56752=>"011011110",
  56753=>"111010111",
  56754=>"010001110",
  56755=>"100110101",
  56756=>"111001100",
  56757=>"110111111",
  56758=>"000001101",
  56759=>"110110000",
  56760=>"100001101",
  56761=>"010100000",
  56762=>"011101010",
  56763=>"001100111",
  56764=>"101110111",
  56765=>"101001100",
  56766=>"001100000",
  56767=>"011000110",
  56768=>"000111111",
  56769=>"110100101",
  56770=>"111101100",
  56771=>"001011111",
  56772=>"101110101",
  56773=>"110101101",
  56774=>"001010111",
  56775=>"001100111",
  56776=>"111100111",
  56777=>"101000101",
  56778=>"100000000",
  56779=>"010010010",
  56780=>"010000000",
  56781=>"011111001",
  56782=>"110111001",
  56783=>"000111101",
  56784=>"101101011",
  56785=>"000111001",
  56786=>"011110001",
  56787=>"101110111",
  56788=>"100000101",
  56789=>"010011110",
  56790=>"011110110",
  56791=>"110000010",
  56792=>"111000000",
  56793=>"100001001",
  56794=>"001000000",
  56795=>"110101001",
  56796=>"110000010",
  56797=>"011111011",
  56798=>"001110111",
  56799=>"100101100",
  56800=>"111000100",
  56801=>"011000001",
  56802=>"101110100",
  56803=>"101110111",
  56804=>"101101100",
  56805=>"110100111",
  56806=>"110000110",
  56807=>"100011011",
  56808=>"001000001",
  56809=>"011011111",
  56810=>"010001001",
  56811=>"111110111",
  56812=>"011001011",
  56813=>"101000100",
  56814=>"110011010",
  56815=>"010110100",
  56816=>"101100010",
  56817=>"111101111",
  56818=>"111100010",
  56819=>"010011111",
  56820=>"010100110",
  56821=>"010000100",
  56822=>"100111011",
  56823=>"100111011",
  56824=>"011101010",
  56825=>"001001010",
  56826=>"000101111",
  56827=>"101010100",
  56828=>"001001011",
  56829=>"111001101",
  56830=>"111001110",
  56831=>"011101111",
  56832=>"111111000",
  56833=>"000010111",
  56834=>"010111110",
  56835=>"111100110",
  56836=>"111101101",
  56837=>"111001110",
  56838=>"011100011",
  56839=>"010010110",
  56840=>"101010111",
  56841=>"000011001",
  56842=>"111110101",
  56843=>"001011001",
  56844=>"111001111",
  56845=>"110110001",
  56846=>"110000011",
  56847=>"100010000",
  56848=>"010101100",
  56849=>"010100110",
  56850=>"011011001",
  56851=>"001101110",
  56852=>"110101110",
  56853=>"011010001",
  56854=>"101010100",
  56855=>"110100110",
  56856=>"010101001",
  56857=>"101110001",
  56858=>"101111011",
  56859=>"001101100",
  56860=>"100101111",
  56861=>"101001001",
  56862=>"101001100",
  56863=>"111001010",
  56864=>"100101011",
  56865=>"011011110",
  56866=>"000101000",
  56867=>"010111101",
  56868=>"011101000",
  56869=>"001101101",
  56870=>"100010001",
  56871=>"000111100",
  56872=>"001000010",
  56873=>"110111011",
  56874=>"001000000",
  56875=>"010100111",
  56876=>"101101000",
  56877=>"001111011",
  56878=>"101111001",
  56879=>"110100001",
  56880=>"001000001",
  56881=>"101111111",
  56882=>"001000010",
  56883=>"001100000",
  56884=>"010000100",
  56885=>"110000010",
  56886=>"110010001",
  56887=>"110101100",
  56888=>"000100011",
  56889=>"011100110",
  56890=>"011000111",
  56891=>"000001110",
  56892=>"001111000",
  56893=>"111011101",
  56894=>"011111000",
  56895=>"100000110",
  56896=>"000111111",
  56897=>"111010111",
  56898=>"100000000",
  56899=>"111001101",
  56900=>"001110001",
  56901=>"101111101",
  56902=>"001001010",
  56903=>"001100001",
  56904=>"111111011",
  56905=>"001001110",
  56906=>"111011111",
  56907=>"101110101",
  56908=>"000001100",
  56909=>"011001100",
  56910=>"100001111",
  56911=>"101001110",
  56912=>"100101110",
  56913=>"000101011",
  56914=>"111100110",
  56915=>"110110011",
  56916=>"001010010",
  56917=>"011101010",
  56918=>"001010110",
  56919=>"111010011",
  56920=>"001100101",
  56921=>"000001011",
  56922=>"100110101",
  56923=>"101110011",
  56924=>"000101010",
  56925=>"111001101",
  56926=>"110111111",
  56927=>"010100000",
  56928=>"001011010",
  56929=>"000101111",
  56930=>"101111111",
  56931=>"011010000",
  56932=>"001001100",
  56933=>"010100101",
  56934=>"000100110",
  56935=>"000000110",
  56936=>"000100101",
  56937=>"010011010",
  56938=>"011010001",
  56939=>"110011110",
  56940=>"111010110",
  56941=>"000011001",
  56942=>"010110101",
  56943=>"100011111",
  56944=>"100001010",
  56945=>"010001000",
  56946=>"011111010",
  56947=>"000001100",
  56948=>"001000101",
  56949=>"111011110",
  56950=>"001001010",
  56951=>"110000011",
  56952=>"100111111",
  56953=>"001011111",
  56954=>"110111101",
  56955=>"000101011",
  56956=>"110011100",
  56957=>"000110011",
  56958=>"011000100",
  56959=>"000001101",
  56960=>"001110111",
  56961=>"111101101",
  56962=>"111000000",
  56963=>"111111111",
  56964=>"110110011",
  56965=>"100000111",
  56966=>"001111000",
  56967=>"101111101",
  56968=>"000001110",
  56969=>"000100100",
  56970=>"001100010",
  56971=>"011111000",
  56972=>"001000101",
  56973=>"111000100",
  56974=>"010010000",
  56975=>"101001000",
  56976=>"011111110",
  56977=>"010001010",
  56978=>"010110011",
  56979=>"011111011",
  56980=>"111111101",
  56981=>"010110101",
  56982=>"010000000",
  56983=>"000101001",
  56984=>"111001010",
  56985=>"110011000",
  56986=>"001101000",
  56987=>"001101101",
  56988=>"011110001",
  56989=>"101010111",
  56990=>"111110000",
  56991=>"000000101",
  56992=>"100100101",
  56993=>"101101101",
  56994=>"111110101",
  56995=>"010010011",
  56996=>"001100110",
  56997=>"000011001",
  56998=>"111001000",
  56999=>"100001010",
  57000=>"111100001",
  57001=>"010010000",
  57002=>"111000110",
  57003=>"000010010",
  57004=>"001011110",
  57005=>"110101000",
  57006=>"000000000",
  57007=>"110100011",
  57008=>"010001101",
  57009=>"000100100",
  57010=>"011100111",
  57011=>"001100010",
  57012=>"100011110",
  57013=>"011000110",
  57014=>"001101100",
  57015=>"101001110",
  57016=>"000101011",
  57017=>"111011010",
  57018=>"000100000",
  57019=>"101110101",
  57020=>"111100111",
  57021=>"101101001",
  57022=>"010110000",
  57023=>"101010010",
  57024=>"001101111",
  57025=>"111100101",
  57026=>"010010000",
  57027=>"101100000",
  57028=>"100110000",
  57029=>"011101000",
  57030=>"001110111",
  57031=>"111110111",
  57032=>"000100000",
  57033=>"100011111",
  57034=>"101110110",
  57035=>"011010000",
  57036=>"001100011",
  57037=>"011111011",
  57038=>"000011000",
  57039=>"011100001",
  57040=>"111010001",
  57041=>"111001010",
  57042=>"011001010",
  57043=>"000011001",
  57044=>"101000011",
  57045=>"100001111",
  57046=>"011001111",
  57047=>"100011000",
  57048=>"011010000",
  57049=>"000100001",
  57050=>"010101010",
  57051=>"111101101",
  57052=>"011111110",
  57053=>"110010110",
  57054=>"010111110",
  57055=>"101010101",
  57056=>"011011101",
  57057=>"101011110",
  57058=>"111100000",
  57059=>"010100111",
  57060=>"000001111",
  57061=>"000111100",
  57062=>"110100110",
  57063=>"110101011",
  57064=>"111000001",
  57065=>"011000110",
  57066=>"000101100",
  57067=>"001010110",
  57068=>"000100111",
  57069=>"100000110",
  57070=>"010110011",
  57071=>"011011110",
  57072=>"001100111",
  57073=>"010100111",
  57074=>"010110101",
  57075=>"100101111",
  57076=>"001101011",
  57077=>"111000010",
  57078=>"000001011",
  57079=>"110110011",
  57080=>"011101101",
  57081=>"110101001",
  57082=>"111011001",
  57083=>"110001101",
  57084=>"010011010",
  57085=>"000111101",
  57086=>"011100111",
  57087=>"110100101",
  57088=>"101101011",
  57089=>"001110110",
  57090=>"100110011",
  57091=>"010000100",
  57092=>"111011100",
  57093=>"011010000",
  57094=>"111010001",
  57095=>"010000111",
  57096=>"110101110",
  57097=>"001010010",
  57098=>"100100101",
  57099=>"010000000",
  57100=>"100000010",
  57101=>"110100111",
  57102=>"111010011",
  57103=>"000100101",
  57104=>"010111110",
  57105=>"000111001",
  57106=>"111111101",
  57107=>"000111111",
  57108=>"101110100",
  57109=>"110011100",
  57110=>"100010110",
  57111=>"111000000",
  57112=>"001110101",
  57113=>"111000111",
  57114=>"001000101",
  57115=>"100101011",
  57116=>"011011000",
  57117=>"011010110",
  57118=>"110010010",
  57119=>"000111001",
  57120=>"111111111",
  57121=>"101001001",
  57122=>"111111001",
  57123=>"001101010",
  57124=>"101010111",
  57125=>"100001111",
  57126=>"000010100",
  57127=>"010110011",
  57128=>"111001000",
  57129=>"101010010",
  57130=>"011101110",
  57131=>"111111011",
  57132=>"101100011",
  57133=>"000110000",
  57134=>"100100111",
  57135=>"010111100",
  57136=>"111111000",
  57137=>"000001100",
  57138=>"010100001",
  57139=>"110111000",
  57140=>"111111111",
  57141=>"010110111",
  57142=>"100000100",
  57143=>"111111000",
  57144=>"010011100",
  57145=>"011100011",
  57146=>"110011011",
  57147=>"101100110",
  57148=>"110110101",
  57149=>"011010010",
  57150=>"001101110",
  57151=>"011001100",
  57152=>"011100100",
  57153=>"011000110",
  57154=>"100100110",
  57155=>"111100100",
  57156=>"000001101",
  57157=>"001010110",
  57158=>"100011111",
  57159=>"010110111",
  57160=>"011110010",
  57161=>"001100100",
  57162=>"010001110",
  57163=>"000110000",
  57164=>"110111111",
  57165=>"110100110",
  57166=>"001000100",
  57167=>"111100000",
  57168=>"011010001",
  57169=>"110110101",
  57170=>"110011100",
  57171=>"100010011",
  57172=>"111111100",
  57173=>"010010010",
  57174=>"101001000",
  57175=>"010000101",
  57176=>"010101100",
  57177=>"000000001",
  57178=>"000111110",
  57179=>"110000010",
  57180=>"111011001",
  57181=>"000001001",
  57182=>"110001111",
  57183=>"101001111",
  57184=>"011000000",
  57185=>"111000011",
  57186=>"001011111",
  57187=>"100010010",
  57188=>"011111000",
  57189=>"000011101",
  57190=>"000011000",
  57191=>"101011101",
  57192=>"001010000",
  57193=>"101111011",
  57194=>"111110111",
  57195=>"110001001",
  57196=>"111100110",
  57197=>"010000001",
  57198=>"011000010",
  57199=>"111000000",
  57200=>"011001111",
  57201=>"010101111",
  57202=>"010111100",
  57203=>"111111101",
  57204=>"000000001",
  57205=>"110010101",
  57206=>"011100101",
  57207=>"011101000",
  57208=>"100001101",
  57209=>"100011000",
  57210=>"110011110",
  57211=>"111100110",
  57212=>"101011010",
  57213=>"001011011",
  57214=>"011111001",
  57215=>"001111000",
  57216=>"010100000",
  57217=>"011111001",
  57218=>"110110111",
  57219=>"010000100",
  57220=>"001000100",
  57221=>"100011011",
  57222=>"111111100",
  57223=>"100101001",
  57224=>"001011111",
  57225=>"111000010",
  57226=>"110101101",
  57227=>"000010101",
  57228=>"111100010",
  57229=>"011110000",
  57230=>"000111110",
  57231=>"010111000",
  57232=>"101111101",
  57233=>"111010110",
  57234=>"011011110",
  57235=>"000011010",
  57236=>"101001010",
  57237=>"110101101",
  57238=>"011101000",
  57239=>"111000011",
  57240=>"101111111",
  57241=>"101110111",
  57242=>"111010111",
  57243=>"000110000",
  57244=>"001100001",
  57245=>"000010001",
  57246=>"011111011",
  57247=>"100110101",
  57248=>"110110000",
  57249=>"100110110",
  57250=>"011010111",
  57251=>"111101101",
  57252=>"011011001",
  57253=>"010110101",
  57254=>"110100000",
  57255=>"001101110",
  57256=>"000011001",
  57257=>"110111100",
  57258=>"100000001",
  57259=>"110000001",
  57260=>"000111000",
  57261=>"110011100",
  57262=>"011010010",
  57263=>"101101101",
  57264=>"101001101",
  57265=>"110001000",
  57266=>"111001101",
  57267=>"100110000",
  57268=>"001101000",
  57269=>"110111100",
  57270=>"001011011",
  57271=>"111000000",
  57272=>"000001011",
  57273=>"011101011",
  57274=>"110011010",
  57275=>"000000000",
  57276=>"110111101",
  57277=>"110110001",
  57278=>"000001111",
  57279=>"100001001",
  57280=>"000111000",
  57281=>"010111010",
  57282=>"001110101",
  57283=>"000000001",
  57284=>"011111010",
  57285=>"000000000",
  57286=>"010101111",
  57287=>"010101011",
  57288=>"101000001",
  57289=>"111111111",
  57290=>"001001101",
  57291=>"111111010",
  57292=>"101010110",
  57293=>"110011000",
  57294=>"110101110",
  57295=>"001011011",
  57296=>"011101111",
  57297=>"010011110",
  57298=>"100100110",
  57299=>"100011111",
  57300=>"100010101",
  57301=>"100001000",
  57302=>"110100111",
  57303=>"110000001",
  57304=>"100110011",
  57305=>"000011110",
  57306=>"100110001",
  57307=>"111000001",
  57308=>"111111110",
  57309=>"001000000",
  57310=>"100000001",
  57311=>"011000101",
  57312=>"101110111",
  57313=>"100111011",
  57314=>"010101100",
  57315=>"110100010",
  57316=>"101100100",
  57317=>"110000010",
  57318=>"101000111",
  57319=>"000001011",
  57320=>"011001111",
  57321=>"110011111",
  57322=>"111011101",
  57323=>"111101001",
  57324=>"010110010",
  57325=>"000001111",
  57326=>"110011000",
  57327=>"100100001",
  57328=>"111101110",
  57329=>"100111100",
  57330=>"100100111",
  57331=>"101110001",
  57332=>"011101110",
  57333=>"111000100",
  57334=>"110000101",
  57335=>"000011100",
  57336=>"000011000",
  57337=>"010100100",
  57338=>"011110010",
  57339=>"111111010",
  57340=>"111100011",
  57341=>"011010101",
  57342=>"011100001",
  57343=>"100000000",
  57344=>"110100000",
  57345=>"001001011",
  57346=>"010111110",
  57347=>"011010010",
  57348=>"010000011",
  57349=>"111101100",
  57350=>"011001101",
  57351=>"010010100",
  57352=>"010100101",
  57353=>"011100111",
  57354=>"011011000",
  57355=>"010111010",
  57356=>"000100110",
  57357=>"001001000",
  57358=>"111010110",
  57359=>"000010100",
  57360=>"100001011",
  57361=>"110110010",
  57362=>"101101010",
  57363=>"011101001",
  57364=>"000100000",
  57365=>"001101010",
  57366=>"000111000",
  57367=>"101000000",
  57368=>"110101011",
  57369=>"011111100",
  57370=>"101000101",
  57371=>"101000010",
  57372=>"000011100",
  57373=>"001110011",
  57374=>"101100100",
  57375=>"110010001",
  57376=>"110000001",
  57377=>"011100100",
  57378=>"111011011",
  57379=>"001000001",
  57380=>"111110011",
  57381=>"111101110",
  57382=>"011001111",
  57383=>"000111100",
  57384=>"101110011",
  57385=>"110101100",
  57386=>"101100101",
  57387=>"010111111",
  57388=>"010011110",
  57389=>"100111101",
  57390=>"100111100",
  57391=>"011111010",
  57392=>"100011111",
  57393=>"001001010",
  57394=>"111000000",
  57395=>"101000100",
  57396=>"111000100",
  57397=>"000001110",
  57398=>"010100110",
  57399=>"111110000",
  57400=>"001100001",
  57401=>"000000001",
  57402=>"110000101",
  57403=>"110000001",
  57404=>"011010000",
  57405=>"101100001",
  57406=>"010010001",
  57407=>"100110011",
  57408=>"010011101",
  57409=>"000011111",
  57410=>"100110100",
  57411=>"000110111",
  57412=>"111010000",
  57413=>"011011001",
  57414=>"101001000",
  57415=>"001011010",
  57416=>"000110111",
  57417=>"101110010",
  57418=>"111111100",
  57419=>"000010101",
  57420=>"101111101",
  57421=>"100111011",
  57422=>"101010000",
  57423=>"111111111",
  57424=>"101110100",
  57425=>"101110111",
  57426=>"101111001",
  57427=>"010110001",
  57428=>"100110110",
  57429=>"101100111",
  57430=>"000101010",
  57431=>"000010010",
  57432=>"101110110",
  57433=>"001100011",
  57434=>"111011110",
  57435=>"001100000",
  57436=>"000100000",
  57437=>"111011111",
  57438=>"000111000",
  57439=>"010101000",
  57440=>"111111000",
  57441=>"010001000",
  57442=>"010101000",
  57443=>"111001000",
  57444=>"010100101",
  57445=>"111001010",
  57446=>"001110010",
  57447=>"111011011",
  57448=>"111001001",
  57449=>"111101011",
  57450=>"101100100",
  57451=>"011100111",
  57452=>"010011001",
  57453=>"011100100",
  57454=>"110110000",
  57455=>"100010011",
  57456=>"010011110",
  57457=>"100000101",
  57458=>"110011111",
  57459=>"101110011",
  57460=>"011010010",
  57461=>"111001110",
  57462=>"001000101",
  57463=>"000101000",
  57464=>"111100001",
  57465=>"101011100",
  57466=>"010110010",
  57467=>"101001011",
  57468=>"010001000",
  57469=>"010010000",
  57470=>"000100010",
  57471=>"111000000",
  57472=>"010001000",
  57473=>"011000111",
  57474=>"000000001",
  57475=>"011100111",
  57476=>"011001011",
  57477=>"101101000",
  57478=>"100101011",
  57479=>"110000010",
  57480=>"110110001",
  57481=>"001001110",
  57482=>"000101010",
  57483=>"101101110",
  57484=>"011000111",
  57485=>"110000001",
  57486=>"001011000",
  57487=>"101001111",
  57488=>"101001001",
  57489=>"111110001",
  57490=>"000010100",
  57491=>"011110110",
  57492=>"000110101",
  57493=>"110000000",
  57494=>"101010111",
  57495=>"001011101",
  57496=>"010011101",
  57497=>"110001110",
  57498=>"010010110",
  57499=>"101101111",
  57500=>"001000101",
  57501=>"000100100",
  57502=>"000101100",
  57503=>"101011101",
  57504=>"010000100",
  57505=>"100010111",
  57506=>"110100110",
  57507=>"010000000",
  57508=>"011100111",
  57509=>"011010001",
  57510=>"101100110",
  57511=>"001110111",
  57512=>"010000101",
  57513=>"010110001",
  57514=>"100101010",
  57515=>"100011110",
  57516=>"010110000",
  57517=>"001100011",
  57518=>"100011100",
  57519=>"010101111",
  57520=>"110001001",
  57521=>"011111011",
  57522=>"101011001",
  57523=>"101111101",
  57524=>"100101100",
  57525=>"001000001",
  57526=>"110000010",
  57527=>"110100000",
  57528=>"111001100",
  57529=>"100111000",
  57530=>"011001000",
  57531=>"101000100",
  57532=>"100101001",
  57533=>"000011010",
  57534=>"110001111",
  57535=>"000001111",
  57536=>"000100110",
  57537=>"110111011",
  57538=>"000010000",
  57539=>"011001000",
  57540=>"101111110",
  57541=>"011101100",
  57542=>"000100000",
  57543=>"100001110",
  57544=>"000011000",
  57545=>"100000001",
  57546=>"100100110",
  57547=>"000111110",
  57548=>"111010110",
  57549=>"101111001",
  57550=>"010000011",
  57551=>"111001010",
  57552=>"010100111",
  57553=>"100110010",
  57554=>"000001100",
  57555=>"100101111",
  57556=>"011011001",
  57557=>"111011001",
  57558=>"100011010",
  57559=>"110010110",
  57560=>"100010010",
  57561=>"001011011",
  57562=>"000000010",
  57563=>"001001011",
  57564=>"101001101",
  57565=>"111001100",
  57566=>"011011001",
  57567=>"111101110",
  57568=>"001100000",
  57569=>"000001000",
  57570=>"100100100",
  57571=>"101110111",
  57572=>"000101011",
  57573=>"110110011",
  57574=>"000101010",
  57575=>"111111110",
  57576=>"011011011",
  57577=>"100111111",
  57578=>"011110010",
  57579=>"000110010",
  57580=>"001110101",
  57581=>"000010100",
  57582=>"010000101",
  57583=>"101101100",
  57584=>"111000011",
  57585=>"001001010",
  57586=>"000101000",
  57587=>"010110100",
  57588=>"101001010",
  57589=>"000000100",
  57590=>"101111110",
  57591=>"100001101",
  57592=>"101000011",
  57593=>"010001101",
  57594=>"101010000",
  57595=>"001101000",
  57596=>"110011110",
  57597=>"110010010",
  57598=>"010111011",
  57599=>"000111101",
  57600=>"011110011",
  57601=>"010000010",
  57602=>"111100111",
  57603=>"001011111",
  57604=>"011010000",
  57605=>"000000110",
  57606=>"100010000",
  57607=>"101000100",
  57608=>"111000110",
  57609=>"100011000",
  57610=>"111001101",
  57611=>"010111100",
  57612=>"111000111",
  57613=>"010011111",
  57614=>"110011000",
  57615=>"101100001",
  57616=>"100000011",
  57617=>"011000000",
  57618=>"001111011",
  57619=>"101011101",
  57620=>"010101001",
  57621=>"100100000",
  57622=>"111101111",
  57623=>"001101101",
  57624=>"111111101",
  57625=>"110000111",
  57626=>"100001000",
  57627=>"001010101",
  57628=>"010010010",
  57629=>"111001110",
  57630=>"101101001",
  57631=>"011001101",
  57632=>"000101100",
  57633=>"011001110",
  57634=>"110000010",
  57635=>"100011010",
  57636=>"011110011",
  57637=>"000011100",
  57638=>"101101001",
  57639=>"111000111",
  57640=>"000100100",
  57641=>"110111110",
  57642=>"010100101",
  57643=>"101101011",
  57644=>"010100001",
  57645=>"110110010",
  57646=>"001101000",
  57647=>"111110101",
  57648=>"001000101",
  57649=>"110011010",
  57650=>"111110100",
  57651=>"101010010",
  57652=>"100000101",
  57653=>"101001100",
  57654=>"010111000",
  57655=>"110011101",
  57656=>"000110000",
  57657=>"101101111",
  57658=>"001101111",
  57659=>"000000010",
  57660=>"110010101",
  57661=>"001101110",
  57662=>"101010000",
  57663=>"001001101",
  57664=>"010100001",
  57665=>"110100100",
  57666=>"100011101",
  57667=>"101101100",
  57668=>"000100100",
  57669=>"111010010",
  57670=>"010001000",
  57671=>"110010011",
  57672=>"101101110",
  57673=>"110101100",
  57674=>"000100100",
  57675=>"001101011",
  57676=>"000001000",
  57677=>"010000110",
  57678=>"111100100",
  57679=>"010010001",
  57680=>"011010001",
  57681=>"110110111",
  57682=>"101110010",
  57683=>"110000111",
  57684=>"010100001",
  57685=>"110011110",
  57686=>"010100000",
  57687=>"001011100",
  57688=>"001001100",
  57689=>"101001001",
  57690=>"000110101",
  57691=>"001010100",
  57692=>"000011000",
  57693=>"111110111",
  57694=>"001000010",
  57695=>"000111101",
  57696=>"001100010",
  57697=>"011000011",
  57698=>"111101000",
  57699=>"111000010",
  57700=>"010100000",
  57701=>"100101010",
  57702=>"010110000",
  57703=>"100111010",
  57704=>"000111001",
  57705=>"111011010",
  57706=>"101011001",
  57707=>"100110010",
  57708=>"011010110",
  57709=>"001111010",
  57710=>"001000000",
  57711=>"100110011",
  57712=>"111011001",
  57713=>"101001011",
  57714=>"011100101",
  57715=>"011101110",
  57716=>"011011110",
  57717=>"111111000",
  57718=>"101100001",
  57719=>"111000111",
  57720=>"101111100",
  57721=>"110000111",
  57722=>"111111110",
  57723=>"110001001",
  57724=>"100111110",
  57725=>"001001000",
  57726=>"111000001",
  57727=>"001100001",
  57728=>"101011100",
  57729=>"111110010",
  57730=>"001000101",
  57731=>"000101001",
  57732=>"000100011",
  57733=>"000010111",
  57734=>"010111011",
  57735=>"111101011",
  57736=>"111000101",
  57737=>"101000110",
  57738=>"111101001",
  57739=>"001011001",
  57740=>"010000100",
  57741=>"010010100",
  57742=>"111100000",
  57743=>"010010001",
  57744=>"110001000",
  57745=>"101101111",
  57746=>"100001110",
  57747=>"101101101",
  57748=>"011100110",
  57749=>"100000111",
  57750=>"000101011",
  57751=>"100010011",
  57752=>"001100100",
  57753=>"011100110",
  57754=>"000001101",
  57755=>"100011001",
  57756=>"000010010",
  57757=>"011000100",
  57758=>"101010001",
  57759=>"000000111",
  57760=>"110010010",
  57761=>"010010111",
  57762=>"101100000",
  57763=>"001001100",
  57764=>"100010011",
  57765=>"010000001",
  57766=>"010011011",
  57767=>"101000001",
  57768=>"111010001",
  57769=>"101001110",
  57770=>"000101101",
  57771=>"110001101",
  57772=>"001111000",
  57773=>"011111101",
  57774=>"111001111",
  57775=>"100001000",
  57776=>"010000001",
  57777=>"100011100",
  57778=>"111111100",
  57779=>"000111001",
  57780=>"000111100",
  57781=>"110010010",
  57782=>"100111101",
  57783=>"001101101",
  57784=>"000101010",
  57785=>"011110101",
  57786=>"011010111",
  57787=>"100011001",
  57788=>"000000000",
  57789=>"010001111",
  57790=>"000101100",
  57791=>"100010001",
  57792=>"000011010",
  57793=>"111100010",
  57794=>"010000101",
  57795=>"011000000",
  57796=>"001001001",
  57797=>"111110001",
  57798=>"010100101",
  57799=>"101100010",
  57800=>"101111110",
  57801=>"010000100",
  57802=>"100001000",
  57803=>"100011001",
  57804=>"110110110",
  57805=>"011010111",
  57806=>"100011010",
  57807=>"010100011",
  57808=>"111010001",
  57809=>"111110111",
  57810=>"101100011",
  57811=>"001011000",
  57812=>"101001010",
  57813=>"111001100",
  57814=>"010000011",
  57815=>"111011001",
  57816=>"111011001",
  57817=>"010001011",
  57818=>"111001111",
  57819=>"010010000",
  57820=>"100100101",
  57821=>"100011101",
  57822=>"011011000",
  57823=>"000000101",
  57824=>"011111000",
  57825=>"101111010",
  57826=>"100000100",
  57827=>"001100110",
  57828=>"001101000",
  57829=>"011100011",
  57830=>"000010000",
  57831=>"010001100",
  57832=>"011110000",
  57833=>"111110111",
  57834=>"000000110",
  57835=>"011000010",
  57836=>"000001111",
  57837=>"100101000",
  57838=>"000100000",
  57839=>"100110000",
  57840=>"010111001",
  57841=>"101010010",
  57842=>"000100110",
  57843=>"001110101",
  57844=>"000101101",
  57845=>"111101110",
  57846=>"110010101",
  57847=>"100101101",
  57848=>"100011100",
  57849=>"100110111",
  57850=>"010100000",
  57851=>"101111101",
  57852=>"010110100",
  57853=>"100101000",
  57854=>"101111011",
  57855=>"101111110",
  57856=>"100001001",
  57857=>"010010111",
  57858=>"101010100",
  57859=>"111100111",
  57860=>"011010000",
  57861=>"010000001",
  57862=>"100101101",
  57863=>"110010001",
  57864=>"101100001",
  57865=>"001101101",
  57866=>"011011110",
  57867=>"101101000",
  57868=>"000001001",
  57869=>"100011000",
  57870=>"110010111",
  57871=>"101100000",
  57872=>"010000011",
  57873=>"011011101",
  57874=>"000010011",
  57875=>"000010110",
  57876=>"000000111",
  57877=>"110001101",
  57878=>"010111000",
  57879=>"010100100",
  57880=>"101111001",
  57881=>"110100101",
  57882=>"000010000",
  57883=>"010010001",
  57884=>"100110000",
  57885=>"000011011",
  57886=>"011001100",
  57887=>"110111110",
  57888=>"101011001",
  57889=>"101111110",
  57890=>"101110111",
  57891=>"010001011",
  57892=>"101110010",
  57893=>"010100000",
  57894=>"100101010",
  57895=>"101111111",
  57896=>"100001010",
  57897=>"101001100",
  57898=>"000000110",
  57899=>"001101001",
  57900=>"010011100",
  57901=>"100000010",
  57902=>"100010001",
  57903=>"111000101",
  57904=>"001000001",
  57905=>"111011101",
  57906=>"100011110",
  57907=>"000011000",
  57908=>"001001001",
  57909=>"010001111",
  57910=>"111100001",
  57911=>"000110000",
  57912=>"101000111",
  57913=>"111001101",
  57914=>"100111100",
  57915=>"000100001",
  57916=>"110101000",
  57917=>"000010010",
  57918=>"111111011",
  57919=>"010010101",
  57920=>"000000100",
  57921=>"010111000",
  57922=>"100110001",
  57923=>"011001010",
  57924=>"101011000",
  57925=>"101110100",
  57926=>"110111111",
  57927=>"101100100",
  57928=>"011110000",
  57929=>"001000000",
  57930=>"100101001",
  57931=>"111100001",
  57932=>"010001111",
  57933=>"001110100",
  57934=>"000010010",
  57935=>"100100000",
  57936=>"110111111",
  57937=>"000001111",
  57938=>"100010111",
  57939=>"110000011",
  57940=>"110110011",
  57941=>"110110000",
  57942=>"111101001",
  57943=>"011100010",
  57944=>"011110100",
  57945=>"010001010",
  57946=>"111110110",
  57947=>"111101010",
  57948=>"011000100",
  57949=>"100101100",
  57950=>"100001011",
  57951=>"011111001",
  57952=>"100011010",
  57953=>"100010000",
  57954=>"011010000",
  57955=>"100100100",
  57956=>"001000101",
  57957=>"110101101",
  57958=>"001011100",
  57959=>"101110110",
  57960=>"101000000",
  57961=>"101000011",
  57962=>"000111010",
  57963=>"100000111",
  57964=>"001110100",
  57965=>"101100001",
  57966=>"111110010",
  57967=>"001110110",
  57968=>"100011000",
  57969=>"000100011",
  57970=>"101101101",
  57971=>"110001100",
  57972=>"011111101",
  57973=>"000010101",
  57974=>"100000100",
  57975=>"010111100",
  57976=>"001101010",
  57977=>"111111100",
  57978=>"010100110",
  57979=>"100111100",
  57980=>"011101010",
  57981=>"010010100",
  57982=>"101101111",
  57983=>"000011001",
  57984=>"111010000",
  57985=>"000111110",
  57986=>"001100000",
  57987=>"010011111",
  57988=>"001011101",
  57989=>"111111110",
  57990=>"011000000",
  57991=>"101000011",
  57992=>"000100000",
  57993=>"011001110",
  57994=>"001010011",
  57995=>"000001000",
  57996=>"110101100",
  57997=>"001111000",
  57998=>"100010100",
  57999=>"110100010",
  58000=>"101000111",
  58001=>"001010101",
  58002=>"110001111",
  58003=>"111010010",
  58004=>"010010100",
  58005=>"101110100",
  58006=>"010010000",
  58007=>"100111011",
  58008=>"001101001",
  58009=>"000111101",
  58010=>"001010000",
  58011=>"110001011",
  58012=>"101111111",
  58013=>"111111010",
  58014=>"010010010",
  58015=>"110011000",
  58016=>"001110001",
  58017=>"010101100",
  58018=>"000001011",
  58019=>"111011111",
  58020=>"011100011",
  58021=>"111010011",
  58022=>"110101101",
  58023=>"001101111",
  58024=>"110010101",
  58025=>"011100100",
  58026=>"110101011",
  58027=>"110100110",
  58028=>"101100001",
  58029=>"101001011",
  58030=>"101100011",
  58031=>"100001100",
  58032=>"010011011",
  58033=>"000001111",
  58034=>"110011010",
  58035=>"101011100",
  58036=>"000110111",
  58037=>"011001100",
  58038=>"011100100",
  58039=>"010100100",
  58040=>"010111010",
  58041=>"011010111",
  58042=>"011011001",
  58043=>"000001100",
  58044=>"010111011",
  58045=>"011010000",
  58046=>"001001010",
  58047=>"101000110",
  58048=>"110010001",
  58049=>"110110010",
  58050=>"000111001",
  58051=>"101010000",
  58052=>"101010000",
  58053=>"000010000",
  58054=>"110101000",
  58055=>"100011001",
  58056=>"111110110",
  58057=>"010011000",
  58058=>"110011111",
  58059=>"000111111",
  58060=>"000000100",
  58061=>"111110011",
  58062=>"001011011",
  58063=>"000111010",
  58064=>"111101100",
  58065=>"101110111",
  58066=>"110010011",
  58067=>"011010110",
  58068=>"101101011",
  58069=>"110000000",
  58070=>"011010000",
  58071=>"011100010",
  58072=>"001000101",
  58073=>"011001111",
  58074=>"011100011",
  58075=>"000001001",
  58076=>"101100001",
  58077=>"011101001",
  58078=>"111101110",
  58079=>"000010100",
  58080=>"001000100",
  58081=>"001001111",
  58082=>"111111000",
  58083=>"101011110",
  58084=>"101011010",
  58085=>"101010100",
  58086=>"010110011",
  58087=>"101101000",
  58088=>"101101111",
  58089=>"011011100",
  58090=>"011101111",
  58091=>"110110001",
  58092=>"000000011",
  58093=>"100000101",
  58094=>"110100111",
  58095=>"001001110",
  58096=>"111110011",
  58097=>"011101010",
  58098=>"011001110",
  58099=>"111011101",
  58100=>"100011010",
  58101=>"110110101",
  58102=>"000011110",
  58103=>"111110001",
  58104=>"001110101",
  58105=>"010100110",
  58106=>"110001100",
  58107=>"100111001",
  58108=>"100110000",
  58109=>"101110101",
  58110=>"110010111",
  58111=>"100011000",
  58112=>"000100000",
  58113=>"001100000",
  58114=>"001011111",
  58115=>"001010101",
  58116=>"000101011",
  58117=>"000000011",
  58118=>"011010101",
  58119=>"000011111",
  58120=>"011011000",
  58121=>"011011111",
  58122=>"110010100",
  58123=>"111011111",
  58124=>"010101100",
  58125=>"110011001",
  58126=>"101000110",
  58127=>"100010000",
  58128=>"000100100",
  58129=>"110000001",
  58130=>"010101111",
  58131=>"100001101",
  58132=>"000010101",
  58133=>"100110001",
  58134=>"110000111",
  58135=>"110010110",
  58136=>"010010000",
  58137=>"100000111",
  58138=>"011000000",
  58139=>"000001110",
  58140=>"000000111",
  58141=>"110111110",
  58142=>"000010000",
  58143=>"011000011",
  58144=>"000010011",
  58145=>"001010111",
  58146=>"101101100",
  58147=>"011101001",
  58148=>"100011000",
  58149=>"001101101",
  58150=>"100101001",
  58151=>"111100001",
  58152=>"101101101",
  58153=>"010101000",
  58154=>"000000110",
  58155=>"001110110",
  58156=>"101111100",
  58157=>"010000001",
  58158=>"001001001",
  58159=>"001011000",
  58160=>"100010001",
  58161=>"101110100",
  58162=>"111101111",
  58163=>"101000100",
  58164=>"010110001",
  58165=>"100101110",
  58166=>"001100100",
  58167=>"101001110",
  58168=>"101010110",
  58169=>"100111101",
  58170=>"100000100",
  58171=>"010111101",
  58172=>"010001000",
  58173=>"110110010",
  58174=>"010100011",
  58175=>"010011100",
  58176=>"011110110",
  58177=>"001011101",
  58178=>"011001010",
  58179=>"100000101",
  58180=>"011001011",
  58181=>"111110100",
  58182=>"000000101",
  58183=>"010011100",
  58184=>"110011101",
  58185=>"111011011",
  58186=>"010001001",
  58187=>"110101101",
  58188=>"000010000",
  58189=>"010001001",
  58190=>"010101011",
  58191=>"110100100",
  58192=>"011011001",
  58193=>"001011010",
  58194=>"111100111",
  58195=>"110010000",
  58196=>"000011000",
  58197=>"000001000",
  58198=>"100001101",
  58199=>"110011000",
  58200=>"011111111",
  58201=>"101110110",
  58202=>"101001101",
  58203=>"111010011",
  58204=>"101110000",
  58205=>"111000111",
  58206=>"101101111",
  58207=>"101110101",
  58208=>"010011111",
  58209=>"110011000",
  58210=>"110011110",
  58211=>"101100001",
  58212=>"101100011",
  58213=>"011101100",
  58214=>"001001100",
  58215=>"001010011",
  58216=>"010101111",
  58217=>"001010001",
  58218=>"101010111",
  58219=>"111101101",
  58220=>"110001110",
  58221=>"011111010",
  58222=>"100000010",
  58223=>"110100101",
  58224=>"100000101",
  58225=>"111110101",
  58226=>"100101100",
  58227=>"011001110",
  58228=>"100110101",
  58229=>"000110010",
  58230=>"010011011",
  58231=>"010000100",
  58232=>"011101001",
  58233=>"100100111",
  58234=>"101000111",
  58235=>"010011010",
  58236=>"000001000",
  58237=>"001100111",
  58238=>"001111011",
  58239=>"000011110",
  58240=>"001100100",
  58241=>"000000001",
  58242=>"101001111",
  58243=>"000011000",
  58244=>"010100111",
  58245=>"001111100",
  58246=>"101010101",
  58247=>"010000101",
  58248=>"010100100",
  58249=>"110101111",
  58250=>"010111000",
  58251=>"000111010",
  58252=>"100111110",
  58253=>"011110111",
  58254=>"110100101",
  58255=>"101111111",
  58256=>"101000001",
  58257=>"000000011",
  58258=>"001000101",
  58259=>"111111000",
  58260=>"001111011",
  58261=>"101010011",
  58262=>"011101000",
  58263=>"000001100",
  58264=>"000001001",
  58265=>"101101101",
  58266=>"110110001",
  58267=>"011000111",
  58268=>"000000001",
  58269=>"100011111",
  58270=>"011010000",
  58271=>"100110011",
  58272=>"010111011",
  58273=>"001111001",
  58274=>"011010000",
  58275=>"111111110",
  58276=>"011000010",
  58277=>"111010011",
  58278=>"101111000",
  58279=>"100010010",
  58280=>"000001101",
  58281=>"110100100",
  58282=>"000100101",
  58283=>"011011100",
  58284=>"000000110",
  58285=>"010111110",
  58286=>"011010100",
  58287=>"111101011",
  58288=>"011110110",
  58289=>"100111111",
  58290=>"100010110",
  58291=>"010001111",
  58292=>"110000001",
  58293=>"010110010",
  58294=>"010110100",
  58295=>"110010011",
  58296=>"101101011",
  58297=>"100011001",
  58298=>"001111000",
  58299=>"010100101",
  58300=>"000011000",
  58301=>"001111111",
  58302=>"001010100",
  58303=>"000011010",
  58304=>"001110011",
  58305=>"000111101",
  58306=>"000101110",
  58307=>"100101010",
  58308=>"000001000",
  58309=>"001011000",
  58310=>"001111000",
  58311=>"010010001",
  58312=>"000010011",
  58313=>"111010110",
  58314=>"100000011",
  58315=>"111110110",
  58316=>"110110111",
  58317=>"100100011",
  58318=>"001000010",
  58319=>"111110101",
  58320=>"101010111",
  58321=>"010000111",
  58322=>"111000101",
  58323=>"000010000",
  58324=>"101001110",
  58325=>"101000111",
  58326=>"101011111",
  58327=>"010000001",
  58328=>"110001100",
  58329=>"011111101",
  58330=>"110111101",
  58331=>"001000100",
  58332=>"000100001",
  58333=>"001110000",
  58334=>"111111010",
  58335=>"111001100",
  58336=>"101111001",
  58337=>"100000111",
  58338=>"101111100",
  58339=>"000101111",
  58340=>"000100000",
  58341=>"000010010",
  58342=>"100111110",
  58343=>"001011011",
  58344=>"010000100",
  58345=>"101000110",
  58346=>"110100110",
  58347=>"001001111",
  58348=>"101000110",
  58349=>"011001000",
  58350=>"111100110",
  58351=>"010011110",
  58352=>"101010010",
  58353=>"101101100",
  58354=>"110001000",
  58355=>"001000001",
  58356=>"100001101",
  58357=>"011000001",
  58358=>"110010100",
  58359=>"111001100",
  58360=>"110100000",
  58361=>"011101111",
  58362=>"000001111",
  58363=>"000101110",
  58364=>"101000001",
  58365=>"000101111",
  58366=>"000001010",
  58367=>"011011100",
  58368=>"100001001",
  58369=>"111100000",
  58370=>"101111110",
  58371=>"110101000",
  58372=>"101111111",
  58373=>"110101110",
  58374=>"000111111",
  58375=>"110110010",
  58376=>"111011010",
  58377=>"001110101",
  58378=>"010111011",
  58379=>"010111101",
  58380=>"000011000",
  58381=>"001111110",
  58382=>"011101010",
  58383=>"100101000",
  58384=>"101010111",
  58385=>"000000101",
  58386=>"101111110",
  58387=>"110000011",
  58388=>"010011111",
  58389=>"011101011",
  58390=>"110010111",
  58391=>"101000101",
  58392=>"010110100",
  58393=>"110110010",
  58394=>"000000110",
  58395=>"100110010",
  58396=>"101000111",
  58397=>"011001001",
  58398=>"001100010",
  58399=>"000000011",
  58400=>"011010101",
  58401=>"001000110",
  58402=>"111001111",
  58403=>"010000100",
  58404=>"010101111",
  58405=>"100100100",
  58406=>"011101100",
  58407=>"100100101",
  58408=>"110101000",
  58409=>"110100101",
  58410=>"111100101",
  58411=>"110010101",
  58412=>"011010001",
  58413=>"111001001",
  58414=>"011101111",
  58415=>"101101010",
  58416=>"110101011",
  58417=>"110011000",
  58418=>"001100111",
  58419=>"010111000",
  58420=>"111100110",
  58421=>"000101101",
  58422=>"000000010",
  58423=>"010000010",
  58424=>"111101011",
  58425=>"110001111",
  58426=>"101011111",
  58427=>"111100000",
  58428=>"000110101",
  58429=>"110110111",
  58430=>"000010111",
  58431=>"011111101",
  58432=>"101111111",
  58433=>"010001101",
  58434=>"011100111",
  58435=>"100000110",
  58436=>"011101011",
  58437=>"101101001",
  58438=>"111100101",
  58439=>"000110100",
  58440=>"001001000",
  58441=>"001011111",
  58442=>"100010100",
  58443=>"111001100",
  58444=>"100011111",
  58445=>"100110101",
  58446=>"010010111",
  58447=>"001101000",
  58448=>"011110110",
  58449=>"100110101",
  58450=>"111010010",
  58451=>"111110100",
  58452=>"101011011",
  58453=>"101011100",
  58454=>"101010110",
  58455=>"011011111",
  58456=>"111001101",
  58457=>"000001001",
  58458=>"111110111",
  58459=>"000100111",
  58460=>"001110100",
  58461=>"010100001",
  58462=>"111101111",
  58463=>"000001010",
  58464=>"000100101",
  58465=>"110111100",
  58466=>"001100010",
  58467=>"000101111",
  58468=>"111001000",
  58469=>"001001001",
  58470=>"101010110",
  58471=>"000111100",
  58472=>"001011001",
  58473=>"101110100",
  58474=>"111001001",
  58475=>"111010101",
  58476=>"110100010",
  58477=>"100100110",
  58478=>"110010101",
  58479=>"000011000",
  58480=>"010101000",
  58481=>"111101101",
  58482=>"111110011",
  58483=>"101011000",
  58484=>"100011001",
  58485=>"100100100",
  58486=>"101100101",
  58487=>"001000010",
  58488=>"011010000",
  58489=>"011011011",
  58490=>"000101110",
  58491=>"011001000",
  58492=>"011111100",
  58493=>"010001011",
  58494=>"010000111",
  58495=>"011111010",
  58496=>"101000010",
  58497=>"100100011",
  58498=>"100001111",
  58499=>"001101101",
  58500=>"100001110",
  58501=>"001110010",
  58502=>"010101011",
  58503=>"000101010",
  58504=>"001110101",
  58505=>"010110000",
  58506=>"111100111",
  58507=>"110111100",
  58508=>"111001100",
  58509=>"111110100",
  58510=>"001111011",
  58511=>"110001010",
  58512=>"000100101",
  58513=>"001100010",
  58514=>"000010100",
  58515=>"001110001",
  58516=>"000100111",
  58517=>"110000010",
  58518=>"000011000",
  58519=>"100110100",
  58520=>"001111010",
  58521=>"111110010",
  58522=>"101000101",
  58523=>"111101111",
  58524=>"111100101",
  58525=>"100100110",
  58526=>"100010010",
  58527=>"000010001",
  58528=>"011000110",
  58529=>"101110001",
  58530=>"100011101",
  58531=>"101111011",
  58532=>"100100100",
  58533=>"100111001",
  58534=>"011101110",
  58535=>"001010110",
  58536=>"000001111",
  58537=>"001010101",
  58538=>"001100001",
  58539=>"101001000",
  58540=>"001110111",
  58541=>"001100100",
  58542=>"101101000",
  58543=>"001001000",
  58544=>"000100101",
  58545=>"101010011",
  58546=>"010010011",
  58547=>"110000101",
  58548=>"100100000",
  58549=>"000000110",
  58550=>"111111100",
  58551=>"010010010",
  58552=>"101110111",
  58553=>"110100111",
  58554=>"110101011",
  58555=>"101111110",
  58556=>"100001100",
  58557=>"000010010",
  58558=>"000010110",
  58559=>"001000000",
  58560=>"110000000",
  58561=>"010100100",
  58562=>"110101111",
  58563=>"011111010",
  58564=>"111101010",
  58565=>"100001111",
  58566=>"011101110",
  58567=>"011101111",
  58568=>"011011011",
  58569=>"111110000",
  58570=>"100101001",
  58571=>"001110100",
  58572=>"010000000",
  58573=>"001110101",
  58574=>"001000100",
  58575=>"010000001",
  58576=>"011110101",
  58577=>"111110010",
  58578=>"101111001",
  58579=>"110111101",
  58580=>"110000010",
  58581=>"100011010",
  58582=>"101100010",
  58583=>"100110101",
  58584=>"111011011",
  58585=>"001101000",
  58586=>"101101011",
  58587=>"010100111",
  58588=>"001000100",
  58589=>"110101001",
  58590=>"000010010",
  58591=>"001011010",
  58592=>"000111001",
  58593=>"110111010",
  58594=>"000010001",
  58595=>"100110110",
  58596=>"111110000",
  58597=>"100000010",
  58598=>"010011111",
  58599=>"011010001",
  58600=>"011000101",
  58601=>"000001000",
  58602=>"011111000",
  58603=>"001010000",
  58604=>"011110000",
  58605=>"011010010",
  58606=>"011001110",
  58607=>"011101001",
  58608=>"111110010",
  58609=>"001100001",
  58610=>"010110000",
  58611=>"101110001",
  58612=>"101100000",
  58613=>"100001110",
  58614=>"101001000",
  58615=>"000010011",
  58616=>"011110100",
  58617=>"010010100",
  58618=>"100110011",
  58619=>"010000101",
  58620=>"101001010",
  58621=>"110001000",
  58622=>"000000000",
  58623=>"111100000",
  58624=>"000110011",
  58625=>"101010111",
  58626=>"000001010",
  58627=>"000110001",
  58628=>"011100110",
  58629=>"110010000",
  58630=>"001001111",
  58631=>"100101100",
  58632=>"101000011",
  58633=>"100101011",
  58634=>"001111010",
  58635=>"101010100",
  58636=>"110110111",
  58637=>"100111001",
  58638=>"101000001",
  58639=>"000001100",
  58640=>"101111000",
  58641=>"100101101",
  58642=>"110111010",
  58643=>"110010111",
  58644=>"101110111",
  58645=>"000001100",
  58646=>"100101101",
  58647=>"111101100",
  58648=>"011000100",
  58649=>"001110010",
  58650=>"100100000",
  58651=>"111110101",
  58652=>"111001111",
  58653=>"110000000",
  58654=>"001111110",
  58655=>"001001000",
  58656=>"011111010",
  58657=>"000011100",
  58658=>"000001011",
  58659=>"111001101",
  58660=>"001111011",
  58661=>"010010001",
  58662=>"100100100",
  58663=>"001011000",
  58664=>"111010000",
  58665=>"010101011",
  58666=>"101110111",
  58667=>"011000000",
  58668=>"101100011",
  58669=>"111001111",
  58670=>"010011101",
  58671=>"100011111",
  58672=>"010000111",
  58673=>"101110110",
  58674=>"000000100",
  58675=>"001011010",
  58676=>"110010100",
  58677=>"010001111",
  58678=>"010101100",
  58679=>"010100101",
  58680=>"001011010",
  58681=>"101100001",
  58682=>"111000111",
  58683=>"010111101",
  58684=>"110100101",
  58685=>"001111000",
  58686=>"111111010",
  58687=>"111010001",
  58688=>"111011001",
  58689=>"111101101",
  58690=>"000110101",
  58691=>"110000001",
  58692=>"100100110",
  58693=>"110001001",
  58694=>"011000110",
  58695=>"110111001",
  58696=>"001000110",
  58697=>"011100011",
  58698=>"110100011",
  58699=>"010101111",
  58700=>"001111010",
  58701=>"000011010",
  58702=>"111101001",
  58703=>"011011011",
  58704=>"011001100",
  58705=>"111101101",
  58706=>"101011110",
  58707=>"101101011",
  58708=>"100011101",
  58709=>"110000001",
  58710=>"100101111",
  58711=>"000000101",
  58712=>"101111000",
  58713=>"101010111",
  58714=>"001001011",
  58715=>"100110010",
  58716=>"101011001",
  58717=>"100011111",
  58718=>"100000000",
  58719=>"100011100",
  58720=>"011101100",
  58721=>"000110011",
  58722=>"000100010",
  58723=>"111000111",
  58724=>"001011010",
  58725=>"010101100",
  58726=>"011111011",
  58727=>"010111001",
  58728=>"010000111",
  58729=>"111110000",
  58730=>"010110101",
  58731=>"111011000",
  58732=>"001011100",
  58733=>"100101000",
  58734=>"001010111",
  58735=>"110110111",
  58736=>"011001000",
  58737=>"110101000",
  58738=>"000010110",
  58739=>"111101000",
  58740=>"000101101",
  58741=>"000110110",
  58742=>"000001000",
  58743=>"100101010",
  58744=>"000011011",
  58745=>"001101100",
  58746=>"000000101",
  58747=>"100101001",
  58748=>"100010100",
  58749=>"101100000",
  58750=>"111001101",
  58751=>"100101100",
  58752=>"100011011",
  58753=>"010111000",
  58754=>"111110100",
  58755=>"110110100",
  58756=>"001111100",
  58757=>"100100101",
  58758=>"110110001",
  58759=>"010100011",
  58760=>"010011111",
  58761=>"111101100",
  58762=>"000010001",
  58763=>"101100111",
  58764=>"100101100",
  58765=>"111100101",
  58766=>"111100011",
  58767=>"011010000",
  58768=>"010100001",
  58769=>"011010001",
  58770=>"000010111",
  58771=>"110011000",
  58772=>"010000001",
  58773=>"101010011",
  58774=>"110110111",
  58775=>"100111010",
  58776=>"000101111",
  58777=>"111110101",
  58778=>"100111100",
  58779=>"101010111",
  58780=>"101001100",
  58781=>"011111010",
  58782=>"011111010",
  58783=>"000111101",
  58784=>"100001101",
  58785=>"110010111",
  58786=>"010001001",
  58787=>"101110110",
  58788=>"111110001",
  58789=>"000010101",
  58790=>"001001101",
  58791=>"001000101",
  58792=>"100110100",
  58793=>"110111100",
  58794=>"010101000",
  58795=>"100001100",
  58796=>"100100110",
  58797=>"100100000",
  58798=>"110011001",
  58799=>"101000001",
  58800=>"001101000",
  58801=>"101100000",
  58802=>"100001001",
  58803=>"110111111",
  58804=>"110001011",
  58805=>"100111001",
  58806=>"110101010",
  58807=>"110101111",
  58808=>"001111011",
  58809=>"100101001",
  58810=>"000011011",
  58811=>"100000000",
  58812=>"001100100",
  58813=>"011011111",
  58814=>"100010110",
  58815=>"011010111",
  58816=>"000011000",
  58817=>"111010001",
  58818=>"010010101",
  58819=>"000101110",
  58820=>"000100111",
  58821=>"000011111",
  58822=>"111110000",
  58823=>"001011010",
  58824=>"000011001",
  58825=>"011110110",
  58826=>"111000000",
  58827=>"101011000",
  58828=>"001111011",
  58829=>"000101101",
  58830=>"101011001",
  58831=>"100001010",
  58832=>"101111100",
  58833=>"110110000",
  58834=>"100001010",
  58835=>"010100001",
  58836=>"000110100",
  58837=>"000100011",
  58838=>"100111100",
  58839=>"000010000",
  58840=>"001011101",
  58841=>"101010111",
  58842=>"110111010",
  58843=>"101001111",
  58844=>"101000111",
  58845=>"001011100",
  58846=>"011111100",
  58847=>"100110010",
  58848=>"010010001",
  58849=>"010100000",
  58850=>"010001010",
  58851=>"110000000",
  58852=>"110010110",
  58853=>"001000110",
  58854=>"011100010",
  58855=>"001000010",
  58856=>"010011010",
  58857=>"111101000",
  58858=>"101000001",
  58859=>"011100011",
  58860=>"100100011",
  58861=>"001011010",
  58862=>"001100000",
  58863=>"101111011",
  58864=>"100000010",
  58865=>"001101000",
  58866=>"111010000",
  58867=>"000000100",
  58868=>"000010000",
  58869=>"011101001",
  58870=>"001000001",
  58871=>"001100100",
  58872=>"100001001",
  58873=>"110001011",
  58874=>"010011011",
  58875=>"100101111",
  58876=>"111100111",
  58877=>"111001111",
  58878=>"110110110",
  58879=>"110101000",
  58880=>"100010000",
  58881=>"000101111",
  58882=>"011100001",
  58883=>"001001111",
  58884=>"111101011",
  58885=>"100110111",
  58886=>"011111100",
  58887=>"101011111",
  58888=>"011001111",
  58889=>"100001101",
  58890=>"100110100",
  58891=>"111100001",
  58892=>"000110111",
  58893=>"110110100",
  58894=>"100000110",
  58895=>"000100001",
  58896=>"101111110",
  58897=>"000001111",
  58898=>"101011011",
  58899=>"011010001",
  58900=>"101110010",
  58901=>"001100000",
  58902=>"000110111",
  58903=>"100101110",
  58904=>"100101101",
  58905=>"101010110",
  58906=>"110110010",
  58907=>"100111111",
  58908=>"110001011",
  58909=>"100101111",
  58910=>"000010100",
  58911=>"011101010",
  58912=>"001000000",
  58913=>"010110000",
  58914=>"010010010",
  58915=>"101000111",
  58916=>"001001000",
  58917=>"001010000",
  58918=>"011010011",
  58919=>"110011000",
  58920=>"111010101",
  58921=>"010001011",
  58922=>"100110000",
  58923=>"101000100",
  58924=>"001010010",
  58925=>"010000111",
  58926=>"111110010",
  58927=>"110111010",
  58928=>"101111010",
  58929=>"000111100",
  58930=>"010000110",
  58931=>"001110111",
  58932=>"011011011",
  58933=>"000110001",
  58934=>"011001011",
  58935=>"000001111",
  58936=>"101000000",
  58937=>"000111000",
  58938=>"000111100",
  58939=>"100110010",
  58940=>"101110101",
  58941=>"101010011",
  58942=>"000000001",
  58943=>"001101101",
  58944=>"110010011",
  58945=>"001000000",
  58946=>"011000101",
  58947=>"010000010",
  58948=>"010101000",
  58949=>"001111111",
  58950=>"111010001",
  58951=>"111001011",
  58952=>"010001000",
  58953=>"110001001",
  58954=>"001010110",
  58955=>"100111100",
  58956=>"010101101",
  58957=>"101101011",
  58958=>"111111101",
  58959=>"111011011",
  58960=>"011110101",
  58961=>"000001101",
  58962=>"100100100",
  58963=>"100110111",
  58964=>"100111001",
  58965=>"111111101",
  58966=>"110111000",
  58967=>"010110111",
  58968=>"111011000",
  58969=>"110100100",
  58970=>"111110100",
  58971=>"001100101",
  58972=>"000001001",
  58973=>"011111000",
  58974=>"101101001",
  58975=>"101000001",
  58976=>"101001000",
  58977=>"001101001",
  58978=>"000101110",
  58979=>"001011010",
  58980=>"110001100",
  58981=>"101000100",
  58982=>"000100110",
  58983=>"111111010",
  58984=>"011011001",
  58985=>"010000010",
  58986=>"111101110",
  58987=>"100001101",
  58988=>"001001011",
  58989=>"111101101",
  58990=>"011010011",
  58991=>"001111010",
  58992=>"100001110",
  58993=>"000010001",
  58994=>"011111101",
  58995=>"000011001",
  58996=>"011100110",
  58997=>"100100101",
  58998=>"001010100",
  58999=>"000010000",
  59000=>"110111010",
  59001=>"001111111",
  59002=>"111000000",
  59003=>"010000010",
  59004=>"101100001",
  59005=>"011010110",
  59006=>"011100101",
  59007=>"011111001",
  59008=>"111101000",
  59009=>"111001110",
  59010=>"001010100",
  59011=>"011000110",
  59012=>"111001011",
  59013=>"100011010",
  59014=>"011100101",
  59015=>"010100011",
  59016=>"010001011",
  59017=>"001000000",
  59018=>"111100011",
  59019=>"000011110",
  59020=>"101100011",
  59021=>"101111011",
  59022=>"001011000",
  59023=>"000111101",
  59024=>"001011101",
  59025=>"110001001",
  59026=>"010100010",
  59027=>"100111001",
  59028=>"001011101",
  59029=>"010000111",
  59030=>"011111001",
  59031=>"110010000",
  59032=>"111101011",
  59033=>"100000101",
  59034=>"100000101",
  59035=>"010001101",
  59036=>"000101011",
  59037=>"100000110",
  59038=>"100100111",
  59039=>"010001000",
  59040=>"101110100",
  59041=>"101010110",
  59042=>"110101101",
  59043=>"101000111",
  59044=>"110010110",
  59045=>"011101101",
  59046=>"011010011",
  59047=>"011010110",
  59048=>"111010011",
  59049=>"101111110",
  59050=>"100001111",
  59051=>"011011011",
  59052=>"001010111",
  59053=>"011111011",
  59054=>"010101001",
  59055=>"100010000",
  59056=>"011101100",
  59057=>"100101000",
  59058=>"001100010",
  59059=>"010100110",
  59060=>"010011111",
  59061=>"011110011",
  59062=>"110100110",
  59063=>"000011101",
  59064=>"010100010",
  59065=>"111000110",
  59066=>"110111101",
  59067=>"011110010",
  59068=>"001011000",
  59069=>"010010000",
  59070=>"000010111",
  59071=>"010001010",
  59072=>"011001010",
  59073=>"000001110",
  59074=>"101101011",
  59075=>"101001110",
  59076=>"011001110",
  59077=>"111101000",
  59078=>"001011101",
  59079=>"010100001",
  59080=>"011000111",
  59081=>"011100001",
  59082=>"011101011",
  59083=>"000001100",
  59084=>"001111101",
  59085=>"111111110",
  59086=>"111011010",
  59087=>"000011010",
  59088=>"101100101",
  59089=>"011000001",
  59090=>"000011110",
  59091=>"011110000",
  59092=>"110010100",
  59093=>"001100010",
  59094=>"101111111",
  59095=>"011101111",
  59096=>"000010000",
  59097=>"010001010",
  59098=>"001011111",
  59099=>"101000111",
  59100=>"010101110",
  59101=>"010101000",
  59102=>"111110001",
  59103=>"000000010",
  59104=>"001111110",
  59105=>"010011000",
  59106=>"011101001",
  59107=>"010101111",
  59108=>"000110111",
  59109=>"110010010",
  59110=>"011100010",
  59111=>"000110111",
  59112=>"100111011",
  59113=>"000000100",
  59114=>"010011100",
  59115=>"101111011",
  59116=>"110111100",
  59117=>"110001110",
  59118=>"001101001",
  59119=>"000100011",
  59120=>"000000110",
  59121=>"101110100",
  59122=>"011011111",
  59123=>"101001000",
  59124=>"001110011",
  59125=>"001111010",
  59126=>"000010001",
  59127=>"010001010",
  59128=>"100011100",
  59129=>"010111010",
  59130=>"100000110",
  59131=>"000000111",
  59132=>"010101110",
  59133=>"010000111",
  59134=>"111001000",
  59135=>"111111011",
  59136=>"101111101",
  59137=>"011110000",
  59138=>"011111010",
  59139=>"001100001",
  59140=>"100101001",
  59141=>"111111000",
  59142=>"111010001",
  59143=>"011001000",
  59144=>"011010001",
  59145=>"100010100",
  59146=>"000100110",
  59147=>"001100011",
  59148=>"011010010",
  59149=>"110110010",
  59150=>"000110011",
  59151=>"111101110",
  59152=>"100111011",
  59153=>"000111000",
  59154=>"100110011",
  59155=>"100001000",
  59156=>"000111010",
  59157=>"010100101",
  59158=>"000101010",
  59159=>"100001000",
  59160=>"001001000",
  59161=>"010011110",
  59162=>"011110110",
  59163=>"111111111",
  59164=>"010001001",
  59165=>"010000111",
  59166=>"000111111",
  59167=>"001000001",
  59168=>"111110010",
  59169=>"011110011",
  59170=>"010111011",
  59171=>"111010000",
  59172=>"110110111",
  59173=>"000000101",
  59174=>"011101010",
  59175=>"011000001",
  59176=>"101101101",
  59177=>"010011001",
  59178=>"011001000",
  59179=>"000010100",
  59180=>"011000111",
  59181=>"000010111",
  59182=>"111111111",
  59183=>"010111111",
  59184=>"111011101",
  59185=>"010010001",
  59186=>"101001100",
  59187=>"010100010",
  59188=>"110110000",
  59189=>"011001010",
  59190=>"011011000",
  59191=>"100001111",
  59192=>"000011010",
  59193=>"001110011",
  59194=>"101000011",
  59195=>"100100111",
  59196=>"101111001",
  59197=>"101001101",
  59198=>"011011100",
  59199=>"100011100",
  59200=>"100011110",
  59201=>"111000100",
  59202=>"110001010",
  59203=>"100001111",
  59204=>"001101111",
  59205=>"000000001",
  59206=>"110011110",
  59207=>"100001001",
  59208=>"110111111",
  59209=>"110100011",
  59210=>"000001001",
  59211=>"010111001",
  59212=>"111111010",
  59213=>"011110010",
  59214=>"101100100",
  59215=>"100010110",
  59216=>"101110111",
  59217=>"001010001",
  59218=>"101111001",
  59219=>"010110000",
  59220=>"001001011",
  59221=>"100011010",
  59222=>"010100111",
  59223=>"100110101",
  59224=>"100001001",
  59225=>"100010011",
  59226=>"010011000",
  59227=>"101010110",
  59228=>"101010011",
  59229=>"111010011",
  59230=>"100010111",
  59231=>"111100111",
  59232=>"101000100",
  59233=>"010000111",
  59234=>"101110110",
  59235=>"110000010",
  59236=>"111000000",
  59237=>"010010110",
  59238=>"110001001",
  59239=>"011111111",
  59240=>"110000000",
  59241=>"111011011",
  59242=>"111100010",
  59243=>"011001011",
  59244=>"001001000",
  59245=>"111011000",
  59246=>"100100001",
  59247=>"111110000",
  59248=>"001001000",
  59249=>"011011000",
  59250=>"111100000",
  59251=>"000111111",
  59252=>"101100101",
  59253=>"111111110",
  59254=>"110111010",
  59255=>"110110010",
  59256=>"011101100",
  59257=>"111101100",
  59258=>"001100110",
  59259=>"110001101",
  59260=>"011111101",
  59261=>"110000111",
  59262=>"111100011",
  59263=>"101110010",
  59264=>"000111110",
  59265=>"111011101",
  59266=>"001111011",
  59267=>"100100100",
  59268=>"100111110",
  59269=>"000000010",
  59270=>"001110000",
  59271=>"000100101",
  59272=>"100111010",
  59273=>"001010011",
  59274=>"011101110",
  59275=>"000000100",
  59276=>"000001000",
  59277=>"000011000",
  59278=>"100101001",
  59279=>"101100110",
  59280=>"001111101",
  59281=>"110110111",
  59282=>"011001000",
  59283=>"000000000",
  59284=>"010110111",
  59285=>"100010011",
  59286=>"001101110",
  59287=>"101101010",
  59288=>"111001111",
  59289=>"100001010",
  59290=>"000100010",
  59291=>"101111111",
  59292=>"111101110",
  59293=>"011010000",
  59294=>"110100101",
  59295=>"010000101",
  59296=>"110111101",
  59297=>"110011010",
  59298=>"000010111",
  59299=>"011110010",
  59300=>"100001011",
  59301=>"011001110",
  59302=>"001101000",
  59303=>"000101000",
  59304=>"100100010",
  59305=>"101110101",
  59306=>"111010111",
  59307=>"111111100",
  59308=>"001010011",
  59309=>"010101111",
  59310=>"100001100",
  59311=>"100101000",
  59312=>"111010111",
  59313=>"000101100",
  59314=>"101000011",
  59315=>"101010100",
  59316=>"001100010",
  59317=>"011011111",
  59318=>"011001101",
  59319=>"000100100",
  59320=>"100110001",
  59321=>"010100000",
  59322=>"001111110",
  59323=>"011010111",
  59324=>"011011111",
  59325=>"100000100",
  59326=>"000101110",
  59327=>"101111011",
  59328=>"110111111",
  59329=>"000010111",
  59330=>"010111100",
  59331=>"010111000",
  59332=>"100000101",
  59333=>"011001010",
  59334=>"011111100",
  59335=>"100001101",
  59336=>"101100110",
  59337=>"001100010",
  59338=>"011010101",
  59339=>"111011101",
  59340=>"111000011",
  59341=>"000000010",
  59342=>"110011110",
  59343=>"110000010",
  59344=>"010001110",
  59345=>"010001110",
  59346=>"000001010",
  59347=>"111000001",
  59348=>"011111111",
  59349=>"000101110",
  59350=>"011000010",
  59351=>"000010001",
  59352=>"111101010",
  59353=>"001011110",
  59354=>"001101111",
  59355=>"111111010",
  59356=>"011110001",
  59357=>"101100110",
  59358=>"111101111",
  59359=>"110111101",
  59360=>"111110100",
  59361=>"100001101",
  59362=>"101010111",
  59363=>"100001000",
  59364=>"000110111",
  59365=>"010010010",
  59366=>"111100111",
  59367=>"011001101",
  59368=>"011101011",
  59369=>"011110011",
  59370=>"000010110",
  59371=>"110010011",
  59372=>"110100111",
  59373=>"110001100",
  59374=>"100001011",
  59375=>"111011101",
  59376=>"111011111",
  59377=>"000010010",
  59378=>"000000011",
  59379=>"100101001",
  59380=>"110100101",
  59381=>"011000011",
  59382=>"110011001",
  59383=>"000100001",
  59384=>"001001010",
  59385=>"001111010",
  59386=>"110111011",
  59387=>"011111001",
  59388=>"000100100",
  59389=>"100111000",
  59390=>"011010011",
  59391=>"000010100",
  59392=>"000001101",
  59393=>"000011101",
  59394=>"111100111",
  59395=>"110011100",
  59396=>"000011011",
  59397=>"000001100",
  59398=>"100000000",
  59399=>"000011111",
  59400=>"100001000",
  59401=>"001011100",
  59402=>"111001001",
  59403=>"010011111",
  59404=>"100100110",
  59405=>"001001000",
  59406=>"111001100",
  59407=>"111001111",
  59408=>"000001101",
  59409=>"000001101",
  59410=>"101011011",
  59411=>"101100010",
  59412=>"001100101",
  59413=>"100010001",
  59414=>"110011100",
  59415=>"101000110",
  59416=>"111011001",
  59417=>"111110010",
  59418=>"110011111",
  59419=>"000101000",
  59420=>"111000011",
  59421=>"000001000",
  59422=>"100101111",
  59423=>"001011111",
  59424=>"011101011",
  59425=>"111111000",
  59426=>"110000000",
  59427=>"101100100",
  59428=>"010001010",
  59429=>"001010011",
  59430=>"000111111",
  59431=>"100000000",
  59432=>"010110101",
  59433=>"101001011",
  59434=>"100100001",
  59435=>"000000111",
  59436=>"111100100",
  59437=>"000001011",
  59438=>"111100001",
  59439=>"011110100",
  59440=>"001010101",
  59441=>"000110100",
  59442=>"000100000",
  59443=>"111011111",
  59444=>"001111111",
  59445=>"001000101",
  59446=>"010001100",
  59447=>"001100111",
  59448=>"010011010",
  59449=>"011011101",
  59450=>"010001111",
  59451=>"100100001",
  59452=>"100000111",
  59453=>"000001011",
  59454=>"011111101",
  59455=>"100100101",
  59456=>"000011011",
  59457=>"000100100",
  59458=>"010001011",
  59459=>"110110001",
  59460=>"100100000",
  59461=>"100111100",
  59462=>"110001011",
  59463=>"001010000",
  59464=>"100110010",
  59465=>"000000000",
  59466=>"110001000",
  59467=>"010001101",
  59468=>"110110000",
  59469=>"001110001",
  59470=>"000100011",
  59471=>"011011110",
  59472=>"110001011",
  59473=>"111101101",
  59474=>"000111110",
  59475=>"010011101",
  59476=>"001110000",
  59477=>"000101100",
  59478=>"010010001",
  59479=>"101100111",
  59480=>"000000011",
  59481=>"011101101",
  59482=>"101101101",
  59483=>"111001100",
  59484=>"010011000",
  59485=>"100000011",
  59486=>"111101011",
  59487=>"000101101",
  59488=>"100101111",
  59489=>"011000000",
  59490=>"000000001",
  59491=>"011000010",
  59492=>"010101100",
  59493=>"100011000",
  59494=>"110010110",
  59495=>"001110100",
  59496=>"111011011",
  59497=>"010001100",
  59498=>"100011100",
  59499=>"101011110",
  59500=>"100001110",
  59501=>"111100101",
  59502=>"111011011",
  59503=>"101010101",
  59504=>"101100110",
  59505=>"010010111",
  59506=>"100101111",
  59507=>"100111010",
  59508=>"001011111",
  59509=>"111111101",
  59510=>"110111110",
  59511=>"011010001",
  59512=>"110111100",
  59513=>"001001010",
  59514=>"100001101",
  59515=>"111111110",
  59516=>"111001101",
  59517=>"011101100",
  59518=>"001000111",
  59519=>"111000101",
  59520=>"110101001",
  59521=>"110000100",
  59522=>"000001000",
  59523=>"011100101",
  59524=>"001001100",
  59525=>"110011101",
  59526=>"111111111",
  59527=>"010001100",
  59528=>"110110010",
  59529=>"011100100",
  59530=>"110111011",
  59531=>"010010101",
  59532=>"111110011",
  59533=>"101111110",
  59534=>"100010001",
  59535=>"100011101",
  59536=>"000001001",
  59537=>"111000101",
  59538=>"110100010",
  59539=>"010110011",
  59540=>"010011101",
  59541=>"100110101",
  59542=>"000010100",
  59543=>"101111000",
  59544=>"011000000",
  59545=>"101000001",
  59546=>"010011100",
  59547=>"010110011",
  59548=>"101111100",
  59549=>"100010101",
  59550=>"011001100",
  59551=>"011110110",
  59552=>"101100011",
  59553=>"001101110",
  59554=>"011110110",
  59555=>"111111011",
  59556=>"000000001",
  59557=>"001010101",
  59558=>"001000011",
  59559=>"101101110",
  59560=>"011111000",
  59561=>"000001011",
  59562=>"011011010",
  59563=>"101001001",
  59564=>"111000110",
  59565=>"111111000",
  59566=>"001011000",
  59567=>"100001011",
  59568=>"110100100",
  59569=>"000010110",
  59570=>"110011000",
  59571=>"000011111",
  59572=>"001000001",
  59573=>"000110001",
  59574=>"110011000",
  59575=>"100100000",
  59576=>"001101001",
  59577=>"101110100",
  59578=>"001101100",
  59579=>"010010011",
  59580=>"001111101",
  59581=>"001010001",
  59582=>"001101110",
  59583=>"111000111",
  59584=>"010111100",
  59585=>"111010000",
  59586=>"110010010",
  59587=>"010111011",
  59588=>"010001001",
  59589=>"000110011",
  59590=>"011010010",
  59591=>"011111000",
  59592=>"010111110",
  59593=>"111010101",
  59594=>"001000100",
  59595=>"011110010",
  59596=>"111001111",
  59597=>"111010101",
  59598=>"000010101",
  59599=>"000001000",
  59600=>"110100110",
  59601=>"110110001",
  59602=>"101000101",
  59603=>"001101110",
  59604=>"110100101",
  59605=>"010100100",
  59606=>"110101111",
  59607=>"001000101",
  59608=>"100100100",
  59609=>"110110000",
  59610=>"110011001",
  59611=>"100100011",
  59612=>"011110010",
  59613=>"010110101",
  59614=>"000001111",
  59615=>"011101110",
  59616=>"001001101",
  59617=>"110100000",
  59618=>"110110010",
  59619=>"000101011",
  59620=>"001101001",
  59621=>"110100000",
  59622=>"001110000",
  59623=>"110111100",
  59624=>"111000001",
  59625=>"001110001",
  59626=>"001000010",
  59627=>"111100101",
  59628=>"111100001",
  59629=>"111000000",
  59630=>"110100010",
  59631=>"010000000",
  59632=>"011101011",
  59633=>"010110001",
  59634=>"010000100",
  59635=>"011010001",
  59636=>"111001110",
  59637=>"111000100",
  59638=>"101000010",
  59639=>"110110000",
  59640=>"010010000",
  59641=>"001111000",
  59642=>"101011100",
  59643=>"110010001",
  59644=>"000000110",
  59645=>"100000101",
  59646=>"010111011",
  59647=>"110100111",
  59648=>"001000000",
  59649=>"100010111",
  59650=>"111000011",
  59651=>"110111100",
  59652=>"000110000",
  59653=>"000110101",
  59654=>"000100111",
  59655=>"100110000",
  59656=>"010111010",
  59657=>"011111001",
  59658=>"001011000",
  59659=>"101000100",
  59660=>"101100011",
  59661=>"001001110",
  59662=>"101010110",
  59663=>"011001101",
  59664=>"111011100",
  59665=>"100010010",
  59666=>"110001100",
  59667=>"011010011",
  59668=>"100000010",
  59669=>"100100000",
  59670=>"101111001",
  59671=>"001000101",
  59672=>"110001101",
  59673=>"101100000",
  59674=>"000011111",
  59675=>"001101100",
  59676=>"101011110",
  59677=>"000101001",
  59678=>"100001010",
  59679=>"011001110",
  59680=>"111010000",
  59681=>"011101010",
  59682=>"110101100",
  59683=>"000001101",
  59684=>"110011010",
  59685=>"010000000",
  59686=>"010000111",
  59687=>"110001101",
  59688=>"110011000",
  59689=>"001010101",
  59690=>"011010010",
  59691=>"100001110",
  59692=>"111100011",
  59693=>"101011000",
  59694=>"011110101",
  59695=>"010000101",
  59696=>"110110000",
  59697=>"101010000",
  59698=>"000110010",
  59699=>"011101100",
  59700=>"001011001",
  59701=>"100110101",
  59702=>"111011000",
  59703=>"100010101",
  59704=>"001011000",
  59705=>"100101100",
  59706=>"011110110",
  59707=>"000110000",
  59708=>"001100010",
  59709=>"101011011",
  59710=>"110111110",
  59711=>"101010110",
  59712=>"110000101",
  59713=>"001010000",
  59714=>"110010111",
  59715=>"011110110",
  59716=>"111110111",
  59717=>"100000011",
  59718=>"100110000",
  59719=>"011111111",
  59720=>"100111111",
  59721=>"100101011",
  59722=>"101011001",
  59723=>"000110011",
  59724=>"100100011",
  59725=>"000111110",
  59726=>"001001111",
  59727=>"111110010",
  59728=>"100001100",
  59729=>"011000010",
  59730=>"011011111",
  59731=>"111101111",
  59732=>"100010000",
  59733=>"000010010",
  59734=>"011110101",
  59735=>"000011010",
  59736=>"010100010",
  59737=>"000001111",
  59738=>"001101000",
  59739=>"110101000",
  59740=>"000010110",
  59741=>"000001100",
  59742=>"011101101",
  59743=>"000000011",
  59744=>"101111010",
  59745=>"011000011",
  59746=>"111100101",
  59747=>"011010100",
  59748=>"000001111",
  59749=>"111111110",
  59750=>"011000001",
  59751=>"010100111",
  59752=>"011011111",
  59753=>"000110100",
  59754=>"100110111",
  59755=>"100111111",
  59756=>"000011001",
  59757=>"010111111",
  59758=>"001111010",
  59759=>"111010111",
  59760=>"111110101",
  59761=>"100000101",
  59762=>"011100010",
  59763=>"000010100",
  59764=>"111111100",
  59765=>"011000111",
  59766=>"100111100",
  59767=>"011011101",
  59768=>"101100101",
  59769=>"000111110",
  59770=>"001111001",
  59771=>"101011010",
  59772=>"000101000",
  59773=>"000101000",
  59774=>"101001110",
  59775=>"111100001",
  59776=>"101001100",
  59777=>"000101001",
  59778=>"101010000",
  59779=>"010011000",
  59780=>"111111011",
  59781=>"110110001",
  59782=>"100011100",
  59783=>"101010011",
  59784=>"101011000",
  59785=>"011000101",
  59786=>"110100000",
  59787=>"001001101",
  59788=>"010000100",
  59789=>"101100101",
  59790=>"100110111",
  59791=>"100111111",
  59792=>"011000111",
  59793=>"010111000",
  59794=>"101001011",
  59795=>"110111000",
  59796=>"110101100",
  59797=>"001110010",
  59798=>"010110110",
  59799=>"100110111",
  59800=>"100001000",
  59801=>"100010110",
  59802=>"111101101",
  59803=>"100001001",
  59804=>"101010001",
  59805=>"101101111",
  59806=>"010011001",
  59807=>"110000010",
  59808=>"000111111",
  59809=>"101110011",
  59810=>"000010011",
  59811=>"001110011",
  59812=>"110110011",
  59813=>"000100000",
  59814=>"000001111",
  59815=>"110111001",
  59816=>"111010111",
  59817=>"011100000",
  59818=>"100100000",
  59819=>"000110100",
  59820=>"101101101",
  59821=>"100010001",
  59822=>"010111111",
  59823=>"111101100",
  59824=>"001010001",
  59825=>"111000110",
  59826=>"110010001",
  59827=>"000101100",
  59828=>"000001000",
  59829=>"010110011",
  59830=>"000100111",
  59831=>"000001011",
  59832=>"101101000",
  59833=>"100010010",
  59834=>"100000111",
  59835=>"101001010",
  59836=>"101010001",
  59837=>"101001011",
  59838=>"100001011",
  59839=>"101001100",
  59840=>"000101100",
  59841=>"110100011",
  59842=>"110011101",
  59843=>"001000101",
  59844=>"011101101",
  59845=>"101001011",
  59846=>"111010001",
  59847=>"111001110",
  59848=>"001001100",
  59849=>"001000010",
  59850=>"011100001",
  59851=>"001011111",
  59852=>"111001100",
  59853=>"001111000",
  59854=>"101001110",
  59855=>"110110110",
  59856=>"111000011",
  59857=>"110000011",
  59858=>"011101001",
  59859=>"000110100",
  59860=>"101101001",
  59861=>"010000101",
  59862=>"011101011",
  59863=>"010000101",
  59864=>"001011100",
  59865=>"010100100",
  59866=>"100001010",
  59867=>"110001000",
  59868=>"111111100",
  59869=>"100010001",
  59870=>"011011101",
  59871=>"000001010",
  59872=>"101001011",
  59873=>"110110001",
  59874=>"101101101",
  59875=>"000000001",
  59876=>"010000010",
  59877=>"011011111",
  59878=>"100011000",
  59879=>"100000100",
  59880=>"111101000",
  59881=>"001011001",
  59882=>"001100110",
  59883=>"111001101",
  59884=>"100000110",
  59885=>"100001111",
  59886=>"101110110",
  59887=>"010010111",
  59888=>"110010000",
  59889=>"101101111",
  59890=>"001011000",
  59891=>"000001001",
  59892=>"111010100",
  59893=>"110101110",
  59894=>"110111110",
  59895=>"001011010",
  59896=>"001101101",
  59897=>"100010011",
  59898=>"000000000",
  59899=>"111010100",
  59900=>"101001101",
  59901=>"110010100",
  59902=>"011111010",
  59903=>"010111111",
  59904=>"000111000",
  59905=>"001111100",
  59906=>"000000010",
  59907=>"000100100",
  59908=>"110010001",
  59909=>"101000000",
  59910=>"100001001",
  59911=>"100111000",
  59912=>"100000001",
  59913=>"010110011",
  59914=>"001111000",
  59915=>"110011001",
  59916=>"100001111",
  59917=>"001101000",
  59918=>"111101100",
  59919=>"110010000",
  59920=>"001100000",
  59921=>"101100010",
  59922=>"011000000",
  59923=>"111101100",
  59924=>"101000101",
  59925=>"111011111",
  59926=>"000010110",
  59927=>"111001110",
  59928=>"000101101",
  59929=>"000000100",
  59930=>"000101000",
  59931=>"001001110",
  59932=>"010110001",
  59933=>"011000011",
  59934=>"011001100",
  59935=>"110111011",
  59936=>"101011001",
  59937=>"000000000",
  59938=>"101111110",
  59939=>"100010101",
  59940=>"001100000",
  59941=>"010110010",
  59942=>"100000000",
  59943=>"000001101",
  59944=>"101111001",
  59945=>"110101101",
  59946=>"011011100",
  59947=>"000001000",
  59948=>"111100110",
  59949=>"011101101",
  59950=>"110001001",
  59951=>"010111001",
  59952=>"011001101",
  59953=>"100010100",
  59954=>"010011000",
  59955=>"001011011",
  59956=>"110110100",
  59957=>"110100001",
  59958=>"110000001",
  59959=>"101000110",
  59960=>"100011010",
  59961=>"010000111",
  59962=>"111110000",
  59963=>"110110010",
  59964=>"001011111",
  59965=>"111011110",
  59966=>"100010111",
  59967=>"010011100",
  59968=>"000000000",
  59969=>"111101111",
  59970=>"001101010",
  59971=>"010000111",
  59972=>"100101111",
  59973=>"000010100",
  59974=>"010110100",
  59975=>"011010000",
  59976=>"101101000",
  59977=>"001001010",
  59978=>"111111110",
  59979=>"111110101",
  59980=>"000110110",
  59981=>"101111100",
  59982=>"001111110",
  59983=>"110000000",
  59984=>"110000011",
  59985=>"010000010",
  59986=>"101101111",
  59987=>"001101101",
  59988=>"001110000",
  59989=>"100001001",
  59990=>"101010000",
  59991=>"111000101",
  59992=>"000101111",
  59993=>"000100111",
  59994=>"110110110",
  59995=>"010011000",
  59996=>"101100100",
  59997=>"011110111",
  59998=>"010110110",
  59999=>"001101011",
  60000=>"011010101",
  60001=>"001100010",
  60002=>"010000111",
  60003=>"000010110",
  60004=>"011000111",
  60005=>"100000010",
  60006=>"111001100",
  60007=>"000100001",
  60008=>"010011111",
  60009=>"100100000",
  60010=>"100000111",
  60011=>"111000100",
  60012=>"010111001",
  60013=>"000101101",
  60014=>"001111101",
  60015=>"010001111",
  60016=>"100111101",
  60017=>"000000000",
  60018=>"111000010",
  60019=>"010001010",
  60020=>"111101000",
  60021=>"110101010",
  60022=>"000100011",
  60023=>"101011110",
  60024=>"111000000",
  60025=>"001101000",
  60026=>"000100000",
  60027=>"101011100",
  60028=>"010100111",
  60029=>"000100100",
  60030=>"011011101",
  60031=>"101100111",
  60032=>"100110110",
  60033=>"011111010",
  60034=>"110000001",
  60035=>"010111011",
  60036=>"100111001",
  60037=>"110010101",
  60038=>"101000100",
  60039=>"101000111",
  60040=>"000101000",
  60041=>"000111100",
  60042=>"010111111",
  60043=>"001111100",
  60044=>"100000111",
  60045=>"111111110",
  60046=>"010010111",
  60047=>"110111011",
  60048=>"011000111",
  60049=>"011101110",
  60050=>"010101000",
  60051=>"100111010",
  60052=>"110101100",
  60053=>"000101101",
  60054=>"000101101",
  60055=>"111110111",
  60056=>"000101100",
  60057=>"010001100",
  60058=>"100010101",
  60059=>"010101100",
  60060=>"100110000",
  60061=>"101111010",
  60062=>"011000001",
  60063=>"010000010",
  60064=>"110010110",
  60065=>"011001101",
  60066=>"010011000",
  60067=>"111111011",
  60068=>"000000010",
  60069=>"011000000",
  60070=>"101110100",
  60071=>"111110101",
  60072=>"111010100",
  60073=>"100001100",
  60074=>"001010010",
  60075=>"000100011",
  60076=>"001100000",
  60077=>"101001111",
  60078=>"010010101",
  60079=>"100111110",
  60080=>"111111010",
  60081=>"111100110",
  60082=>"100111001",
  60083=>"001011000",
  60084=>"110010100",
  60085=>"001000111",
  60086=>"001001110",
  60087=>"111111011",
  60088=>"011011011",
  60089=>"001011110",
  60090=>"011111101",
  60091=>"000100001",
  60092=>"001011000",
  60093=>"111001110",
  60094=>"000011111",
  60095=>"111000001",
  60096=>"000100100",
  60097=>"000001001",
  60098=>"010110000",
  60099=>"001000010",
  60100=>"001000000",
  60101=>"101010100",
  60102=>"110001110",
  60103=>"001111111",
  60104=>"100011110",
  60105=>"010000000",
  60106=>"101100101",
  60107=>"001000111",
  60108=>"001100100",
  60109=>"011010011",
  60110=>"001100111",
  60111=>"100111001",
  60112=>"100000011",
  60113=>"010000001",
  60114=>"011000111",
  60115=>"000001000",
  60116=>"101101001",
  60117=>"100111000",
  60118=>"001010100",
  60119=>"111111100",
  60120=>"110000010",
  60121=>"000000011",
  60122=>"111101110",
  60123=>"001000110",
  60124=>"100100111",
  60125=>"101100111",
  60126=>"000111011",
  60127=>"000101110",
  60128=>"010000001",
  60129=>"011001110",
  60130=>"010001000",
  60131=>"100001010",
  60132=>"101101010",
  60133=>"001101110",
  60134=>"110110111",
  60135=>"100110101",
  60136=>"011110011",
  60137=>"011000110",
  60138=>"101011111",
  60139=>"000111101",
  60140=>"011110010",
  60141=>"101100010",
  60142=>"001100000",
  60143=>"000000010",
  60144=>"110101001",
  60145=>"100111111",
  60146=>"010000100",
  60147=>"111111000",
  60148=>"010111010",
  60149=>"110110010",
  60150=>"010100110",
  60151=>"101100000",
  60152=>"111000001",
  60153=>"001110001",
  60154=>"101111011",
  60155=>"111010111",
  60156=>"011011110",
  60157=>"011110010",
  60158=>"111010010",
  60159=>"110101101",
  60160=>"100100100",
  60161=>"111111111",
  60162=>"000010100",
  60163=>"010100011",
  60164=>"100101001",
  60165=>"111110100",
  60166=>"111000001",
  60167=>"100110001",
  60168=>"111111001",
  60169=>"010010110",
  60170=>"100100100",
  60171=>"101000010",
  60172=>"010100110",
  60173=>"100001011",
  60174=>"010000011",
  60175=>"100100000",
  60176=>"010110011",
  60177=>"101001010",
  60178=>"010110001",
  60179=>"010100000",
  60180=>"100010001",
  60181=>"011011010",
  60182=>"111000011",
  60183=>"110101110",
  60184=>"101100101",
  60185=>"011110000",
  60186=>"100010101",
  60187=>"000111010",
  60188=>"010110100",
  60189=>"110001011",
  60190=>"110011100",
  60191=>"000000001",
  60192=>"111110111",
  60193=>"101011000",
  60194=>"010001101",
  60195=>"000100110",
  60196=>"010101111",
  60197=>"101101111",
  60198=>"001110100",
  60199=>"001000001",
  60200=>"100000000",
  60201=>"000011100",
  60202=>"010000000",
  60203=>"111111100",
  60204=>"000110100",
  60205=>"110000010",
  60206=>"101001110",
  60207=>"110111011",
  60208=>"110100001",
  60209=>"011101001",
  60210=>"111000100",
  60211=>"001110010",
  60212=>"101110001",
  60213=>"011111010",
  60214=>"010100010",
  60215=>"000110001",
  60216=>"111111110",
  60217=>"010011101",
  60218=>"000010101",
  60219=>"111100011",
  60220=>"110000011",
  60221=>"001001010",
  60222=>"001110111",
  60223=>"110110110",
  60224=>"011100010",
  60225=>"101001101",
  60226=>"110010000",
  60227=>"101101100",
  60228=>"010100101",
  60229=>"001011100",
  60230=>"001011111",
  60231=>"001111100",
  60232=>"011101111",
  60233=>"001100100",
  60234=>"100010101",
  60235=>"100111010",
  60236=>"111100000",
  60237=>"111000011",
  60238=>"010001011",
  60239=>"001000010",
  60240=>"101011101",
  60241=>"111011010",
  60242=>"001000100",
  60243=>"111000100",
  60244=>"010001101",
  60245=>"111111110",
  60246=>"101100100",
  60247=>"000010010",
  60248=>"000101011",
  60249=>"001100001",
  60250=>"000100101",
  60251=>"111000110",
  60252=>"100011101",
  60253=>"001111101",
  60254=>"010110010",
  60255=>"100010011",
  60256=>"111000010",
  60257=>"110110010",
  60258=>"000111110",
  60259=>"000010000",
  60260=>"100101111",
  60261=>"000110100",
  60262=>"000111110",
  60263=>"000010000",
  60264=>"000100111",
  60265=>"001111100",
  60266=>"010010001",
  60267=>"110110111",
  60268=>"100111000",
  60269=>"010000100",
  60270=>"111110110",
  60271=>"000101010",
  60272=>"000100001",
  60273=>"111110100",
  60274=>"001000100",
  60275=>"011111000",
  60276=>"100100011",
  60277=>"010101111",
  60278=>"101010100",
  60279=>"001000100",
  60280=>"100010110",
  60281=>"111001000",
  60282=>"100101011",
  60283=>"010001011",
  60284=>"010001001",
  60285=>"101011101",
  60286=>"101101101",
  60287=>"011011101",
  60288=>"001001111",
  60289=>"001010000",
  60290=>"101111010",
  60291=>"100000011",
  60292=>"010111111",
  60293=>"010110111",
  60294=>"101101100",
  60295=>"110001110",
  60296=>"010101110",
  60297=>"000010010",
  60298=>"111001011",
  60299=>"101111111",
  60300=>"110011111",
  60301=>"010011000",
  60302=>"010101000",
  60303=>"100001100",
  60304=>"101001110",
  60305=>"110110010",
  60306=>"101111001",
  60307=>"100110100",
  60308=>"000011011",
  60309=>"001111110",
  60310=>"111000100",
  60311=>"001111101",
  60312=>"100100000",
  60313=>"101011101",
  60314=>"000100010",
  60315=>"110000101",
  60316=>"100100101",
  60317=>"100000000",
  60318=>"100001000",
  60319=>"110011011",
  60320=>"000000011",
  60321=>"001100101",
  60322=>"110011110",
  60323=>"001101000",
  60324=>"011000110",
  60325=>"011111111",
  60326=>"001011010",
  60327=>"111011011",
  60328=>"010001010",
  60329=>"111100111",
  60330=>"010011111",
  60331=>"011111001",
  60332=>"111000100",
  60333=>"011110011",
  60334=>"011111110",
  60335=>"001100001",
  60336=>"111111100",
  60337=>"100111100",
  60338=>"000101000",
  60339=>"011000100",
  60340=>"011110111",
  60341=>"001101110",
  60342=>"001101111",
  60343=>"110011110",
  60344=>"100000001",
  60345=>"011111111",
  60346=>"001011001",
  60347=>"011110100",
  60348=>"111100110",
  60349=>"000111111",
  60350=>"001101110",
  60351=>"101000111",
  60352=>"001010110",
  60353=>"111010010",
  60354=>"101000110",
  60355=>"100111011",
  60356=>"011101001",
  60357=>"001100100",
  60358=>"101110001",
  60359=>"110011100",
  60360=>"111100011",
  60361=>"000111111",
  60362=>"011000010",
  60363=>"001000010",
  60364=>"010111001",
  60365=>"101100111",
  60366=>"100111001",
  60367=>"101000011",
  60368=>"111010101",
  60369=>"011100001",
  60370=>"111101000",
  60371=>"010111101",
  60372=>"101101111",
  60373=>"110111110",
  60374=>"111100100",
  60375=>"111000000",
  60376=>"100100111",
  60377=>"110110111",
  60378=>"011000110",
  60379=>"000101111",
  60380=>"101110000",
  60381=>"001110011",
  60382=>"111010100",
  60383=>"001010110",
  60384=>"110100101",
  60385=>"011010110",
  60386=>"101111111",
  60387=>"110110010",
  60388=>"111110110",
  60389=>"110011010",
  60390=>"001001001",
  60391=>"100101110",
  60392=>"000100101",
  60393=>"000000001",
  60394=>"110000001",
  60395=>"000111000",
  60396=>"011111010",
  60397=>"111101110",
  60398=>"001001100",
  60399=>"000110111",
  60400=>"011110010",
  60401=>"101010111",
  60402=>"100111010",
  60403=>"000001111",
  60404=>"000000000",
  60405=>"001010000",
  60406=>"011100100",
  60407=>"010010000",
  60408=>"110100000",
  60409=>"111000000",
  60410=>"000100110",
  60411=>"110001000",
  60412=>"110100000",
  60413=>"110010001",
  60414=>"110111000",
  60415=>"011000001",
  60416=>"101111101",
  60417=>"111101101",
  60418=>"100100001",
  60419=>"110010000",
  60420=>"000101111",
  60421=>"001100000",
  60422=>"000100000",
  60423=>"011001001",
  60424=>"110101110",
  60425=>"100010100",
  60426=>"011011010",
  60427=>"000000100",
  60428=>"110110111",
  60429=>"110101111",
  60430=>"101111000",
  60431=>"000100111",
  60432=>"011001001",
  60433=>"101110110",
  60434=>"010000100",
  60435=>"100000001",
  60436=>"110000000",
  60437=>"111101111",
  60438=>"000100010",
  60439=>"111111110",
  60440=>"111110101",
  60441=>"000001001",
  60442=>"011110000",
  60443=>"000100001",
  60444=>"010000101",
  60445=>"000100000",
  60446=>"111111010",
  60447=>"110100000",
  60448=>"110111110",
  60449=>"000011101",
  60450=>"110101111",
  60451=>"100001010",
  60452=>"110110011",
  60453=>"110000100",
  60454=>"100100101",
  60455=>"000101100",
  60456=>"100110011",
  60457=>"001000110",
  60458=>"110101110",
  60459=>"010110100",
  60460=>"011110100",
  60461=>"110010000",
  60462=>"110001111",
  60463=>"011111110",
  60464=>"101000000",
  60465=>"110110001",
  60466=>"101100010",
  60467=>"001010100",
  60468=>"010001101",
  60469=>"100100110",
  60470=>"000101010",
  60471=>"000010000",
  60472=>"011111100",
  60473=>"101001111",
  60474=>"000001111",
  60475=>"101000010",
  60476=>"111001011",
  60477=>"110111001",
  60478=>"100001011",
  60479=>"111110011",
  60480=>"111010110",
  60481=>"010010001",
  60482=>"000010101",
  60483=>"100110000",
  60484=>"111101000",
  60485=>"111100001",
  60486=>"011110010",
  60487=>"111100101",
  60488=>"000111000",
  60489=>"110011001",
  60490=>"010100011",
  60491=>"101011001",
  60492=>"010000001",
  60493=>"010001011",
  60494=>"110001110",
  60495=>"110000010",
  60496=>"101100111",
  60497=>"111000111",
  60498=>"000110101",
  60499=>"110000001",
  60500=>"100010001",
  60501=>"110001010",
  60502=>"100000011",
  60503=>"011001001",
  60504=>"111011111",
  60505=>"010001100",
  60506=>"001011010",
  60507=>"001111100",
  60508=>"001011111",
  60509=>"100100010",
  60510=>"000000100",
  60511=>"110101101",
  60512=>"000001011",
  60513=>"111101010",
  60514=>"110001101",
  60515=>"010101000",
  60516=>"000001011",
  60517=>"111001011",
  60518=>"001001001",
  60519=>"010011001",
  60520=>"000100101",
  60521=>"000110111",
  60522=>"000011001",
  60523=>"000100000",
  60524=>"111001100",
  60525=>"111101111",
  60526=>"001001110",
  60527=>"101000111",
  60528=>"100000010",
  60529=>"110101011",
  60530=>"011001110",
  60531=>"100000100",
  60532=>"111010000",
  60533=>"110111011",
  60534=>"110001110",
  60535=>"001101000",
  60536=>"011100111",
  60537=>"001000010",
  60538=>"001000110",
  60539=>"010001010",
  60540=>"100110111",
  60541=>"100111111",
  60542=>"110100110",
  60543=>"001110110",
  60544=>"000010011",
  60545=>"110000000",
  60546=>"011110000",
  60547=>"001111100",
  60548=>"000110101",
  60549=>"110011000",
  60550=>"001010101",
  60551=>"101000010",
  60552=>"010001010",
  60553=>"110011110",
  60554=>"111101101",
  60555=>"101010100",
  60556=>"011011110",
  60557=>"000100110",
  60558=>"011000110",
  60559=>"000001010",
  60560=>"110001101",
  60561=>"111100101",
  60562=>"101111000",
  60563=>"011111111",
  60564=>"101010110",
  60565=>"001010110",
  60566=>"111111010",
  60567=>"001010111",
  60568=>"110100000",
  60569=>"110100000",
  60570=>"100111111",
  60571=>"100111101",
  60572=>"010100101",
  60573=>"100100001",
  60574=>"011100011",
  60575=>"010011000",
  60576=>"100011111",
  60577=>"101111110",
  60578=>"111111110",
  60579=>"101111101",
  60580=>"011011011",
  60581=>"110101111",
  60582=>"001010000",
  60583=>"000110101",
  60584=>"101000001",
  60585=>"010001111",
  60586=>"000001001",
  60587=>"011000100",
  60588=>"010000100",
  60589=>"100100101",
  60590=>"101010011",
  60591=>"010011100",
  60592=>"100010001",
  60593=>"001000101",
  60594=>"101000011",
  60595=>"000010100",
  60596=>"111011101",
  60597=>"000100111",
  60598=>"100101111",
  60599=>"101110001",
  60600=>"000100101",
  60601=>"010101000",
  60602=>"011011111",
  60603=>"100100111",
  60604=>"011111010",
  60605=>"100110111",
  60606=>"101001001",
  60607=>"111011011",
  60608=>"110111110",
  60609=>"101101000",
  60610=>"110010000",
  60611=>"101011001",
  60612=>"100101001",
  60613=>"111110000",
  60614=>"000010000",
  60615=>"011101000",
  60616=>"110101001",
  60617=>"000000100",
  60618=>"101110000",
  60619=>"001101100",
  60620=>"100100010",
  60621=>"010101000",
  60622=>"111000110",
  60623=>"111111010",
  60624=>"100011010",
  60625=>"010010100",
  60626=>"111011000",
  60627=>"101000100",
  60628=>"110110110",
  60629=>"111010101",
  60630=>"100101011",
  60631=>"100111100",
  60632=>"000101000",
  60633=>"101100100",
  60634=>"111001011",
  60635=>"011110110",
  60636=>"010110101",
  60637=>"101010100",
  60638=>"110011001",
  60639=>"011011010",
  60640=>"100001000",
  60641=>"111100100",
  60642=>"101110100",
  60643=>"110000100",
  60644=>"111000000",
  60645=>"000001110",
  60646=>"010100110",
  60647=>"010111010",
  60648=>"110100011",
  60649=>"111010001",
  60650=>"100010001",
  60651=>"110000001",
  60652=>"110111010",
  60653=>"001111010",
  60654=>"010111000",
  60655=>"000100000",
  60656=>"111000101",
  60657=>"001010010",
  60658=>"010001101",
  60659=>"100001000",
  60660=>"010001110",
  60661=>"110001000",
  60662=>"000101010",
  60663=>"000010010",
  60664=>"000100101",
  60665=>"110010111",
  60666=>"110110011",
  60667=>"010110010",
  60668=>"101000000",
  60669=>"110011001",
  60670=>"100010101",
  60671=>"111001111",
  60672=>"001110101",
  60673=>"010001111",
  60674=>"111100000",
  60675=>"001010100",
  60676=>"110111000",
  60677=>"111111001",
  60678=>"110111101",
  60679=>"100100010",
  60680=>"110111010",
  60681=>"100110010",
  60682=>"100001100",
  60683=>"001011001",
  60684=>"101111110",
  60685=>"111010000",
  60686=>"000100101",
  60687=>"000001101",
  60688=>"010111110",
  60689=>"101111001",
  60690=>"001010100",
  60691=>"011100011",
  60692=>"000111011",
  60693=>"111100010",
  60694=>"000100000",
  60695=>"110001110",
  60696=>"100000111",
  60697=>"000101000",
  60698=>"010100000",
  60699=>"100001101",
  60700=>"111110100",
  60701=>"000111101",
  60702=>"011101101",
  60703=>"000010001",
  60704=>"110100011",
  60705=>"010010100",
  60706=>"001011001",
  60707=>"100111110",
  60708=>"101101010",
  60709=>"100010010",
  60710=>"100111101",
  60711=>"111111010",
  60712=>"000110110",
  60713=>"010010101",
  60714=>"000111111",
  60715=>"000110101",
  60716=>"000000001",
  60717=>"101001001",
  60718=>"011101101",
  60719=>"001111010",
  60720=>"101011101",
  60721=>"110010111",
  60722=>"010110011",
  60723=>"000011001",
  60724=>"101110010",
  60725=>"000001010",
  60726=>"010000110",
  60727=>"110000000",
  60728=>"100011111",
  60729=>"001101011",
  60730=>"010110001",
  60731=>"101100011",
  60732=>"001101110",
  60733=>"000111000",
  60734=>"000111110",
  60735=>"011001110",
  60736=>"011100101",
  60737=>"101111011",
  60738=>"011010010",
  60739=>"110100110",
  60740=>"111100001",
  60741=>"101110010",
  60742=>"111000001",
  60743=>"100000000",
  60744=>"001001001",
  60745=>"100010101",
  60746=>"010100010",
  60747=>"111100001",
  60748=>"011111011",
  60749=>"011101110",
  60750=>"001011011",
  60751=>"000111101",
  60752=>"110010000",
  60753=>"100100100",
  60754=>"110110110",
  60755=>"111000101",
  60756=>"100111110",
  60757=>"011111111",
  60758=>"000011100",
  60759=>"111111001",
  60760=>"001010000",
  60761=>"100001111",
  60762=>"001001100",
  60763=>"101010111",
  60764=>"000010111",
  60765=>"000100111",
  60766=>"111000010",
  60767=>"000000110",
  60768=>"001110111",
  60769=>"001000001",
  60770=>"100111101",
  60771=>"010010010",
  60772=>"001010100",
  60773=>"001010101",
  60774=>"110110001",
  60775=>"111110000",
  60776=>"100000110",
  60777=>"001010010",
  60778=>"000001101",
  60779=>"110110011",
  60780=>"110110010",
  60781=>"100100011",
  60782=>"000101100",
  60783=>"100001000",
  60784=>"110000011",
  60785=>"101001001",
  60786=>"011111101",
  60787=>"011110011",
  60788=>"100100011",
  60789=>"001001010",
  60790=>"000010011",
  60791=>"011111010",
  60792=>"000000111",
  60793=>"011110001",
  60794=>"100010000",
  60795=>"100011000",
  60796=>"110001101",
  60797=>"111100011",
  60798=>"100101000",
  60799=>"110000001",
  60800=>"001000001",
  60801=>"100111111",
  60802=>"101101101",
  60803=>"100001000",
  60804=>"111011101",
  60805=>"000011111",
  60806=>"001010101",
  60807=>"000001101",
  60808=>"110001100",
  60809=>"111001010",
  60810=>"001000010",
  60811=>"110001001",
  60812=>"000001010",
  60813=>"011001111",
  60814=>"000111111",
  60815=>"110000011",
  60816=>"011011110",
  60817=>"110010010",
  60818=>"011001001",
  60819=>"111010010",
  60820=>"100001001",
  60821=>"010010010",
  60822=>"110101000",
  60823=>"110111111",
  60824=>"111000100",
  60825=>"111111000",
  60826=>"011001100",
  60827=>"111111001",
  60828=>"111010111",
  60829=>"101100011",
  60830=>"001011001",
  60831=>"011111011",
  60832=>"010011101",
  60833=>"010100111",
  60834=>"110000111",
  60835=>"111111011",
  60836=>"111001111",
  60837=>"110110100",
  60838=>"100110100",
  60839=>"011100000",
  60840=>"000100011",
  60841=>"010110101",
  60842=>"010100000",
  60843=>"110111001",
  60844=>"011010001",
  60845=>"000011000",
  60846=>"110011000",
  60847=>"011010110",
  60848=>"001011011",
  60849=>"000010101",
  60850=>"010110110",
  60851=>"111001101",
  60852=>"111001011",
  60853=>"001110110",
  60854=>"000101000",
  60855=>"111101011",
  60856=>"000001001",
  60857=>"010100101",
  60858=>"101001010",
  60859=>"101000111",
  60860=>"101111010",
  60861=>"110011011",
  60862=>"111001111",
  60863=>"111101100",
  60864=>"101110001",
  60865=>"001100001",
  60866=>"001001111",
  60867=>"011100001",
  60868=>"101100111",
  60869=>"001001101",
  60870=>"010100110",
  60871=>"100100111",
  60872=>"010110011",
  60873=>"101011010",
  60874=>"111101010",
  60875=>"001110001",
  60876=>"000101111",
  60877=>"010001011",
  60878=>"001000001",
  60879=>"100101110",
  60880=>"110110111",
  60881=>"100000000",
  60882=>"000010001",
  60883=>"101110001",
  60884=>"001111111",
  60885=>"010100000",
  60886=>"001011111",
  60887=>"110100010",
  60888=>"011011001",
  60889=>"111001101",
  60890=>"100000110",
  60891=>"000101011",
  60892=>"110111000",
  60893=>"100011001",
  60894=>"111101010",
  60895=>"011111000",
  60896=>"100100000",
  60897=>"011101101",
  60898=>"111111100",
  60899=>"001100000",
  60900=>"111010011",
  60901=>"101010011",
  60902=>"010010000",
  60903=>"011110011",
  60904=>"001111101",
  60905=>"001110110",
  60906=>"000110001",
  60907=>"111111111",
  60908=>"010011011",
  60909=>"110101111",
  60910=>"100100101",
  60911=>"101010100",
  60912=>"110010110",
  60913=>"100101001",
  60914=>"011010100",
  60915=>"000111001",
  60916=>"011101100",
  60917=>"100100000",
  60918=>"001011100",
  60919=>"111010001",
  60920=>"101011000",
  60921=>"000101110",
  60922=>"001110001",
  60923=>"000001101",
  60924=>"110111011",
  60925=>"100011111",
  60926=>"001010000",
  60927=>"001110100",
  60928=>"011001010",
  60929=>"010100101",
  60930=>"110010111",
  60931=>"100101100",
  60932=>"111100011",
  60933=>"110000000",
  60934=>"111010111",
  60935=>"101001010",
  60936=>"110001001",
  60937=>"110000011",
  60938=>"101000010",
  60939=>"010010000",
  60940=>"101010101",
  60941=>"111100000",
  60942=>"111110000",
  60943=>"000101011",
  60944=>"100001011",
  60945=>"000110111",
  60946=>"111110000",
  60947=>"011100011",
  60948=>"110111000",
  60949=>"010000000",
  60950=>"011110111",
  60951=>"100001101",
  60952=>"000100010",
  60953=>"011010101",
  60954=>"000010000",
  60955=>"011001000",
  60956=>"001101101",
  60957=>"001011111",
  60958=>"100010110",
  60959=>"110000101",
  60960=>"010101100",
  60961=>"110100111",
  60962=>"110000001",
  60963=>"101011111",
  60964=>"101001111",
  60965=>"111110011",
  60966=>"100011110",
  60967=>"100100101",
  60968=>"011011110",
  60969=>"011101001",
  60970=>"100001010",
  60971=>"110110000",
  60972=>"101100100",
  60973=>"000001101",
  60974=>"101110000",
  60975=>"010000100",
  60976=>"000011000",
  60977=>"110101001",
  60978=>"000101010",
  60979=>"111110001",
  60980=>"001001111",
  60981=>"001010010",
  60982=>"100010011",
  60983=>"000101111",
  60984=>"000011000",
  60985=>"000100000",
  60986=>"001001000",
  60987=>"101000110",
  60988=>"010100110",
  60989=>"001000111",
  60990=>"101100110",
  60991=>"111111101",
  60992=>"001101000",
  60993=>"101100110",
  60994=>"111010001",
  60995=>"010111001",
  60996=>"010011011",
  60997=>"011110001",
  60998=>"000001100",
  60999=>"010011101",
  61000=>"001001110",
  61001=>"000111011",
  61002=>"110101100",
  61003=>"100011010",
  61004=>"111111010",
  61005=>"110100000",
  61006=>"111000101",
  61007=>"001011011",
  61008=>"000000111",
  61009=>"111011110",
  61010=>"011101101",
  61011=>"111011101",
  61012=>"001101000",
  61013=>"110110000",
  61014=>"001100001",
  61015=>"000101010",
  61016=>"011010111",
  61017=>"111110000",
  61018=>"010011111",
  61019=>"101101001",
  61020=>"110011100",
  61021=>"011011001",
  61022=>"101011000",
  61023=>"101010011",
  61024=>"011110110",
  61025=>"011011001",
  61026=>"110010111",
  61027=>"001100101",
  61028=>"011100000",
  61029=>"001100101",
  61030=>"001000101",
  61031=>"111000010",
  61032=>"001100001",
  61033=>"101001000",
  61034=>"000000111",
  61035=>"000100101",
  61036=>"101101000",
  61037=>"000011011",
  61038=>"000010010",
  61039=>"011010110",
  61040=>"101101010",
  61041=>"111000000",
  61042=>"100111000",
  61043=>"101100110",
  61044=>"100110101",
  61045=>"010111100",
  61046=>"011000010",
  61047=>"010000100",
  61048=>"111110001",
  61049=>"110101000",
  61050=>"101100111",
  61051=>"001001101",
  61052=>"001011001",
  61053=>"001000000",
  61054=>"010001100",
  61055=>"010110110",
  61056=>"001010111",
  61057=>"011001011",
  61058=>"110111011",
  61059=>"011101100",
  61060=>"100000000",
  61061=>"010111011",
  61062=>"110101101",
  61063=>"110110000",
  61064=>"011111110",
  61065=>"011110011",
  61066=>"011111011",
  61067=>"010111000",
  61068=>"111100111",
  61069=>"111111010",
  61070=>"111001010",
  61071=>"111011101",
  61072=>"001101110",
  61073=>"001110111",
  61074=>"000111001",
  61075=>"010110110",
  61076=>"000110000",
  61077=>"100100000",
  61078=>"001110110",
  61079=>"000010000",
  61080=>"111001000",
  61081=>"000000100",
  61082=>"011110101",
  61083=>"010010010",
  61084=>"101100010",
  61085=>"000100110",
  61086=>"100011100",
  61087=>"100001110",
  61088=>"101010111",
  61089=>"000011100",
  61090=>"000011001",
  61091=>"001011001",
  61092=>"100000010",
  61093=>"001101001",
  61094=>"011101100",
  61095=>"000010001",
  61096=>"011100010",
  61097=>"101111011",
  61098=>"001110111",
  61099=>"000001101",
  61100=>"001110011",
  61101=>"100000100",
  61102=>"100110111",
  61103=>"111010000",
  61104=>"000010111",
  61105=>"010010111",
  61106=>"111100010",
  61107=>"110101111",
  61108=>"100000011",
  61109=>"101001110",
  61110=>"000011111",
  61111=>"000110010",
  61112=>"000010101",
  61113=>"101111010",
  61114=>"111010011",
  61115=>"011000001",
  61116=>"100110011",
  61117=>"011100000",
  61118=>"101101011",
  61119=>"100100100",
  61120=>"001000001",
  61121=>"000110111",
  61122=>"001000010",
  61123=>"000111010",
  61124=>"111111001",
  61125=>"001011001",
  61126=>"011100111",
  61127=>"001101100",
  61128=>"101000011",
  61129=>"010101110",
  61130=>"100110000",
  61131=>"001011000",
  61132=>"000010011",
  61133=>"000011000",
  61134=>"000001110",
  61135=>"111010111",
  61136=>"000100010",
  61137=>"110101101",
  61138=>"000100100",
  61139=>"000100011",
  61140=>"010011101",
  61141=>"100000101",
  61142=>"000101101",
  61143=>"001101010",
  61144=>"110110111",
  61145=>"111010100",
  61146=>"000000001",
  61147=>"101000000",
  61148=>"111001000",
  61149=>"000101001",
  61150=>"010111100",
  61151=>"010001111",
  61152=>"010100111",
  61153=>"000111101",
  61154=>"011110101",
  61155=>"110100110",
  61156=>"000011000",
  61157=>"001010110",
  61158=>"000000111",
  61159=>"110001100",
  61160=>"011100001",
  61161=>"100101010",
  61162=>"001101001",
  61163=>"100011101",
  61164=>"010100001",
  61165=>"001011011",
  61166=>"110110111",
  61167=>"010011111",
  61168=>"001010110",
  61169=>"011011001",
  61170=>"101100100",
  61171=>"010001100",
  61172=>"010100011",
  61173=>"000000111",
  61174=>"010111010",
  61175=>"000010100",
  61176=>"110101011",
  61177=>"101011001",
  61178=>"000011000",
  61179=>"111001000",
  61180=>"100101010",
  61181=>"110100001",
  61182=>"011000011",
  61183=>"000000111",
  61184=>"011111111",
  61185=>"011111100",
  61186=>"011011011",
  61187=>"000000110",
  61188=>"111010010",
  61189=>"010011010",
  61190=>"010000101",
  61191=>"010110010",
  61192=>"010011100",
  61193=>"000110011",
  61194=>"011001111",
  61195=>"110000011",
  61196=>"100010110",
  61197=>"010101101",
  61198=>"110100010",
  61199=>"001100011",
  61200=>"111100110",
  61201=>"010001000",
  61202=>"101100001",
  61203=>"001011101",
  61204=>"101010011",
  61205=>"000110111",
  61206=>"110100110",
  61207=>"001000101",
  61208=>"111011001",
  61209=>"110000101",
  61210=>"110001001",
  61211=>"001100011",
  61212=>"000111000",
  61213=>"101100101",
  61214=>"101001000",
  61215=>"000010110",
  61216=>"011110000",
  61217=>"100011100",
  61218=>"101110101",
  61219=>"010100010",
  61220=>"101111000",
  61221=>"000011000",
  61222=>"101000110",
  61223=>"000010110",
  61224=>"000010000",
  61225=>"110001111",
  61226=>"001001101",
  61227=>"110011011",
  61228=>"000001010",
  61229=>"001011000",
  61230=>"101101101",
  61231=>"100010001",
  61232=>"111110001",
  61233=>"010110001",
  61234=>"000111101",
  61235=>"011000110",
  61236=>"101000101",
  61237=>"110010100",
  61238=>"111000000",
  61239=>"110110101",
  61240=>"011010001",
  61241=>"110101010",
  61242=>"011101000",
  61243=>"000001001",
  61244=>"111000001",
  61245=>"000111010",
  61246=>"111001010",
  61247=>"010010110",
  61248=>"001010101",
  61249=>"011011010",
  61250=>"101001010",
  61251=>"000101000",
  61252=>"001011000",
  61253=>"101000001",
  61254=>"110000010",
  61255=>"100110101",
  61256=>"001000000",
  61257=>"000100100",
  61258=>"010101100",
  61259=>"110111110",
  61260=>"101000001",
  61261=>"000101010",
  61262=>"100010100",
  61263=>"100110101",
  61264=>"011111011",
  61265=>"001110001",
  61266=>"011001001",
  61267=>"000001101",
  61268=>"101101010",
  61269=>"011000010",
  61270=>"100101010",
  61271=>"000110001",
  61272=>"111001001",
  61273=>"111111100",
  61274=>"011011001",
  61275=>"110000000",
  61276=>"000101000",
  61277=>"011010100",
  61278=>"110000100",
  61279=>"010101101",
  61280=>"011110000",
  61281=>"111100111",
  61282=>"011000110",
  61283=>"010001111",
  61284=>"001101010",
  61285=>"000110100",
  61286=>"100011111",
  61287=>"111101001",
  61288=>"011111111",
  61289=>"100101110",
  61290=>"100111001",
  61291=>"001000111",
  61292=>"101111110",
  61293=>"011100110",
  61294=>"111101001",
  61295=>"011011101",
  61296=>"000111000",
  61297=>"001011001",
  61298=>"111111011",
  61299=>"001110001",
  61300=>"111110101",
  61301=>"000011001",
  61302=>"001110101",
  61303=>"010111111",
  61304=>"100111000",
  61305=>"100111010",
  61306=>"101110101",
  61307=>"100100010",
  61308=>"010011001",
  61309=>"100111100",
  61310=>"011011001",
  61311=>"111111010",
  61312=>"111011010",
  61313=>"011011100",
  61314=>"001011010",
  61315=>"010111111",
  61316=>"001000100",
  61317=>"000111101",
  61318=>"000100111",
  61319=>"101110010",
  61320=>"101000001",
  61321=>"001110101",
  61322=>"000100010",
  61323=>"101110111",
  61324=>"101100110",
  61325=>"110001111",
  61326=>"010010110",
  61327=>"000110011",
  61328=>"101101011",
  61329=>"111011111",
  61330=>"010010111",
  61331=>"100101111",
  61332=>"001011100",
  61333=>"100100010",
  61334=>"001100100",
  61335=>"010000000",
  61336=>"111111100",
  61337=>"010000011",
  61338=>"110111001",
  61339=>"001101010",
  61340=>"011110101",
  61341=>"110101010",
  61342=>"011001110",
  61343=>"100001101",
  61344=>"000110100",
  61345=>"010100111",
  61346=>"001101100",
  61347=>"101011100",
  61348=>"001010111",
  61349=>"010110010",
  61350=>"011100001",
  61351=>"101000110",
  61352=>"010010010",
  61353=>"000011101",
  61354=>"100011011",
  61355=>"111101001",
  61356=>"000101100",
  61357=>"010011101",
  61358=>"001000110",
  61359=>"101110000",
  61360=>"000110001",
  61361=>"111011000",
  61362=>"111011101",
  61363=>"111110011",
  61364=>"011111000",
  61365=>"101111110",
  61366=>"111110110",
  61367=>"111110111",
  61368=>"101110100",
  61369=>"001011110",
  61370=>"111011110",
  61371=>"100110111",
  61372=>"111100100",
  61373=>"110101100",
  61374=>"000000111",
  61375=>"110111111",
  61376=>"100110101",
  61377=>"100001010",
  61378=>"010001110",
  61379=>"000010010",
  61380=>"111001100",
  61381=>"110101101",
  61382=>"001000110",
  61383=>"011100101",
  61384=>"100111101",
  61385=>"000000001",
  61386=>"110101111",
  61387=>"000110000",
  61388=>"000110001",
  61389=>"111001101",
  61390=>"111111111",
  61391=>"011110111",
  61392=>"000010000",
  61393=>"110100001",
  61394=>"000110100",
  61395=>"100110010",
  61396=>"000110010",
  61397=>"001010111",
  61398=>"011111101",
  61399=>"111011101",
  61400=>"111111100",
  61401=>"100011100",
  61402=>"101110011",
  61403=>"110010110",
  61404=>"101011000",
  61405=>"101000111",
  61406=>"100100111",
  61407=>"010000000",
  61408=>"011110110",
  61409=>"101000011",
  61410=>"111000111",
  61411=>"000000001",
  61412=>"110101001",
  61413=>"111000011",
  61414=>"001001110",
  61415=>"100110110",
  61416=>"000010100",
  61417=>"000110001",
  61418=>"110011010",
  61419=>"000111001",
  61420=>"101010001",
  61421=>"011101011",
  61422=>"100111101",
  61423=>"001111110",
  61424=>"101010001",
  61425=>"000111010",
  61426=>"100001001",
  61427=>"001011100",
  61428=>"110101011",
  61429=>"101111111",
  61430=>"010010000",
  61431=>"111011111",
  61432=>"001001011",
  61433=>"100001011",
  61434=>"111011011",
  61435=>"100001010",
  61436=>"111111111",
  61437=>"000101110",
  61438=>"010111101",
  61439=>"100101111",
  61440=>"000111011",
  61441=>"111111111",
  61442=>"010101001",
  61443=>"011110111",
  61444=>"110011101",
  61445=>"111111010",
  61446=>"100111111",
  61447=>"111110101",
  61448=>"001011011",
  61449=>"101101010",
  61450=>"010101011",
  61451=>"000000110",
  61452=>"110010100",
  61453=>"011010010",
  61454=>"011001000",
  61455=>"001111110",
  61456=>"001100111",
  61457=>"110000101",
  61458=>"101110001",
  61459=>"011011100",
  61460=>"001011111",
  61461=>"101011000",
  61462=>"000100000",
  61463=>"001010000",
  61464=>"111011101",
  61465=>"100010111",
  61466=>"110001110",
  61467=>"011000000",
  61468=>"000111010",
  61469=>"111011111",
  61470=>"010110000",
  61471=>"001101001",
  61472=>"011100011",
  61473=>"011010000",
  61474=>"110101011",
  61475=>"000001111",
  61476=>"011010100",
  61477=>"010000110",
  61478=>"000010010",
  61479=>"101111111",
  61480=>"001010111",
  61481=>"110011010",
  61482=>"011100100",
  61483=>"101000001",
  61484=>"100001111",
  61485=>"000000011",
  61486=>"001100111",
  61487=>"110101011",
  61488=>"100101111",
  61489=>"111010000",
  61490=>"011111100",
  61491=>"011111110",
  61492=>"111001100",
  61493=>"011011011",
  61494=>"000000001",
  61495=>"001010001",
  61496=>"000101111",
  61497=>"100001010",
  61498=>"101111111",
  61499=>"000110101",
  61500=>"101110011",
  61501=>"001001000",
  61502=>"110101110",
  61503=>"001000001",
  61504=>"001101110",
  61505=>"010110000",
  61506=>"110111100",
  61507=>"000000001",
  61508=>"001110111",
  61509=>"010001011",
  61510=>"001010001",
  61511=>"101110001",
  61512=>"010010001",
  61513=>"110010010",
  61514=>"000100111",
  61515=>"101001100",
  61516=>"011100001",
  61517=>"011111010",
  61518=>"001000010",
  61519=>"101111000",
  61520=>"001010100",
  61521=>"000100110",
  61522=>"101000001",
  61523=>"111010111",
  61524=>"010110111",
  61525=>"011110010",
  61526=>"101111101",
  61527=>"101111000",
  61528=>"000101110",
  61529=>"111110110",
  61530=>"110000101",
  61531=>"000110111",
  61532=>"001100100",
  61533=>"011001111",
  61534=>"100111001",
  61535=>"101011000",
  61536=>"000100000",
  61537=>"011011010",
  61538=>"111000010",
  61539=>"000011111",
  61540=>"100000101",
  61541=>"100100110",
  61542=>"010011001",
  61543=>"110011010",
  61544=>"001000001",
  61545=>"001101101",
  61546=>"001110011",
  61547=>"100100111",
  61548=>"111100000",
  61549=>"000000010",
  61550=>"010010100",
  61551=>"001000100",
  61552=>"011011000",
  61553=>"001011110",
  61554=>"111000001",
  61555=>"100111010",
  61556=>"000001000",
  61557=>"010000000",
  61558=>"111000011",
  61559=>"100011111",
  61560=>"011000000",
  61561=>"111000001",
  61562=>"011011110",
  61563=>"111001101",
  61564=>"110000010",
  61565=>"111110011",
  61566=>"111000010",
  61567=>"001000111",
  61568=>"100101110",
  61569=>"111100110",
  61570=>"010100001",
  61571=>"011000001",
  61572=>"100001000",
  61573=>"001101111",
  61574=>"011101111",
  61575=>"111011100",
  61576=>"001000000",
  61577=>"011011110",
  61578=>"111100110",
  61579=>"000100011",
  61580=>"110101101",
  61581=>"000101000",
  61582=>"101110100",
  61583=>"011001011",
  61584=>"000110111",
  61585=>"111100111",
  61586=>"101010010",
  61587=>"100101101",
  61588=>"100111011",
  61589=>"111010111",
  61590=>"101101110",
  61591=>"110010100",
  61592=>"110001010",
  61593=>"010111111",
  61594=>"010100001",
  61595=>"010100110",
  61596=>"110011011",
  61597=>"000011111",
  61598=>"110110011",
  61599=>"011100101",
  61600=>"101001011",
  61601=>"111010001",
  61602=>"110011001",
  61603=>"001010001",
  61604=>"011101000",
  61605=>"111101000",
  61606=>"111101111",
  61607=>"011100000",
  61608=>"010001101",
  61609=>"100001011",
  61610=>"011111001",
  61611=>"011110101",
  61612=>"101001000",
  61613=>"010011110",
  61614=>"001000100",
  61615=>"110100011",
  61616=>"011101100",
  61617=>"011000000",
  61618=>"100100010",
  61619=>"101101110",
  61620=>"100100100",
  61621=>"100000000",
  61622=>"100110111",
  61623=>"110101011",
  61624=>"111010011",
  61625=>"101111101",
  61626=>"101010010",
  61627=>"011100101",
  61628=>"011111000",
  61629=>"000111000",
  61630=>"110010111",
  61631=>"011010110",
  61632=>"000101011",
  61633=>"101110100",
  61634=>"001001000",
  61635=>"110100010",
  61636=>"000110110",
  61637=>"111011101",
  61638=>"011001100",
  61639=>"101011011",
  61640=>"011111010",
  61641=>"011110101",
  61642=>"100111001",
  61643=>"001011110",
  61644=>"110111010",
  61645=>"100000010",
  61646=>"000111111",
  61647=>"110110110",
  61648=>"001111101",
  61649=>"110000110",
  61650=>"110101011",
  61651=>"110111000",
  61652=>"100000100",
  61653=>"100011011",
  61654=>"011111001",
  61655=>"110101011",
  61656=>"001101101",
  61657=>"100101111",
  61658=>"001111110",
  61659=>"011100100",
  61660=>"000111010",
  61661=>"000110111",
  61662=>"000110011",
  61663=>"001110110",
  61664=>"111100111",
  61665=>"011111001",
  61666=>"000011011",
  61667=>"000000110",
  61668=>"011110011",
  61669=>"011101000",
  61670=>"001010010",
  61671=>"010010010",
  61672=>"011000011",
  61673=>"111100101",
  61674=>"010011100",
  61675=>"101101101",
  61676=>"001110111",
  61677=>"110111011",
  61678=>"111011110",
  61679=>"111111001",
  61680=>"110011110",
  61681=>"110010001",
  61682=>"111111000",
  61683=>"000110010",
  61684=>"001011100",
  61685=>"111000111",
  61686=>"101100010",
  61687=>"000001010",
  61688=>"110001111",
  61689=>"001001000",
  61690=>"100100111",
  61691=>"100001001",
  61692=>"001001101",
  61693=>"111111100",
  61694=>"000010100",
  61695=>"111111000",
  61696=>"111110110",
  61697=>"000111101",
  61698=>"011000000",
  61699=>"010000101",
  61700=>"001010000",
  61701=>"001111101",
  61702=>"100101010",
  61703=>"010011101",
  61704=>"111010000",
  61705=>"011000100",
  61706=>"100010001",
  61707=>"001100110",
  61708=>"101100111",
  61709=>"110101001",
  61710=>"110100000",
  61711=>"100100010",
  61712=>"001000000",
  61713=>"011100101",
  61714=>"000010110",
  61715=>"111010100",
  61716=>"101000101",
  61717=>"001001011",
  61718=>"000101001",
  61719=>"001100001",
  61720=>"011101001",
  61721=>"000101000",
  61722=>"000011011",
  61723=>"000110010",
  61724=>"100101001",
  61725=>"011000111",
  61726=>"010001011",
  61727=>"110110111",
  61728=>"100011010",
  61729=>"010010100",
  61730=>"001011111",
  61731=>"100011100",
  61732=>"000101111",
  61733=>"111101100",
  61734=>"101010110",
  61735=>"000000010",
  61736=>"111010101",
  61737=>"100010001",
  61738=>"000000001",
  61739=>"101100111",
  61740=>"011001010",
  61741=>"101011111",
  61742=>"010100001",
  61743=>"110100000",
  61744=>"111000110",
  61745=>"101110001",
  61746=>"111011111",
  61747=>"110011110",
  61748=>"010110000",
  61749=>"000100000",
  61750=>"101100100",
  61751=>"001100100",
  61752=>"000010111",
  61753=>"001100010",
  61754=>"111101101",
  61755=>"111110111",
  61756=>"110010001",
  61757=>"011100000",
  61758=>"010100101",
  61759=>"011000000",
  61760=>"111111110",
  61761=>"010000001",
  61762=>"010110000",
  61763=>"001000100",
  61764=>"101101010",
  61765=>"110001111",
  61766=>"101000010",
  61767=>"001100100",
  61768=>"101011110",
  61769=>"111011110",
  61770=>"010001010",
  61771=>"000111110",
  61772=>"000001000",
  61773=>"100100111",
  61774=>"110101110",
  61775=>"100111111",
  61776=>"001111100",
  61777=>"001111010",
  61778=>"111100001",
  61779=>"100111101",
  61780=>"101100111",
  61781=>"010100100",
  61782=>"111100011",
  61783=>"001111110",
  61784=>"111101000",
  61785=>"111110100",
  61786=>"010101100",
  61787=>"110111100",
  61788=>"010100001",
  61789=>"101100011",
  61790=>"111101100",
  61791=>"001011110",
  61792=>"100110010",
  61793=>"010110000",
  61794=>"010000001",
  61795=>"111111000",
  61796=>"100000001",
  61797=>"011111100",
  61798=>"101000000",
  61799=>"110001101",
  61800=>"011011011",
  61801=>"000001100",
  61802=>"010011110",
  61803=>"000111111",
  61804=>"010011100",
  61805=>"011111000",
  61806=>"110100000",
  61807=>"100011001",
  61808=>"010001001",
  61809=>"000001000",
  61810=>"100001011",
  61811=>"001000011",
  61812=>"000101011",
  61813=>"010001111",
  61814=>"000110011",
  61815=>"000010111",
  61816=>"111010010",
  61817=>"111010110",
  61818=>"000011101",
  61819=>"010001001",
  61820=>"011100010",
  61821=>"001011001",
  61822=>"101011110",
  61823=>"010100010",
  61824=>"100101111",
  61825=>"010111100",
  61826=>"110000100",
  61827=>"111001010",
  61828=>"000101100",
  61829=>"001001001",
  61830=>"011000010",
  61831=>"000110110",
  61832=>"000011100",
  61833=>"000110101",
  61834=>"001110011",
  61835=>"111100001",
  61836=>"101110010",
  61837=>"110000001",
  61838=>"000011100",
  61839=>"011101101",
  61840=>"010101110",
  61841=>"110101110",
  61842=>"111010111",
  61843=>"100011001",
  61844=>"000001010",
  61845=>"111010001",
  61846=>"100111101",
  61847=>"001000110",
  61848=>"100101111",
  61849=>"111111110",
  61850=>"000100100",
  61851=>"001111111",
  61852=>"000011000",
  61853=>"001010011",
  61854=>"010000110",
  61855=>"001001001",
  61856=>"101111100",
  61857=>"010111110",
  61858=>"010000011",
  61859=>"110110110",
  61860=>"000001001",
  61861=>"101000001",
  61862=>"000000101",
  61863=>"011011110",
  61864=>"000000100",
  61865=>"011000111",
  61866=>"111110000",
  61867=>"010000111",
  61868=>"101010101",
  61869=>"010100100",
  61870=>"111010011",
  61871=>"100011001",
  61872=>"010001101",
  61873=>"110111001",
  61874=>"000001111",
  61875=>"101111101",
  61876=>"111011011",
  61877=>"000110010",
  61878=>"111010000",
  61879=>"100000010",
  61880=>"001100001",
  61881=>"000101011",
  61882=>"110000001",
  61883=>"111110100",
  61884=>"111111000",
  61885=>"011100001",
  61886=>"111110111",
  61887=>"110111001",
  61888=>"000001100",
  61889=>"001001110",
  61890=>"001010111",
  61891=>"001010000",
  61892=>"100001101",
  61893=>"011110100",
  61894=>"111101101",
  61895=>"101000000",
  61896=>"011001010",
  61897=>"010111111",
  61898=>"110111111",
  61899=>"111001101",
  61900=>"010111111",
  61901=>"101110111",
  61902=>"000100001",
  61903=>"101011100",
  61904=>"111011101",
  61905=>"011001010",
  61906=>"100011000",
  61907=>"110000000",
  61908=>"000100010",
  61909=>"011011111",
  61910=>"100001101",
  61911=>"000100101",
  61912=>"000110100",
  61913=>"001010010",
  61914=>"011011000",
  61915=>"000001111",
  61916=>"001011010",
  61917=>"000111011",
  61918=>"111000011",
  61919=>"111111100",
  61920=>"000110100",
  61921=>"001011110",
  61922=>"000101101",
  61923=>"111100110",
  61924=>"011000000",
  61925=>"000010001",
  61926=>"111000101",
  61927=>"100100000",
  61928=>"110100011",
  61929=>"111011100",
  61930=>"001111010",
  61931=>"001100111",
  61932=>"010000010",
  61933=>"011111011",
  61934=>"011101010",
  61935=>"111101000",
  61936=>"111111110",
  61937=>"011011011",
  61938=>"001111101",
  61939=>"001101101",
  61940=>"111101111",
  61941=>"110111000",
  61942=>"111000010",
  61943=>"100010010",
  61944=>"111101111",
  61945=>"010110011",
  61946=>"100110000",
  61947=>"010101010",
  61948=>"111101011",
  61949=>"010000110",
  61950=>"000101111",
  61951=>"001000001",
  61952=>"001110101",
  61953=>"000010101",
  61954=>"100011000",
  61955=>"110111010",
  61956=>"111010111",
  61957=>"000101000",
  61958=>"011011011",
  61959=>"010001011",
  61960=>"000000100",
  61961=>"011111111",
  61962=>"000000111",
  61963=>"101011010",
  61964=>"111110111",
  61965=>"101111000",
  61966=>"111110001",
  61967=>"111000110",
  61968=>"111100001",
  61969=>"001101011",
  61970=>"110011011",
  61971=>"111100101",
  61972=>"110101111",
  61973=>"000010001",
  61974=>"011101110",
  61975=>"000000001",
  61976=>"110011000",
  61977=>"101110110",
  61978=>"101100000",
  61979=>"111001111",
  61980=>"001110001",
  61981=>"010010001",
  61982=>"010101000",
  61983=>"111110001",
  61984=>"000111111",
  61985=>"011101111",
  61986=>"010110110",
  61987=>"100101111",
  61988=>"010110110",
  61989=>"011001001",
  61990=>"010100000",
  61991=>"000111011",
  61992=>"001000001",
  61993=>"011001000",
  61994=>"111111111",
  61995=>"110011100",
  61996=>"011111100",
  61997=>"101010111",
  61998=>"101010101",
  61999=>"011100100",
  62000=>"110101001",
  62001=>"000011000",
  62002=>"110100110",
  62003=>"111010111",
  62004=>"001110001",
  62005=>"101011011",
  62006=>"100111001",
  62007=>"011110111",
  62008=>"101111011",
  62009=>"000110100",
  62010=>"000110110",
  62011=>"101110010",
  62012=>"000100010",
  62013=>"111100111",
  62014=>"111111101",
  62015=>"000010011",
  62016=>"100001110",
  62017=>"110111110",
  62018=>"001111011",
  62019=>"011111011",
  62020=>"000001000",
  62021=>"111111010",
  62022=>"110101000",
  62023=>"001101100",
  62024=>"111110111",
  62025=>"111110000",
  62026=>"110111011",
  62027=>"010111110",
  62028=>"100100000",
  62029=>"000110000",
  62030=>"011010001",
  62031=>"010001101",
  62032=>"101010111",
  62033=>"100001111",
  62034=>"101111011",
  62035=>"101100101",
  62036=>"011001000",
  62037=>"001000111",
  62038=>"011101101",
  62039=>"000011000",
  62040=>"111101101",
  62041=>"011110111",
  62042=>"111110100",
  62043=>"010101001",
  62044=>"000001101",
  62045=>"101111111",
  62046=>"111100011",
  62047=>"000101100",
  62048=>"110111010",
  62049=>"010111000",
  62050=>"110110011",
  62051=>"001001101",
  62052=>"010111011",
  62053=>"110011100",
  62054=>"010111100",
  62055=>"110101101",
  62056=>"101011000",
  62057=>"100101101",
  62058=>"110100110",
  62059=>"110011101",
  62060=>"111110111",
  62061=>"111100100",
  62062=>"100010111",
  62063=>"011101110",
  62064=>"110011110",
  62065=>"001001111",
  62066=>"000110100",
  62067=>"000010101",
  62068=>"110111100",
  62069=>"001000001",
  62070=>"110111000",
  62071=>"000100110",
  62072=>"001101000",
  62073=>"010010000",
  62074=>"111001000",
  62075=>"001011001",
  62076=>"011011110",
  62077=>"001110010",
  62078=>"110011000",
  62079=>"001100111",
  62080=>"111111101",
  62081=>"001000100",
  62082=>"000000100",
  62083=>"000000100",
  62084=>"111101111",
  62085=>"100000011",
  62086=>"110011011",
  62087=>"110001101",
  62088=>"011010011",
  62089=>"000010011",
  62090=>"001010000",
  62091=>"010010010",
  62092=>"100010101",
  62093=>"111111010",
  62094=>"100000001",
  62095=>"011000011",
  62096=>"100111010",
  62097=>"100010000",
  62098=>"010011100",
  62099=>"111000110",
  62100=>"101101111",
  62101=>"011111110",
  62102=>"100001010",
  62103=>"000110011",
  62104=>"110101100",
  62105=>"110010111",
  62106=>"010101011",
  62107=>"110111110",
  62108=>"010111101",
  62109=>"010100011",
  62110=>"111100111",
  62111=>"110110100",
  62112=>"010010101",
  62113=>"010101000",
  62114=>"001011111",
  62115=>"000000110",
  62116=>"001010111",
  62117=>"110110101",
  62118=>"111011001",
  62119=>"100111111",
  62120=>"100111111",
  62121=>"101111010",
  62122=>"101110001",
  62123=>"011100011",
  62124=>"101111000",
  62125=>"010100000",
  62126=>"100110010",
  62127=>"111011111",
  62128=>"010100111",
  62129=>"010001111",
  62130=>"000000110",
  62131=>"111111001",
  62132=>"000011001",
  62133=>"101101000",
  62134=>"100111011",
  62135=>"101010110",
  62136=>"110010001",
  62137=>"101110100",
  62138=>"100011000",
  62139=>"110100001",
  62140=>"100011011",
  62141=>"111111101",
  62142=>"100000000",
  62143=>"110010100",
  62144=>"000011001",
  62145=>"101011011",
  62146=>"101110110",
  62147=>"100010011",
  62148=>"000100111",
  62149=>"111001011",
  62150=>"010111010",
  62151=>"000001000",
  62152=>"010000100",
  62153=>"110011011",
  62154=>"110000000",
  62155=>"000000111",
  62156=>"110011111",
  62157=>"010010011",
  62158=>"101100101",
  62159=>"101110001",
  62160=>"110100010",
  62161=>"011000100",
  62162=>"111111011",
  62163=>"010010111",
  62164=>"000000001",
  62165=>"001110000",
  62166=>"001110101",
  62167=>"110011100",
  62168=>"100100010",
  62169=>"010011011",
  62170=>"110111111",
  62171=>"101111000",
  62172=>"111001101",
  62173=>"100111100",
  62174=>"111011010",
  62175=>"010010101",
  62176=>"111000010",
  62177=>"010000001",
  62178=>"110000110",
  62179=>"110001000",
  62180=>"100101111",
  62181=>"110111010",
  62182=>"001101111",
  62183=>"111000110",
  62184=>"011011000",
  62185=>"001010000",
  62186=>"101101000",
  62187=>"010011000",
  62188=>"111111001",
  62189=>"100011001",
  62190=>"101110100",
  62191=>"111001011",
  62192=>"010010010",
  62193=>"001111010",
  62194=>"111010011",
  62195=>"110101101",
  62196=>"011011001",
  62197=>"111110100",
  62198=>"111111101",
  62199=>"110011101",
  62200=>"110000100",
  62201=>"011011000",
  62202=>"111100100",
  62203=>"100010001",
  62204=>"001100011",
  62205=>"111010101",
  62206=>"000100010",
  62207=>"010001111",
  62208=>"111010100",
  62209=>"010100110",
  62210=>"011101000",
  62211=>"000010101",
  62212=>"101011001",
  62213=>"000010011",
  62214=>"011011011",
  62215=>"001000101",
  62216=>"101000000",
  62217=>"110011101",
  62218=>"111010010",
  62219=>"011111110",
  62220=>"111011000",
  62221=>"010011100",
  62222=>"000110011",
  62223=>"011110010",
  62224=>"100000111",
  62225=>"001110000",
  62226=>"110101010",
  62227=>"100110100",
  62228=>"111101001",
  62229=>"010101111",
  62230=>"001101101",
  62231=>"001001010",
  62232=>"100111101",
  62233=>"011000110",
  62234=>"001011001",
  62235=>"001000011",
  62236=>"110101110",
  62237=>"101010000",
  62238=>"110110110",
  62239=>"100000010",
  62240=>"011110010",
  62241=>"111110101",
  62242=>"010010001",
  62243=>"111100111",
  62244=>"100111010",
  62245=>"010100001",
  62246=>"110010100",
  62247=>"100110110",
  62248=>"101000100",
  62249=>"111100011",
  62250=>"000001101",
  62251=>"110000111",
  62252=>"000100001",
  62253=>"001011111",
  62254=>"000001010",
  62255=>"000000011",
  62256=>"101001100",
  62257=>"010101101",
  62258=>"010001110",
  62259=>"000110010",
  62260=>"010010110",
  62261=>"000000101",
  62262=>"111111100",
  62263=>"111011101",
  62264=>"100001010",
  62265=>"101010101",
  62266=>"000011111",
  62267=>"101101011",
  62268=>"110111110",
  62269=>"110110111",
  62270=>"111000110",
  62271=>"101010001",
  62272=>"111100101",
  62273=>"100011010",
  62274=>"110010110",
  62275=>"011010111",
  62276=>"011001000",
  62277=>"110101101",
  62278=>"010000000",
  62279=>"001110111",
  62280=>"001100100",
  62281=>"100000100",
  62282=>"011011110",
  62283=>"011110101",
  62284=>"101011100",
  62285=>"100000111",
  62286=>"011110110",
  62287=>"111111111",
  62288=>"000000101",
  62289=>"010000000",
  62290=>"011011110",
  62291=>"101110100",
  62292=>"001100101",
  62293=>"000100111",
  62294=>"110011101",
  62295=>"110001101",
  62296=>"000110001",
  62297=>"011110011",
  62298=>"011111010",
  62299=>"010111111",
  62300=>"000111011",
  62301=>"111111111",
  62302=>"110100111",
  62303=>"000110111",
  62304=>"110110010",
  62305=>"010001110",
  62306=>"111101100",
  62307=>"011110011",
  62308=>"111010001",
  62309=>"001111011",
  62310=>"110110010",
  62311=>"111111101",
  62312=>"110110000",
  62313=>"111000101",
  62314=>"010000001",
  62315=>"000101010",
  62316=>"000111001",
  62317=>"110010100",
  62318=>"110111111",
  62319=>"010000110",
  62320=>"010011101",
  62321=>"000111011",
  62322=>"111011010",
  62323=>"100110110",
  62324=>"101111110",
  62325=>"010001101",
  62326=>"100111110",
  62327=>"011000101",
  62328=>"011110011",
  62329=>"111100110",
  62330=>"111110110",
  62331=>"110100001",
  62332=>"101100000",
  62333=>"110101010",
  62334=>"000010100",
  62335=>"010011011",
  62336=>"101010001",
  62337=>"010000000",
  62338=>"101101010",
  62339=>"100110010",
  62340=>"101000110",
  62341=>"001010011",
  62342=>"100100010",
  62343=>"010110011",
  62344=>"100001110",
  62345=>"110000100",
  62346=>"100000011",
  62347=>"000011011",
  62348=>"100011100",
  62349=>"011110111",
  62350=>"010100100",
  62351=>"011000110",
  62352=>"010100011",
  62353=>"100010100",
  62354=>"001001000",
  62355=>"000111001",
  62356=>"011000100",
  62357=>"111001001",
  62358=>"100110101",
  62359=>"110101100",
  62360=>"111110110",
  62361=>"010010000",
  62362=>"000001011",
  62363=>"111010111",
  62364=>"100010101",
  62365=>"111110010",
  62366=>"001111000",
  62367=>"001101001",
  62368=>"001010110",
  62369=>"100011001",
  62370=>"000110111",
  62371=>"011000111",
  62372=>"001100111",
  62373=>"011101011",
  62374=>"110010111",
  62375=>"000011110",
  62376=>"111110000",
  62377=>"000000000",
  62378=>"110011111",
  62379=>"011001111",
  62380=>"001101100",
  62381=>"101000001",
  62382=>"010101000",
  62383=>"001111101",
  62384=>"100111011",
  62385=>"000000100",
  62386=>"011010010",
  62387=>"000011111",
  62388=>"001011001",
  62389=>"110101110",
  62390=>"010000101",
  62391=>"001001011",
  62392=>"101111111",
  62393=>"010110101",
  62394=>"001110111",
  62395=>"010010101",
  62396=>"111000010",
  62397=>"110010010",
  62398=>"011111111",
  62399=>"011101101",
  62400=>"001000110",
  62401=>"110111011",
  62402=>"101000100",
  62403=>"001000101",
  62404=>"000000000",
  62405=>"110011111",
  62406=>"010001000",
  62407=>"110000001",
  62408=>"011100010",
  62409=>"000111101",
  62410=>"000110010",
  62411=>"101101011",
  62412=>"111000010",
  62413=>"010001111",
  62414=>"100110001",
  62415=>"110100101",
  62416=>"111000100",
  62417=>"011111011",
  62418=>"111101111",
  62419=>"100110010",
  62420=>"101111111",
  62421=>"111000010",
  62422=>"000000110",
  62423=>"000001110",
  62424=>"111100001",
  62425=>"100100101",
  62426=>"000010101",
  62427=>"110010101",
  62428=>"000011101",
  62429=>"100101010",
  62430=>"100000101",
  62431=>"111000000",
  62432=>"011101000",
  62433=>"111100010",
  62434=>"010000100",
  62435=>"010000111",
  62436=>"100111110",
  62437=>"111100111",
  62438=>"001011111",
  62439=>"101111100",
  62440=>"110101010",
  62441=>"111010111",
  62442=>"010010100",
  62443=>"111110100",
  62444=>"111000001",
  62445=>"001101110",
  62446=>"001011111",
  62447=>"010011010",
  62448=>"110100010",
  62449=>"101000101",
  62450=>"111001010",
  62451=>"001001110",
  62452=>"101000101",
  62453=>"101111000",
  62454=>"110110110",
  62455=>"100100000",
  62456=>"101000010",
  62457=>"100000001",
  62458=>"101010011",
  62459=>"100111111",
  62460=>"110110000",
  62461=>"000010010",
  62462=>"001001000",
  62463=>"110011111",
  62464=>"011000011",
  62465=>"001011010",
  62466=>"101001000",
  62467=>"000101010",
  62468=>"110110001",
  62469=>"001110000",
  62470=>"000000001",
  62471=>"111100111",
  62472=>"001100100",
  62473=>"010110101",
  62474=>"101010001",
  62475=>"000101100",
  62476=>"000001001",
  62477=>"001000011",
  62478=>"110011110",
  62479=>"011010111",
  62480=>"101111011",
  62481=>"001000011",
  62482=>"011101010",
  62483=>"110010001",
  62484=>"101111101",
  62485=>"110101011",
  62486=>"101010001",
  62487=>"001000001",
  62488=>"010000101",
  62489=>"110001011",
  62490=>"000010000",
  62491=>"001000011",
  62492=>"111001110",
  62493=>"110100111",
  62494=>"111001100",
  62495=>"010000011",
  62496=>"011100101",
  62497=>"010110010",
  62498=>"011101100",
  62499=>"011001000",
  62500=>"010001111",
  62501=>"100010101",
  62502=>"000000001",
  62503=>"011001101",
  62504=>"010001110",
  62505=>"101011000",
  62506=>"001101111",
  62507=>"001110011",
  62508=>"100001011",
  62509=>"000000111",
  62510=>"000000101",
  62511=>"000101011",
  62512=>"110110000",
  62513=>"000110111",
  62514=>"101101000",
  62515=>"101000110",
  62516=>"011101100",
  62517=>"011110011",
  62518=>"011010000",
  62519=>"110110000",
  62520=>"000000000",
  62521=>"111011001",
  62522=>"101111011",
  62523=>"100100011",
  62524=>"111000111",
  62525=>"100010001",
  62526=>"111001010",
  62527=>"000010101",
  62528=>"101110100",
  62529=>"001010100",
  62530=>"100010000",
  62531=>"110010110",
  62532=>"110111010",
  62533=>"000111101",
  62534=>"011101011",
  62535=>"000101010",
  62536=>"100111011",
  62537=>"001110011",
  62538=>"010101111",
  62539=>"010101100",
  62540=>"001110100",
  62541=>"011111001",
  62542=>"111000011",
  62543=>"111100111",
  62544=>"010101001",
  62545=>"001101011",
  62546=>"110110110",
  62547=>"101101111",
  62548=>"101011000",
  62549=>"011010000",
  62550=>"011001000",
  62551=>"010111110",
  62552=>"011001010",
  62553=>"110100011",
  62554=>"001001100",
  62555=>"000010101",
  62556=>"000101010",
  62557=>"000100011",
  62558=>"001000010",
  62559=>"000001011",
  62560=>"010101110",
  62561=>"001100111",
  62562=>"101110010",
  62563=>"111001001",
  62564=>"001000001",
  62565=>"010010110",
  62566=>"101111111",
  62567=>"000001000",
  62568=>"010110010",
  62569=>"110100111",
  62570=>"001001100",
  62571=>"101110011",
  62572=>"011110101",
  62573=>"001010110",
  62574=>"111101001",
  62575=>"000000001",
  62576=>"100010101",
  62577=>"000010111",
  62578=>"111011100",
  62579=>"101011010",
  62580=>"011011101",
  62581=>"110100010",
  62582=>"000010000",
  62583=>"110101101",
  62584=>"011010101",
  62585=>"011001001",
  62586=>"110101100",
  62587=>"110000110",
  62588=>"011010111",
  62589=>"100111000",
  62590=>"000000101",
  62591=>"101010110",
  62592=>"010100001",
  62593=>"100111011",
  62594=>"110110111",
  62595=>"100110011",
  62596=>"011011000",
  62597=>"001010011",
  62598=>"100011011",
  62599=>"110010001",
  62600=>"010010000",
  62601=>"101011011",
  62602=>"011100100",
  62603=>"100111101",
  62604=>"011100000",
  62605=>"010001111",
  62606=>"111010001",
  62607=>"001011011",
  62608=>"000111110",
  62609=>"001101100",
  62610=>"111001000",
  62611=>"100011000",
  62612=>"010010010",
  62613=>"101011101",
  62614=>"101001011",
  62615=>"101010000",
  62616=>"111010111",
  62617=>"010111111",
  62618=>"010111100",
  62619=>"001000001",
  62620=>"001001100",
  62621=>"011111010",
  62622=>"111010110",
  62623=>"000110101",
  62624=>"011010010",
  62625=>"110011010",
  62626=>"110010111",
  62627=>"000001011",
  62628=>"010111011",
  62629=>"101111100",
  62630=>"001010011",
  62631=>"011001110",
  62632=>"111001000",
  62633=>"100001010",
  62634=>"010010101",
  62635=>"100110000",
  62636=>"111011111",
  62637=>"111100000",
  62638=>"101010111",
  62639=>"110011100",
  62640=>"011000100",
  62641=>"001001011",
  62642=>"010110110",
  62643=>"110001110",
  62644=>"010101010",
  62645=>"001011100",
  62646=>"110110010",
  62647=>"101010001",
  62648=>"010001000",
  62649=>"110010011",
  62650=>"010110010",
  62651=>"001110010",
  62652=>"100110011",
  62653=>"000100111",
  62654=>"011011100",
  62655=>"000010111",
  62656=>"111111110",
  62657=>"100111000",
  62658=>"011001101",
  62659=>"111110001",
  62660=>"000001010",
  62661=>"100000111",
  62662=>"101101011",
  62663=>"001000110",
  62664=>"100000101",
  62665=>"001110100",
  62666=>"000111100",
  62667=>"100010010",
  62668=>"100111000",
  62669=>"011100010",
  62670=>"010010000",
  62671=>"110011100",
  62672=>"011100000",
  62673=>"100100110",
  62674=>"000010001",
  62675=>"110001111",
  62676=>"111000111",
  62677=>"110011011",
  62678=>"001000000",
  62679=>"110111110",
  62680=>"110101011",
  62681=>"110001101",
  62682=>"000101111",
  62683=>"100001000",
  62684=>"001111011",
  62685=>"110101111",
  62686=>"110101110",
  62687=>"010010000",
  62688=>"010001001",
  62689=>"111000101",
  62690=>"110011101",
  62691=>"010001000",
  62692=>"010101110",
  62693=>"000001110",
  62694=>"001000000",
  62695=>"111010010",
  62696=>"000011100",
  62697=>"011100101",
  62698=>"000100111",
  62699=>"111010101",
  62700=>"010001010",
  62701=>"000011000",
  62702=>"011111011",
  62703=>"001101111",
  62704=>"111110011",
  62705=>"010100011",
  62706=>"101011101",
  62707=>"001110011",
  62708=>"100000010",
  62709=>"100010110",
  62710=>"011001110",
  62711=>"000100000",
  62712=>"010101000",
  62713=>"110100000",
  62714=>"010000100",
  62715=>"101000101",
  62716=>"010100110",
  62717=>"101000010",
  62718=>"001101110",
  62719=>"000010100",
  62720=>"001100000",
  62721=>"100111111",
  62722=>"010111000",
  62723=>"010011101",
  62724=>"101010011",
  62725=>"100001111",
  62726=>"011111001",
  62727=>"110111101",
  62728=>"100101010",
  62729=>"011001111",
  62730=>"101101111",
  62731=>"011001101",
  62732=>"001010010",
  62733=>"010100101",
  62734=>"011110111",
  62735=>"001110001",
  62736=>"111000101",
  62737=>"111101000",
  62738=>"000001101",
  62739=>"010010110",
  62740=>"000100111",
  62741=>"001101000",
  62742=>"100100101",
  62743=>"111000111",
  62744=>"100110111",
  62745=>"110111001",
  62746=>"100100000",
  62747=>"111010010",
  62748=>"100110101",
  62749=>"010000010",
  62750=>"001010010",
  62751=>"111111000",
  62752=>"001000000",
  62753=>"110110101",
  62754=>"100010110",
  62755=>"000100101",
  62756=>"111000000",
  62757=>"110011111",
  62758=>"000011001",
  62759=>"010011111",
  62760=>"101100001",
  62761=>"100101010",
  62762=>"001001000",
  62763=>"110001001",
  62764=>"010011000",
  62765=>"001011011",
  62766=>"011100011",
  62767=>"111100001",
  62768=>"110011100",
  62769=>"011111110",
  62770=>"110111110",
  62771=>"010111010",
  62772=>"101110110",
  62773=>"001000100",
  62774=>"011111110",
  62775=>"110001100",
  62776=>"110101111",
  62777=>"011101010",
  62778=>"101001101",
  62779=>"010010010",
  62780=>"000010010",
  62781=>"101000010",
  62782=>"100110100",
  62783=>"000110010",
  62784=>"010010111",
  62785=>"010001111",
  62786=>"011110111",
  62787=>"010010101",
  62788=>"010100100",
  62789=>"100010110",
  62790=>"101110000",
  62791=>"110010110",
  62792=>"000011101",
  62793=>"111110001",
  62794=>"110100010",
  62795=>"010010100",
  62796=>"110011111",
  62797=>"100111110",
  62798=>"110110001",
  62799=>"100110111",
  62800=>"100000000",
  62801=>"001101101",
  62802=>"111101001",
  62803=>"010111010",
  62804=>"011111010",
  62805=>"000100000",
  62806=>"000000001",
  62807=>"001110000",
  62808=>"101000010",
  62809=>"001111010",
  62810=>"000001011",
  62811=>"100100000",
  62812=>"000111100",
  62813=>"000101001",
  62814=>"011101010",
  62815=>"000100101",
  62816=>"110001011",
  62817=>"110101110",
  62818=>"111101110",
  62819=>"011000100",
  62820=>"010010110",
  62821=>"011001001",
  62822=>"011111001",
  62823=>"111100110",
  62824=>"110001110",
  62825=>"111100010",
  62826=>"100110111",
  62827=>"100000010",
  62828=>"101001010",
  62829=>"001011111",
  62830=>"001110100",
  62831=>"101000011",
  62832=>"010000010",
  62833=>"010110110",
  62834=>"100001001",
  62835=>"100000010",
  62836=>"110101110",
  62837=>"000000100",
  62838=>"001100001",
  62839=>"010000100",
  62840=>"000100110",
  62841=>"001110001",
  62842=>"110000111",
  62843=>"101110100",
  62844=>"100011100",
  62845=>"011000010",
  62846=>"001110101",
  62847=>"110011000",
  62848=>"100100000",
  62849=>"011100110",
  62850=>"010100000",
  62851=>"100100001",
  62852=>"110110110",
  62853=>"110101000",
  62854=>"001000101",
  62855=>"001111001",
  62856=>"101101001",
  62857=>"001010000",
  62858=>"010001100",
  62859=>"101101110",
  62860=>"100000000",
  62861=>"000110000",
  62862=>"110011001",
  62863=>"111110011",
  62864=>"101110110",
  62865=>"010100001",
  62866=>"010000001",
  62867=>"000011101",
  62868=>"000001110",
  62869=>"001100101",
  62870=>"101010010",
  62871=>"110011101",
  62872=>"001101001",
  62873=>"000101110",
  62874=>"010011111",
  62875=>"000010111",
  62876=>"110100110",
  62877=>"001110010",
  62878=>"111110111",
  62879=>"011001010",
  62880=>"111100100",
  62881=>"001000010",
  62882=>"110001010",
  62883=>"001001010",
  62884=>"110010000",
  62885=>"100011000",
  62886=>"010011010",
  62887=>"110001011",
  62888=>"101001001",
  62889=>"011110101",
  62890=>"000100101",
  62891=>"111000000",
  62892=>"011100010",
  62893=>"000001110",
  62894=>"010010100",
  62895=>"001001001",
  62896=>"100011110",
  62897=>"000101000",
  62898=>"001110001",
  62899=>"100001110",
  62900=>"100110101",
  62901=>"110011100",
  62902=>"100000101",
  62903=>"111010100",
  62904=>"001010111",
  62905=>"010001011",
  62906=>"110111001",
  62907=>"011001101",
  62908=>"110011110",
  62909=>"010011001",
  62910=>"000100100",
  62911=>"101000011",
  62912=>"011011000",
  62913=>"110111111",
  62914=>"001011000",
  62915=>"001001011",
  62916=>"101000110",
  62917=>"011000000",
  62918=>"010001001",
  62919=>"101001001",
  62920=>"011100000",
  62921=>"111101001",
  62922=>"011000011",
  62923=>"100110000",
  62924=>"110010000",
  62925=>"100010001",
  62926=>"100001010",
  62927=>"001011110",
  62928=>"100111001",
  62929=>"011000110",
  62930=>"000110100",
  62931=>"000010111",
  62932=>"000011110",
  62933=>"101010011",
  62934=>"101101111",
  62935=>"111001100",
  62936=>"000111101",
  62937=>"100000011",
  62938=>"001001111",
  62939=>"101011011",
  62940=>"000110100",
  62941=>"000011011",
  62942=>"100011001",
  62943=>"010110000",
  62944=>"000000000",
  62945=>"110001111",
  62946=>"011110010",
  62947=>"110111111",
  62948=>"010001101",
  62949=>"110010011",
  62950=>"111111101",
  62951=>"100011001",
  62952=>"010110001",
  62953=>"101011010",
  62954=>"100111110",
  62955=>"010010111",
  62956=>"110111110",
  62957=>"011000110",
  62958=>"001011101",
  62959=>"101110110",
  62960=>"000100110",
  62961=>"110001111",
  62962=>"110010101",
  62963=>"100100001",
  62964=>"011111111",
  62965=>"001010000",
  62966=>"011011110",
  62967=>"010001101",
  62968=>"100011010",
  62969=>"001000010",
  62970=>"101001000",
  62971=>"010100111",
  62972=>"001101010",
  62973=>"111110111",
  62974=>"010011011",
  62975=>"100000000",
  62976=>"010001000",
  62977=>"011111001",
  62978=>"110000110",
  62979=>"000101100",
  62980=>"110011011",
  62981=>"111110100",
  62982=>"000100100",
  62983=>"101010001",
  62984=>"001000011",
  62985=>"000110001",
  62986=>"001101001",
  62987=>"001001101",
  62988=>"000010000",
  62989=>"110011101",
  62990=>"000100000",
  62991=>"000000110",
  62992=>"001010110",
  62993=>"001000000",
  62994=>"111100011",
  62995=>"011111000",
  62996=>"010001000",
  62997=>"011101100",
  62998=>"101111000",
  62999=>"110111001",
  63000=>"000011000",
  63001=>"101011111",
  63002=>"010000100",
  63003=>"111111000",
  63004=>"101001101",
  63005=>"110001010",
  63006=>"011010101",
  63007=>"001100000",
  63008=>"000110101",
  63009=>"111010111",
  63010=>"100011010",
  63011=>"101101010",
  63012=>"110011110",
  63013=>"101100110",
  63014=>"110110100",
  63015=>"000010001",
  63016=>"111110100",
  63017=>"101111000",
  63018=>"000101010",
  63019=>"011010111",
  63020=>"110000101",
  63021=>"100010110",
  63022=>"010100000",
  63023=>"111111111",
  63024=>"011010011",
  63025=>"010110010",
  63026=>"000010010",
  63027=>"100011011",
  63028=>"101010111",
  63029=>"110010000",
  63030=>"001110100",
  63031=>"110001110",
  63032=>"011011110",
  63033=>"000110100",
  63034=>"010001010",
  63035=>"100111111",
  63036=>"001011110",
  63037=>"000000010",
  63038=>"011010001",
  63039=>"101000111",
  63040=>"011111110",
  63041=>"111001010",
  63042=>"001011100",
  63043=>"110101010",
  63044=>"111111111",
  63045=>"001101010",
  63046=>"000110100",
  63047=>"000001001",
  63048=>"111101010",
  63049=>"101011100",
  63050=>"111000010",
  63051=>"011011101",
  63052=>"001000101",
  63053=>"011101010",
  63054=>"101011010",
  63055=>"111110101",
  63056=>"101011100",
  63057=>"110111010",
  63058=>"010011000",
  63059=>"111011011",
  63060=>"111001010",
  63061=>"100000001",
  63062=>"010100111",
  63063=>"011000100",
  63064=>"010111010",
  63065=>"001011100",
  63066=>"001000001",
  63067=>"000111101",
  63068=>"000101010",
  63069=>"000010100",
  63070=>"000111110",
  63071=>"101000101",
  63072=>"101101001",
  63073=>"000001001",
  63074=>"111001110",
  63075=>"110101011",
  63076=>"000101000",
  63077=>"001110011",
  63078=>"010001111",
  63079=>"000101000",
  63080=>"100010100",
  63081=>"010111100",
  63082=>"010100000",
  63083=>"001000001",
  63084=>"100000000",
  63085=>"010000011",
  63086=>"100001100",
  63087=>"110111110",
  63088=>"110111001",
  63089=>"101110100",
  63090=>"011111100",
  63091=>"100001101",
  63092=>"010000000",
  63093=>"000010000",
  63094=>"000111111",
  63095=>"100011011",
  63096=>"101000110",
  63097=>"001000110",
  63098=>"011001010",
  63099=>"100100011",
  63100=>"010111110",
  63101=>"100011111",
  63102=>"101000010",
  63103=>"100111011",
  63104=>"100111111",
  63105=>"011110010",
  63106=>"000100010",
  63107=>"011101001",
  63108=>"001111101",
  63109=>"001111110",
  63110=>"000001111",
  63111=>"101000001",
  63112=>"111100011",
  63113=>"011101101",
  63114=>"001101110",
  63115=>"110111001",
  63116=>"001000011",
  63117=>"100110011",
  63118=>"010001010",
  63119=>"100111010",
  63120=>"110011100",
  63121=>"011111111",
  63122=>"101110011",
  63123=>"110110100",
  63124=>"010111111",
  63125=>"000000110",
  63126=>"101011101",
  63127=>"101111100",
  63128=>"100101001",
  63129=>"100111100",
  63130=>"101011001",
  63131=>"110110110",
  63132=>"110000100",
  63133=>"001110001",
  63134=>"011101000",
  63135=>"001100010",
  63136=>"111001011",
  63137=>"111001000",
  63138=>"010011000",
  63139=>"011011101",
  63140=>"100010001",
  63141=>"101100011",
  63142=>"110101101",
  63143=>"001000110",
  63144=>"010100101",
  63145=>"100100011",
  63146=>"000110111",
  63147=>"110101100",
  63148=>"011110010",
  63149=>"100001001",
  63150=>"010001000",
  63151=>"001101101",
  63152=>"110000011",
  63153=>"101000101",
  63154=>"111101110",
  63155=>"100000100",
  63156=>"001101111",
  63157=>"110100100",
  63158=>"110111011",
  63159=>"011110000",
  63160=>"000111010",
  63161=>"000111010",
  63162=>"110111100",
  63163=>"101001111",
  63164=>"000001101",
  63165=>"000101110",
  63166=>"100000010",
  63167=>"000110101",
  63168=>"001010000",
  63169=>"000101100",
  63170=>"001100100",
  63171=>"111100001",
  63172=>"010111011",
  63173=>"101010100",
  63174=>"011110001",
  63175=>"010011010",
  63176=>"010110110",
  63177=>"110000010",
  63178=>"001011010",
  63179=>"001111100",
  63180=>"001001101",
  63181=>"111111100",
  63182=>"010011001",
  63183=>"100100111",
  63184=>"110001101",
  63185=>"011010011",
  63186=>"110110011",
  63187=>"100011001",
  63188=>"010011000",
  63189=>"111001100",
  63190=>"001101001",
  63191=>"111110000",
  63192=>"110000111",
  63193=>"011010110",
  63194=>"111010100",
  63195=>"011110011",
  63196=>"001110000",
  63197=>"101111010",
  63198=>"110101110",
  63199=>"010110100",
  63200=>"010000010",
  63201=>"111011110",
  63202=>"100110010",
  63203=>"010000100",
  63204=>"101011111",
  63205=>"111000000",
  63206=>"001011101",
  63207=>"110011010",
  63208=>"110011011",
  63209=>"011110000",
  63210=>"110111101",
  63211=>"001010101",
  63212=>"001000110",
  63213=>"010010110",
  63214=>"100010100",
  63215=>"010001101",
  63216=>"000100010",
  63217=>"101010000",
  63218=>"111000000",
  63219=>"100101010",
  63220=>"001110110",
  63221=>"000010010",
  63222=>"101111001",
  63223=>"101101101",
  63224=>"110111000",
  63225=>"011101000",
  63226=>"110110111",
  63227=>"111001001",
  63228=>"011110001",
  63229=>"010011101",
  63230=>"010101100",
  63231=>"111100100",
  63232=>"001111000",
  63233=>"010100001",
  63234=>"011011000",
  63235=>"010110110",
  63236=>"000110000",
  63237=>"010110111",
  63238=>"100110110",
  63239=>"000010101",
  63240=>"100111100",
  63241=>"110100001",
  63242=>"011101110",
  63243=>"001010001",
  63244=>"000000001",
  63245=>"101111011",
  63246=>"011111101",
  63247=>"111010111",
  63248=>"101010110",
  63249=>"011010100",
  63250=>"000110101",
  63251=>"011101111",
  63252=>"001010000",
  63253=>"001111000",
  63254=>"001110000",
  63255=>"110100010",
  63256=>"011001010",
  63257=>"110011110",
  63258=>"011101110",
  63259=>"010111001",
  63260=>"101100010",
  63261=>"110011101",
  63262=>"110001010",
  63263=>"011010111",
  63264=>"011011001",
  63265=>"111011111",
  63266=>"001101110",
  63267=>"000100010",
  63268=>"010110011",
  63269=>"001011100",
  63270=>"011110111",
  63271=>"100101001",
  63272=>"010011100",
  63273=>"111101010",
  63274=>"110010001",
  63275=>"010111011",
  63276=>"011101001",
  63277=>"111000111",
  63278=>"010011011",
  63279=>"000101100",
  63280=>"100000010",
  63281=>"100101001",
  63282=>"110111100",
  63283=>"100000011",
  63284=>"000001010",
  63285=>"001100111",
  63286=>"111100100",
  63287=>"011100000",
  63288=>"100100100",
  63289=>"100111011",
  63290=>"000011110",
  63291=>"100111010",
  63292=>"011100110",
  63293=>"001001010",
  63294=>"000010110",
  63295=>"110011011",
  63296=>"011110101",
  63297=>"000110111",
  63298=>"000111111",
  63299=>"001000010",
  63300=>"010111101",
  63301=>"000101011",
  63302=>"001011100",
  63303=>"010010100",
  63304=>"000000101",
  63305=>"010001101",
  63306=>"101110110",
  63307=>"001011110",
  63308=>"001110010",
  63309=>"011111100",
  63310=>"000001110",
  63311=>"110011100",
  63312=>"010110011",
  63313=>"000100100",
  63314=>"100011000",
  63315=>"111010001",
  63316=>"110011001",
  63317=>"010000010",
  63318=>"001100100",
  63319=>"110100111",
  63320=>"100011011",
  63321=>"100010100",
  63322=>"011000111",
  63323=>"111101101",
  63324=>"101000101",
  63325=>"010011010",
  63326=>"111001000",
  63327=>"011101011",
  63328=>"110011000",
  63329=>"000010000",
  63330=>"000000001",
  63331=>"011000011",
  63332=>"011000001",
  63333=>"110010001",
  63334=>"001001101",
  63335=>"010000111",
  63336=>"111010110",
  63337=>"001011010",
  63338=>"111011101",
  63339=>"010010011",
  63340=>"111011100",
  63341=>"100011001",
  63342=>"101001101",
  63343=>"110110001",
  63344=>"011110101",
  63345=>"000000010",
  63346=>"001100010",
  63347=>"000000010",
  63348=>"000011001",
  63349=>"000101000",
  63350=>"011001100",
  63351=>"111001001",
  63352=>"011101000",
  63353=>"001010010",
  63354=>"011000101",
  63355=>"111010111",
  63356=>"000110001",
  63357=>"101100000",
  63358=>"001011011",
  63359=>"010001111",
  63360=>"101100011",
  63361=>"010110000",
  63362=>"000111011",
  63363=>"001101001",
  63364=>"011100110",
  63365=>"000010001",
  63366=>"110111011",
  63367=>"000010100",
  63368=>"000111110",
  63369=>"111100010",
  63370=>"101001101",
  63371=>"100010000",
  63372=>"110111001",
  63373=>"111111110",
  63374=>"110010000",
  63375=>"100101110",
  63376=>"001000101",
  63377=>"110100000",
  63378=>"001000110",
  63379=>"110001100",
  63380=>"000101001",
  63381=>"000111001",
  63382=>"101111011",
  63383=>"110111101",
  63384=>"101010101",
  63385=>"010010000",
  63386=>"101010110",
  63387=>"101010001",
  63388=>"001011100",
  63389=>"101111101",
  63390=>"011001111",
  63391=>"010101110",
  63392=>"010110010",
  63393=>"000000111",
  63394=>"010010111",
  63395=>"011010101",
  63396=>"011001000",
  63397=>"101111011",
  63398=>"100000110",
  63399=>"101100000",
  63400=>"110111100",
  63401=>"001111100",
  63402=>"011111000",
  63403=>"001101000",
  63404=>"111110001",
  63405=>"000001110",
  63406=>"101101000",
  63407=>"100000110",
  63408=>"111110000",
  63409=>"011101001",
  63410=>"001000011",
  63411=>"110010000",
  63412=>"010111000",
  63413=>"101101100",
  63414=>"111000101",
  63415=>"110010000",
  63416=>"010000110",
  63417=>"011100010",
  63418=>"111000011",
  63419=>"111110001",
  63420=>"000110000",
  63421=>"000111000",
  63422=>"000100000",
  63423=>"011111000",
  63424=>"001111101",
  63425=>"011000110",
  63426=>"011011100",
  63427=>"001000011",
  63428=>"110010001",
  63429=>"000100111",
  63430=>"000111010",
  63431=>"001010000",
  63432=>"000000001",
  63433=>"100101010",
  63434=>"110100100",
  63435=>"001000101",
  63436=>"001011110",
  63437=>"010001100",
  63438=>"101000110",
  63439=>"101010011",
  63440=>"001110101",
  63441=>"010100001",
  63442=>"000111100",
  63443=>"101100011",
  63444=>"101011110",
  63445=>"010101100",
  63446=>"110111100",
  63447=>"000101111",
  63448=>"000000000",
  63449=>"101010111",
  63450=>"000111111",
  63451=>"111011000",
  63452=>"000100000",
  63453=>"100110100",
  63454=>"100011110",
  63455=>"101110010",
  63456=>"011110000",
  63457=>"001110101",
  63458=>"011100101",
  63459=>"000110001",
  63460=>"000100000",
  63461=>"001011011",
  63462=>"000000101",
  63463=>"101110111",
  63464=>"101101010",
  63465=>"001010011",
  63466=>"001011011",
  63467=>"000010111",
  63468=>"101011110",
  63469=>"001111011",
  63470=>"011100101",
  63471=>"001101000",
  63472=>"100000111",
  63473=>"101101010",
  63474=>"011011011",
  63475=>"111111010",
  63476=>"010000000",
  63477=>"110100000",
  63478=>"111101100",
  63479=>"100110101",
  63480=>"000101001",
  63481=>"000001001",
  63482=>"111000101",
  63483=>"100101110",
  63484=>"010001000",
  63485=>"110100100",
  63486=>"111101101",
  63487=>"110100000",
  63488=>"011110010",
  63489=>"001110001",
  63490=>"001001101",
  63491=>"011111000",
  63492=>"101011111",
  63493=>"010100000",
  63494=>"011110101",
  63495=>"110111000",
  63496=>"001001001",
  63497=>"011111111",
  63498=>"100001101",
  63499=>"111000100",
  63500=>"000010101",
  63501=>"110110011",
  63502=>"001001101",
  63503=>"011011101",
  63504=>"111111100",
  63505=>"000010010",
  63506=>"110010000",
  63507=>"110000011",
  63508=>"011110100",
  63509=>"101011000",
  63510=>"000000000",
  63511=>"110101011",
  63512=>"001110011",
  63513=>"100010101",
  63514=>"110011110",
  63515=>"001011011",
  63516=>"101000111",
  63517=>"100000001",
  63518=>"101111010",
  63519=>"100110001",
  63520=>"110000110",
  63521=>"000110001",
  63522=>"001001001",
  63523=>"111000011",
  63524=>"111011011",
  63525=>"101000101",
  63526=>"001110100",
  63527=>"100101001",
  63528=>"010001111",
  63529=>"001110111",
  63530=>"100001111",
  63531=>"100110111",
  63532=>"010110011",
  63533=>"101101111",
  63534=>"001100111",
  63535=>"011010010",
  63536=>"111100111",
  63537=>"000111111",
  63538=>"100001001",
  63539=>"111110110",
  63540=>"001100101",
  63541=>"010101000",
  63542=>"001110111",
  63543=>"111111101",
  63544=>"111111010",
  63545=>"110010110",
  63546=>"001111010",
  63547=>"110000001",
  63548=>"001000111",
  63549=>"001001001",
  63550=>"111111010",
  63551=>"001011101",
  63552=>"111111000",
  63553=>"001101010",
  63554=>"000000111",
  63555=>"001001101",
  63556=>"111010110",
  63557=>"110100111",
  63558=>"000111110",
  63559=>"011000100",
  63560=>"101011011",
  63561=>"000101001",
  63562=>"000010110",
  63563=>"001010011",
  63564=>"010111010",
  63565=>"001101001",
  63566=>"000111000",
  63567=>"001001100",
  63568=>"110001111",
  63569=>"100111100",
  63570=>"110100111",
  63571=>"000100000",
  63572=>"100000011",
  63573=>"101100101",
  63574=>"010101001",
  63575=>"000010001",
  63576=>"000101111",
  63577=>"011011111",
  63578=>"001000001",
  63579=>"010110111",
  63580=>"010000100",
  63581=>"010000000",
  63582=>"001010000",
  63583=>"100001111",
  63584=>"100010000",
  63585=>"000111000",
  63586=>"000001000",
  63587=>"001001001",
  63588=>"111110000",
  63589=>"110011111",
  63590=>"000111011",
  63591=>"001110110",
  63592=>"011100111",
  63593=>"101000110",
  63594=>"001101101",
  63595=>"101001100",
  63596=>"011111101",
  63597=>"111011001",
  63598=>"010010101",
  63599=>"001001000",
  63600=>"010111000",
  63601=>"100100110",
  63602=>"100001010",
  63603=>"101110101",
  63604=>"101000110",
  63605=>"000000111",
  63606=>"011001100",
  63607=>"001000110",
  63608=>"110111111",
  63609=>"111010001",
  63610=>"101001001",
  63611=>"001100111",
  63612=>"101110001",
  63613=>"000000000",
  63614=>"011011000",
  63615=>"100010001",
  63616=>"010000000",
  63617=>"110011011",
  63618=>"010000110",
  63619=>"000000101",
  63620=>"010001111",
  63621=>"110011011",
  63622=>"001101110",
  63623=>"111111100",
  63624=>"011101000",
  63625=>"100110110",
  63626=>"100111100",
  63627=>"000000001",
  63628=>"101000111",
  63629=>"111101000",
  63630=>"110000100",
  63631=>"101000000",
  63632=>"010011110",
  63633=>"010100110",
  63634=>"101001101",
  63635=>"010010110",
  63636=>"001100001",
  63637=>"111111111",
  63638=>"110001001",
  63639=>"100010001",
  63640=>"111001111",
  63641=>"111011001",
  63642=>"011101111",
  63643=>"011000011",
  63644=>"101011111",
  63645=>"000111100",
  63646=>"101001010",
  63647=>"111100011",
  63648=>"010001000",
  63649=>"010010001",
  63650=>"100111110",
  63651=>"000100010",
  63652=>"011010100",
  63653=>"001111011",
  63654=>"001101000",
  63655=>"010111100",
  63656=>"010111010",
  63657=>"011100011",
  63658=>"110001010",
  63659=>"111001100",
  63660=>"010111010",
  63661=>"000011110",
  63662=>"001100100",
  63663=>"011001011",
  63664=>"110111111",
  63665=>"101111011",
  63666=>"100110100",
  63667=>"111001110",
  63668=>"000001010",
  63669=>"100010010",
  63670=>"110011110",
  63671=>"111000011",
  63672=>"011011101",
  63673=>"001010101",
  63674=>"001010110",
  63675=>"001101111",
  63676=>"000000110",
  63677=>"101011011",
  63678=>"100101111",
  63679=>"111000101",
  63680=>"001110100",
  63681=>"101111001",
  63682=>"111110110",
  63683=>"101111001",
  63684=>"001001000",
  63685=>"111001101",
  63686=>"010011100",
  63687=>"100110001",
  63688=>"000111101",
  63689=>"000101100",
  63690=>"000000101",
  63691=>"110111111",
  63692=>"001001001",
  63693=>"010001100",
  63694=>"110110001",
  63695=>"100001111",
  63696=>"110011100",
  63697=>"100100001",
  63698=>"000010011",
  63699=>"000011001",
  63700=>"110000101",
  63701=>"101111111",
  63702=>"001100000",
  63703=>"100100100",
  63704=>"010110101",
  63705=>"010110011",
  63706=>"110110111",
  63707=>"101011001",
  63708=>"111101000",
  63709=>"110100111",
  63710=>"111101101",
  63711=>"110010100",
  63712=>"001001001",
  63713=>"001110001",
  63714=>"011111111",
  63715=>"111100100",
  63716=>"011111000",
  63717=>"100100101",
  63718=>"011110001",
  63719=>"100000101",
  63720=>"011000100",
  63721=>"110100010",
  63722=>"100001000",
  63723=>"100010101",
  63724=>"011011101",
  63725=>"011100110",
  63726=>"101110101",
  63727=>"001101000",
  63728=>"000100110",
  63729=>"110010110",
  63730=>"010100110",
  63731=>"001111000",
  63732=>"010110110",
  63733=>"010010010",
  63734=>"111000111",
  63735=>"110000011",
  63736=>"100001111",
  63737=>"100101101",
  63738=>"100110100",
  63739=>"010100001",
  63740=>"111101111",
  63741=>"010011100",
  63742=>"000001101",
  63743=>"000101101",
  63744=>"011111110",
  63745=>"000001111",
  63746=>"011010010",
  63747=>"000100111",
  63748=>"000000111",
  63749=>"001010011",
  63750=>"001001000",
  63751=>"011100011",
  63752=>"110010001",
  63753=>"001010110",
  63754=>"011011001",
  63755=>"001110100",
  63756=>"000111110",
  63757=>"110001000",
  63758=>"111100010",
  63759=>"000111011",
  63760=>"000100110",
  63761=>"110001110",
  63762=>"101010011",
  63763=>"011101010",
  63764=>"111000011",
  63765=>"001001011",
  63766=>"100100100",
  63767=>"110101100",
  63768=>"011110100",
  63769=>"101111100",
  63770=>"011110011",
  63771=>"111011110",
  63772=>"000110001",
  63773=>"001101100",
  63774=>"000101000",
  63775=>"101101010",
  63776=>"111111101",
  63777=>"000110010",
  63778=>"100001001",
  63779=>"100010100",
  63780=>"111001100",
  63781=>"100100011",
  63782=>"111100110",
  63783=>"011000000",
  63784=>"011011010",
  63785=>"001110111",
  63786=>"111110010",
  63787=>"100010011",
  63788=>"000010000",
  63789=>"111110010",
  63790=>"101010011",
  63791=>"001110011",
  63792=>"111101110",
  63793=>"000010010",
  63794=>"011100001",
  63795=>"111110111",
  63796=>"111001011",
  63797=>"010110011",
  63798=>"011111111",
  63799=>"111100100",
  63800=>"101110001",
  63801=>"100111111",
  63802=>"000001100",
  63803=>"110001001",
  63804=>"000011110",
  63805=>"110010010",
  63806=>"100100010",
  63807=>"110101111",
  63808=>"001110101",
  63809=>"111000100",
  63810=>"000000110",
  63811=>"111111001",
  63812=>"111111000",
  63813=>"100001011",
  63814=>"111010101",
  63815=>"110000010",
  63816=>"000011111",
  63817=>"000100001",
  63818=>"001010011",
  63819=>"101101011",
  63820=>"100001101",
  63821=>"111101111",
  63822=>"000111110",
  63823=>"001111000",
  63824=>"100100010",
  63825=>"001111101",
  63826=>"011011011",
  63827=>"110110000",
  63828=>"100100001",
  63829=>"010001111",
  63830=>"110110101",
  63831=>"110000011",
  63832=>"100000110",
  63833=>"001101011",
  63834=>"100000110",
  63835=>"111110101",
  63836=>"011110010",
  63837=>"001110001",
  63838=>"000110011",
  63839=>"100111101",
  63840=>"110011010",
  63841=>"001011000",
  63842=>"111110111",
  63843=>"011010110",
  63844=>"010100000",
  63845=>"010001110",
  63846=>"010110011",
  63847=>"111111111",
  63848=>"010011000",
  63849=>"100001101",
  63850=>"111111001",
  63851=>"110000100",
  63852=>"000100110",
  63853=>"111001001",
  63854=>"101011011",
  63855=>"100110101",
  63856=>"000111000",
  63857=>"110000001",
  63858=>"111100101",
  63859=>"011101101",
  63860=>"111100000",
  63861=>"101001011",
  63862=>"011011100",
  63863=>"100000000",
  63864=>"000101111",
  63865=>"001001010",
  63866=>"011110101",
  63867=>"111001111",
  63868=>"010001010",
  63869=>"110001110",
  63870=>"001100000",
  63871=>"000110100",
  63872=>"000011010",
  63873=>"011001110",
  63874=>"000011111",
  63875=>"101000010",
  63876=>"000011101",
  63877=>"101100001",
  63878=>"000101100",
  63879=>"001111010",
  63880=>"011001001",
  63881=>"000010010",
  63882=>"001010000",
  63883=>"001110001",
  63884=>"011110011",
  63885=>"101000101",
  63886=>"011111111",
  63887=>"100010011",
  63888=>"111101000",
  63889=>"001001111",
  63890=>"001101010",
  63891=>"011000111",
  63892=>"110100101",
  63893=>"001000010",
  63894=>"101101001",
  63895=>"101111111",
  63896=>"100110010",
  63897=>"111101110",
  63898=>"011000010",
  63899=>"101101001",
  63900=>"010100000",
  63901=>"011100000",
  63902=>"110011101",
  63903=>"101011110",
  63904=>"100100001",
  63905=>"010001000",
  63906=>"000111101",
  63907=>"110110001",
  63908=>"111011000",
  63909=>"011011111",
  63910=>"110000100",
  63911=>"111100111",
  63912=>"110001111",
  63913=>"101010101",
  63914=>"110001111",
  63915=>"100100000",
  63916=>"011100101",
  63917=>"000011011",
  63918=>"111110110",
  63919=>"101001110",
  63920=>"100110110",
  63921=>"100000010",
  63922=>"010101010",
  63923=>"101100011",
  63924=>"111000111",
  63925=>"110000011",
  63926=>"110100000",
  63927=>"110000000",
  63928=>"011101111",
  63929=>"110100101",
  63930=>"011000101",
  63931=>"110010101",
  63932=>"000000010",
  63933=>"001101110",
  63934=>"011011110",
  63935=>"111110100",
  63936=>"100001000",
  63937=>"110101101",
  63938=>"001110110",
  63939=>"111000111",
  63940=>"001101110",
  63941=>"110110010",
  63942=>"111110111",
  63943=>"111100010",
  63944=>"010001111",
  63945=>"000111011",
  63946=>"101110100",
  63947=>"110011010",
  63948=>"010110100",
  63949=>"111110011",
  63950=>"000101000",
  63951=>"000111111",
  63952=>"010001001",
  63953=>"001011010",
  63954=>"000101101",
  63955=>"110001010",
  63956=>"000010110",
  63957=>"101101000",
  63958=>"110110111",
  63959=>"000000100",
  63960=>"000010111",
  63961=>"110110001",
  63962=>"000111000",
  63963=>"101101101",
  63964=>"010001011",
  63965=>"011100110",
  63966=>"000011111",
  63967=>"101111111",
  63968=>"101111110",
  63969=>"010000101",
  63970=>"000000111",
  63971=>"111111010",
  63972=>"010111111",
  63973=>"101110110",
  63974=>"000011111",
  63975=>"010100011",
  63976=>"001100111",
  63977=>"111010100",
  63978=>"010000011",
  63979=>"000000000",
  63980=>"110111001",
  63981=>"111101000",
  63982=>"010100111",
  63983=>"110000111",
  63984=>"110011100",
  63985=>"111110110",
  63986=>"011101101",
  63987=>"110100101",
  63988=>"000110110",
  63989=>"001011001",
  63990=>"101101011",
  63991=>"100110100",
  63992=>"001100011",
  63993=>"110111100",
  63994=>"010000000",
  63995=>"011001010",
  63996=>"001000110",
  63997=>"001110111",
  63998=>"011101011",
  63999=>"011000110",
  64000=>"000111000",
  64001=>"100010010",
  64002=>"110101100",
  64003=>"111100011",
  64004=>"100011001",
  64005=>"100100100",
  64006=>"111000101",
  64007=>"011001101",
  64008=>"011111010",
  64009=>"010001100",
  64010=>"001010100",
  64011=>"000011010",
  64012=>"010001010",
  64013=>"011111010",
  64014=>"010011111",
  64015=>"011001101",
  64016=>"010100110",
  64017=>"001000110",
  64018=>"101111010",
  64019=>"101011111",
  64020=>"110111101",
  64021=>"011111001",
  64022=>"101010001",
  64023=>"101110011",
  64024=>"011001111",
  64025=>"101101011",
  64026=>"101001110",
  64027=>"110000000",
  64028=>"110011101",
  64029=>"011111101",
  64030=>"010110000",
  64031=>"010001100",
  64032=>"010011111",
  64033=>"111111110",
  64034=>"101010010",
  64035=>"001111001",
  64036=>"010100110",
  64037=>"000100010",
  64038=>"111100100",
  64039=>"010111110",
  64040=>"000111011",
  64041=>"011001001",
  64042=>"110101110",
  64043=>"110010110",
  64044=>"011001111",
  64045=>"111011001",
  64046=>"101000000",
  64047=>"111001001",
  64048=>"110011010",
  64049=>"101101110",
  64050=>"111111111",
  64051=>"011111110",
  64052=>"101001111",
  64053=>"100000111",
  64054=>"011101110",
  64055=>"010010110",
  64056=>"110111011",
  64057=>"000010010",
  64058=>"010010111",
  64059=>"011010110",
  64060=>"011000100",
  64061=>"010010100",
  64062=>"110100011",
  64063=>"100110110",
  64064=>"110111101",
  64065=>"111111101",
  64066=>"101110101",
  64067=>"111011110",
  64068=>"000110111",
  64069=>"101100000",
  64070=>"111011000",
  64071=>"111100000",
  64072=>"001111110",
  64073=>"010000001",
  64074=>"110000011",
  64075=>"001100000",
  64076=>"001001011",
  64077=>"100000001",
  64078=>"101000011",
  64079=>"000000100",
  64080=>"100010110",
  64081=>"011100111",
  64082=>"011001000",
  64083=>"000110001",
  64084=>"011000111",
  64085=>"010110100",
  64086=>"111010011",
  64087=>"000010110",
  64088=>"010111011",
  64089=>"001100000",
  64090=>"100000100",
  64091=>"101100100",
  64092=>"011000010",
  64093=>"111111001",
  64094=>"110101110",
  64095=>"111010000",
  64096=>"000100000",
  64097=>"110101000",
  64098=>"111110010",
  64099=>"011001100",
  64100=>"001011000",
  64101=>"000000010",
  64102=>"110000110",
  64103=>"001101101",
  64104=>"010010011",
  64105=>"011100000",
  64106=>"010100011",
  64107=>"011010000",
  64108=>"101001011",
  64109=>"110000010",
  64110=>"111000001",
  64111=>"110110110",
  64112=>"100110110",
  64113=>"101101100",
  64114=>"111110011",
  64115=>"001001111",
  64116=>"100111111",
  64117=>"011010000",
  64118=>"011000011",
  64119=>"000111011",
  64120=>"101110000",
  64121=>"001010001",
  64122=>"000101100",
  64123=>"000000000",
  64124=>"110111000",
  64125=>"101001001",
  64126=>"101000011",
  64127=>"110110001",
  64128=>"100100011",
  64129=>"010010100",
  64130=>"001101100",
  64131=>"011101001",
  64132=>"011000001",
  64133=>"101000000",
  64134=>"001000101",
  64135=>"100010111",
  64136=>"111101000",
  64137=>"100100101",
  64138=>"111101001",
  64139=>"010110101",
  64140=>"111100000",
  64141=>"110110010",
  64142=>"010100010",
  64143=>"001110011",
  64144=>"111111011",
  64145=>"000010100",
  64146=>"001000001",
  64147=>"010111100",
  64148=>"000000011",
  64149=>"010000001",
  64150=>"010110000",
  64151=>"100011011",
  64152=>"101110100",
  64153=>"000011010",
  64154=>"110110110",
  64155=>"011011000",
  64156=>"100011000",
  64157=>"101000010",
  64158=>"110001010",
  64159=>"010011111",
  64160=>"001001000",
  64161=>"110101000",
  64162=>"100000101",
  64163=>"001101111",
  64164=>"010101100",
  64165=>"001101101",
  64166=>"110101001",
  64167=>"000110000",
  64168=>"111000100",
  64169=>"101100011",
  64170=>"101100111",
  64171=>"000110111",
  64172=>"011100000",
  64173=>"000101110",
  64174=>"100111100",
  64175=>"010101100",
  64176=>"110011111",
  64177=>"011001110",
  64178=>"110011010",
  64179=>"000011001",
  64180=>"111110000",
  64181=>"010110111",
  64182=>"100100010",
  64183=>"111110110",
  64184=>"101100010",
  64185=>"011011110",
  64186=>"010110001",
  64187=>"110100001",
  64188=>"110010101",
  64189=>"111010001",
  64190=>"010000101",
  64191=>"010011111",
  64192=>"111110010",
  64193=>"110001100",
  64194=>"010100101",
  64195=>"101000001",
  64196=>"100100110",
  64197=>"100000001",
  64198=>"100100110",
  64199=>"110111000",
  64200=>"011110011",
  64201=>"110001101",
  64202=>"110010101",
  64203=>"111111110",
  64204=>"110111000",
  64205=>"110111110",
  64206=>"001100010",
  64207=>"111010001",
  64208=>"001001110",
  64209=>"110111011",
  64210=>"000110011",
  64211=>"100000011",
  64212=>"100000001",
  64213=>"111001011",
  64214=>"010101110",
  64215=>"001101100",
  64216=>"001010010",
  64217=>"000100001",
  64218=>"001011101",
  64219=>"100110100",
  64220=>"111000000",
  64221=>"000010010",
  64222=>"000011011",
  64223=>"100101111",
  64224=>"100100010",
  64225=>"101111011",
  64226=>"001110111",
  64227=>"100010111",
  64228=>"000001100",
  64229=>"110110010",
  64230=>"111010010",
  64231=>"110111111",
  64232=>"100111000",
  64233=>"100011011",
  64234=>"000101111",
  64235=>"000001001",
  64236=>"101110110",
  64237=>"110001011",
  64238=>"010111111",
  64239=>"111010100",
  64240=>"000010100",
  64241=>"010111100",
  64242=>"111010111",
  64243=>"010011001",
  64244=>"011001011",
  64245=>"010010100",
  64246=>"100101001",
  64247=>"100000110",
  64248=>"101000110",
  64249=>"000101101",
  64250=>"111101010",
  64251=>"000000010",
  64252=>"001110000",
  64253=>"101000010",
  64254=>"010000101",
  64255=>"100111110",
  64256=>"011101011",
  64257=>"101001011",
  64258=>"101010011",
  64259=>"011010101",
  64260=>"111111011",
  64261=>"100110110",
  64262=>"111100000",
  64263=>"000111001",
  64264=>"111011100",
  64265=>"111011111",
  64266=>"010000000",
  64267=>"001100010",
  64268=>"100010101",
  64269=>"110101100",
  64270=>"010011011",
  64271=>"111110100",
  64272=>"100110100",
  64273=>"101101110",
  64274=>"111001111",
  64275=>"110000000",
  64276=>"110111101",
  64277=>"010000000",
  64278=>"110111010",
  64279=>"101111010",
  64280=>"101100001",
  64281=>"010101110",
  64282=>"100010101",
  64283=>"000011001",
  64284=>"110011001",
  64285=>"000100101",
  64286=>"110010101",
  64287=>"000001010",
  64288=>"101110000",
  64289=>"110111101",
  64290=>"111110110",
  64291=>"110110101",
  64292=>"100110101",
  64293=>"111001100",
  64294=>"000010111",
  64295=>"100101110",
  64296=>"110100111",
  64297=>"011110001",
  64298=>"010011100",
  64299=>"111001110",
  64300=>"111101100",
  64301=>"100010111",
  64302=>"100100100",
  64303=>"100100110",
  64304=>"000000111",
  64305=>"011110100",
  64306=>"000011111",
  64307=>"101011000",
  64308=>"111110111",
  64309=>"110011101",
  64310=>"010011100",
  64311=>"111100100",
  64312=>"010001100",
  64313=>"000110010",
  64314=>"011101100",
  64315=>"000101100",
  64316=>"011000100",
  64317=>"001010101",
  64318=>"100100010",
  64319=>"011011101",
  64320=>"011010001",
  64321=>"000000000",
  64322=>"000001010",
  64323=>"100110100",
  64324=>"100101111",
  64325=>"010000111",
  64326=>"010111101",
  64327=>"111101100",
  64328=>"001001011",
  64329=>"101110101",
  64330=>"011111111",
  64331=>"000010011",
  64332=>"110110011",
  64333=>"001011111",
  64334=>"000001110",
  64335=>"101001110",
  64336=>"111100100",
  64337=>"101010001",
  64338=>"110001001",
  64339=>"010010001",
  64340=>"101100111",
  64341=>"111011110",
  64342=>"100001111",
  64343=>"010111001",
  64344=>"110101011",
  64345=>"111101101",
  64346=>"110011010",
  64347=>"100011000",
  64348=>"000011101",
  64349=>"010010110",
  64350=>"001011101",
  64351=>"111000001",
  64352=>"111101100",
  64353=>"110000110",
  64354=>"110000000",
  64355=>"000000011",
  64356=>"010010010",
  64357=>"100111000",
  64358=>"001010111",
  64359=>"001010000",
  64360=>"001000000",
  64361=>"101011110",
  64362=>"010101100",
  64363=>"010000001",
  64364=>"011100000",
  64365=>"101000000",
  64366=>"100100110",
  64367=>"001010001",
  64368=>"000111011",
  64369=>"001111110",
  64370=>"101010011",
  64371=>"011111011",
  64372=>"101001001",
  64373=>"111100101",
  64374=>"111010110",
  64375=>"111110101",
  64376=>"001110111",
  64377=>"100011001",
  64378=>"000010011",
  64379=>"111001011",
  64380=>"001001011",
  64381=>"011101011",
  64382=>"010000110",
  64383=>"110011010",
  64384=>"000100110",
  64385=>"101011111",
  64386=>"110000111",
  64387=>"110110111",
  64388=>"000011000",
  64389=>"011101010",
  64390=>"001111011",
  64391=>"111011101",
  64392=>"011100011",
  64393=>"111100100",
  64394=>"101001100",
  64395=>"101000010",
  64396=>"100111010",
  64397=>"110100010",
  64398=>"001101011",
  64399=>"101111011",
  64400=>"010000011",
  64401=>"100111101",
  64402=>"000011111",
  64403=>"100001100",
  64404=>"000111110",
  64405=>"100111011",
  64406=>"111011011",
  64407=>"111100110",
  64408=>"111100011",
  64409=>"010110001",
  64410=>"011101101",
  64411=>"111100101",
  64412=>"110011110",
  64413=>"101100001",
  64414=>"011011110",
  64415=>"111111110",
  64416=>"001100010",
  64417=>"000110110",
  64418=>"010001110",
  64419=>"011100010",
  64420=>"110100000",
  64421=>"010100011",
  64422=>"100011100",
  64423=>"101011000",
  64424=>"010100000",
  64425=>"101100000",
  64426=>"000001010",
  64427=>"111100011",
  64428=>"001101100",
  64429=>"010011010",
  64430=>"000010011",
  64431=>"101111010",
  64432=>"001000111",
  64433=>"111111001",
  64434=>"101100011",
  64435=>"010111001",
  64436=>"110110000",
  64437=>"010001010",
  64438=>"001101000",
  64439=>"010000111",
  64440=>"100111011",
  64441=>"011010001",
  64442=>"110001000",
  64443=>"111110101",
  64444=>"001000110",
  64445=>"011010011",
  64446=>"000011001",
  64447=>"000010110",
  64448=>"011011010",
  64449=>"101001001",
  64450=>"101011000",
  64451=>"110100011",
  64452=>"001001010",
  64453=>"100111010",
  64454=>"110000101",
  64455=>"101110110",
  64456=>"111100001",
  64457=>"101001111",
  64458=>"010011110",
  64459=>"101001000",
  64460=>"000001100",
  64461=>"000011010",
  64462=>"110110111",
  64463=>"111011001",
  64464=>"010111101",
  64465=>"100011010",
  64466=>"001110000",
  64467=>"000010100",
  64468=>"100010010",
  64469=>"110100000",
  64470=>"100111011",
  64471=>"010000000",
  64472=>"111001011",
  64473=>"101100101",
  64474=>"101100111",
  64475=>"000100011",
  64476=>"110111000",
  64477=>"001001110",
  64478=>"000100011",
  64479=>"001111100",
  64480=>"011111011",
  64481=>"010001010",
  64482=>"100101110",
  64483=>"000111001",
  64484=>"000010010",
  64485=>"000110111",
  64486=>"010001000",
  64487=>"010111011",
  64488=>"001001101",
  64489=>"001100101",
  64490=>"011010110",
  64491=>"011010101",
  64492=>"100000000",
  64493=>"100000110",
  64494=>"111100110",
  64495=>"001011001",
  64496=>"000111111",
  64497=>"010010100",
  64498=>"011010111",
  64499=>"000001110",
  64500=>"010101100",
  64501=>"001001000",
  64502=>"110000001",
  64503=>"110010010",
  64504=>"001001101",
  64505=>"000010000",
  64506=>"010100100",
  64507=>"111010011",
  64508=>"001000001",
  64509=>"110111010",
  64510=>"100100010",
  64511=>"001001100",
  64512=>"100101101",
  64513=>"101100011",
  64514=>"110001101",
  64515=>"000111010",
  64516=>"010001101",
  64517=>"000100001",
  64518=>"100110110",
  64519=>"101100001",
  64520=>"101100110",
  64521=>"011111101",
  64522=>"110111100",
  64523=>"011111100",
  64524=>"110011111",
  64525=>"111101000",
  64526=>"100001101",
  64527=>"010110010",
  64528=>"010001100",
  64529=>"100000001",
  64530=>"011100111",
  64531=>"001110101",
  64532=>"101110110",
  64533=>"100000011",
  64534=>"110111010",
  64535=>"101111100",
  64536=>"100010111",
  64537=>"100010101",
  64538=>"111101010",
  64539=>"101011010",
  64540=>"100000110",
  64541=>"111110010",
  64542=>"011111010",
  64543=>"100010000",
  64544=>"111011101",
  64545=>"110110010",
  64546=>"100010010",
  64547=>"110010111",
  64548=>"000001011",
  64549=>"101110001",
  64550=>"001011100",
  64551=>"110101011",
  64552=>"001111111",
  64553=>"010101010",
  64554=>"101001000",
  64555=>"111101111",
  64556=>"001011011",
  64557=>"101011100",
  64558=>"000001000",
  64559=>"100101111",
  64560=>"110110110",
  64561=>"000101011",
  64562=>"111110000",
  64563=>"111011000",
  64564=>"010111010",
  64565=>"010010011",
  64566=>"100001110",
  64567=>"001000101",
  64568=>"100010110",
  64569=>"011011100",
  64570=>"111011101",
  64571=>"001110000",
  64572=>"111001110",
  64573=>"110110110",
  64574=>"100010011",
  64575=>"000110000",
  64576=>"000010101",
  64577=>"001011001",
  64578=>"100010000",
  64579=>"100010101",
  64580=>"100100100",
  64581=>"111000001",
  64582=>"100110111",
  64583=>"000110001",
  64584=>"101001101",
  64585=>"100110100",
  64586=>"001001001",
  64587=>"001110010",
  64588=>"111111110",
  64589=>"011011110",
  64590=>"110000000",
  64591=>"101110001",
  64592=>"100000111",
  64593=>"110000001",
  64594=>"000010100",
  64595=>"111111000",
  64596=>"010011101",
  64597=>"011111101",
  64598=>"100100011",
  64599=>"001001001",
  64600=>"001111010",
  64601=>"010011001",
  64602=>"001001010",
  64603=>"001000111",
  64604=>"000011110",
  64605=>"000101010",
  64606=>"100001101",
  64607=>"101010111",
  64608=>"000100111",
  64609=>"101110101",
  64610=>"111010001",
  64611=>"000101011",
  64612=>"111111101",
  64613=>"101011010",
  64614=>"111100001",
  64615=>"101101100",
  64616=>"010000010",
  64617=>"001001000",
  64618=>"111001001",
  64619=>"011000110",
  64620=>"001101110",
  64621=>"010101100",
  64622=>"010110001",
  64623=>"100111101",
  64624=>"110110000",
  64625=>"010011011",
  64626=>"100000101",
  64627=>"011100000",
  64628=>"001001111",
  64629=>"101001101",
  64630=>"001111100",
  64631=>"001111100",
  64632=>"111100010",
  64633=>"001111110",
  64634=>"000111001",
  64635=>"101000011",
  64636=>"010111110",
  64637=>"001100010",
  64638=>"001100100",
  64639=>"010100100",
  64640=>"111000001",
  64641=>"001111110",
  64642=>"010010100",
  64643=>"100010001",
  64644=>"101010000",
  64645=>"000010111",
  64646=>"010010110",
  64647=>"110000010",
  64648=>"101110010",
  64649=>"010010001",
  64650=>"011110001",
  64651=>"111010101",
  64652=>"000000100",
  64653=>"110100000",
  64654=>"111111011",
  64655=>"010110000",
  64656=>"101000101",
  64657=>"110000011",
  64658=>"111101101",
  64659=>"011000110",
  64660=>"001001001",
  64661=>"101001111",
  64662=>"011100111",
  64663=>"100010110",
  64664=>"111100111",
  64665=>"100111110",
  64666=>"011100010",
  64667=>"100011001",
  64668=>"100010110",
  64669=>"101100101",
  64670=>"010001111",
  64671=>"100001011",
  64672=>"000101110",
  64673=>"011110101",
  64674=>"000000110",
  64675=>"011000000",
  64676=>"100101001",
  64677=>"110000001",
  64678=>"000011010",
  64679=>"001111110",
  64680=>"100110010",
  64681=>"111010001",
  64682=>"011111010",
  64683=>"010000000",
  64684=>"101010111",
  64685=>"111110101",
  64686=>"011010101",
  64687=>"010110010",
  64688=>"000000100",
  64689=>"100110000",
  64690=>"110100101",
  64691=>"010001000",
  64692=>"101001010",
  64693=>"011000100",
  64694=>"001001110",
  64695=>"010110010",
  64696=>"110001110",
  64697=>"011111111",
  64698=>"000000000",
  64699=>"110000010",
  64700=>"111011101",
  64701=>"110001101",
  64702=>"010011010",
  64703=>"111101101",
  64704=>"000111000",
  64705=>"001100010",
  64706=>"111111001",
  64707=>"000100100",
  64708=>"101111011",
  64709=>"011100111",
  64710=>"001000000",
  64711=>"000000001",
  64712=>"100110000",
  64713=>"010001000",
  64714=>"011111000",
  64715=>"000101010",
  64716=>"001101101",
  64717=>"110101000",
  64718=>"100001001",
  64719=>"011100111",
  64720=>"000001010",
  64721=>"001101000",
  64722=>"110100000",
  64723=>"100011110",
  64724=>"001110100",
  64725=>"000000000",
  64726=>"011110101",
  64727=>"111100100",
  64728=>"101010001",
  64729=>"000111100",
  64730=>"000100100",
  64731=>"101000000",
  64732=>"110000001",
  64733=>"101001000",
  64734=>"100010001",
  64735=>"110100111",
  64736=>"111110111",
  64737=>"100100010",
  64738=>"000101000",
  64739=>"010101111",
  64740=>"010010111",
  64741=>"111110010",
  64742=>"001111100",
  64743=>"000000001",
  64744=>"011111111",
  64745=>"100000011",
  64746=>"000000101",
  64747=>"100110111",
  64748=>"000100001",
  64749=>"110111110",
  64750=>"100101100",
  64751=>"100101111",
  64752=>"000011101",
  64753=>"010011100",
  64754=>"001011101",
  64755=>"001011111",
  64756=>"011011110",
  64757=>"001011011",
  64758=>"100111110",
  64759=>"100000111",
  64760=>"000001011",
  64761=>"110110001",
  64762=>"111000101",
  64763=>"001101000",
  64764=>"100000001",
  64765=>"101111110",
  64766=>"111011000",
  64767=>"110001101",
  64768=>"111000001",
  64769=>"010001100",
  64770=>"111001111",
  64771=>"011100101",
  64772=>"110010110",
  64773=>"111100111",
  64774=>"001011011",
  64775=>"000101011",
  64776=>"111111111",
  64777=>"011000001",
  64778=>"110011011",
  64779=>"001110011",
  64780=>"011011111",
  64781=>"100011111",
  64782=>"000001101",
  64783=>"111110100",
  64784=>"010010101",
  64785=>"010100110",
  64786=>"000001101",
  64787=>"111111110",
  64788=>"000100010",
  64789=>"111110010",
  64790=>"001111110",
  64791=>"000010101",
  64792=>"111001000",
  64793=>"001101001",
  64794=>"111100010",
  64795=>"001100011",
  64796=>"000010001",
  64797=>"111111100",
  64798=>"010001001",
  64799=>"000101111",
  64800=>"011110011",
  64801=>"100010001",
  64802=>"100101110",
  64803=>"110010111",
  64804=>"011010101",
  64805=>"111111110",
  64806=>"011110010",
  64807=>"000010110",
  64808=>"100001010",
  64809=>"011010000",
  64810=>"110111011",
  64811=>"111110000",
  64812=>"100011111",
  64813=>"010101111",
  64814=>"101010010",
  64815=>"110111100",
  64816=>"111000011",
  64817=>"011110001",
  64818=>"111001101",
  64819=>"001010011",
  64820=>"000001000",
  64821=>"011010111",
  64822=>"000110111",
  64823=>"111101010",
  64824=>"111100100",
  64825=>"000010011",
  64826=>"011011101",
  64827=>"001101001",
  64828=>"010111101",
  64829=>"011011111",
  64830=>"001000010",
  64831=>"100110100",
  64832=>"000001000",
  64833=>"100110101",
  64834=>"101001111",
  64835=>"111100100",
  64836=>"001101101",
  64837=>"011110010",
  64838=>"100000000",
  64839=>"001010001",
  64840=>"001101000",
  64841=>"110111010",
  64842=>"000111100",
  64843=>"000001000",
  64844=>"011101000",
  64845=>"111011110",
  64846=>"000101010",
  64847=>"100101000",
  64848=>"011111001",
  64849=>"001011101",
  64850=>"100100100",
  64851=>"111100110",
  64852=>"101001101",
  64853=>"100011100",
  64854=>"001110010",
  64855=>"000010100",
  64856=>"011010001",
  64857=>"001001000",
  64858=>"010011000",
  64859=>"000100000",
  64860=>"010010000",
  64861=>"001110010",
  64862=>"100011100",
  64863=>"010000000",
  64864=>"100001101",
  64865=>"101111000",
  64866=>"010011110",
  64867=>"000001100",
  64868=>"110111011",
  64869=>"001000101",
  64870=>"000001010",
  64871=>"110000111",
  64872=>"000000110",
  64873=>"001111000",
  64874=>"110111111",
  64875=>"011010110",
  64876=>"110111111",
  64877=>"000111100",
  64878=>"000011001",
  64879=>"010100100",
  64880=>"011000001",
  64881=>"000110011",
  64882=>"110101110",
  64883=>"000010101",
  64884=>"111101111",
  64885=>"110110000",
  64886=>"011100001",
  64887=>"101100111",
  64888=>"001011000",
  64889=>"000000000",
  64890=>"111010010",
  64891=>"100111010",
  64892=>"101010101",
  64893=>"010101110",
  64894=>"001100111",
  64895=>"011011000",
  64896=>"100001000",
  64897=>"001100110",
  64898=>"101001011",
  64899=>"011001110",
  64900=>"101100110",
  64901=>"110100010",
  64902=>"010111110",
  64903=>"110100100",
  64904=>"111010010",
  64905=>"000101000",
  64906=>"111010010",
  64907=>"010110011",
  64908=>"011101001",
  64909=>"100100100",
  64910=>"110000010",
  64911=>"101101000",
  64912=>"100101111",
  64913=>"000001100",
  64914=>"110010001",
  64915=>"101100010",
  64916=>"101100110",
  64917=>"101101100",
  64918=>"000101100",
  64919=>"101000010",
  64920=>"010100001",
  64921=>"000011101",
  64922=>"011110110",
  64923=>"111000011",
  64924=>"111011010",
  64925=>"111100010",
  64926=>"101101101",
  64927=>"111100011",
  64928=>"001010111",
  64929=>"110000000",
  64930=>"010100100",
  64931=>"011111001",
  64932=>"000110101",
  64933=>"001101000",
  64934=>"000000000",
  64935=>"011110011",
  64936=>"011010001",
  64937=>"111111001",
  64938=>"111111111",
  64939=>"000111001",
  64940=>"100111000",
  64941=>"011000001",
  64942=>"100111111",
  64943=>"001001000",
  64944=>"010111100",
  64945=>"101101111",
  64946=>"010000100",
  64947=>"011010010",
  64948=>"100011100",
  64949=>"011001001",
  64950=>"111011011",
  64951=>"110110010",
  64952=>"110011100",
  64953=>"000100111",
  64954=>"000011000",
  64955=>"110010010",
  64956=>"011000101",
  64957=>"101111000",
  64958=>"010111111",
  64959=>"001101110",
  64960=>"100000000",
  64961=>"110010001",
  64962=>"010000101",
  64963=>"110110100",
  64964=>"100101100",
  64965=>"101101001",
  64966=>"011101010",
  64967=>"110101011",
  64968=>"111111001",
  64969=>"010011010",
  64970=>"111101101",
  64971=>"000000011",
  64972=>"001100010",
  64973=>"010000001",
  64974=>"101110011",
  64975=>"100111010",
  64976=>"101111111",
  64977=>"111010010",
  64978=>"000010100",
  64979=>"100110110",
  64980=>"010111101",
  64981=>"000000100",
  64982=>"110001001",
  64983=>"011100100",
  64984=>"101101010",
  64985=>"100101000",
  64986=>"010010111",
  64987=>"011001000",
  64988=>"011000010",
  64989=>"001000100",
  64990=>"000111111",
  64991=>"010011000",
  64992=>"101010100",
  64993=>"011000010",
  64994=>"101000110",
  64995=>"010001000",
  64996=>"000100110",
  64997=>"110100000",
  64998=>"011101000",
  64999=>"111110000",
  65000=>"101111110",
  65001=>"010000000",
  65002=>"100100001",
  65003=>"111011110",
  65004=>"011110111",
  65005=>"001011111",
  65006=>"110100101",
  65007=>"111000001",
  65008=>"111001011",
  65009=>"000101001",
  65010=>"000001111",
  65011=>"000101110",
  65012=>"101010001",
  65013=>"010011001",
  65014=>"100000110",
  65015=>"100101100",
  65016=>"111000000",
  65017=>"100000100",
  65018=>"110001000",
  65019=>"001011111",
  65020=>"100111100",
  65021=>"000000111",
  65022=>"100101100",
  65023=>"111001101",
  65024=>"110000111",
  65025=>"100100001",
  65026=>"100001000",
  65027=>"001010001",
  65028=>"110111011",
  65029=>"111100111",
  65030=>"111111011",
  65031=>"100001011",
  65032=>"111111101",
  65033=>"101110111",
  65034=>"111010011",
  65035=>"010100010",
  65036=>"000000011",
  65037=>"000000000",
  65038=>"110110011",
  65039=>"101110000",
  65040=>"001001100",
  65041=>"111111010",
  65042=>"110010001",
  65043=>"001011000",
  65044=>"001011001",
  65045=>"100010001",
  65046=>"010010000",
  65047=>"011011100",
  65048=>"110001111",
  65049=>"010001111",
  65050=>"001000110",
  65051=>"111110001",
  65052=>"001100011",
  65053=>"101001011",
  65054=>"011100001",
  65055=>"111011110",
  65056=>"011011010",
  65057=>"011101011",
  65058=>"101000000",
  65059=>"111010111",
  65060=>"111100100",
  65061=>"010101111",
  65062=>"010011111",
  65063=>"011101000",
  65064=>"111001100",
  65065=>"011000111",
  65066=>"011011110",
  65067=>"100010010",
  65068=>"100110110",
  65069=>"111111000",
  65070=>"000011101",
  65071=>"100000001",
  65072=>"011010010",
  65073=>"101101000",
  65074=>"011111010",
  65075=>"101110010",
  65076=>"101011100",
  65077=>"011111010",
  65078=>"000000101",
  65079=>"011111011",
  65080=>"111000110",
  65081=>"001111000",
  65082=>"100101111",
  65083=>"111011111",
  65084=>"011000110",
  65085=>"000101010",
  65086=>"111111110",
  65087=>"010010000",
  65088=>"011110101",
  65089=>"101101110",
  65090=>"110101001",
  65091=>"011111110",
  65092=>"011000101",
  65093=>"101010010",
  65094=>"010010010",
  65095=>"000111011",
  65096=>"110010111",
  65097=>"100100000",
  65098=>"111010001",
  65099=>"111101100",
  65100=>"011101000",
  65101=>"110101111",
  65102=>"110111111",
  65103=>"110011110",
  65104=>"101010011",
  65105=>"000110110",
  65106=>"101111100",
  65107=>"111011101",
  65108=>"110010110",
  65109=>"100101111",
  65110=>"011001011",
  65111=>"001100110",
  65112=>"001000101",
  65113=>"011101110",
  65114=>"011101001",
  65115=>"000101111",
  65116=>"001101101",
  65117=>"010100011",
  65118=>"001110010",
  65119=>"101100101",
  65120=>"000110010",
  65121=>"010010111",
  65122=>"100000011",
  65123=>"000000001",
  65124=>"000100110",
  65125=>"101101100",
  65126=>"011101100",
  65127=>"110010111",
  65128=>"000011000",
  65129=>"001001110",
  65130=>"111110010",
  65131=>"111010110",
  65132=>"101100100",
  65133=>"100101101",
  65134=>"100101101",
  65135=>"001001101",
  65136=>"111011110",
  65137=>"010000001",
  65138=>"000100001",
  65139=>"001101010",
  65140=>"001001100",
  65141=>"001000000",
  65142=>"010110110",
  65143=>"000111011",
  65144=>"110100100",
  65145=>"111011011",
  65146=>"000010111",
  65147=>"111100100",
  65148=>"000010101",
  65149=>"000010001",
  65150=>"001011110",
  65151=>"001101011",
  65152=>"010000110",
  65153=>"011011111",
  65154=>"000110100",
  65155=>"010010001",
  65156=>"001100010",
  65157=>"101000000",
  65158=>"010111101",
  65159=>"010000001",
  65160=>"010001011",
  65161=>"111011000",
  65162=>"010100000",
  65163=>"111000111",
  65164=>"010101010",
  65165=>"010010100",
  65166=>"001111001",
  65167=>"110111010",
  65168=>"101011111",
  65169=>"110001010",
  65170=>"100101110",
  65171=>"111111110",
  65172=>"001000010",
  65173=>"000010010",
  65174=>"000101110",
  65175=>"110000001",
  65176=>"111011001",
  65177=>"010101111",
  65178=>"000100000",
  65179=>"100101101",
  65180=>"011110001",
  65181=>"100011111",
  65182=>"110011011",
  65183=>"001100100",
  65184=>"101011101",
  65185=>"000000001",
  65186=>"111101101",
  65187=>"111011101",
  65188=>"010100010",
  65189=>"111010101",
  65190=>"011011011",
  65191=>"010110010",
  65192=>"001101001",
  65193=>"100001001",
  65194=>"111010010",
  65195=>"110100100",
  65196=>"010100101",
  65197=>"110110010",
  65198=>"111101111",
  65199=>"000010011",
  65200=>"111110001",
  65201=>"111101101",
  65202=>"001000000",
  65203=>"011111010",
  65204=>"010100001",
  65205=>"011000011",
  65206=>"001001111",
  65207=>"001010111",
  65208=>"010101110",
  65209=>"011101110",
  65210=>"100110011",
  65211=>"010010001",
  65212=>"000000000",
  65213=>"010011110",
  65214=>"100111101",
  65215=>"000111011",
  65216=>"001100111",
  65217=>"000110100",
  65218=>"000011010",
  65219=>"111000110",
  65220=>"011001011",
  65221=>"111101010",
  65222=>"110111110",
  65223=>"100011010",
  65224=>"011111011",
  65225=>"101000010",
  65226=>"011000001",
  65227=>"000000001",
  65228=>"100101001",
  65229=>"100101111",
  65230=>"100101100",
  65231=>"010011000",
  65232=>"110110100",
  65233=>"010010000",
  65234=>"101111010",
  65235=>"001011001",
  65236=>"010110000",
  65237=>"000001001",
  65238=>"100001110",
  65239=>"101110010",
  65240=>"110010001",
  65241=>"011010011",
  65242=>"001000100",
  65243=>"101001011",
  65244=>"101011010",
  65245=>"000011010",
  65246=>"110100101",
  65247=>"010101110",
  65248=>"110001000",
  65249=>"010001100",
  65250=>"101010111",
  65251=>"011001110",
  65252=>"000111110",
  65253=>"001001000",
  65254=>"000100110",
  65255=>"111101101",
  65256=>"110101000",
  65257=>"101010011",
  65258=>"000000110",
  65259=>"111101101",
  65260=>"000000001",
  65261=>"001100010",
  65262=>"100101110",
  65263=>"110001000",
  65264=>"110111011",
  65265=>"000111110",
  65266=>"101101010",
  65267=>"001010100",
  65268=>"111000011",
  65269=>"111011101",
  65270=>"111111000",
  65271=>"011000100",
  65272=>"110101001",
  65273=>"001110000",
  65274=>"001010011",
  65275=>"001000110",
  65276=>"101100101",
  65277=>"110010110",
  65278=>"101000010",
  65279=>"011100000",
  65280=>"100010011",
  65281=>"100000000",
  65282=>"000111101",
  65283=>"000110000",
  65284=>"000101100",
  65285=>"010111110",
  65286=>"011001000",
  65287=>"110111110",
  65288=>"001010000",
  65289=>"011111000",
  65290=>"000011011",
  65291=>"101000101",
  65292=>"010010100",
  65293=>"110111101",
  65294=>"100101010",
  65295=>"000011011",
  65296=>"110111011",
  65297=>"100101000",
  65298=>"001010001",
  65299=>"001101011",
  65300=>"010110001",
  65301=>"111110000",
  65302=>"110101001",
  65303=>"100000001",
  65304=>"010010110",
  65305=>"010011100",
  65306=>"011110011",
  65307=>"010011110",
  65308=>"010000110",
  65309=>"011101010",
  65310=>"111000010",
  65311=>"001001111",
  65312=>"100010100",
  65313=>"011110010",
  65314=>"110111111",
  65315=>"111100001",
  65316=>"010100011",
  65317=>"101000001",
  65318=>"111111000",
  65319=>"000010100",
  65320=>"110001001",
  65321=>"011001110",
  65322=>"100101010",
  65323=>"111101000",
  65324=>"001010010",
  65325=>"100000111",
  65326=>"110001001",
  65327=>"100111001",
  65328=>"101000010",
  65329=>"110010000",
  65330=>"001011000",
  65331=>"101011110",
  65332=>"001001111",
  65333=>"001101001",
  65334=>"100011101",
  65335=>"111101001",
  65336=>"010000111",
  65337=>"101011100",
  65338=>"010010110",
  65339=>"001001111",
  65340=>"000111100",
  65341=>"010000101",
  65342=>"000101000",
  65343=>"001101001",
  65344=>"100101000",
  65345=>"111001000",
  65346=>"011011001",
  65347=>"111100101",
  65348=>"111011100",
  65349=>"110011101",
  65350=>"000100110",
  65351=>"010101000",
  65352=>"001000100",
  65353=>"110011011",
  65354=>"111001000",
  65355=>"000111001",
  65356=>"111101011",
  65357=>"101100101",
  65358=>"000000100",
  65359=>"000010111",
  65360=>"000100101",
  65361=>"100100010",
  65362=>"110001011",
  65363=>"100000101",
  65364=>"011010100",
  65365=>"010000000",
  65366=>"110000111",
  65367=>"100000001",
  65368=>"110101000",
  65369=>"001101110",
  65370=>"011000010",
  65371=>"011001011",
  65372=>"100001110",
  65373=>"111111011",
  65374=>"111100111",
  65375=>"100101010",
  65376=>"111100111",
  65377=>"001010111",
  65378=>"010111000",
  65379=>"011001101",
  65380=>"011001101",
  65381=>"001101100",
  65382=>"100111000",
  65383=>"100000010",
  65384=>"101111000",
  65385=>"100111001",
  65386=>"010011100",
  65387=>"101100111",
  65388=>"101100110",
  65389=>"101110111",
  65390=>"011100100",
  65391=>"010001011",
  65392=>"011001110",
  65393=>"111101110",
  65394=>"100111111",
  65395=>"111000100",
  65396=>"101100001",
  65397=>"010111100",
  65398=>"011001101",
  65399=>"110001010",
  65400=>"100000011",
  65401=>"111101101",
  65402=>"011011100",
  65403=>"000110011",
  65404=>"010011010",
  65405=>"100010001",
  65406=>"001000011",
  65407=>"111010100",
  65408=>"101110101",
  65409=>"110110111",
  65410=>"100111101",
  65411=>"011011100",
  65412=>"001011010",
  65413=>"001011000",
  65414=>"000001111",
  65415=>"110011010",
  65416=>"111001111",
  65417=>"010000101",
  65418=>"101111110",
  65419=>"010010000",
  65420=>"001011100",
  65421=>"101111110",
  65422=>"001101101",
  65423=>"100000011",
  65424=>"001101101",
  65425=>"010101110",
  65426=>"100011100",
  65427=>"101001010",
  65428=>"010101011",
  65429=>"011011100",
  65430=>"011001000",
  65431=>"000011001",
  65432=>"010010101",
  65433=>"010101010",
  65434=>"111100111",
  65435=>"010001111",
  65436=>"101111011",
  65437=>"001011101",
  65438=>"100010111",
  65439=>"111011010",
  65440=>"110111010",
  65441=>"111101010",
  65442=>"111111000",
  65443=>"001101011",
  65444=>"101100001",
  65445=>"101111111",
  65446=>"010000000",
  65447=>"000110011",
  65448=>"011001000",
  65449=>"011010101",
  65450=>"010111110",
  65451=>"011100100",
  65452=>"010100011",
  65453=>"110011000",
  65454=>"111011101",
  65455=>"101001110",
  65456=>"100101000",
  65457=>"100000001",
  65458=>"010010011",
  65459=>"011011010",
  65460=>"011111111",
  65461=>"011111010",
  65462=>"110110001",
  65463=>"010010101",
  65464=>"001011011",
  65465=>"111001110",
  65466=>"111010010",
  65467=>"110101001",
  65468=>"010011000",
  65469=>"101001101",
  65470=>"010010000",
  65471=>"011001010",
  65472=>"101111110",
  65473=>"010110010",
  65474=>"100000011",
  65475=>"111001100",
  65476=>"000101100",
  65477=>"010010011",
  65478=>"110010110",
  65479=>"000110000",
  65480=>"001101110",
  65481=>"001001111",
  65482=>"111100100",
  65483=>"101011010",
  65484=>"010100001",
  65485=>"101100111",
  65486=>"011010100",
  65487=>"100001001",
  65488=>"100101001",
  65489=>"101000001",
  65490=>"100100101",
  65491=>"111110110",
  65492=>"000011111",
  65493=>"010011011",
  65494=>"100001011",
  65495=>"110010110",
  65496=>"001011000",
  65497=>"001100000",
  65498=>"110101000",
  65499=>"001000000",
  65500=>"000001001",
  65501=>"000101110",
  65502=>"111001110",
  65503=>"101000000",
  65504=>"010111111",
  65505=>"000100000",
  65506=>"000011000",
  65507=>"011111001",
  65508=>"110001101",
  65509=>"010100010",
  65510=>"101001110",
  65511=>"000110101",
  65512=>"101101110",
  65513=>"110111001",
  65514=>"001100101",
  65515=>"000000100",
  65516=>"000110111",
  65517=>"100011011",
  65518=>"010000001",
  65519=>"110101011",
  65520=>"010100111",
  65521=>"011100101",
  65522=>"011111001",
  65523=>"111110011",
  65524=>"000000100",
  65525=>"001101111",
  65526=>"110111000",
  65527=>"000110001",
  65528=>"000100101",
  65529=>"101010001",
  65530=>"000111011",
  65531=>"011001010",
  65532=>"111101101",
  65533=>"011000011",
  65534=>"000010010",
  65535=>"000111000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;