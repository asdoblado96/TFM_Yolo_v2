LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L9_1_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L9_1_BNROM;

ARCHITECTURE RTL OF L9_1_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 62) OF STD_LOGIC_VECTOR(15 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0 => "0000000000000111",
  1 => "0000000000101001",
  2 => "1111111111001101",
  3 => "0000011010000111",
  4 => "1111001111010101",
  5 => "1111111101101101",
  6 => "1111111111111001",
  7 => "0000000011100000",
  8 => "0000000000001010",
  9 => "0000000010011110",
  10 => "1111111010111101",
  11 => "0000000100111100",
  12 => "1111111110100110",
  13 => "0000000101010101",
  14 => "1111111110011111",
  15 => "1111111110010000",
  16 => "1111111111010110",
  17 => "1111111101110010",
  18 => "1111111101001011",
  19 => "0000001001100010",
  20 => "0000000001110001",
  21 => "1111111110101110",
  22 => "1111111101001011",
  23 => "1111111011001100",
  24 => "1111111111000101",
  25 => "1111111101110011",
  26 => "1111111111001010",
  27 => "1111100000101101",
  28 => "1111111100101000",
  29 => "1110110111011100",
  30 => "1111111110000011",
  31 => "1111111110101101",
  32 => "0000000000111110",
  33 => "1111111111100100",
  34 => "1111111111011110",
  35 => "1111111101111011",
  36 => "0000000001010000",
  37 => "1111111110101110",
  38 => "0000000101101011",
  39 => "1111111100010010",
  40 => "1111111110111110",
  41 => "0000000000100111",
  42 => "1111111100001011",
  43 => "1111111110110011",
  44 => "0000001100001000",
  45 => "0000000001000110",
  46 => "1111111110011001",
  47 => "1111111111011100",
  48 => "1111111100011011",
  49 => "0000000001011010",
  50 => "0000000000111011",
  51 => "1111111101000100",
  52 => "1111110011010111",
  53 => "1111110110100100",
  54 => "1110111101011010",
  55 => "1111111101101011",
  56 => "1111111110111111",
  57 => "1111111110110101",
  58 => "1111111111011110",
  59 => "1111111111100100",
  60 => "1111111110101001",
  61 => "1111111111100100",
  62 => "0000000010100100");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;