LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_7_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(6 DOWNTO 0));
END L7_7_BNROM;

ARCHITECTURE RTL OF L7_7_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"1111011111100100"&"0010000101010010",
  1=>"1110001010001101"&"0010100110101010",
  2=>"1110110001111101"&"0010100011011000",
  3=>"1101101000001000"&"0010101010001011",
  4=>"1111000111101100"&"0010010011011111",
  5=>"1111001101001000"&"0010000011010110",
  6=>"1110111010000011"&"0010100111011100",
  7=>"1110001001100110"&"0010100111001110",
  8=>"1110101101100101"&"0010010000000110",
  9=>"1110110100111001"&"0010101010010001",
  10=>"1111110000011101"&"0010100000000001",
  11=>"1110011110111100"&"0010011001010011",
  12=>"1110100110111101"&"0010001100000101",
  13=>"1110101010111111"&"0010101001001001",
  14=>"1111101000001100"&"0010001011011011",
  15=>"1111011100110111"&"0010001101011110",
  16=>"1110101101110010"&"0010111101111010",
  17=>"1110011001101101"&"0001111110101111",
  18=>"1111011011101110"&"0010001101110000",
  19=>"1111110010100100"&"0010110000101001",
  20=>"0000000001110100"&"0010010010101111",
  21=>"1111011000011011"&"0010011011000011",
  22=>"1110100101011110"&"0001111111010100",
  23=>"1110101011000010"&"0010001101111101",
  24=>"1110110110011110"&"0010011001010010",
  25=>"1110011111000101"&"0010010100111101",
  26=>"1110011000111101"&"0010110010000110",
  27=>"1110011000100011"&"0010101101010010",
  28=>"1110111101011101"&"0010010000111010",
  29=>"1111011001100101"&"0010001001010111",
  30=>"1111100110111011"&"0001011100100110",
  31=>"1111110110001100"&"0010010101110010",
  32=>"1111000101001000"&"0010001101001011",
  33=>"1111010001101011"&"0010101100100110",
  34=>"1101101110011010"&"0010101100010100",
  35=>"1110000100111011"&"0010011110110000",
  36=>"1110111011101110"&"0010011101101010",
  37=>"1101100010110100"&"0010011110110111",
  38=>"1110000111001111"&"0011000011001111",
  39=>"1111000010011100"&"0010101010110010",
  40=>"1111110001100000"&"0010010000100011",
  41=>"1110100001011100"&"0010110100011101",
  42=>"1111111001010010"&"0010011100001010",
  43=>"1110010110101111"&"0010010011011101",
  44=>"1101111010000111"&"0010100100001011",
  45=>"1110010110101101"&"0010001111110010",
  46=>"1101111101111010"&"0001111011110100",
  47=>"1110010101101001"&"0010011001101010",
  48=>"1111000101000011"&"0010001010000011",
  49=>"1110010110110010"&"0010111000110000",
  50=>"1110011100111101"&"0010011100001001",
  51=>"1111010010111110"&"0010000110010000",
  52=>"1111000011011001"&"0010011010100100",
  53=>"1110101011101110"&"0010011001100110",
  54=>"1111001100101001"&"0010001100111001",
  55=>"1111001111001101"&"0010010011100100",
  56=>"1111001101010101"&"0010011100001111",
  57=>"1111011011011111"&"0010010001000011",
  58=>"1110010101110010"&"0011000111101100",
  59=>"1111011111101010"&"0010001111110110",
  60=>"1110111101101111"&"0010100010011011",
  61=>"1110110010110101"&"0010010110101110",
  62=>"1111011101100110"&"0010001101111101",
  63=>"1111100100000101"&"0010101101111011",
  64=>"1111011011111100"&"0010001000110011",
  65=>"1110010011110110"&"0010101100110000",
  66=>"1110011100100111"&"0010010111000000",
  67=>"1111000101010111"&"0001111111010101",
  68=>"1110100010011010"&"0010100010101001",
  69=>"0000001100001110"&"0010010100111110",
  70=>"1110000101100101"&"0010001110110000",
  71=>"1111001011101001"&"0010011000011001",
  72=>"1111001100100010"&"0010000110010111",
  73=>"1110111000100011"&"0010011100110100",
  74=>"1111000011110101"&"0010010100011110",
  75=>"1111010001111000"&"0010010110101011",
  76=>"1110011100100101"&"0010011011011100",
  77=>"0000000100011101"&"0010000101110100",
  78=>"1110110100110011"&"0010000010011101",
  79=>"1110101000000111"&"0010011110100110",
  80=>"1110011010100101"&"0010011110000010",
  81=>"1110010010110010"&"0010010100100111",
  82=>"1111001010001101"&"0010011111110010",
  83=>"1111010001010110"&"0001111111000011",
  84=>"1111100101101011"&"0010001101010000",
  85=>"1111010000110101"&"0010010010000111",
  86=>"1110000011000101"&"0010110000110110",
  87=>"1111001111100100"&"0010100001000111",
  88=>"1110111000110001"&"0010010100110001",
  89=>"1110110111010010"&"0010101111110010",
  90=>"1111101101000001"&"0010001000000110",
  91=>"1110001110101000"&"0010110100001111",
  92=>"1110010000110010"&"0010011100101111",
  93=>"1110001001100010"&"0010101010101101",
  94=>"1110101000011101"&"0010001011101000",
  95=>"1101101010111010"&"0010001010111000",
  96=>"1111101101110110"&"0010001100100000",
  97=>"1110111010110000"&"0010010010111011",
  98=>"1110100101111000"&"0010001110000101",
  99=>"1111000001001010"&"0010010101101110",
  100=>"1111011011101001"&"0010000110010000",
  101=>"1110100010111110"&"0010010110001101",
  102=>"1110010100100000"&"0010100111000011",
  103=>"1111001010101011"&"0010011101000111",
  104=>"1101101010000111"&"0010011100100101",
  105=>"0000001000100101"&"0010001100000011",
  106=>"1111110010001100"&"0010001001010000",
  107=>"1111010101101011"&"0010101001110001",
  108=>"1101100011111111"&"0010101011010000",
  109=>"1111110000110010"&"0010111010100000",
  110=>"1110101111110101"&"0010001110100011",
  111=>"1111101001000111"&"0010100000010110",
  112=>"1110001010010010"&"0010101110111011",
  113=>"1111000010110010"&"0010001101011001",
  114=>"1110111111000010"&"0010100011110111",
  115=>"1110011110011011"&"0010010011100001",
  116=>"1110100011001101"&"0010001110000100",
  117=>"1110101000011111"&"0010010111101001",
  118=>"1111001001011001"&"0001111011110010",
  119=>"1110000110001000"&"0010111011110001",
  120=>"1111001011101111"&"0010101001011101",
  121=>"1111100000111011"&"0010001011010101",
  122=>"1111111011001100"&"0010001101111111",
  123=>"1110001001011000"&"0010110011001000",
  124=>"1111001001000010"&"0000110000110100",
  125=>"1110010001111101"&"0010011010001110",
  126=>"1110111001000100"&"0010100001000111",
  127=>"1110110110110011"&"0010010010001101");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;