LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_4_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_4_WROM;

ARCHITECTURE RTL OF L7_4_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"000000111",
  1=>"100110010",
  2=>"111111010",
  3=>"001101011",
  4=>"000110110",
  5=>"000100000",
  6=>"110110111",
  7=>"111111111",
  8=>"111001000",
  9=>"111111111",
  10=>"011111111",
  11=>"101000000",
  12=>"100100100",
  13=>"111100101",
  14=>"101111111",
  15=>"000110000",
  16=>"000000001",
  17=>"100100111",
  18=>"000000100",
  19=>"100000000",
  20=>"000000000",
  21=>"100000000",
  22=>"111101001",
  23=>"100100100",
  24=>"111111000",
  25=>"000110110",
  26=>"111001000",
  27=>"001000011",
  28=>"000100111",
  29=>"001000000",
  30=>"001010000",
  31=>"111001000",
  32=>"111001001",
  33=>"000000000",
  34=>"000110110",
  35=>"000000000",
  36=>"000100110",
  37=>"111111111",
  38=>"000000000",
  39=>"000000000",
  40=>"011111111",
  41=>"000000000",
  42=>"000001000",
  43=>"010111000",
  44=>"001111111",
  45=>"110101111",
  46=>"000000000",
  47=>"000000000",
  48=>"110110000",
  49=>"010000000",
  50=>"000000001",
  51=>"111111011",
  52=>"101001101",
  53=>"000001111",
  54=>"101100000",
  55=>"000100111",
  56=>"111111111",
  57=>"000000001",
  58=>"000000000",
  59=>"000000000",
  60=>"001001000",
  61=>"111111111",
  62=>"110101001",
  63=>"011111111",
  64=>"000011111",
  65=>"000000000",
  66=>"000101101",
  67=>"000000000",
  68=>"111111111",
  69=>"111111110",
  70=>"000000111",
  71=>"000000000",
  72=>"011011001",
  73=>"111111000",
  74=>"111111111",
  75=>"000000000",
  76=>"111111111",
  77=>"100000000",
  78=>"111000000",
  79=>"000000101",
  80=>"000000101",
  81=>"111001100",
  82=>"100111111",
  83=>"111111111",
  84=>"000000000",
  85=>"111111111",
  86=>"000000000",
  87=>"100100100",
  88=>"110010000",
  89=>"111101001",
  90=>"111000001",
  91=>"100100100",
  92=>"000000001",
  93=>"111111111",
  94=>"111000000",
  95=>"000001111",
  96=>"100000000",
  97=>"110000000",
  98=>"111111111",
  99=>"000000100",
  100=>"010110110",
  101=>"000000011",
  102=>"001001001",
  103=>"101101101",
  104=>"111000000",
  105=>"111111111",
  106=>"000000111",
  107=>"111111111",
  108=>"110111111",
  109=>"100100111",
  110=>"111111111",
  111=>"111111111",
  112=>"111111111",
  113=>"000000111",
  114=>"111111111",
  115=>"011000000",
  116=>"110111011",
  117=>"000000000",
  118=>"111111000",
  119=>"000000000",
  120=>"111111111",
  121=>"001000001",
  122=>"111101111",
  123=>"100000000",
  124=>"000101111",
  125=>"111111101",
  126=>"000000111",
  127=>"000000000",
  128=>"000000000",
  129=>"110000000",
  130=>"111001001",
  131=>"011011111",
  132=>"111111100",
  133=>"000000111",
  134=>"111111110",
  135=>"000110110",
  136=>"111101000",
  137=>"111001101",
  138=>"000000000",
  139=>"111111111",
  140=>"111111011",
  141=>"100000000",
  142=>"000111111",
  143=>"101100111",
  144=>"111001000",
  145=>"000000111",
  146=>"111101111",
  147=>"000000000",
  148=>"000000110",
  149=>"000000000",
  150=>"111111111",
  151=>"111001001",
  152=>"000000000",
  153=>"001100110",
  154=>"111100000",
  155=>"111111010",
  156=>"111111000",
  157=>"111001001",
  158=>"000000111",
  159=>"111000000",
  160=>"111100111",
  161=>"101001011",
  162=>"000000000",
  163=>"111111111",
  164=>"000000000",
  165=>"000010110",
  166=>"000000111",
  167=>"110110110",
  168=>"111000000",
  169=>"000000000",
  170=>"111100110",
  171=>"000010111",
  172=>"110111111",
  173=>"111111000",
  174=>"001000000",
  175=>"110111011",
  176=>"000000000",
  177=>"001000000",
  178=>"000000111",
  179=>"111101000",
  180=>"000101101",
  181=>"000000000",
  182=>"000000001",
  183=>"101101000",
  184=>"010111111",
  185=>"001000000",
  186=>"110111001",
  187=>"100101111",
  188=>"111111111",
  189=>"111111100",
  190=>"000000000",
  191=>"011001000",
  192=>"111001000",
  193=>"001111111",
  194=>"111001001",
  195=>"111111111",
  196=>"110111111",
  197=>"000000000",
  198=>"000000000",
  199=>"111111000",
  200=>"110000000",
  201=>"010110100",
  202=>"010000000",
  203=>"111111111",
  204=>"111111000",
  205=>"011011011",
  206=>"100000000",
  207=>"111100000",
  208=>"110011000",
  209=>"000000000",
  210=>"101101111",
  211=>"110110000",
  212=>"011000000",
  213=>"111111111",
  214=>"011001011",
  215=>"000000110",
  216=>"000000011",
  217=>"000100111",
  218=>"000000000",
  219=>"111111000",
  220=>"111111111",
  221=>"011011011",
  222=>"000111111",
  223=>"000000000",
  224=>"111111111",
  225=>"010010111",
  226=>"111000110",
  227=>"111000010",
  228=>"000110111",
  229=>"011001001",
  230=>"100100111",
  231=>"000000001",
  232=>"101101111",
  233=>"000010011",
  234=>"110000000",
  235=>"111111101",
  236=>"000000001",
  237=>"101000111",
  238=>"111110010",
  239=>"000001111",
  240=>"111111110",
  241=>"111111111",
  242=>"101000100",
  243=>"111101101",
  244=>"000000000",
  245=>"110110100",
  246=>"110110000",
  247=>"000000101",
  248=>"000000111",
  249=>"110101101",
  250=>"010000000",
  251=>"000000000",
  252=>"011001011",
  253=>"100110111",
  254=>"111001001",
  255=>"001001000",
  256=>"011000001",
  257=>"111111000",
  258=>"111001111",
  259=>"111001000",
  260=>"111111111",
  261=>"000100110",
  262=>"000000000",
  263=>"111111011",
  264=>"110100001",
  265=>"111111111",
  266=>"000000001",
  267=>"000001011",
  268=>"000000110",
  269=>"111111110",
  270=>"111001001",
  271=>"111111111",
  272=>"000001001",
  273=>"111000101",
  274=>"000000000",
  275=>"001100100",
  276=>"000101111",
  277=>"000000111",
  278=>"100000000",
  279=>"101111000",
  280=>"011110111",
  281=>"000000000",
  282=>"001001000",
  283=>"111110001",
  284=>"000000000",
  285=>"000000110",
  286=>"111111000",
  287=>"001000111",
  288=>"111111111",
  289=>"111001001",
  290=>"000000000",
  291=>"111111111",
  292=>"000100000",
  293=>"111111100",
  294=>"111111111",
  295=>"010000010",
  296=>"100110110",
  297=>"000000000",
  298=>"011001100",
  299=>"001111001",
  300=>"000000000",
  301=>"111011001",
  302=>"000000000",
  303=>"000011111",
  304=>"000000000",
  305=>"111111111",
  306=>"111111111",
  307=>"100100111",
  308=>"111111000",
  309=>"101000101",
  310=>"111110000",
  311=>"000000000",
  312=>"111111000",
  313=>"000000111",
  314=>"101000000",
  315=>"000000000",
  316=>"001001011",
  317=>"111111011",
  318=>"010010010",
  319=>"000111111",
  320=>"000010000",
  321=>"111111111",
  322=>"111111000",
  323=>"111111000",
  324=>"111111111",
  325=>"000000000",
  326=>"111111100",
  327=>"111111110",
  328=>"111000000",
  329=>"000000000",
  330=>"110111000",
  331=>"011011011",
  332=>"000001101",
  333=>"100111111",
  334=>"100100111",
  335=>"000010110",
  336=>"011001001",
  337=>"000000111",
  338=>"111111111",
  339=>"111110010",
  340=>"000000000",
  341=>"001000001",
  342=>"111001000",
  343=>"000000000",
  344=>"000000000",
  345=>"000000000",
  346=>"111111100",
  347=>"001111111",
  348=>"000000000",
  349=>"111111111",
  350=>"000000000",
  351=>"111111111",
  352=>"000011000",
  353=>"110000110",
  354=>"100111110",
  355=>"000111111",
  356=>"111001000",
  357=>"001000111",
  358=>"001111100",
  359=>"101111000",
  360=>"111101100",
  361=>"000110111",
  362=>"000000000",
  363=>"000010000",
  364=>"111110110",
  365=>"111111100",
  366=>"000000000",
  367=>"111111111",
  368=>"110111111",
  369=>"110000000",
  370=>"011000000",
  371=>"011011011",
  372=>"111000000",
  373=>"111111010",
  374=>"111110000",
  375=>"111010000",
  376=>"000000011",
  377=>"011000110",
  378=>"110000000",
  379=>"111100000",
  380=>"000000000",
  381=>"001000000",
  382=>"111111111",
  383=>"111110000",
  384=>"001001110",
  385=>"111111111",
  386=>"111111111",
  387=>"000000100",
  388=>"000000000",
  389=>"110111111",
  390=>"111110000",
  391=>"111110100",
  392=>"011111111",
  393=>"111101000",
  394=>"000100000",
  395=>"110111111",
  396=>"111101001",
  397=>"000001001",
  398=>"011001001",
  399=>"011111000",
  400=>"111111111",
  401=>"000000000",
  402=>"111111101",
  403=>"111111110",
  404=>"001101111",
  405=>"000000000",
  406=>"111110110",
  407=>"011001001",
  408=>"000000000",
  409=>"000000111",
  410=>"011000010",
  411=>"110100100",
  412=>"100101111",
  413=>"111111000",
  414=>"000000000",
  415=>"000000100",
  416=>"111100000",
  417=>"111111111",
  418=>"001001101",
  419=>"000000000",
  420=>"010111111",
  421=>"110110000",
  422=>"000001111",
  423=>"111111000",
  424=>"111000000",
  425=>"110010000",
  426=>"111110100",
  427=>"111010000",
  428=>"000000000",
  429=>"111101101",
  430=>"110110000",
  431=>"111110000",
  432=>"111111100",
  433=>"111111010",
  434=>"111110100",
  435=>"111100110",
  436=>"110111111",
  437=>"000000000",
  438=>"100111111",
  439=>"111111101",
  440=>"000111111",
  441=>"111111111",
  442=>"111111010",
  443=>"111111001",
  444=>"100000000",
  445=>"011111111",
  446=>"000000010",
  447=>"101111100",
  448=>"011111111",
  449=>"000000000",
  450=>"111111011",
  451=>"111111000",
  452=>"010000010",
  453=>"000110110",
  454=>"111010010",
  455=>"000000000",
  456=>"010000000",
  457=>"111000000",
  458=>"000000010",
  459=>"000001001",
  460=>"000000000",
  461=>"111111111",
  462=>"100000000",
  463=>"110010000",
  464=>"000000000",
  465=>"111111111",
  466=>"000011111",
  467=>"000000000",
  468=>"100100111",
  469=>"000100110",
  470=>"000000000",
  471=>"001001001",
  472=>"100111111",
  473=>"000000110",
  474=>"111111100",
  475=>"111011001",
  476=>"000000000",
  477=>"000001111",
  478=>"100100000",
  479=>"000111001",
  480=>"000000111",
  481=>"000000000",
  482=>"001000000",
  483=>"001111111",
  484=>"111111111",
  485=>"001101111",
  486=>"111001001",
  487=>"000000000",
  488=>"000000111",
  489=>"001101111",
  490=>"000110111",
  491=>"000001111",
  492=>"111111101",
  493=>"111000000",
  494=>"100111000",
  495=>"111111111",
  496=>"100000100",
  497=>"111100000",
  498=>"000000000",
  499=>"110100111",
  500=>"000011111",
  501=>"000000000",
  502=>"000000111",
  503=>"101001001",
  504=>"000000000",
  505=>"011000001",
  506=>"110111111",
  507=>"111111011",
  508=>"111110000",
  509=>"110110111",
  510=>"111111111",
  511=>"000011000",
  512=>"011001000",
  513=>"111111011",
  514=>"000000000",
  515=>"011111110",
  516=>"001001111",
  517=>"110101000",
  518=>"001001001",
  519=>"000111111",
  520=>"000000000",
  521=>"101001001",
  522=>"111111001",
  523=>"000011111",
  524=>"111110000",
  525=>"111001000",
  526=>"001111111",
  527=>"110000000",
  528=>"111000000",
  529=>"100100111",
  530=>"111111111",
  531=>"010100100",
  532=>"111011000",
  533=>"101100110",
  534=>"110111111",
  535=>"111110011",
  536=>"111111111",
  537=>"000001011",
  538=>"000000000",
  539=>"000000000",
  540=>"001001111",
  541=>"110000001",
  542=>"011011110",
  543=>"100111111",
  544=>"100000000",
  545=>"011111111",
  546=>"000000000",
  547=>"000000000",
  548=>"011010000",
  549=>"111101100",
  550=>"011011010",
  551=>"011111000",
  552=>"111110000",
  553=>"000000011",
  554=>"000000100",
  555=>"000001000",
  556=>"000000000",
  557=>"000100111",
  558=>"011111111",
  559=>"000000000",
  560=>"011110011",
  561=>"000011111",
  562=>"111101111",
  563=>"000111110",
  564=>"110100000",
  565=>"000011011",
  566=>"110110111",
  567=>"111011110",
  568=>"001000101",
  569=>"001111111",
  570=>"000000000",
  571=>"111111000",
  572=>"111111111",
  573=>"100001111",
  574=>"000000000",
  575=>"000111001",
  576=>"111111011",
  577=>"110111111",
  578=>"111001000",
  579=>"111111110",
  580=>"001001111",
  581=>"001000000",
  582=>"000110100",
  583=>"000000000",
  584=>"111111111",
  585=>"100000100",
  586=>"000000100",
  587=>"001101000",
  588=>"111011001",
  589=>"001000011",
  590=>"111111111",
  591=>"101111111",
  592=>"100000000",
  593=>"010111011",
  594=>"111100111",
  595=>"110110110",
  596=>"100000001",
  597=>"000001111",
  598=>"100000111",
  599=>"101001000",
  600=>"111111110",
  601=>"000000111",
  602=>"111111111",
  603=>"111011111",
  604=>"111111111",
  605=>"000000000",
  606=>"111100100",
  607=>"111111111",
  608=>"111110110",
  609=>"111111111",
  610=>"000010000",
  611=>"110000111",
  612=>"000100111",
  613=>"000100111",
  614=>"000000010",
  615=>"000110110",
  616=>"111111111",
  617=>"100000001",
  618=>"111111111",
  619=>"111111111",
  620=>"000000000",
  621=>"000000000",
  622=>"111111111",
  623=>"111111010",
  624=>"000001111",
  625=>"011111111",
  626=>"111110010",
  627=>"111111000",
  628=>"111111111",
  629=>"111111110",
  630=>"001000111",
  631=>"101000000",
  632=>"111101100",
  633=>"111111111",
  634=>"011011111",
  635=>"101001111",
  636=>"001011001",
  637=>"010000000",
  638=>"111011111",
  639=>"000000000",
  640=>"000000000",
  641=>"101000000",
  642=>"111111111",
  643=>"011111111",
  644=>"111111011",
  645=>"000100001",
  646=>"111111111",
  647=>"111111111",
  648=>"111001111",
  649=>"000000001",
  650=>"111001101",
  651=>"000000001",
  652=>"000010000",
  653=>"101000000",
  654=>"011111111",
  655=>"111111111",
  656=>"001001101",
  657=>"000000000",
  658=>"111101101",
  659=>"001101001",
  660=>"001000000",
  661=>"110011000",
  662=>"011000000",
  663=>"111111111",
  664=>"111110111",
  665=>"111011011",
  666=>"110111111",
  667=>"111111111",
  668=>"111110110",
  669=>"111111101",
  670=>"111111001",
  671=>"000011110",
  672=>"100100111",
  673=>"111111111",
  674=>"000000000",
  675=>"111100111",
  676=>"111011000",
  677=>"001001001",
  678=>"000000000",
  679=>"100000000",
  680=>"000000000",
  681=>"000000000",
  682=>"111111111",
  683=>"000000000",
  684=>"000100000",
  685=>"011011011",
  686=>"001001000",
  687=>"000000000",
  688=>"000110110",
  689=>"000100100",
  690=>"000000000",
  691=>"000000000",
  692=>"111111111",
  693=>"010011001",
  694=>"000000000",
  695=>"011001100",
  696=>"100000011",
  697=>"000000111",
  698=>"111111111",
  699=>"001011011",
  700=>"000000000",
  701=>"000101000",
  702=>"111001011",
  703=>"111101000",
  704=>"000000000",
  705=>"000001001",
  706=>"111111100",
  707=>"111111111",
  708=>"000000000",
  709=>"011111010",
  710=>"111111000",
  711=>"000000111",
  712=>"010110010",
  713=>"000110110",
  714=>"111111111",
  715=>"000001000",
  716=>"111111000",
  717=>"111111111",
  718=>"111111111",
  719=>"001111111",
  720=>"111101001",
  721=>"111010111",
  722=>"111011001",
  723=>"000000000",
  724=>"101001011",
  725=>"001001100",
  726=>"000000000",
  727=>"000000000",
  728=>"001111111",
  729=>"000000001",
  730=>"111111111",
  731=>"000001011",
  732=>"000010000",
  733=>"000000001",
  734=>"101110110",
  735=>"001011011",
  736=>"100100111",
  737=>"000000000",
  738=>"111010000",
  739=>"000000000",
  740=>"111011011",
  741=>"110111111",
  742=>"000000001",
  743=>"001001000",
  744=>"111111111",
  745=>"100000011",
  746=>"010111001",
  747=>"000000000",
  748=>"100100100",
  749=>"111110111",
  750=>"111000000",
  751=>"011000000",
  752=>"111000000",
  753=>"011011011",
  754=>"010000011",
  755=>"000011111",
  756=>"111001000",
  757=>"111111111",
  758=>"001101111",
  759=>"111010011",
  760=>"111111000",
  761=>"100111111",
  762=>"000000000",
  763=>"111111110",
  764=>"101001001",
  765=>"000111101",
  766=>"101111111",
  767=>"011110110",
  768=>"000000000",
  769=>"001001001",
  770=>"101000001",
  771=>"100011111",
  772=>"111111111",
  773=>"000001101",
  774=>"000000000",
  775=>"011111101",
  776=>"000000000",
  777=>"111111111",
  778=>"111110110",
  779=>"111111111",
  780=>"000000001",
  781=>"000100111",
  782=>"111101111",
  783=>"111100110",
  784=>"000101101",
  785=>"000000000",
  786=>"110111111",
  787=>"000000001",
  788=>"000000000",
  789=>"111111111",
  790=>"001001000",
  791=>"011111111",
  792=>"100101000",
  793=>"000000000",
  794=>"101001000",
  795=>"111111111",
  796=>"000001111",
  797=>"111111111",
  798=>"001011011",
  799=>"100111011",
  800=>"011111111",
  801=>"010011111",
  802=>"111100111",
  803=>"000100110",
  804=>"000010111",
  805=>"111111111",
  806=>"111111001",
  807=>"001000000",
  808=>"000000000",
  809=>"001111111",
  810=>"001011110",
  811=>"000000100",
  812=>"010111011",
  813=>"101011000",
  814=>"111010111",
  815=>"111111111",
  816=>"000000000",
  817=>"111010110",
  818=>"100000000",
  819=>"110100000",
  820=>"000000111",
  821=>"111111000",
  822=>"001011011",
  823=>"110010000",
  824=>"000100111",
  825=>"011111111",
  826=>"000000000",
  827=>"101111111",
  828=>"000000000",
  829=>"011111000",
  830=>"101001101",
  831=>"001111010",
  832=>"000000000",
  833=>"111000000",
  834=>"011111111",
  835=>"000000010",
  836=>"111111111",
  837=>"000001000",
  838=>"000000000",
  839=>"111111111",
  840=>"000000000",
  841=>"111010011",
  842=>"110111111",
  843=>"101100110",
  844=>"101100010",
  845=>"111111000",
  846=>"101100001",
  847=>"100100100",
  848=>"000000000",
  849=>"000000011",
  850=>"000000000",
  851=>"000000000",
  852=>"111000000",
  853=>"111111111",
  854=>"111000001",
  855=>"000001000",
  856=>"111101100",
  857=>"000000000",
  858=>"000000101",
  859=>"110011111",
  860=>"110010011",
  861=>"000000000",
  862=>"000000000",
  863=>"011000000",
  864=>"111011111",
  865=>"001011001",
  866=>"111001001",
  867=>"000000000",
  868=>"000000000",
  869=>"101111111",
  870=>"100100111",
  871=>"111011111",
  872=>"111011011",
  873=>"000010000",
  874=>"101111001",
  875=>"001011111",
  876=>"000110110",
  877=>"011000000",
  878=>"011000000",
  879=>"001011111",
  880=>"111000100",
  881=>"111111111",
  882=>"110100111",
  883=>"011001100",
  884=>"101101100",
  885=>"000111111",
  886=>"111111101",
  887=>"111000110",
  888=>"111111111",
  889=>"011011000",
  890=>"111101100",
  891=>"111111111",
  892=>"000110110",
  893=>"000000111",
  894=>"111000101",
  895=>"111111100",
  896=>"000100110",
  897=>"110110111",
  898=>"000000001",
  899=>"000000000",
  900=>"010111111",
  901=>"110111111",
  902=>"111111111",
  903=>"011011011",
  904=>"001001001",
  905=>"100000011",
  906=>"111111111",
  907=>"110110000",
  908=>"000000000",
  909=>"000000100",
  910=>"011111111",
  911=>"100111000",
  912=>"111111111",
  913=>"000001011",
  914=>"011001000",
  915=>"000000000",
  916=>"000111111",
  917=>"111111111",
  918=>"100111111",
  919=>"000001111",
  920=>"111001000",
  921=>"111001111",
  922=>"000000011",
  923=>"001011000",
  924=>"000000000",
  925=>"000000001",
  926=>"100100000",
  927=>"111111111",
  928=>"111111011",
  929=>"011000000",
  930=>"100111111",
  931=>"011011011",
  932=>"111111111",
  933=>"000000000",
  934=>"000110111",
  935=>"011000000",
  936=>"110000000",
  937=>"010010010",
  938=>"000000000",
  939=>"000000110",
  940=>"010001000",
  941=>"110110111",
  942=>"101101111",
  943=>"000000000",
  944=>"000000000",
  945=>"111111111",
  946=>"111111000",
  947=>"001001111",
  948=>"110111111",
  949=>"001111011",
  950=>"110111111",
  951=>"011111111",
  952=>"011111001",
  953=>"111111111",
  954=>"000010010",
  955=>"100000000",
  956=>"100110000",
  957=>"000000100",
  958=>"110111101",
  959=>"001011010",
  960=>"001001111",
  961=>"001100000",
  962=>"001000000",
  963=>"000000000",
  964=>"000010010",
  965=>"000001001",
  966=>"011111011",
  967=>"110111111",
  968=>"111011111",
  969=>"101011111",
  970=>"000010111",
  971=>"000000000",
  972=>"000011000",
  973=>"000000000",
  974=>"111011111",
  975=>"101111011",
  976=>"000101111",
  977=>"000111010",
  978=>"000000000",
  979=>"000010000",
  980=>"110111111",
  981=>"001011011",
  982=>"101101000",
  983=>"100000110",
  984=>"000110110",
  985=>"001001001",
  986=>"101100100",
  987=>"000000011",
  988=>"111111111",
  989=>"000001111",
  990=>"000000000",
  991=>"111111111",
  992=>"100001111",
  993=>"110000000",
  994=>"011010000",
  995=>"000000010",
  996=>"000010111",
  997=>"100110111",
  998=>"011111100",
  999=>"101000000",
  1000=>"000001001",
  1001=>"011010011",
  1002=>"000000000",
  1003=>"010010000",
  1004=>"111011100",
  1005=>"000000000",
  1006=>"110000000",
  1007=>"000110010",
  1008=>"100101000",
  1009=>"111111110",
  1010=>"111111111",
  1011=>"000011011",
  1012=>"011001000",
  1013=>"001111111",
  1014=>"001000000",
  1015=>"000000001",
  1016=>"010010000",
  1017=>"100110000",
  1018=>"110111111",
  1019=>"111111111",
  1020=>"111111111",
  1021=>"111110000",
  1022=>"000000111",
  1023=>"000000111",
  1024=>"001000001",
  1025=>"110111000",
  1026=>"000000000",
  1027=>"000000000",
  1028=>"100101111",
  1029=>"011000000",
  1030=>"100110000",
  1031=>"000000000",
  1032=>"011010111",
  1033=>"111111111",
  1034=>"100100000",
  1035=>"111000110",
  1036=>"100111110",
  1037=>"001001111",
  1038=>"000000000",
  1039=>"100100100",
  1040=>"110000000",
  1041=>"000010111",
  1042=>"001001001",
  1043=>"000000100",
  1044=>"000000000",
  1045=>"111111111",
  1046=>"001111111",
  1047=>"111011000",
  1048=>"000000110",
  1049=>"000100010",
  1050=>"000000000",
  1051=>"100000000",
  1052=>"110110110",
  1053=>"011011111",
  1054=>"101101001",
  1055=>"011111011",
  1056=>"111011000",
  1057=>"100000000",
  1058=>"110000000",
  1059=>"000000000",
  1060=>"000000000",
  1061=>"001001001",
  1062=>"111111000",
  1063=>"111111111",
  1064=>"111000000",
  1065=>"111100000",
  1066=>"000000000",
  1067=>"110110110",
  1068=>"111001111",
  1069=>"111111111",
  1070=>"000101001",
  1071=>"110111111",
  1072=>"000111111",
  1073=>"000100100",
  1074=>"001001000",
  1075=>"000000000",
  1076=>"000001001",
  1077=>"111111110",
  1078=>"000011001",
  1079=>"011011111",
  1080=>"111111111",
  1081=>"000000000",
  1082=>"111111000",
  1083=>"111111111",
  1084=>"000000000",
  1085=>"000000011",
  1086=>"001111111",
  1087=>"000000000",
  1088=>"000010010",
  1089=>"011111001",
  1090=>"111110000",
  1091=>"110000000",
  1092=>"000000000",
  1093=>"100110100",
  1094=>"010000000",
  1095=>"111111111",
  1096=>"011010110",
  1097=>"001001011",
  1098=>"000010110",
  1099=>"001000111",
  1100=>"000000111",
  1101=>"111111111",
  1102=>"111111101",
  1103=>"111111111",
  1104=>"000000000",
  1105=>"000011011",
  1106=>"000000000",
  1107=>"100111010",
  1108=>"111111101",
  1109=>"000010010",
  1110=>"111100000",
  1111=>"000001000",
  1112=>"111010001",
  1113=>"011100111",
  1114=>"001011111",
  1115=>"000000001",
  1116=>"100100000",
  1117=>"001111000",
  1118=>"010100111",
  1119=>"010000000",
  1120=>"000000000",
  1121=>"111001001",
  1122=>"000000000",
  1123=>"000000000",
  1124=>"100000000",
  1125=>"000000000",
  1126=>"000000000",
  1127=>"111111111",
  1128=>"000000000",
  1129=>"111111111",
  1130=>"000000000",
  1131=>"111111111",
  1132=>"000100111",
  1133=>"111111111",
  1134=>"111111111",
  1135=>"000000000",
  1136=>"111111011",
  1137=>"000111111",
  1138=>"011011011",
  1139=>"111111000",
  1140=>"000000000",
  1141=>"110000100",
  1142=>"110111111",
  1143=>"011000111",
  1144=>"111110101",
  1145=>"110111111",
  1146=>"111010000",
  1147=>"001000001",
  1148=>"111100100",
  1149=>"000000000",
  1150=>"000111011",
  1151=>"111000000",
  1152=>"000010000",
  1153=>"000000000",
  1154=>"000000000",
  1155=>"111010010",
  1156=>"111111111",
  1157=>"000000000",
  1158=>"000010000",
  1159=>"000000001",
  1160=>"000100100",
  1161=>"000011111",
  1162=>"000000000",
  1163=>"000000000",
  1164=>"000000111",
  1165=>"000000000",
  1166=>"000011111",
  1167=>"111111111",
  1168=>"001000111",
  1169=>"101000000",
  1170=>"000011000",
  1171=>"000111110",
  1172=>"000000000",
  1173=>"110110000",
  1174=>"000100111",
  1175=>"010000110",
  1176=>"110000010",
  1177=>"111111111",
  1178=>"100000000",
  1179=>"000111010",
  1180=>"111111111",
  1181=>"011111000",
  1182=>"111111111",
  1183=>"000110111",
  1184=>"111111111",
  1185=>"101001000",
  1186=>"111111001",
  1187=>"000000010",
  1188=>"100011011",
  1189=>"100000110",
  1190=>"101000000",
  1191=>"111111001",
  1192=>"111000000",
  1193=>"000000000",
  1194=>"010000000",
  1195=>"111001001",
  1196=>"111111111",
  1197=>"011000111",
  1198=>"000000000",
  1199=>"000000111",
  1200=>"000000000",
  1201=>"000011011",
  1202=>"101000000",
  1203=>"111000100",
  1204=>"111111111",
  1205=>"111010110",
  1206=>"000000000",
  1207=>"000000111",
  1208=>"111111101",
  1209=>"000000000",
  1210=>"010111111",
  1211=>"111111111",
  1212=>"000000000",
  1213=>"000000000",
  1214=>"111111111",
  1215=>"111111110",
  1216=>"000000011",
  1217=>"000000000",
  1218=>"000000000",
  1219=>"000000000",
  1220=>"111111111",
  1221=>"011001000",
  1222=>"111111011",
  1223=>"111111000",
  1224=>"011111111",
  1225=>"111111000",
  1226=>"111001000",
  1227=>"000110111",
  1228=>"001011111",
  1229=>"000000000",
  1230=>"110100000",
  1231=>"000000000",
  1232=>"000000000",
  1233=>"000001000",
  1234=>"100100000",
  1235=>"000000000",
  1236=>"000111111",
  1237=>"001011000",
  1238=>"000001001",
  1239=>"110000011",
  1240=>"111111111",
  1241=>"100110000",
  1242=>"111011000",
  1243=>"111111110",
  1244=>"111111111",
  1245=>"000000111",
  1246=>"000000000",
  1247=>"111111110",
  1248=>"000000010",
  1249=>"001001111",
  1250=>"000000010",
  1251=>"111011110",
  1252=>"110111111",
  1253=>"100110010",
  1254=>"010001001",
  1255=>"111111110",
  1256=>"111111111",
  1257=>"101111011",
  1258=>"111111111",
  1259=>"011111110",
  1260=>"111111111",
  1261=>"000000000",
  1262=>"000100001",
  1263=>"000000000",
  1264=>"001010000",
  1265=>"100010000",
  1266=>"000111111",
  1267=>"111000000",
  1268=>"011011010",
  1269=>"110000001",
  1270=>"111111111",
  1271=>"111011111",
  1272=>"000000000",
  1273=>"000110111",
  1274=>"100100110",
  1275=>"111011011",
  1276=>"001011011",
  1277=>"110000000",
  1278=>"111111111",
  1279=>"011111111",
  1280=>"111111011",
  1281=>"000000000",
  1282=>"111111111",
  1283=>"000000000",
  1284=>"111111111",
  1285=>"011000000",
  1286=>"000000000",
  1287=>"110110110",
  1288=>"111111111",
  1289=>"111111111",
  1290=>"111110000",
  1291=>"111111110",
  1292=>"000000001",
  1293=>"000000000",
  1294=>"111111000",
  1295=>"000000000",
  1296=>"111111011",
  1297=>"000010000",
  1298=>"001001011",
  1299=>"010101100",
  1300=>"000000000",
  1301=>"100000000",
  1302=>"001011001",
  1303=>"000000000",
  1304=>"000000000",
  1305=>"010110111",
  1306=>"111101111",
  1307=>"111000000",
  1308=>"111111111",
  1309=>"111000000",
  1310=>"111111010",
  1311=>"100101000",
  1312=>"111111000",
  1313=>"100000000",
  1314=>"000000000",
  1315=>"111110110",
  1316=>"011001101",
  1317=>"000000000",
  1318=>"000011111",
  1319=>"000000000",
  1320=>"111111111",
  1321=>"111000000",
  1322=>"011000000",
  1323=>"000000000",
  1324=>"011111010",
  1325=>"110000000",
  1326=>"000000000",
  1327=>"111111000",
  1328=>"111111111",
  1329=>"111111111",
  1330=>"101000101",
  1331=>"000001111",
  1332=>"001001101",
  1333=>"111111111",
  1334=>"111111111",
  1335=>"110100100",
  1336=>"000000000",
  1337=>"000000100",
  1338=>"001100000",
  1339=>"011010000",
  1340=>"000000000",
  1341=>"011111011",
  1342=>"111011101",
  1343=>"000000000",
  1344=>"010010001",
  1345=>"111111111",
  1346=>"000000000",
  1347=>"000000101",
  1348=>"001000000",
  1349=>"111111111",
  1350=>"001000000",
  1351=>"101000001",
  1352=>"000000000",
  1353=>"000000000",
  1354=>"111111111",
  1355=>"110110100",
  1356=>"000000000",
  1357=>"001000000",
  1358=>"111000000",
  1359=>"011111111",
  1360=>"001100100",
  1361=>"000000000",
  1362=>"100000000",
  1363=>"111111111",
  1364=>"000000000",
  1365=>"011001001",
  1366=>"000000000",
  1367=>"000111111",
  1368=>"001111110",
  1369=>"111111001",
  1370=>"000100010",
  1371=>"000000111",
  1372=>"001001111",
  1373=>"111111111",
  1374=>"101100000",
  1375=>"111100000",
  1376=>"011111111",
  1377=>"111111111",
  1378=>"001101011",
  1379=>"000000000",
  1380=>"111111110",
  1381=>"000000000",
  1382=>"000000000",
  1383=>"111111111",
  1384=>"110011001",
  1385=>"000000000",
  1386=>"000110110",
  1387=>"111011010",
  1388=>"111110000",
  1389=>"110110000",
  1390=>"000000000",
  1391=>"000000000",
  1392=>"000000000",
  1393=>"000000100",
  1394=>"000000000",
  1395=>"111010011",
  1396=>"000110111",
  1397=>"111111111",
  1398=>"000000000",
  1399=>"010010001",
  1400=>"000001001",
  1401=>"111111111",
  1402=>"000000000",
  1403=>"111110111",
  1404=>"111011111",
  1405=>"110010010",
  1406=>"111011000",
  1407=>"111000000",
  1408=>"100111110",
  1409=>"000000000",
  1410=>"000111111",
  1411=>"111111110",
  1412=>"111111111",
  1413=>"000000011",
  1414=>"111011111",
  1415=>"000111111",
  1416=>"101111111",
  1417=>"011000111",
  1418=>"110111111",
  1419=>"011111001",
  1420=>"111111111",
  1421=>"000000010",
  1422=>"101111111",
  1423=>"000000000",
  1424=>"000000000",
  1425=>"101000010",
  1426=>"000100000",
  1427=>"000110000",
  1428=>"111111111",
  1429=>"000000000",
  1430=>"000111111",
  1431=>"110000011",
  1432=>"010111000",
  1433=>"111111101",
  1434=>"111111011",
  1435=>"111111111",
  1436=>"111111011",
  1437=>"001101111",
  1438=>"000011001",
  1439=>"110111111",
  1440=>"000000000",
  1441=>"011001011",
  1442=>"111111111",
  1443=>"111111111",
  1444=>"001000000",
  1445=>"111111111",
  1446=>"000000000",
  1447=>"111111111",
  1448=>"001100000",
  1449=>"111111000",
  1450=>"000000000",
  1451=>"000001111",
  1452=>"111000000",
  1453=>"001111000",
  1454=>"111111101",
  1455=>"000000100",
  1456=>"111011111",
  1457=>"000000101",
  1458=>"100000111",
  1459=>"000000000",
  1460=>"000100111",
  1461=>"111111111",
  1462=>"000000010",
  1463=>"000000000",
  1464=>"000000000",
  1465=>"111111111",
  1466=>"111010000",
  1467=>"111010000",
  1468=>"111111111",
  1469=>"110110110",
  1470=>"000000000",
  1471=>"000000000",
  1472=>"111111111",
  1473=>"100000000",
  1474=>"101000000",
  1475=>"000000000",
  1476=>"111111110",
  1477=>"001000000",
  1478=>"111111111",
  1479=>"000000000",
  1480=>"111111001",
  1481=>"000000000",
  1482=>"111111111",
  1483=>"111111001",
  1484=>"111011101",
  1485=>"000000000",
  1486=>"000001000",
  1487=>"111000000",
  1488=>"111111000",
  1489=>"010010111",
  1490=>"000000000",
  1491=>"111000000",
  1492=>"000001001",
  1493=>"111110111",
  1494=>"010011011",
  1495=>"111011011",
  1496=>"000000000",
  1497=>"111000000",
  1498=>"010000000",
  1499=>"100000000",
  1500=>"000111111",
  1501=>"100110010",
  1502=>"111110100",
  1503=>"001101110",
  1504=>"000000100",
  1505=>"111101101",
  1506=>"111000000",
  1507=>"111111111",
  1508=>"000000001",
  1509=>"000000000",
  1510=>"111000000",
  1511=>"111011000",
  1512=>"000000000",
  1513=>"000000000",
  1514=>"111000000",
  1515=>"100110100",
  1516=>"000111111",
  1517=>"111111111",
  1518=>"100000000",
  1519=>"111001001",
  1520=>"100100111",
  1521=>"111110111",
  1522=>"000000000",
  1523=>"000000000",
  1524=>"001000000",
  1525=>"000000000",
  1526=>"111011011",
  1527=>"000000000",
  1528=>"111111111",
  1529=>"000000000",
  1530=>"110111111",
  1531=>"001000000",
  1532=>"111111111",
  1533=>"111101000",
  1534=>"000011011",
  1535=>"100000000",
  1536=>"101101100",
  1537=>"000000000",
  1538=>"100100000",
  1539=>"001000000",
  1540=>"111111110",
  1541=>"111111001",
  1542=>"000000000",
  1543=>"111111111",
  1544=>"000101000",
  1545=>"111101000",
  1546=>"100100000",
  1547=>"111111111",
  1548=>"000111100",
  1549=>"111111011",
  1550=>"110110111",
  1551=>"000000000",
  1552=>"111111111",
  1553=>"100100100",
  1554=>"000111000",
  1555=>"000001000",
  1556=>"000010111",
  1557=>"011001001",
  1558=>"000000000",
  1559=>"111001111",
  1560=>"100100100",
  1561=>"100100000",
  1562=>"000000000",
  1563=>"000010000",
  1564=>"110000000",
  1565=>"000000000",
  1566=>"111110100",
  1567=>"111101001",
  1568=>"000000110",
  1569=>"101001000",
  1570=>"001011111",
  1571=>"111111111",
  1572=>"111111111",
  1573=>"111000001",
  1574=>"111000010",
  1575=>"111100111",
  1576=>"111111111",
  1577=>"000000000",
  1578=>"101111111",
  1579=>"111111111",
  1580=>"111111111",
  1581=>"100111111",
  1582=>"111111111",
  1583=>"000110111",
  1584=>"000000000",
  1585=>"001000000",
  1586=>"001000000",
  1587=>"111111011",
  1588=>"010111000",
  1589=>"100110110",
  1590=>"000110010",
  1591=>"110110110",
  1592=>"011111100",
  1593=>"111011111",
  1594=>"000000001",
  1595=>"111000000",
  1596=>"000000000",
  1597=>"000000000",
  1598=>"000000000",
  1599=>"000000000",
  1600=>"111111000",
  1601=>"111111111",
  1602=>"000000000",
  1603=>"111000000",
  1604=>"111111001",
  1605=>"000111111",
  1606=>"111111000",
  1607=>"000000101",
  1608=>"000000001",
  1609=>"001001111",
  1610=>"000000000",
  1611=>"001001000",
  1612=>"110011000",
  1613=>"111111110",
  1614=>"000000000",
  1615=>"111111000",
  1616=>"000000000",
  1617=>"000100111",
  1618=>"000000000",
  1619=>"000110110",
  1620=>"111111111",
  1621=>"111111010",
  1622=>"101001111",
  1623=>"000000111",
  1624=>"000000000",
  1625=>"001000000",
  1626=>"000000000",
  1627=>"100000000",
  1628=>"111000000",
  1629=>"111111111",
  1630=>"111001001",
  1631=>"011111111",
  1632=>"001000000",
  1633=>"000000000",
  1634=>"000001001",
  1635=>"110110010",
  1636=>"111111000",
  1637=>"001001001",
  1638=>"110110111",
  1639=>"111111111",
  1640=>"000000000",
  1641=>"010000110",
  1642=>"000000000",
  1643=>"001001101",
  1644=>"000000000",
  1645=>"111111111",
  1646=>"111111111",
  1647=>"100100000",
  1648=>"111110110",
  1649=>"000100111",
  1650=>"111011000",
  1651=>"110101111",
  1652=>"111111011",
  1653=>"110111011",
  1654=>"000000000",
  1655=>"111111110",
  1656=>"000110011",
  1657=>"111111111",
  1658=>"101000101",
  1659=>"000111111",
  1660=>"111110000",
  1661=>"000001000",
  1662=>"111111111",
  1663=>"111111111",
  1664=>"111111111",
  1665=>"000000000",
  1666=>"010111111",
  1667=>"100011111",
  1668=>"000000000",
  1669=>"101000000",
  1670=>"001001000",
  1671=>"000000110",
  1672=>"000010011",
  1673=>"100000111",
  1674=>"000000000",
  1675=>"111111111",
  1676=>"001111111",
  1677=>"010000000",
  1678=>"000000000",
  1679=>"111011011",
  1680=>"001000000",
  1681=>"000000000",
  1682=>"000000100",
  1683=>"100000000",
  1684=>"001111001",
  1685=>"110100100",
  1686=>"000111111",
  1687=>"000000000",
  1688=>"000010011",
  1689=>"111111111",
  1690=>"000000111",
  1691=>"000000000",
  1692=>"011111111",
  1693=>"000000000",
  1694=>"111111011",
  1695=>"111111111",
  1696=>"000000000",
  1697=>"111110000",
  1698=>"111111110",
  1699=>"000000011",
  1700=>"001001001",
  1701=>"110110111",
  1702=>"110100000",
  1703=>"001000000",
  1704=>"111111000",
  1705=>"111111111",
  1706=>"000111111",
  1707=>"111111111",
  1708=>"111111111",
  1709=>"100100100",
  1710=>"111111011",
  1711=>"111111111",
  1712=>"111111110",
  1713=>"110111001",
  1714=>"111111000",
  1715=>"010000000",
  1716=>"111110111",
  1717=>"011011111",
  1718=>"000000000",
  1719=>"111101000",
  1720=>"000000000",
  1721=>"000000011",
  1722=>"111000000",
  1723=>"000000000",
  1724=>"111111111",
  1725=>"111111111",
  1726=>"111000111",
  1727=>"110000000",
  1728=>"010110010",
  1729=>"000000000",
  1730=>"000001001",
  1731=>"001000000",
  1732=>"000000000",
  1733=>"000001111",
  1734=>"001000000",
  1735=>"000000000",
  1736=>"110011001",
  1737=>"111111111",
  1738=>"111101001",
  1739=>"001111011",
  1740=>"111111111",
  1741=>"000000000",
  1742=>"010110111",
  1743=>"101100110",
  1744=>"000110011",
  1745=>"000010011",
  1746=>"101111110",
  1747=>"000000000",
  1748=>"000000000",
  1749=>"111111111",
  1750=>"000000000",
  1751=>"000000000",
  1752=>"000000000",
  1753=>"110100000",
  1754=>"000000000",
  1755=>"111011111",
  1756=>"000011011",
  1757=>"111001001",
  1758=>"111111111",
  1759=>"000010110",
  1760=>"000000000",
  1761=>"001001000",
  1762=>"000011001",
  1763=>"111111111",
  1764=>"110110111",
  1765=>"001000000",
  1766=>"000000000",
  1767=>"000000000",
  1768=>"000000111",
  1769=>"111111111",
  1770=>"111111011",
  1771=>"001001011",
  1772=>"110110111",
  1773=>"000000000",
  1774=>"111111111",
  1775=>"111001000",
  1776=>"111011011",
  1777=>"000000000",
  1778=>"111111111",
  1779=>"000000000",
  1780=>"011111111",
  1781=>"110110110",
  1782=>"111111111",
  1783=>"000000000",
  1784=>"111111110",
  1785=>"000010000",
  1786=>"111111111",
  1787=>"000000000",
  1788=>"100000000",
  1789=>"001001111",
  1790=>"101001000",
  1791=>"011001000",
  1792=>"000000000",
  1793=>"011010010",
  1794=>"000000111",
  1795=>"111110111",
  1796=>"000000000",
  1797=>"100110110",
  1798=>"101000000",
  1799=>"111111111",
  1800=>"000000000",
  1801=>"000000101",
  1802=>"111111000",
  1803=>"000000000",
  1804=>"000000000",
  1805=>"000000000",
  1806=>"000000000",
  1807=>"011011111",
  1808=>"000000000",
  1809=>"100110110",
  1810=>"000010000",
  1811=>"001001000",
  1812=>"111111111",
  1813=>"000111111",
  1814=>"110110110",
  1815=>"111011001",
  1816=>"110110100",
  1817=>"111000000",
  1818=>"000010000",
  1819=>"000000000",
  1820=>"111101100",
  1821=>"000000000",
  1822=>"000000001",
  1823=>"110110010",
  1824=>"110100101",
  1825=>"111111011",
  1826=>"000000000",
  1827=>"001001010",
  1828=>"000001000",
  1829=>"000000000",
  1830=>"111111000",
  1831=>"001000000",
  1832=>"110111111",
  1833=>"110111111",
  1834=>"000111111",
  1835=>"011011000",
  1836=>"111111110",
  1837=>"100100100",
  1838=>"000000000",
  1839=>"111111000",
  1840=>"011111011",
  1841=>"000000110",
  1842=>"111111000",
  1843=>"111101000",
  1844=>"000010000",
  1845=>"110110000",
  1846=>"001000000",
  1847=>"000110010",
  1848=>"000000011",
  1849=>"000000000",
  1850=>"111101111",
  1851=>"111111011",
  1852=>"101100000",
  1853=>"000000010",
  1854=>"111111111",
  1855=>"000000000",
  1856=>"111111001",
  1857=>"001000000",
  1858=>"001001011",
  1859=>"110110111",
  1860=>"001111101",
  1861=>"111111000",
  1862=>"010111111",
  1863=>"000000000",
  1864=>"111111111",
  1865=>"000000000",
  1866=>"000000010",
  1867=>"000000010",
  1868=>"000000000",
  1869=>"110111111",
  1870=>"110110010",
  1871=>"110010111",
  1872=>"001101111",
  1873=>"101111111",
  1874=>"011011001",
  1875=>"000000000",
  1876=>"001000000",
  1877=>"111001111",
  1878=>"111110110",
  1879=>"111001001",
  1880=>"000000000",
  1881=>"000000000",
  1882=>"111111000",
  1883=>"100101001",
  1884=>"111111011",
  1885=>"111001000",
  1886=>"000000000",
  1887=>"111111111",
  1888=>"111000000",
  1889=>"111111111",
  1890=>"010011011",
  1891=>"111111111",
  1892=>"010011011",
  1893=>"000000000",
  1894=>"111111111",
  1895=>"000000000",
  1896=>"001011011",
  1897=>"000111111",
  1898=>"111111111",
  1899=>"000000000",
  1900=>"111011011",
  1901=>"111111001",
  1902=>"000000000",
  1903=>"111000000",
  1904=>"110111111",
  1905=>"111011111",
  1906=>"000111011",
  1907=>"101100000",
  1908=>"101001111",
  1909=>"000000000",
  1910=>"111101000",
  1911=>"000000000",
  1912=>"111111111",
  1913=>"111111000",
  1914=>"000110100",
  1915=>"101111111",
  1916=>"010110111",
  1917=>"110110000",
  1918=>"000000000",
  1919=>"111101111",
  1920=>"110111111",
  1921=>"001010010",
  1922=>"000111111",
  1923=>"100111111",
  1924=>"100000111",
  1925=>"000000000",
  1926=>"001010010",
  1927=>"111111011",
  1928=>"000000000",
  1929=>"100101101",
  1930=>"111111011",
  1931=>"000000111",
  1932=>"111111111",
  1933=>"111111111",
  1934=>"110100100",
  1935=>"000000000",
  1936=>"111111111",
  1937=>"111111111",
  1938=>"000000000",
  1939=>"110001000",
  1940=>"000000010",
  1941=>"000110111",
  1942=>"111101111",
  1943=>"001001001",
  1944=>"111111001",
  1945=>"000010000",
  1946=>"000000000",
  1947=>"000000110",
  1948=>"101000111",
  1949=>"100000000",
  1950=>"111001011",
  1951=>"000000000",
  1952=>"111111111",
  1953=>"011011010",
  1954=>"110111111",
  1955=>"000111111",
  1956=>"000000111",
  1957=>"010111111",
  1958=>"000000000",
  1959=>"000000000",
  1960=>"111111111",
  1961=>"001111111",
  1962=>"111111111",
  1963=>"100100110",
  1964=>"000111101",
  1965=>"111111000",
  1966=>"111011011",
  1967=>"000000000",
  1968=>"000000000",
  1969=>"111111111",
  1970=>"001001000",
  1971=>"000000000",
  1972=>"110000000",
  1973=>"110000000",
  1974=>"011111110",
  1975=>"001000000",
  1976=>"001000000",
  1977=>"111101101",
  1978=>"000000000",
  1979=>"000001010",
  1980=>"000000000",
  1981=>"000000111",
  1982=>"100111111",
  1983=>"010011011",
  1984=>"111011011",
  1985=>"000000000",
  1986=>"111111010",
  1987=>"000000000",
  1988=>"001001111",
  1989=>"111111110",
  1990=>"001111111",
  1991=>"000010111",
  1992=>"000000000",
  1993=>"100000000",
  1994=>"101111010",
  1995=>"000000000",
  1996=>"000000000",
  1997=>"111111111",
  1998=>"110111010",
  1999=>"111111111",
  2000=>"100000000",
  2001=>"110000000",
  2002=>"111111111",
  2003=>"011011111",
  2004=>"111000001",
  2005=>"001001111",
  2006=>"111111100",
  2007=>"111111111",
  2008=>"111100000",
  2009=>"000111001",
  2010=>"000000000",
  2011=>"101101111",
  2012=>"000000000",
  2013=>"111110010",
  2014=>"001111000",
  2015=>"101100100",
  2016=>"110110000",
  2017=>"000000000",
  2018=>"100100101",
  2019=>"111100000",
  2020=>"000000111",
  2021=>"111101111",
  2022=>"111111011",
  2023=>"001111110",
  2024=>"100000000",
  2025=>"001001000",
  2026=>"011000001",
  2027=>"001000000",
  2028=>"111111011",
  2029=>"011011001",
  2030=>"000111010",
  2031=>"111111111",
  2032=>"111101100",
  2033=>"000000000",
  2034=>"010010000",
  2035=>"001000000",
  2036=>"111000000",
  2037=>"000110010",
  2038=>"000000100",
  2039=>"011111111",
  2040=>"111111111",
  2041=>"000110110",
  2042=>"000000000",
  2043=>"000000000",
  2044=>"111111111",
  2045=>"010010100",
  2046=>"111111111",
  2047=>"101000001",
  2048=>"001111111",
  2049=>"000110111",
  2050=>"111111111",
  2051=>"001111111",
  2052=>"001001101",
  2053=>"111111111",
  2054=>"000011111",
  2055=>"111111011",
  2056=>"111111111",
  2057=>"100111011",
  2058=>"111000000",
  2059=>"111011111",
  2060=>"000000100",
  2061=>"100000011",
  2062=>"000000001",
  2063=>"111010000",
  2064=>"001000000",
  2065=>"010111111",
  2066=>"000110111",
  2067=>"001001001",
  2068=>"000001111",
  2069=>"001000000",
  2070=>"000000111",
  2071=>"111111111",
  2072=>"111111111",
  2073=>"111110100",
  2074=>"000000000",
  2075=>"111111111",
  2076=>"011000001",
  2077=>"000111001",
  2078=>"110011000",
  2079=>"000000111",
  2080=>"110100011",
  2081=>"000111111",
  2082=>"110111000",
  2083=>"011011111",
  2084=>"001000000",
  2085=>"000000000",
  2086=>"110000000",
  2087=>"111000000",
  2088=>"111101000",
  2089=>"000000000",
  2090=>"111000000",
  2091=>"111111111",
  2092=>"111111111",
  2093=>"000000001",
  2094=>"000000111",
  2095=>"111111001",
  2096=>"000000001",
  2097=>"000000001",
  2098=>"110000000",
  2099=>"110100111",
  2100=>"000000000",
  2101=>"010011111",
  2102=>"000000000",
  2103=>"011000001",
  2104=>"010000011",
  2105=>"111111111",
  2106=>"000000000",
  2107=>"001000000",
  2108=>"011010111",
  2109=>"101000000",
  2110=>"000011000",
  2111=>"111001000",
  2112=>"001000111",
  2113=>"001001001",
  2114=>"011001000",
  2115=>"000111111",
  2116=>"011011111",
  2117=>"001011011",
  2118=>"000000110",
  2119=>"000000000",
  2120=>"001001001",
  2121=>"000000111",
  2122=>"111111111",
  2123=>"100100101",
  2124=>"111111111",
  2125=>"000100001",
  2126=>"000000111",
  2127=>"000000000",
  2128=>"001000000",
  2129=>"000000111",
  2130=>"000100100",
  2131=>"011111110",
  2132=>"100100000",
  2133=>"110000110",
  2134=>"110110111",
  2135=>"011011111",
  2136=>"111111110",
  2137=>"001000111",
  2138=>"011011011",
  2139=>"000000000",
  2140=>"000100000",
  2141=>"111010000",
  2142=>"001000000",
  2143=>"000000000",
  2144=>"011000000",
  2145=>"100000011",
  2146=>"000000000",
  2147=>"000000000",
  2148=>"111100000",
  2149=>"000000000",
  2150=>"111111011",
  2151=>"000000000",
  2152=>"110110000",
  2153=>"000000110",
  2154=>"000000111",
  2155=>"000011101",
  2156=>"001011001",
  2157=>"100110111",
  2158=>"011000111",
  2159=>"011000000",
  2160=>"000000001",
  2161=>"000000111",
  2162=>"001001000",
  2163=>"000111111",
  2164=>"110000000",
  2165=>"000000000",
  2166=>"111111000",
  2167=>"101001111",
  2168=>"000111111",
  2169=>"000000000",
  2170=>"000000000",
  2171=>"111111111",
  2172=>"000000000",
  2173=>"000101111",
  2174=>"100100100",
  2175=>"000000000",
  2176=>"000000000",
  2177=>"001111111",
  2178=>"000000001",
  2179=>"111111011",
  2180=>"110001000",
  2181=>"111101111",
  2182=>"011111100",
  2183=>"000000111",
  2184=>"000000000",
  2185=>"000000111",
  2186=>"000100111",
  2187=>"111111011",
  2188=>"110110111",
  2189=>"000110111",
  2190=>"000000111",
  2191=>"111011001",
  2192=>"001111111",
  2193=>"110110111",
  2194=>"000000000",
  2195=>"111011000",
  2196=>"110111001",
  2197=>"111111111",
  2198=>"001001111",
  2199=>"000000011",
  2200=>"000100111",
  2201=>"011111111",
  2202=>"111111111",
  2203=>"111111000",
  2204=>"001000110",
  2205=>"000000000",
  2206=>"111111111",
  2207=>"000000000",
  2208=>"000000000",
  2209=>"100000000",
  2210=>"000000000",
  2211=>"000001100",
  2212=>"000000111",
  2213=>"111111111",
  2214=>"111111110",
  2215=>"011011011",
  2216=>"111111010",
  2217=>"000000000",
  2218=>"000000111",
  2219=>"111111111",
  2220=>"000000011",
  2221=>"000011111",
  2222=>"000101111",
  2223=>"000000000",
  2224=>"111100111",
  2225=>"101001000",
  2226=>"111111010",
  2227=>"110111111",
  2228=>"001000001",
  2229=>"101111111",
  2230=>"000000001",
  2231=>"011110111",
  2232=>"000110111",
  2233=>"111111111",
  2234=>"000001000",
  2235=>"011010110",
  2236=>"111101111",
  2237=>"000000000",
  2238=>"111111111",
  2239=>"111111110",
  2240=>"111111111",
  2241=>"111101101",
  2242=>"100101101",
  2243=>"111111011",
  2244=>"010000000",
  2245=>"011111011",
  2246=>"100000000",
  2247=>"000000111",
  2248=>"000000010",
  2249=>"000000000",
  2250=>"111101100",
  2251=>"000000000",
  2252=>"000000000",
  2253=>"011011000",
  2254=>"111001000",
  2255=>"000000111",
  2256=>"111000000",
  2257=>"000011111",
  2258=>"111110000",
  2259=>"000000000",
  2260=>"000000011",
  2261=>"111111000",
  2262=>"001000000",
  2263=>"111001000",
  2264=>"111111111",
  2265=>"111111111",
  2266=>"000000011",
  2267=>"000000000",
  2268=>"111011001",
  2269=>"111111111",
  2270=>"110111010",
  2271=>"111000000",
  2272=>"000000000",
  2273=>"000000000",
  2274=>"111111010",
  2275=>"111011000",
  2276=>"111111111",
  2277=>"001000100",
  2278=>"000111111",
  2279=>"110111111",
  2280=>"100110110",
  2281=>"000110111",
  2282=>"111111000",
  2283=>"101010000",
  2284=>"001000000",
  2285=>"000000000",
  2286=>"111000000",
  2287=>"111111111",
  2288=>"111111111",
  2289=>"001001011",
  2290=>"111111011",
  2291=>"101000000",
  2292=>"011111111",
  2293=>"000000000",
  2294=>"011001000",
  2295=>"111100000",
  2296=>"111111111",
  2297=>"111111100",
  2298=>"000000000",
  2299=>"000000000",
  2300=>"001001000",
  2301=>"001000000",
  2302=>"010000001",
  2303=>"111111111",
  2304=>"111111111",
  2305=>"111111000",
  2306=>"111100111",
  2307=>"000111110",
  2308=>"100100100",
  2309=>"111001001",
  2310=>"111111111",
  2311=>"111111111",
  2312=>"001001101",
  2313=>"001000000",
  2314=>"111101111",
  2315=>"111111111",
  2316=>"111101101",
  2317=>"000011111",
  2318=>"111100100",
  2319=>"000000000",
  2320=>"000100100",
  2321=>"000001111",
  2322=>"001001001",
  2323=>"100000000",
  2324=>"000000000",
  2325=>"000000000",
  2326=>"000000000",
  2327=>"000000000",
  2328=>"111111000",
  2329=>"010010000",
  2330=>"110111111",
  2331=>"011000000",
  2332=>"100100111",
  2333=>"000000000",
  2334=>"111111111",
  2335=>"111111000",
  2336=>"000000110",
  2337=>"111100000",
  2338=>"011011111",
  2339=>"111000000",
  2340=>"000000000",
  2341=>"001000001",
  2342=>"000001001",
  2343=>"000000000",
  2344=>"000000111",
  2345=>"010111111",
  2346=>"000000000",
  2347=>"111111111",
  2348=>"000000000",
  2349=>"000000000",
  2350=>"110110111",
  2351=>"111111110",
  2352=>"011111111",
  2353=>"000000111",
  2354=>"001011110",
  2355=>"000000000",
  2356=>"111111111",
  2357=>"111111111",
  2358=>"000000000",
  2359=>"000000001",
  2360=>"000000000",
  2361=>"000000111",
  2362=>"001000000",
  2363=>"111111111",
  2364=>"011111000",
  2365=>"000001101",
  2366=>"000000000",
  2367=>"111111111",
  2368=>"000000011",
  2369=>"111101011",
  2370=>"000000111",
  2371=>"111100111",
  2372=>"000000110",
  2373=>"111011111",
  2374=>"000000001",
  2375=>"000000110",
  2376=>"111110000",
  2377=>"000000000",
  2378=>"000000000",
  2379=>"000000000",
  2380=>"100100000",
  2381=>"111111000",
  2382=>"111111111",
  2383=>"111101100",
  2384=>"000000110",
  2385=>"111111111",
  2386=>"011001000",
  2387=>"111110000",
  2388=>"000110111",
  2389=>"011111011",
  2390=>"111111001",
  2391=>"111000001",
  2392=>"111111111",
  2393=>"000110000",
  2394=>"111000111",
  2395=>"101111111",
  2396=>"111111001",
  2397=>"111111111",
  2398=>"000010111",
  2399=>"111111111",
  2400=>"111111000",
  2401=>"000000011",
  2402=>"111111001",
  2403=>"011011011",
  2404=>"100100000",
  2405=>"111111111",
  2406=>"111111111",
  2407=>"000000000",
  2408=>"001000000",
  2409=>"011011111",
  2410=>"000000001",
  2411=>"000000000",
  2412=>"001001001",
  2413=>"101000101",
  2414=>"000111111",
  2415=>"000000000",
  2416=>"100111000",
  2417=>"100110111",
  2418=>"011010111",
  2419=>"000000000",
  2420=>"000000000",
  2421=>"111101111",
  2422=>"000000000",
  2423=>"111000000",
  2424=>"000001111",
  2425=>"111000000",
  2426=>"110000100",
  2427=>"010001000",
  2428=>"000011011",
  2429=>"110111111",
  2430=>"110000000",
  2431=>"000101111",
  2432=>"111110110",
  2433=>"101000000",
  2434=>"000110110",
  2435=>"111111111",
  2436=>"111111111",
  2437=>"000000000",
  2438=>"000000001",
  2439=>"111111111",
  2440=>"001001000",
  2441=>"111000000",
  2442=>"111111111",
  2443=>"111111000",
  2444=>"111111111",
  2445=>"111111100",
  2446=>"100110110",
  2447=>"000000000",
  2448=>"111111000",
  2449=>"110110110",
  2450=>"011111111",
  2451=>"110111001",
  2452=>"101111001",
  2453=>"010010000",
  2454=>"001000000",
  2455=>"001011010",
  2456=>"111111111",
  2457=>"101111111",
  2458=>"101000000",
  2459=>"000000111",
  2460=>"101111100",
  2461=>"010111111",
  2462=>"000000000",
  2463=>"111010011",
  2464=>"111111000",
  2465=>"001111010",
  2466=>"110110111",
  2467=>"000001111",
  2468=>"000001001",
  2469=>"000111111",
  2470=>"101101111",
  2471=>"111001000",
  2472=>"111111000",
  2473=>"000000000",
  2474=>"111001000",
  2475=>"000000000",
  2476=>"000000000",
  2477=>"111001001",
  2478=>"110100111",
  2479=>"100111111",
  2480=>"000000011",
  2481=>"111111111",
  2482=>"000011001",
  2483=>"111111111",
  2484=>"000000000",
  2485=>"001000000",
  2486=>"111111111",
  2487=>"001001000",
  2488=>"111010111",
  2489=>"000000100",
  2490=>"000011011",
  2491=>"000000000",
  2492=>"000111111",
  2493=>"001111111",
  2494=>"000000000",
  2495=>"000000001",
  2496=>"111000000",
  2497=>"111111111",
  2498=>"111111111",
  2499=>"111011000",
  2500=>"111001101",
  2501=>"111001001",
  2502=>"001011111",
  2503=>"000000000",
  2504=>"111100110",
  2505=>"000000101",
  2506=>"000000011",
  2507=>"000000000",
  2508=>"111010000",
  2509=>"111111011",
  2510=>"110011011",
  2511=>"000010000",
  2512=>"100000000",
  2513=>"111011001",
  2514=>"111111111",
  2515=>"111111011",
  2516=>"100001011",
  2517=>"111111111",
  2518=>"101101111",
  2519=>"001000000",
  2520=>"000000001",
  2521=>"101111111",
  2522=>"011000000",
  2523=>"111000000",
  2524=>"111011010",
  2525=>"000111000",
  2526=>"111000000",
  2527=>"000111111",
  2528=>"000000000",
  2529=>"010001100",
  2530=>"111111111",
  2531=>"011001001",
  2532=>"110000000",
  2533=>"000000101",
  2534=>"001001011",
  2535=>"111111000",
  2536=>"001001000",
  2537=>"111111111",
  2538=>"011011000",
  2539=>"110110100",
  2540=>"111011111",
  2541=>"000000110",
  2542=>"111111111",
  2543=>"000000000",
  2544=>"000000000",
  2545=>"111111111",
  2546=>"100110111",
  2547=>"000000000",
  2548=>"000000010",
  2549=>"111111110",
  2550=>"111111000",
  2551=>"000000001",
  2552=>"000000001",
  2553=>"000000000",
  2554=>"100111111",
  2555=>"001001111",
  2556=>"000000100",
  2557=>"111000000",
  2558=>"111111111",
  2559=>"000000000",
  2560=>"000010010",
  2561=>"001000000",
  2562=>"111111111",
  2563=>"000101101",
  2564=>"101000100",
  2565=>"110111110",
  2566=>"111111100",
  2567=>"000111111",
  2568=>"110000000",
  2569=>"000000000",
  2570=>"000000000",
  2571=>"000000000",
  2572=>"100100100",
  2573=>"111111000",
  2574=>"111011011",
  2575=>"111111000",
  2576=>"110110101",
  2577=>"000111111",
  2578=>"011001000",
  2579=>"000000000",
  2580=>"111111000",
  2581=>"111111111",
  2582=>"000000000",
  2583=>"000000111",
  2584=>"000000111",
  2585=>"101000000",
  2586=>"000000111",
  2587=>"100000110",
  2588=>"111111000",
  2589=>"111011011",
  2590=>"111111011",
  2591=>"100001000",
  2592=>"000101111",
  2593=>"000000111",
  2594=>"111101000",
  2595=>"100101111",
  2596=>"111111111",
  2597=>"110111001",
  2598=>"110000000",
  2599=>"110010000",
  2600=>"111001000",
  2601=>"111000000",
  2602=>"110111111",
  2603=>"100110111",
  2604=>"000000111",
  2605=>"000111110",
  2606=>"000001001",
  2607=>"000000000",
  2608=>"000111100",
  2609=>"001000010",
  2610=>"000000111",
  2611=>"110100110",
  2612=>"000111111",
  2613=>"001001011",
  2614=>"111111101",
  2615=>"001000000",
  2616=>"100101111",
  2617=>"101001110",
  2618=>"100000000",
  2619=>"000110000",
  2620=>"000000111",
  2621=>"111110111",
  2622=>"000101100",
  2623=>"100100111",
  2624=>"100111111",
  2625=>"111111111",
  2626=>"100100000",
  2627=>"111000100",
  2628=>"001000110",
  2629=>"001111011",
  2630=>"111111111",
  2631=>"000000101",
  2632=>"001001111",
  2633=>"000100000",
  2634=>"000000111",
  2635=>"110101111",
  2636=>"000000000",
  2637=>"101001001",
  2638=>"111000000",
  2639=>"100100000",
  2640=>"111011000",
  2641=>"111111010",
  2642=>"000001101",
  2643=>"001011000",
  2644=>"111111010",
  2645=>"100111111",
  2646=>"111000101",
  2647=>"000000111",
  2648=>"111110100",
  2649=>"000101111",
  2650=>"010000000",
  2651=>"111000000",
  2652=>"111111110",
  2653=>"111111111",
  2654=>"010000110",
  2655=>"111111111",
  2656=>"110111000",
  2657=>"001011100",
  2658=>"111111000",
  2659=>"000000111",
  2660=>"000001000",
  2661=>"111111111",
  2662=>"011111001",
  2663=>"111111000",
  2664=>"111111000",
  2665=>"000000000",
  2666=>"111110100",
  2667=>"100111000",
  2668=>"111111101",
  2669=>"111110000",
  2670=>"000000011",
  2671=>"010000001",
  2672=>"111111111",
  2673=>"110110111",
  2674=>"000101111",
  2675=>"111000000",
  2676=>"111111111",
  2677=>"000000001",
  2678=>"000000000",
  2679=>"010000000",
  2680=>"000000111",
  2681=>"100100000",
  2682=>"000000101",
  2683=>"111111000",
  2684=>"011111111",
  2685=>"000101111",
  2686=>"000000100",
  2687=>"100110111",
  2688=>"000001001",
  2689=>"000000110",
  2690=>"111111111",
  2691=>"110111111",
  2692=>"000001000",
  2693=>"110000000",
  2694=>"000011111",
  2695=>"010111000",
  2696=>"111111101",
  2697=>"111111111",
  2698=>"111100000",
  2699=>"000000011",
  2700=>"111101100",
  2701=>"000000000",
  2702=>"111111100",
  2703=>"111110000",
  2704=>"011111111",
  2705=>"111111000",
  2706=>"110000000",
  2707=>"111111000",
  2708=>"011111000",
  2709=>"110000000",
  2710=>"000000000",
  2711=>"000000011",
  2712=>"100100110",
  2713=>"110110000",
  2714=>"111111111",
  2715=>"111111011",
  2716=>"101101111",
  2717=>"111111000",
  2718=>"000000110",
  2719=>"000000000",
  2720=>"000111111",
  2721=>"111111001",
  2722=>"110111111",
  2723=>"111110000",
  2724=>"001101111",
  2725=>"111111100",
  2726=>"000000010",
  2727=>"111011000",
  2728=>"111100111",
  2729=>"101111000",
  2730=>"110110111",
  2731=>"010000110",
  2732=>"000101101",
  2733=>"000000001",
  2734=>"111111111",
  2735=>"011011000",
  2736=>"001000000",
  2737=>"000000110",
  2738=>"110111000",
  2739=>"111111000",
  2740=>"111000000",
  2741=>"000000001",
  2742=>"111111111",
  2743=>"100110011",
  2744=>"001000000",
  2745=>"000111111",
  2746=>"000001111",
  2747=>"000001000",
  2748=>"100100111",
  2749=>"111000000",
  2750=>"100000001",
  2751=>"111111000",
  2752=>"111111100",
  2753=>"000100110",
  2754=>"000000001",
  2755=>"111111000",
  2756=>"000100000",
  2757=>"000111111",
  2758=>"111111000",
  2759=>"000011111",
  2760=>"000000111",
  2761=>"000101111",
  2762=>"000011111",
  2763=>"000000000",
  2764=>"100000000",
  2765=>"101100000",
  2766=>"000000000",
  2767=>"000100101",
  2768=>"111101000",
  2769=>"000000000",
  2770=>"000000000",
  2771=>"000000110",
  2772=>"000000001",
  2773=>"111011000",
  2774=>"001111111",
  2775=>"001111111",
  2776=>"000000000",
  2777=>"111011000",
  2778=>"001011111",
  2779=>"111111111",
  2780=>"111001001",
  2781=>"001001001",
  2782=>"010111000",
  2783=>"111100101",
  2784=>"111111000",
  2785=>"000100111",
  2786=>"111011011",
  2787=>"100000111",
  2788=>"110000000",
  2789=>"111010000",
  2790=>"111100111",
  2791=>"111100000",
  2792=>"110100100",
  2793=>"000001000",
  2794=>"100000000",
  2795=>"001000000",
  2796=>"000000010",
  2797=>"001000000",
  2798=>"000000000",
  2799=>"111011001",
  2800=>"100000000",
  2801=>"111111111",
  2802=>"000000000",
  2803=>"111011011",
  2804=>"000000000",
  2805=>"110111111",
  2806=>"111101000",
  2807=>"110100000",
  2808=>"000000000",
  2809=>"100000000",
  2810=>"111110110",
  2811=>"011111111",
  2812=>"111100111",
  2813=>"110100100",
  2814=>"111111100",
  2815=>"000000000",
  2816=>"000000000",
  2817=>"111111111",
  2818=>"000000111",
  2819=>"000000000",
  2820=>"001001111",
  2821=>"111000000",
  2822=>"111111111",
  2823=>"111000100",
  2824=>"101000000",
  2825=>"111000000",
  2826=>"000000000",
  2827=>"010111011",
  2828=>"111111111",
  2829=>"110000000",
  2830=>"111110000",
  2831=>"000101111",
  2832=>"000000000",
  2833=>"000001011",
  2834=>"111000000",
  2835=>"111111000",
  2836=>"111111111",
  2837=>"000100111",
  2838=>"100011001",
  2839=>"000100110",
  2840=>"111111011",
  2841=>"111111110",
  2842=>"001001011",
  2843=>"111001000",
  2844=>"001000000",
  2845=>"000000000",
  2846=>"111111111",
  2847=>"000000000",
  2848=>"100001000",
  2849=>"111001111",
  2850=>"111111111",
  2851=>"000000000",
  2852=>"110000000",
  2853=>"000000000",
  2854=>"111100000",
  2855=>"111010000",
  2856=>"001000000",
  2857=>"000000000",
  2858=>"101001000",
  2859=>"000000000",
  2860=>"111000000",
  2861=>"011011011",
  2862=>"000000000",
  2863=>"001000000",
  2864=>"111110000",
  2865=>"111111110",
  2866=>"111111111",
  2867=>"000000000",
  2868=>"000000000",
  2869=>"100000000",
  2870=>"110111110",
  2871=>"111100000",
  2872=>"000100000",
  2873=>"111110000",
  2874=>"111111110",
  2875=>"100000111",
  2876=>"001011111",
  2877=>"111111000",
  2878=>"110000000",
  2879=>"111111111",
  2880=>"111110111",
  2881=>"000000000",
  2882=>"111111010",
  2883=>"000000000",
  2884=>"111111101",
  2885=>"000000111",
  2886=>"001111101",
  2887=>"111111000",
  2888=>"111111101",
  2889=>"111000000",
  2890=>"111111111",
  2891=>"000111111",
  2892=>"000000000",
  2893=>"111110100",
  2894=>"100000100",
  2895=>"100111101",
  2896=>"111111100",
  2897=>"111111000",
  2898=>"111110010",
  2899=>"000111111",
  2900=>"000000000",
  2901=>"011111011",
  2902=>"111000000",
  2903=>"111111111",
  2904=>"000000000",
  2905=>"111111101",
  2906=>"111111001",
  2907=>"111000000",
  2908=>"000110111",
  2909=>"001011000",
  2910=>"111111000",
  2911=>"001111111",
  2912=>"101111100",
  2913=>"000000111",
  2914=>"111111110",
  2915=>"001000001",
  2916=>"000000011",
  2917=>"000000001",
  2918=>"010000101",
  2919=>"111111110",
  2920=>"000111111",
  2921=>"000000111",
  2922=>"111001111",
  2923=>"110110111",
  2924=>"010011000",
  2925=>"000000011",
  2926=>"000000111",
  2927=>"111011011",
  2928=>"011000000",
  2929=>"111100111",
  2930=>"000000000",
  2931=>"111111111",
  2932=>"111100111",
  2933=>"101100100",
  2934=>"000000011",
  2935=>"000100110",
  2936=>"101001111",
  2937=>"000000000",
  2938=>"000000000",
  2939=>"110100111",
  2940=>"111111111",
  2941=>"111110000",
  2942=>"000001111",
  2943=>"111000000",
  2944=>"011011111",
  2945=>"000110111",
  2946=>"000000100",
  2947=>"111111111",
  2948=>"100000000",
  2949=>"000000000",
  2950=>"111100000",
  2951=>"111111000",
  2952=>"111111101",
  2953=>"000111101",
  2954=>"111111010",
  2955=>"111111000",
  2956=>"000111111",
  2957=>"000011000",
  2958=>"111111001",
  2959=>"000011011",
  2960=>"001111110",
  2961=>"111000111",
  2962=>"000011011",
  2963=>"000111111",
  2964=>"000101000",
  2965=>"000000000",
  2966=>"001000000",
  2967=>"000000001",
  2968=>"110000111",
  2969=>"000000101",
  2970=>"111101000",
  2971=>"111111111",
  2972=>"000100111",
  2973=>"111111111",
  2974=>"000000000",
  2975=>"111000111",
  2976=>"111000000",
  2977=>"100000011",
  2978=>"111111111",
  2979=>"011000000",
  2980=>"000000100",
  2981=>"111101000",
  2982=>"111111000",
  2983=>"100000000",
  2984=>"000111111",
  2985=>"111100111",
  2986=>"000100101",
  2987=>"011011000",
  2988=>"111001001",
  2989=>"111110110",
  2990=>"111100101",
  2991=>"111111000",
  2992=>"111111111",
  2993=>"111111111",
  2994=>"111111111",
  2995=>"000000000",
  2996=>"111111000",
  2997=>"011000100",
  2998=>"111111111",
  2999=>"000111010",
  3000=>"111000010",
  3001=>"110111001",
  3002=>"001100000",
  3003=>"100110111",
  3004=>"110111000",
  3005=>"111111111",
  3006=>"111001011",
  3007=>"110111001",
  3008=>"000000011",
  3009=>"001001001",
  3010=>"000111111",
  3011=>"101001001",
  3012=>"100000110",
  3013=>"111001111",
  3014=>"110110110",
  3015=>"111100011",
  3016=>"100100100",
  3017=>"111111111",
  3018=>"111000110",
  3019=>"111111000",
  3020=>"000000000",
  3021=>"100111111",
  3022=>"000000000",
  3023=>"000001001",
  3024=>"111111111",
  3025=>"111110110",
  3026=>"000000111",
  3027=>"000010100",
  3028=>"000000111",
  3029=>"111001100",
  3030=>"000000110",
  3031=>"000110001",
  3032=>"000000011",
  3033=>"110111111",
  3034=>"011011000",
  3035=>"011000000",
  3036=>"111110000",
  3037=>"111111100",
  3038=>"110000000",
  3039=>"111000000",
  3040=>"111111111",
  3041=>"110101111",
  3042=>"111101000",
  3043=>"111101000",
  3044=>"110111111",
  3045=>"000000111",
  3046=>"111111000",
  3047=>"101111111",
  3048=>"000000111",
  3049=>"100111111",
  3050=>"111011000",
  3051=>"000000000",
  3052=>"000000111",
  3053=>"000000000",
  3054=>"011000111",
  3055=>"111011111",
  3056=>"111111111",
  3057=>"000100100",
  3058=>"111000101",
  3059=>"000000111",
  3060=>"111000000",
  3061=>"101111111",
  3062=>"111111111",
  3063=>"001001111",
  3064=>"011000111",
  3065=>"111111101",
  3066=>"000111111",
  3067=>"000000111",
  3068=>"111111110",
  3069=>"000000111",
  3070=>"001011111",
  3071=>"111101111",
  3072=>"100111111",
  3073=>"111101001",
  3074=>"111001000",
  3075=>"000111111",
  3076=>"000000001",
  3077=>"111011001",
  3078=>"111101001",
  3079=>"110110000",
  3080=>"110111000",
  3081=>"000000000",
  3082=>"011011111",
  3083=>"111011001",
  3084=>"111001001",
  3085=>"000101111",
  3086=>"100111100",
  3087=>"111111111",
  3088=>"000000000",
  3089=>"010001111",
  3090=>"000000110",
  3091=>"110000000",
  3092=>"001001111",
  3093=>"111011011",
  3094=>"000000010",
  3095=>"001001001",
  3096=>"000000000",
  3097=>"001011111",
  3098=>"011011111",
  3099=>"111111110",
  3100=>"000000100",
  3101=>"000000000",
  3102=>"001111111",
  3103=>"000000000",
  3104=>"000000000",
  3105=>"110111111",
  3106=>"100100110",
  3107=>"000000000",
  3108=>"000000111",
  3109=>"000000000",
  3110=>"000000000",
  3111=>"110010000",
  3112=>"000000000",
  3113=>"001101111",
  3114=>"000001011",
  3115=>"111011000",
  3116=>"000000001",
  3117=>"001011011",
  3118=>"010111111",
  3119=>"111111011",
  3120=>"000000000",
  3121=>"000000001",
  3122=>"000000000",
  3123=>"000000000",
  3124=>"000000000",
  3125=>"100110110",
  3126=>"101101101",
  3127=>"000000100",
  3128=>"001000111",
  3129=>"000001001",
  3130=>"111111000",
  3131=>"010010111",
  3132=>"000000000",
  3133=>"110110100",
  3134=>"000001111",
  3135=>"101001001",
  3136=>"000000000",
  3137=>"000000000",
  3138=>"001001101",
  3139=>"001001111",
  3140=>"111111110",
  3141=>"100100000",
  3142=>"101000000",
  3143=>"111111111",
  3144=>"111111111",
  3145=>"000001001",
  3146=>"111111110",
  3147=>"111111000",
  3148=>"110110110",
  3149=>"000101101",
  3150=>"000001000",
  3151=>"111001001",
  3152=>"011011000",
  3153=>"001111111",
  3154=>"111001011",
  3155=>"011001001",
  3156=>"000001001",
  3157=>"000001001",
  3158=>"000101111",
  3159=>"110110110",
  3160=>"011111111",
  3161=>"111111011",
  3162=>"011110110",
  3163=>"111100000",
  3164=>"001101111",
  3165=>"001011000",
  3166=>"000000000",
  3167=>"000000111",
  3168=>"001011011",
  3169=>"010010101",
  3170=>"110111110",
  3171=>"111010010",
  3172=>"000000000",
  3173=>"111111111",
  3174=>"111110000",
  3175=>"000000000",
  3176=>"000011111",
  3177=>"000000011",
  3178=>"111111111",
  3179=>"000100000",
  3180=>"111110010",
  3181=>"000000111",
  3182=>"100110111",
  3183=>"000110100",
  3184=>"000000001",
  3185=>"111110110",
  3186=>"111111111",
  3187=>"111111111",
  3188=>"000000000",
  3189=>"001001101",
  3190=>"000100101",
  3191=>"001001001",
  3192=>"110111110",
  3193=>"101001001",
  3194=>"101101111",
  3195=>"000010000",
  3196=>"101101101",
  3197=>"110110000",
  3198=>"101000001",
  3199=>"010110010",
  3200=>"001001011",
  3201=>"111111000",
  3202=>"111000000",
  3203=>"100100100",
  3204=>"111001001",
  3205=>"111101101",
  3206=>"000000111",
  3207=>"000001101",
  3208=>"000000001",
  3209=>"010110000",
  3210=>"000000000",
  3211=>"111111001",
  3212=>"000000111",
  3213=>"111110110",
  3214=>"100110101",
  3215=>"110100100",
  3216=>"001111110",
  3217=>"010111110",
  3218=>"001001001",
  3219=>"100100000",
  3220=>"111111001",
  3221=>"110111111",
  3222=>"111111111",
  3223=>"010110111",
  3224=>"110110111",
  3225=>"111111111",
  3226=>"000010000",
  3227=>"100101001",
  3228=>"000000010",
  3229=>"100101111",
  3230=>"101001000",
  3231=>"111111110",
  3232=>"000000000",
  3233=>"000100000",
  3234=>"101101101",
  3235=>"010000000",
  3236=>"111101001",
  3237=>"110111111",
  3238=>"011011000",
  3239=>"111111111",
  3240=>"000110000",
  3241=>"001001001",
  3242=>"101000000",
  3243=>"000000001",
  3244=>"111111110",
  3245=>"101011001",
  3246=>"111111111",
  3247=>"001001001",
  3248=>"000000000",
  3249=>"111111111",
  3250=>"110111111",
  3251=>"010000000",
  3252=>"000000000",
  3253=>"111001001",
  3254=>"111011000",
  3255=>"111001001",
  3256=>"011001101",
  3257=>"001101111",
  3258=>"100100100",
  3259=>"101101001",
  3260=>"000000000",
  3261=>"001111011",
  3262=>"111000000",
  3263=>"010110111",
  3264=>"000100110",
  3265=>"001001101",
  3266=>"111111111",
  3267=>"000000001",
  3268=>"001000000",
  3269=>"111111111",
  3270=>"000000000",
  3271=>"000110001",
  3272=>"000000010",
  3273=>"001010111",
  3274=>"000000000",
  3275=>"000000011",
  3276=>"110110111",
  3277=>"000010000",
  3278=>"101111111",
  3279=>"000000000",
  3280=>"000111011",
  3281=>"111011000",
  3282=>"110110010",
  3283=>"100000000",
  3284=>"011110010",
  3285=>"001000000",
  3286=>"000010000",
  3287=>"111111000",
  3288=>"000000111",
  3289=>"111111111",
  3290=>"000000001",
  3291=>"000000111",
  3292=>"011000000",
  3293=>"000000000",
  3294=>"000000000",
  3295=>"000000100",
  3296=>"000001111",
  3297=>"000001000",
  3298=>"111111111",
  3299=>"111110000",
  3300=>"000000000",
  3301=>"100111111",
  3302=>"110110110",
  3303=>"011011001",
  3304=>"010010110",
  3305=>"110011000",
  3306=>"000100111",
  3307=>"111100000",
  3308=>"111000010",
  3309=>"001001000",
  3310=>"111101101",
  3311=>"001001001",
  3312=>"001011000",
  3313=>"001101100",
  3314=>"001000000",
  3315=>"100111111",
  3316=>"000000000",
  3317=>"000000100",
  3318=>"000101111",
  3319=>"000010110",
  3320=>"000000000",
  3321=>"000000100",
  3322=>"000000000",
  3323=>"111001111",
  3324=>"111110100",
  3325=>"001001111",
  3326=>"001001100",
  3327=>"111111111",
  3328=>"101100000",
  3329=>"000000000",
  3330=>"111111111",
  3331=>"101001101",
  3332=>"010000000",
  3333=>"000001001",
  3334=>"110110000",
  3335=>"001111000",
  3336=>"001001000",
  3337=>"001001001",
  3338=>"111000000",
  3339=>"111111111",
  3340=>"000000000",
  3341=>"010111110",
  3342=>"000000000",
  3343=>"111111001",
  3344=>"011000001",
  3345=>"000000000",
  3346=>"000010010",
  3347=>"000000000",
  3348=>"001000001",
  3349=>"101000111",
  3350=>"001000000",
  3351=>"000000000",
  3352=>"000001001",
  3353=>"100100111",
  3354=>"000110110",
  3355=>"000000110",
  3356=>"111110110",
  3357=>"000000111",
  3358=>"101000000",
  3359=>"111001000",
  3360=>"000000011",
  3361=>"110110110",
  3362=>"011110000",
  3363=>"101111111",
  3364=>"001101111",
  3365=>"110100100",
  3366=>"000001000",
  3367=>"001101100",
  3368=>"000000110",
  3369=>"110110111",
  3370=>"000000000",
  3371=>"000000000",
  3372=>"000000111",
  3373=>"110110110",
  3374=>"000000001",
  3375=>"111111010",
  3376=>"000001001",
  3377=>"000000111",
  3378=>"001101000",
  3379=>"001001000",
  3380=>"010111000",
  3381=>"000000000",
  3382=>"001110110",
  3383=>"101100111",
  3384=>"111011011",
  3385=>"101101111",
  3386=>"111111000",
  3387=>"000010001",
  3388=>"100110010",
  3389=>"111111001",
  3390=>"000000000",
  3391=>"111111000",
  3392=>"100100000",
  3393=>"011110111",
  3394=>"110110111",
  3395=>"000000000",
  3396=>"110010100",
  3397=>"111111111",
  3398=>"000001111",
  3399=>"000000001",
  3400=>"000001100",
  3401=>"000000111",
  3402=>"111101101",
  3403=>"110111111",
  3404=>"001101001",
  3405=>"110111111",
  3406=>"100100111",
  3407=>"110110110",
  3408=>"000000000",
  3409=>"100000001",
  3410=>"000001100",
  3411=>"010110111",
  3412=>"001000000",
  3413=>"001011011",
  3414=>"000000000",
  3415=>"000000000",
  3416=>"000000101",
  3417=>"011011111",
  3418=>"000000000",
  3419=>"000000001",
  3420=>"111111001",
  3421=>"111111111",
  3422=>"111100000",
  3423=>"111111000",
  3424=>"000000000",
  3425=>"101001111",
  3426=>"100100100",
  3427=>"000001001",
  3428=>"000000100",
  3429=>"000110000",
  3430=>"111111011",
  3431=>"111111111",
  3432=>"000000000",
  3433=>"001001001",
  3434=>"010010000",
  3435=>"101001001",
  3436=>"000000100",
  3437=>"110110110",
  3438=>"111000001",
  3439=>"001001000",
  3440=>"000000010",
  3441=>"000000001",
  3442=>"111111110",
  3443=>"111011001",
  3444=>"000111111",
  3445=>"000000000",
  3446=>"111111111",
  3447=>"010111111",
  3448=>"000000011",
  3449=>"111000001",
  3450=>"000000110",
  3451=>"001000000",
  3452=>"001000000",
  3453=>"011011001",
  3454=>"010010000",
  3455=>"111111001",
  3456=>"001001111",
  3457=>"000110111",
  3458=>"011001000",
  3459=>"001000000",
  3460=>"000000000",
  3461=>"010111010",
  3462=>"111101101",
  3463=>"000001000",
  3464=>"111110110",
  3465=>"111111111",
  3466=>"100100111",
  3467=>"010010100",
  3468=>"111111111",
  3469=>"100100100",
  3470=>"111111111",
  3471=>"110111111",
  3472=>"000010010",
  3473=>"001000000",
  3474=>"010110110",
  3475=>"011011000",
  3476=>"001111000",
  3477=>"000010010",
  3478=>"000001000",
  3479=>"001101001",
  3480=>"111111111",
  3481=>"111111110",
  3482=>"001011111",
  3483=>"000001011",
  3484=>"100100111",
  3485=>"000010010",
  3486=>"000000011",
  3487=>"000010101",
  3488=>"100000000",
  3489=>"011111011",
  3490=>"100000010",
  3491=>"111111111",
  3492=>"101111111",
  3493=>"111111110",
  3494=>"000000000",
  3495=>"010010000",
  3496=>"000000001",
  3497=>"001111111",
  3498=>"111000001",
  3499=>"000001111",
  3500=>"001001001",
  3501=>"010000111",
  3502=>"111101001",
  3503=>"000000000",
  3504=>"111111110",
  3505=>"001001001",
  3506=>"011000000",
  3507=>"000000001",
  3508=>"110111111",
  3509=>"101000001",
  3510=>"000000010",
  3511=>"001000001",
  3512=>"001001000",
  3513=>"010111001",
  3514=>"111100101",
  3515=>"000110111",
  3516=>"001111001",
  3517=>"000000100",
  3518=>"111101000",
  3519=>"101001001",
  3520=>"011000000",
  3521=>"111111000",
  3522=>"111111111",
  3523=>"111001000",
  3524=>"001011000",
  3525=>"001100100",
  3526=>"000110000",
  3527=>"111001001",
  3528=>"101100000",
  3529=>"110110111",
  3530=>"001000000",
  3531=>"111101000",
  3532=>"001001001",
  3533=>"000000111",
  3534=>"000000001",
  3535=>"011111111",
  3536=>"000000011",
  3537=>"100101110",
  3538=>"110010000",
  3539=>"111001110",
  3540=>"110111101",
  3541=>"000000000",
  3542=>"000001001",
  3543=>"100100111",
  3544=>"000111111",
  3545=>"000000000",
  3546=>"000000111",
  3547=>"111111000",
  3548=>"010110110",
  3549=>"001001111",
  3550=>"000000010",
  3551=>"011111110",
  3552=>"001001111",
  3553=>"000000000",
  3554=>"000010111",
  3555=>"001010000",
  3556=>"111111111",
  3557=>"111110110",
  3558=>"111111111",
  3559=>"111101001",
  3560=>"001001001",
  3561=>"000000000",
  3562=>"011011000",
  3563=>"010110101",
  3564=>"111111111",
  3565=>"000000000",
  3566=>"110110010",
  3567=>"000000001",
  3568=>"000110111",
  3569=>"111110000",
  3570=>"000000000",
  3571=>"000110111",
  3572=>"101001111",
  3573=>"000010010",
  3574=>"111111111",
  3575=>"100100001",
  3576=>"000000011",
  3577=>"100000110",
  3578=>"001001001",
  3579=>"001001001",
  3580=>"001001000",
  3581=>"111011011",
  3582=>"001111111",
  3583=>"111111111",
  3584=>"111111111",
  3585=>"000000110",
  3586=>"000000000",
  3587=>"000000000",
  3588=>"001000100",
  3589=>"100100100",
  3590=>"111101101",
  3591=>"001001000",
  3592=>"111111000",
  3593=>"000000000",
  3594=>"111111111",
  3595=>"111000000",
  3596=>"001001011",
  3597=>"000000111",
  3598=>"000001000",
  3599=>"100000001",
  3600=>"000110111",
  3601=>"111000000",
  3602=>"111111111",
  3603=>"110000111",
  3604=>"110111111",
  3605=>"000000000",
  3606=>"100111111",
  3607=>"001011011",
  3608=>"000001000",
  3609=>"100111111",
  3610=>"011111111",
  3611=>"000011111",
  3612=>"111111111",
  3613=>"000000000",
  3614=>"111011001",
  3615=>"110111000",
  3616=>"001100000",
  3617=>"111111111",
  3618=>"111111111",
  3619=>"101001000",
  3620=>"111111011",
  3621=>"000000100",
  3622=>"000011111",
  3623=>"000000111",
  3624=>"111111000",
  3625=>"000110110",
  3626=>"000100111",
  3627=>"000011111",
  3628=>"111111111",
  3629=>"000010011",
  3630=>"011110111",
  3631=>"001001001",
  3632=>"011110100",
  3633=>"111101111",
  3634=>"000000111",
  3635=>"010000000",
  3636=>"010010011",
  3637=>"000000000",
  3638=>"000011110",
  3639=>"000110000",
  3640=>"100000000",
  3641=>"000000000",
  3642=>"110000000",
  3643=>"000110000",
  3644=>"111100111",
  3645=>"011001111",
  3646=>"111111111",
  3647=>"000000000",
  3648=>"111110000",
  3649=>"000000000",
  3650=>"111111111",
  3651=>"110110111",
  3652=>"011111111",
  3653=>"000000100",
  3654=>"000000000",
  3655=>"111111111",
  3656=>"001101111",
  3657=>"100000000",
  3658=>"000001001",
  3659=>"111111111",
  3660=>"111110000",
  3661=>"000111111",
  3662=>"000000000",
  3663=>"111111111",
  3664=>"000000010",
  3665=>"000001011",
  3666=>"011000000",
  3667=>"011001001",
  3668=>"000000011",
  3669=>"110000000",
  3670=>"100000000",
  3671=>"001001000",
  3672=>"111110111",
  3673=>"000000000",
  3674=>"000000110",
  3675=>"111111001",
  3676=>"001000000",
  3677=>"000000000",
  3678=>"100000000",
  3679=>"010100100",
  3680=>"001000000",
  3681=>"000001001",
  3682=>"101101100",
  3683=>"111111111",
  3684=>"001001111",
  3685=>"000100101",
  3686=>"110110110",
  3687=>"001111110",
  3688=>"000111111",
  3689=>"000000111",
  3690=>"111111000",
  3691=>"111110110",
  3692=>"111111111",
  3693=>"111111111",
  3694=>"111111111",
  3695=>"111111111",
  3696=>"111111110",
  3697=>"000000100",
  3698=>"000011011",
  3699=>"000000000",
  3700=>"101101111",
  3701=>"111011010",
  3702=>"000000000",
  3703=>"111111111",
  3704=>"000110100",
  3705=>"111111111",
  3706=>"001011111",
  3707=>"000011001",
  3708=>"011011011",
  3709=>"000111110",
  3710=>"000000011",
  3711=>"000110110",
  3712=>"111100100",
  3713=>"110010010",
  3714=>"111111000",
  3715=>"000100111",
  3716=>"111111111",
  3717=>"000000000",
  3718=>"110010000",
  3719=>"001001001",
  3720=>"101111011",
  3721=>"001111111",
  3722=>"111101111",
  3723=>"101101110",
  3724=>"111111110",
  3725=>"110111111",
  3726=>"010001011",
  3727=>"111111111",
  3728=>"001111111",
  3729=>"000010000",
  3730=>"111111111",
  3731=>"111100101",
  3732=>"110110100",
  3733=>"000000110",
  3734=>"000000000",
  3735=>"000000000",
  3736=>"000010111",
  3737=>"111111111",
  3738=>"111111111",
  3739=>"111110000",
  3740=>"000000000",
  3741=>"100110111",
  3742=>"111111110",
  3743=>"111111000",
  3744=>"111110110",
  3745=>"111111011",
  3746=>"111111111",
  3747=>"001000110",
  3748=>"000110110",
  3749=>"000000111",
  3750=>"110110000",
  3751=>"000001001",
  3752=>"000000000",
  3753=>"111111100",
  3754=>"101100101",
  3755=>"000010010",
  3756=>"101111111",
  3757=>"110110100",
  3758=>"001101111",
  3759=>"111111110",
  3760=>"111111111",
  3761=>"111100100",
  3762=>"000011011",
  3763=>"101000000",
  3764=>"011010111",
  3765=>"000111111",
  3766=>"111101000",
  3767=>"000001000",
  3768=>"000000100",
  3769=>"001001001",
  3770=>"000000000",
  3771=>"100110111",
  3772=>"000000000",
  3773=>"111011001",
  3774=>"000000000",
  3775=>"110110111",
  3776=>"000001001",
  3777=>"011111100",
  3778=>"111111111",
  3779=>"100100000",
  3780=>"100000000",
  3781=>"000000000",
  3782=>"101000111",
  3783=>"111110110",
  3784=>"101111111",
  3785=>"111000000",
  3786=>"000000000",
  3787=>"110100000",
  3788=>"000100111",
  3789=>"111110000",
  3790=>"000000000",
  3791=>"110000111",
  3792=>"111111100",
  3793=>"000100101",
  3794=>"111111111",
  3795=>"000000000",
  3796=>"111111000",
  3797=>"000000101",
  3798=>"000000000",
  3799=>"000001000",
  3800=>"111111111",
  3801=>"000011110",
  3802=>"000000000",
  3803=>"000001011",
  3804=>"111111110",
  3805=>"000111000",
  3806=>"000000000",
  3807=>"000000000",
  3808=>"100000001",
  3809=>"000000000",
  3810=>"001000000",
  3811=>"100000000",
  3812=>"001001111",
  3813=>"010011000",
  3814=>"001000000",
  3815=>"000000011",
  3816=>"100111111",
  3817=>"111110000",
  3818=>"111111111",
  3819=>"111111111",
  3820=>"000000000",
  3821=>"000000000",
  3822=>"111110111",
  3823=>"000000000",
  3824=>"111111011",
  3825=>"100000111",
  3826=>"111100101",
  3827=>"000000000",
  3828=>"111000001",
  3829=>"111000000",
  3830=>"011011011",
  3831=>"110111111",
  3832=>"111111111",
  3833=>"000000000",
  3834=>"000111111",
  3835=>"000000000",
  3836=>"110111110",
  3837=>"000000111",
  3838=>"000111111",
  3839=>"000000000",
  3840=>"000000000",
  3841=>"001011001",
  3842=>"111111111",
  3843=>"000010010",
  3844=>"111101101",
  3845=>"010000000",
  3846=>"110100000",
  3847=>"111000111",
  3848=>"010111111",
  3849=>"001000000",
  3850=>"000110100",
  3851=>"001011111",
  3852=>"110110000",
  3853=>"000011011",
  3854=>"111111111",
  3855=>"000111111",
  3856=>"000111111",
  3857=>"001001001",
  3858=>"000000000",
  3859=>"000001101",
  3860=>"111001101",
  3861=>"111101111",
  3862=>"011111111",
  3863=>"011111111",
  3864=>"001001000",
  3865=>"111111111",
  3866=>"000100100",
  3867=>"000000000",
  3868=>"000000100",
  3869=>"000000100",
  3870=>"100100101",
  3871=>"000000000",
  3872=>"000101001",
  3873=>"111111111",
  3874=>"100100110",
  3875=>"000111110",
  3876=>"100100001",
  3877=>"011001000",
  3878=>"111100100",
  3879=>"111111111",
  3880=>"111111111",
  3881=>"000000000",
  3882=>"011111111",
  3883=>"000111000",
  3884=>"010011011",
  3885=>"000100100",
  3886=>"011011000",
  3887=>"000000000",
  3888=>"110111111",
  3889=>"000000110",
  3890=>"001000000",
  3891=>"110000000",
  3892=>"011111111",
  3893=>"100110100",
  3894=>"010110110",
  3895=>"100000000",
  3896=>"000000111",
  3897=>"110010000",
  3898=>"111111111",
  3899=>"000000111",
  3900=>"111000100",
  3901=>"000010110",
  3902=>"111101111",
  3903=>"111000001",
  3904=>"111111111",
  3905=>"010110011",
  3906=>"001001111",
  3907=>"000000110",
  3908=>"011111001",
  3909=>"000011011",
  3910=>"000000100",
  3911=>"001001011",
  3912=>"000000111",
  3913=>"111001000",
  3914=>"110000000",
  3915=>"000000000",
  3916=>"011011000",
  3917=>"111111101",
  3918=>"111001000",
  3919=>"011001111",
  3920=>"110111101",
  3921=>"000100110",
  3922=>"111111001",
  3923=>"000000000",
  3924=>"000000000",
  3925=>"111101111",
  3926=>"111111111",
  3927=>"011001000",
  3928=>"111011000",
  3929=>"000000000",
  3930=>"001001111",
  3931=>"000000000",
  3932=>"000010110",
  3933=>"111000100",
  3934=>"110111100",
  3935=>"110110000",
  3936=>"000000000",
  3937=>"000011011",
  3938=>"001000010",
  3939=>"001001011",
  3940=>"001001111",
  3941=>"000001011",
  3942=>"011001000",
  3943=>"011111011",
  3944=>"001001001",
  3945=>"111111111",
  3946=>"101100111",
  3947=>"000000000",
  3948=>"110110100",
  3949=>"000001111",
  3950=>"001000000",
  3951=>"101101111",
  3952=>"000000100",
  3953=>"111111111",
  3954=>"011111111",
  3955=>"100100100",
  3956=>"111100111",
  3957=>"111111011",
  3958=>"000001001",
  3959=>"000000001",
  3960=>"111101101",
  3961=>"000000111",
  3962=>"111111100",
  3963=>"011000111",
  3964=>"000100111",
  3965=>"111111000",
  3966=>"010000000",
  3967=>"111111111",
  3968=>"001001000",
  3969=>"000000000",
  3970=>"000000111",
  3971=>"000000000",
  3972=>"000000000",
  3973=>"000000000",
  3974=>"110111111",
  3975=>"000101111",
  3976=>"000000000",
  3977=>"110111111",
  3978=>"111110000",
  3979=>"000000000",
  3980=>"011011111",
  3981=>"011101111",
  3982=>"000011000",
  3983=>"000000111",
  3984=>"111000000",
  3985=>"001001001",
  3986=>"111111111",
  3987=>"111001001",
  3988=>"110111001",
  3989=>"000000000",
  3990=>"101101101",
  3991=>"000001111",
  3992=>"000100111",
  3993=>"000110111",
  3994=>"000000000",
  3995=>"011111111",
  3996=>"000000010",
  3997=>"101100101",
  3998=>"000000000",
  3999=>"010100111",
  4000=>"000001000",
  4001=>"011001001",
  4002=>"010111011",
  4003=>"000111111",
  4004=>"010011011",
  4005=>"011111000",
  4006=>"110111001",
  4007=>"000011001",
  4008=>"000000000",
  4009=>"000000000",
  4010=>"011001111",
  4011=>"010110011",
  4012=>"111010000",
  4013=>"110100111",
  4014=>"101111111",
  4015=>"111110111",
  4016=>"111111111",
  4017=>"000000000",
  4018=>"111111111",
  4019=>"001000000",
  4020=>"111111111",
  4021=>"000011111",
  4022=>"111111111",
  4023=>"111111111",
  4024=>"111111111",
  4025=>"000000100",
  4026=>"100100100",
  4027=>"000000000",
  4028=>"000000000",
  4029=>"000000000",
  4030=>"011111110",
  4031=>"001011001",
  4032=>"000000001",
  4033=>"101111001",
  4034=>"000000000",
  4035=>"011001000",
  4036=>"011011000",
  4037=>"111101111",
  4038=>"111110000",
  4039=>"000000111",
  4040=>"000000001",
  4041=>"000001111",
  4042=>"000000000",
  4043=>"000110110",
  4044=>"000000000",
  4045=>"000000000",
  4046=>"010111000",
  4047=>"111111001",
  4048=>"111111111",
  4049=>"110100000",
  4050=>"100111110",
  4051=>"111111111",
  4052=>"001001011",
  4053=>"000000000",
  4054=>"111111011",
  4055=>"101000101",
  4056=>"100100111",
  4057=>"000010011",
  4058=>"001000101",
  4059=>"111110010",
  4060=>"111000111",
  4061=>"110111111",
  4062=>"000000000",
  4063=>"101001101",
  4064=>"000000101",
  4065=>"001001000",
  4066=>"000000110",
  4067=>"110100000",
  4068=>"001001101",
  4069=>"000001111",
  4070=>"001111111",
  4071=>"000000011",
  4072=>"001011011",
  4073=>"111111111",
  4074=>"011000100",
  4075=>"111100111",
  4076=>"000000000",
  4077=>"000000000",
  4078=>"011111111",
  4079=>"110111000",
  4080=>"111111111",
  4081=>"001011001",
  4082=>"111111111",
  4083=>"000111111",
  4084=>"110111001",
  4085=>"000000010",
  4086=>"111011011",
  4087=>"001000100",
  4088=>"111000000",
  4089=>"110101001",
  4090=>"111001111",
  4091=>"000000000",
  4092=>"111111011",
  4093=>"000000001",
  4094=>"000000000",
  4095=>"111111111",
  4096=>"110110000",
  4097=>"111001111",
  4098=>"000000101",
  4099=>"000000111",
  4100=>"111111011",
  4101=>"110000010",
  4102=>"000111111",
  4103=>"111000111",
  4104=>"111000001",
  4105=>"010111111",
  4106=>"000000101",
  4107=>"000000000",
  4108=>"100110110",
  4109=>"111111111",
  4110=>"111111111",
  4111=>"100111111",
  4112=>"001000001",
  4113=>"111100100",
  4114=>"000000001",
  4115=>"000000000",
  4116=>"011000110",
  4117=>"000111111",
  4118=>"111111111",
  4119=>"011011001",
  4120=>"110000000",
  4121=>"110000000",
  4122=>"011011000",
  4123=>"000100111",
  4124=>"111111111",
  4125=>"000010000",
  4126=>"111100101",
  4127=>"001111111",
  4128=>"111111011",
  4129=>"001000100",
  4130=>"110110100",
  4131=>"111010001",
  4132=>"000000000",
  4133=>"001001111",
  4134=>"100100110",
  4135=>"011010011",
  4136=>"011011000",
  4137=>"000111111",
  4138=>"011000000",
  4139=>"000000111",
  4140=>"110110100",
  4141=>"000000000",
  4142=>"111100111",
  4143=>"000010000",
  4144=>"100000111",
  4145=>"011011010",
  4146=>"001001000",
  4147=>"100111000",
  4148=>"010010000",
  4149=>"011000000",
  4150=>"010101111",
  4151=>"000000000",
  4152=>"000000111",
  4153=>"000000000",
  4154=>"111111111",
  4155=>"110111111",
  4156=>"111100101",
  4157=>"011111100",
  4158=>"000000000",
  4159=>"111000101",
  4160=>"000000111",
  4161=>"010101101",
  4162=>"101000100",
  4163=>"000000011",
  4164=>"100010000",
  4165=>"101110110",
  4166=>"111111010",
  4167=>"111101111",
  4168=>"000001000",
  4169=>"110110110",
  4170=>"000010000",
  4171=>"111111111",
  4172=>"111111111",
  4173=>"000000111",
  4174=>"111011111",
  4175=>"111101111",
  4176=>"000000000",
  4177=>"000100111",
  4178=>"111111111",
  4179=>"011101100",
  4180=>"011111111",
  4181=>"110000000",
  4182=>"111111111",
  4183=>"111111000",
  4184=>"111000000",
  4185=>"111000101",
  4186=>"000000111",
  4187=>"010110011",
  4188=>"111000010",
  4189=>"101000001",
  4190=>"111111110",
  4191=>"100111111",
  4192=>"100100100",
  4193=>"101111111",
  4194=>"000111111",
  4195=>"001001101",
  4196=>"111110000",
  4197=>"111111111",
  4198=>"011011111",
  4199=>"001001111",
  4200=>"111111111",
  4201=>"010000000",
  4202=>"000011000",
  4203=>"110110100",
  4204=>"000000000",
  4205=>"010111010",
  4206=>"111101101",
  4207=>"111111111",
  4208=>"001101111",
  4209=>"000001111",
  4210=>"000110110",
  4211=>"101100101",
  4212=>"001111111",
  4213=>"000000111",
  4214=>"010000000",
  4215=>"101111001",
  4216=>"111111111",
  4217=>"000000000",
  4218=>"111101001",
  4219=>"001111011",
  4220=>"111101001",
  4221=>"000000000",
  4222=>"001000000",
  4223=>"000101111",
  4224=>"011011111",
  4225=>"000001000",
  4226=>"111111111",
  4227=>"111000000",
  4228=>"000000000",
  4229=>"111100001",
  4230=>"000000001",
  4231=>"011000000",
  4232=>"111110000",
  4233=>"100000011",
  4234=>"111111111",
  4235=>"000001011",
  4236=>"111001000",
  4237=>"111111010",
  4238=>"100010000",
  4239=>"000001011",
  4240=>"111001101",
  4241=>"110000000",
  4242=>"000010000",
  4243=>"111000100",
  4244=>"001111111",
  4245=>"001000011",
  4246=>"011000000",
  4247=>"110100101",
  4248=>"000001000",
  4249=>"000000011",
  4250=>"000111111",
  4251=>"111111111",
  4252=>"110110010",
  4253=>"111011111",
  4254=>"111111111",
  4255=>"000000000",
  4256=>"000010000",
  4257=>"110111000",
  4258=>"111111111",
  4259=>"000111111",
  4260=>"011001011",
  4261=>"011011111",
  4262=>"110000000",
  4263=>"111100100",
  4264=>"000000000",
  4265=>"101000100",
  4266=>"111111000",
  4267=>"110011111",
  4268=>"100110000",
  4269=>"000101111",
  4270=>"001000000",
  4271=>"111101000",
  4272=>"011111011",
  4273=>"001001100",
  4274=>"010110010",
  4275=>"111101111",
  4276=>"110000011",
  4277=>"000000011",
  4278=>"101000000",
  4279=>"111111010",
  4280=>"000000000",
  4281=>"000111111",
  4282=>"111000000",
  4283=>"001011111",
  4284=>"000000001",
  4285=>"000111010",
  4286=>"000000000",
  4287=>"111111111",
  4288=>"110111111",
  4289=>"001011000",
  4290=>"010111111",
  4291=>"111111111",
  4292=>"111110000",
  4293=>"000000000",
  4294=>"010000000",
  4295=>"111111111",
  4296=>"000010111",
  4297=>"101001111",
  4298=>"001001001",
  4299=>"000000000",
  4300=>"000011111",
  4301=>"100100101",
  4302=>"111111000",
  4303=>"000000000",
  4304=>"110101111",
  4305=>"001111111",
  4306=>"111000000",
  4307=>"000010010",
  4308=>"001100000",
  4309=>"101100000",
  4310=>"001000000",
  4311=>"000000000",
  4312=>"110111000",
  4313=>"111001111",
  4314=>"000110110",
  4315=>"001011111",
  4316=>"100110000",
  4317=>"100000000",
  4318=>"111111110",
  4319=>"000000111",
  4320=>"000000111",
  4321=>"010000111",
  4322=>"000110110",
  4323=>"111111010",
  4324=>"000000000",
  4325=>"011111110",
  4326=>"000000000",
  4327=>"011111010",
  4328=>"111111010",
  4329=>"000010011",
  4330=>"000000100",
  4331=>"000111111",
  4332=>"111000100",
  4333=>"000000000",
  4334=>"101000000",
  4335=>"000001011",
  4336=>"101000000",
  4337=>"111000110",
  4338=>"111001111",
  4339=>"010000111",
  4340=>"111111111",
  4341=>"000100110",
  4342=>"100111111",
  4343=>"001011010",
  4344=>"010110010",
  4345=>"000011011",
  4346=>"000000101",
  4347=>"100100001",
  4348=>"000011001",
  4349=>"001000001",
  4350=>"111001000",
  4351=>"000001111",
  4352=>"001000000",
  4353=>"100100100",
  4354=>"000000000",
  4355=>"111001000",
  4356=>"000000111",
  4357=>"000011111",
  4358=>"111111111",
  4359=>"001011011",
  4360=>"100111111",
  4361=>"000000001",
  4362=>"011011101",
  4363=>"111111111",
  4364=>"000000000",
  4365=>"110100101",
  4366=>"000011011",
  4367=>"010010000",
  4368=>"000010111",
  4369=>"011111110",
  4370=>"111001001",
  4371=>"010111011",
  4372=>"000000111",
  4373=>"001111111",
  4374=>"101100100",
  4375=>"000000101",
  4376=>"110111111",
  4377=>"110110000",
  4378=>"100010000",
  4379=>"000000000",
  4380=>"100100100",
  4381=>"101000001",
  4382=>"000101000",
  4383=>"000000001",
  4384=>"111101000",
  4385=>"000000111",
  4386=>"000000010",
  4387=>"000001111",
  4388=>"111101100",
  4389=>"000111111",
  4390=>"011111111",
  4391=>"111011110",
  4392=>"111000000",
  4393=>"010101000",
  4394=>"110111010",
  4395=>"111100100",
  4396=>"001110100",
  4397=>"111111111",
  4398=>"011011001",
  4399=>"111111110",
  4400=>"110110010",
  4401=>"000000000",
  4402=>"100000111",
  4403=>"111111011",
  4404=>"010111111",
  4405=>"111010000",
  4406=>"010110110",
  4407=>"111011000",
  4408=>"000000000",
  4409=>"100000101",
  4410=>"111000000",
  4411=>"111100111",
  4412=>"100110001",
  4413=>"100011111",
  4414=>"111111001",
  4415=>"110000110",
  4416=>"111100000",
  4417=>"000000001",
  4418=>"110111110",
  4419=>"100000000",
  4420=>"100000110",
  4421=>"001000000",
  4422=>"111011000",
  4423=>"000000100",
  4424=>"101000000",
  4425=>"110000011",
  4426=>"100111111",
  4427=>"000000000",
  4428=>"001000101",
  4429=>"000010000",
  4430=>"111000000",
  4431=>"101000000",
  4432=>"101100000",
  4433=>"000000011",
  4434=>"111110010",
  4435=>"011011010",
  4436=>"111111011",
  4437=>"001001001",
  4438=>"000000000",
  4439=>"100101101",
  4440=>"000000100",
  4441=>"000000000",
  4442=>"000000000",
  4443=>"000000000",
  4444=>"011011011",
  4445=>"111111000",
  4446=>"111011010",
  4447=>"000000000",
  4448=>"011011001",
  4449=>"111000000",
  4450=>"001000000",
  4451=>"111111111",
  4452=>"111111111",
  4453=>"000000111",
  4454=>"000000110",
  4455=>"001000000",
  4456=>"110100100",
  4457=>"000000001",
  4458=>"000000000",
  4459=>"111001111",
  4460=>"011111111",
  4461=>"011011111",
  4462=>"110111111",
  4463=>"100100101",
  4464=>"111111111",
  4465=>"000000010",
  4466=>"111010000",
  4467=>"110111110",
  4468=>"111111010",
  4469=>"111111100",
  4470=>"111101101",
  4471=>"111110100",
  4472=>"100000000",
  4473=>"011001111",
  4474=>"111111111",
  4475=>"000111111",
  4476=>"111111111",
  4477=>"100110111",
  4478=>"011011011",
  4479=>"000111111",
  4480=>"011000000",
  4481=>"110111000",
  4482=>"111011011",
  4483=>"000000000",
  4484=>"000010111",
  4485=>"010010000",
  4486=>"111111111",
  4487=>"111000111",
  4488=>"000100100",
  4489=>"000011001",
  4490=>"000000000",
  4491=>"000110000",
  4492=>"100000111",
  4493=>"110100100",
  4494=>"000011010",
  4495=>"110000000",
  4496=>"101000111",
  4497=>"111000101",
  4498=>"000010000",
  4499=>"001011000",
  4500=>"111111111",
  4501=>"010010000",
  4502=>"111111000",
  4503=>"000001011",
  4504=>"000000111",
  4505=>"111111111",
  4506=>"000000000",
  4507=>"100000000",
  4508=>"011011010",
  4509=>"001000001",
  4510=>"101100110",
  4511=>"000110111",
  4512=>"001000000",
  4513=>"111101111",
  4514=>"010011000",
  4515=>"000011000",
  4516=>"000000000",
  4517=>"111100100",
  4518=>"111000111",
  4519=>"010010110",
  4520=>"111111110",
  4521=>"110111111",
  4522=>"111011111",
  4523=>"000001111",
  4524=>"111111111",
  4525=>"000000110",
  4526=>"000000001",
  4527=>"001000000",
  4528=>"001001101",
  4529=>"001000000",
  4530=>"000000100",
  4531=>"000000111",
  4532=>"111111111",
  4533=>"111000001",
  4534=>"111010000",
  4535=>"111111111",
  4536=>"000000111",
  4537=>"011111011",
  4538=>"111111111",
  4539=>"000000000",
  4540=>"000000000",
  4541=>"010000000",
  4542=>"000111000",
  4543=>"000000111",
  4544=>"111111001",
  4545=>"001001001",
  4546=>"011111011",
  4547=>"100100101",
  4548=>"111111111",
  4549=>"001000100",
  4550=>"011111110",
  4551=>"100100100",
  4552=>"000000000",
  4553=>"001101011",
  4554=>"100101111",
  4555=>"000100000",
  4556=>"000111111",
  4557=>"000000000",
  4558=>"111111111",
  4559=>"100100111",
  4560=>"111111111",
  4561=>"000000000",
  4562=>"011111111",
  4563=>"111001101",
  4564=>"101100100",
  4565=>"000001000",
  4566=>"111010000",
  4567=>"011011111",
  4568=>"000100100",
  4569=>"000000001",
  4570=>"000000101",
  4571=>"001000111",
  4572=>"000111001",
  4573=>"011011111",
  4574=>"110000110",
  4575=>"111111011",
  4576=>"000000111",
  4577=>"000000000",
  4578=>"001111111",
  4579=>"011011010",
  4580=>"111000000",
  4581=>"011000000",
  4582=>"100101111",
  4583=>"111111110",
  4584=>"000001001",
  4585=>"111110111",
  4586=>"000000010",
  4587=>"001011111",
  4588=>"001101111",
  4589=>"000000000",
  4590=>"111101111",
  4591=>"110000000",
  4592=>"100000011",
  4593=>"010110000",
  4594=>"111001101",
  4595=>"000111111",
  4596=>"000000000",
  4597=>"100111111",
  4598=>"111111111",
  4599=>"111111100",
  4600=>"011011101",
  4601=>"000101000",
  4602=>"000111111",
  4603=>"100000000",
  4604=>"111000001",
  4605=>"000101111",
  4606=>"111111111",
  4607=>"111111111",
  4608=>"000000001",
  4609=>"000000000",
  4610=>"000000101",
  4611=>"111111111",
  4612=>"111111111",
  4613=>"000100111",
  4614=>"111111111",
  4615=>"001001000",
  4616=>"110111010",
  4617=>"000000011",
  4618=>"111101101",
  4619=>"000000011",
  4620=>"111111111",
  4621=>"100000000",
  4622=>"000111111",
  4623=>"111111111",
  4624=>"000000000",
  4625=>"000111111",
  4626=>"111111111",
  4627=>"000000000",
  4628=>"000111111",
  4629=>"111111111",
  4630=>"100100100",
  4631=>"000001011",
  4632=>"000100000",
  4633=>"000001011",
  4634=>"000111010",
  4635=>"000010000",
  4636=>"100000000",
  4637=>"111111111",
  4638=>"111111110",
  4639=>"000011011",
  4640=>"100100100",
  4641=>"111110110",
  4642=>"111101111",
  4643=>"000000000",
  4644=>"000000000",
  4645=>"111111110",
  4646=>"000000000",
  4647=>"111011001",
  4648=>"111111011",
  4649=>"000000000",
  4650=>"000000000",
  4651=>"111111111",
  4652=>"000111111",
  4653=>"000110111",
  4654=>"000000110",
  4655=>"111111101",
  4656=>"100000000",
  4657=>"111111111",
  4658=>"100100000",
  4659=>"000000000",
  4660=>"110100100",
  4661=>"110110111",
  4662=>"111001111",
  4663=>"011010000",
  4664=>"111000001",
  4665=>"000000101",
  4666=>"111111111",
  4667=>"000000000",
  4668=>"111000000",
  4669=>"001000000",
  4670=>"000000000",
  4671=>"000000000",
  4672=>"111111110",
  4673=>"110110000",
  4674=>"111000000",
  4675=>"000110000",
  4676=>"111111111",
  4677=>"101101110",
  4678=>"111111111",
  4679=>"111111000",
  4680=>"010000110",
  4681=>"000011111",
  4682=>"011110000",
  4683=>"000110111",
  4684=>"000011111",
  4685=>"110110100",
  4686=>"000000000",
  4687=>"000000000",
  4688=>"101001000",
  4689=>"011111110",
  4690=>"000001111",
  4691=>"110110110",
  4692=>"000000000",
  4693=>"000111111",
  4694=>"111111111",
  4695=>"000001111",
  4696=>"111111011",
  4697=>"000000000",
  4698=>"111111111",
  4699=>"011001001",
  4700=>"000111111",
  4701=>"111111111",
  4702=>"001000000",
  4703=>"111001001",
  4704=>"111101001",
  4705=>"000100111",
  4706=>"000000111",
  4707=>"000100111",
  4708=>"111011000",
  4709=>"000000000",
  4710=>"111110000",
  4711=>"111111111",
  4712=>"000000000",
  4713=>"001000000",
  4714=>"001101111",
  4715=>"000000000",
  4716=>"000000000",
  4717=>"110111110",
  4718=>"111111110",
  4719=>"000000000",
  4720=>"110111111",
  4721=>"000000000",
  4722=>"001111000",
  4723=>"011001111",
  4724=>"000000001",
  4725=>"110010001",
  4726=>"000000000",
  4727=>"000000001",
  4728=>"110111111",
  4729=>"100100000",
  4730=>"000111111",
  4731=>"111111111",
  4732=>"010010110",
  4733=>"000000000",
  4734=>"000000000",
  4735=>"000000100",
  4736=>"111111111",
  4737=>"000110100",
  4738=>"000000000",
  4739=>"001111111",
  4740=>"111111110",
  4741=>"001000111",
  4742=>"001011111",
  4743=>"111111111",
  4744=>"111111111",
  4745=>"001101111",
  4746=>"000000010",
  4747=>"000000100",
  4748=>"111111011",
  4749=>"111001000",
  4750=>"011111000",
  4751=>"000000111",
  4752=>"111111111",
  4753=>"111111111",
  4754=>"000100000",
  4755=>"000000100",
  4756=>"000100111",
  4757=>"100000000",
  4758=>"111111111",
  4759=>"110110110",
  4760=>"001111111",
  4761=>"011000000",
  4762=>"111111111",
  4763=>"010010000",
  4764=>"000000000",
  4765=>"100110000",
  4766=>"111111111",
  4767=>"111111111",
  4768=>"111110111",
  4769=>"111000000",
  4770=>"111111111",
  4771=>"000000011",
  4772=>"110111110",
  4773=>"000000001",
  4774=>"000000000",
  4775=>"011001111",
  4776=>"011011111",
  4777=>"000001001",
  4778=>"000110111",
  4779=>"000000000",
  4780=>"001111111",
  4781=>"110110110",
  4782=>"000001111",
  4783=>"111011011",
  4784=>"000000001",
  4785=>"011011011",
  4786=>"111111011",
  4787=>"000000010",
  4788=>"110110110",
  4789=>"001000000",
  4790=>"000000001",
  4791=>"000000001",
  4792=>"000000000",
  4793=>"111111001",
  4794=>"000000001",
  4795=>"011111000",
  4796=>"000100110",
  4797=>"111111010",
  4798=>"000001000",
  4799=>"111111111",
  4800=>"011011011",
  4801=>"001111111",
  4802=>"000000000",
  4803=>"000000010",
  4804=>"111111111",
  4805=>"101101100",
  4806=>"000111111",
  4807=>"100100000",
  4808=>"111111100",
  4809=>"111111110",
  4810=>"000000000",
  4811=>"111101111",
  4812=>"000000000",
  4813=>"100101111",
  4814=>"000000000",
  4815=>"111111000",
  4816=>"000000000",
  4817=>"111111111",
  4818=>"000000000",
  4819=>"110111111",
  4820=>"111111111",
  4821=>"011111111",
  4822=>"000000000",
  4823=>"010111111",
  4824=>"101111100",
  4825=>"010011000",
  4826=>"000000001",
  4827=>"001011011",
  4828=>"111000000",
  4829=>"111111111",
  4830=>"011000110",
  4831=>"000000001",
  4832=>"000000000",
  4833=>"000000110",
  4834=>"000000000",
  4835=>"111111111",
  4836=>"110111111",
  4837=>"110110111",
  4838=>"000000000",
  4839=>"000000000",
  4840=>"000000000",
  4841=>"101111111",
  4842=>"111111111",
  4843=>"000100100",
  4844=>"111111111",
  4845=>"001100110",
  4846=>"011001101",
  4847=>"101000100",
  4848=>"001000000",
  4849=>"000000001",
  4850=>"000000000",
  4851=>"000000000",
  4852=>"000000011",
  4853=>"111111001",
  4854=>"001111100",
  4855=>"111110110",
  4856=>"100111111",
  4857=>"000000000",
  4858=>"111011000",
  4859=>"111111111",
  4860=>"000001101",
  4861=>"000000000",
  4862=>"001111101",
  4863=>"000000101",
  4864=>"000000000",
  4865=>"001110111",
  4866=>"010000000",
  4867=>"000011000",
  4868=>"111000000",
  4869=>"000000000",
  4870=>"111110000",
  4871=>"110111111",
  4872=>"001000001",
  4873=>"000000000",
  4874=>"100000000",
  4875=>"011010000",
  4876=>"011011011",
  4877=>"101100100",
  4878=>"111111111",
  4879=>"000000000",
  4880=>"100000001",
  4881=>"111100000",
  4882=>"111111000",
  4883=>"000000000",
  4884=>"000000000",
  4885=>"011111000",
  4886=>"111011000",
  4887=>"111111111",
  4888=>"000000000",
  4889=>"111111110",
  4890=>"001110111",
  4891=>"001000000",
  4892=>"111111110",
  4893=>"000000000",
  4894=>"000000111",
  4895=>"111111001",
  4896=>"111111000",
  4897=>"000110111",
  4898=>"000110100",
  4899=>"111111001",
  4900=>"000000000",
  4901=>"111111111",
  4902=>"111100111",
  4903=>"101111011",
  4904=>"000111111",
  4905=>"000000001",
  4906=>"101001000",
  4907=>"000000000",
  4908=>"110110111",
  4909=>"110110111",
  4910=>"000000000",
  4911=>"000010000",
  4912=>"001011010",
  4913=>"000000000",
  4914=>"001100111",
  4915=>"011001100",
  4916=>"000000000",
  4917=>"000000000",
  4918=>"000000000",
  4919=>"000001000",
  4920=>"111100000",
  4921=>"000000000",
  4922=>"000100000",
  4923=>"111111110",
  4924=>"100000000",
  4925=>"000000101",
  4926=>"111111011",
  4927=>"001001100",
  4928=>"000100111",
  4929=>"000000000",
  4930=>"000000000",
  4931=>"010000000",
  4932=>"111111111",
  4933=>"010100000",
  4934=>"100111000",
  4935=>"111101111",
  4936=>"000000111",
  4937=>"011000000",
  4938=>"111111111",
  4939=>"011000000",
  4940=>"111000000",
  4941=>"100000100",
  4942=>"000000001",
  4943=>"011011001",
  4944=>"100000101",
  4945=>"111111011",
  4946=>"111111111",
  4947=>"000000000",
  4948=>"000000000",
  4949=>"011111111",
  4950=>"011000000",
  4951=>"111111111",
  4952=>"000000000",
  4953=>"111110000",
  4954=>"111111111",
  4955=>"000000000",
  4956=>"001101000",
  4957=>"000111111",
  4958=>"111011011",
  4959=>"010000000",
  4960=>"000000000",
  4961=>"000000000",
  4962=>"011001000",
  4963=>"000000100",
  4964=>"001000000",
  4965=>"000000000",
  4966=>"111000001",
  4967=>"001011000",
  4968=>"011001000",
  4969=>"111111000",
  4970=>"000000011",
  4971=>"101110111",
  4972=>"100111000",
  4973=>"000011111",
  4974=>"110010000",
  4975=>"000011111",
  4976=>"000000000",
  4977=>"111001001",
  4978=>"111111111",
  4979=>"110100111",
  4980=>"000000000",
  4981=>"000000000",
  4982=>"000000000",
  4983=>"001111000",
  4984=>"000000000",
  4985=>"111111111",
  4986=>"001000000",
  4987=>"110000111",
  4988=>"001000000",
  4989=>"000000100",
  4990=>"111111111",
  4991=>"000000000",
  4992=>"111111111",
  4993=>"000000000",
  4994=>"000000000",
  4995=>"000000000",
  4996=>"000110111",
  4997=>"000000000",
  4998=>"011000000",
  4999=>"001010011",
  5000=>"111011011",
  5001=>"000100000",
  5002=>"000000110",
  5003=>"011111111",
  5004=>"101000000",
  5005=>"001111111",
  5006=>"111111111",
  5007=>"000000111",
  5008=>"000000000",
  5009=>"111111111",
  5010=>"111111001",
  5011=>"001000000",
  5012=>"111111111",
  5013=>"010000110",
  5014=>"010110000",
  5015=>"000000000",
  5016=>"111111110",
  5017=>"111110000",
  5018=>"111111110",
  5019=>"111111111",
  5020=>"100111000",
  5021=>"000001001",
  5022=>"000000000",
  5023=>"000100111",
  5024=>"101101100",
  5025=>"111111111",
  5026=>"000000000",
  5027=>"111110110",
  5028=>"000000000",
  5029=>"111101111",
  5030=>"001000000",
  5031=>"000100000",
  5032=>"111010111",
  5033=>"001011011",
  5034=>"001001001",
  5035=>"100000110",
  5036=>"000000011",
  5037=>"111001001",
  5038=>"111111111",
  5039=>"100111111",
  5040=>"111111111",
  5041=>"111110000",
  5042=>"111111111",
  5043=>"111111110",
  5044=>"111111111",
  5045=>"000000000",
  5046=>"000011000",
  5047=>"000000000",
  5048=>"100100100",
  5049=>"000000001",
  5050=>"001001000",
  5051=>"111000000",
  5052=>"000000000",
  5053=>"100110110",
  5054=>"000000000",
  5055=>"001011011",
  5056=>"000000000",
  5057=>"111111111",
  5058=>"000000000",
  5059=>"000000000",
  5060=>"100100000",
  5061=>"001001111",
  5062=>"000111100",
  5063=>"000110000",
  5064=>"001000000",
  5065=>"000101001",
  5066=>"011011000",
  5067=>"110110111",
  5068=>"011000000",
  5069=>"000000000",
  5070=>"110111101",
  5071=>"000110000",
  5072=>"000000000",
  5073=>"101001001",
  5074=>"000000010",
  5075=>"111111110",
  5076=>"011111111",
  5077=>"111001011",
  5078=>"110111111",
  5079=>"110111111",
  5080=>"000001011",
  5081=>"001100100",
  5082=>"000100010",
  5083=>"001001000",
  5084=>"000111111",
  5085=>"110001001",
  5086=>"000000000",
  5087=>"011111111",
  5088=>"111111111",
  5089=>"110100000",
  5090=>"000101011",
  5091=>"001001000",
  5092=>"000100110",
  5093=>"010100100",
  5094=>"111111101",
  5095=>"111011011",
  5096=>"111111011",
  5097=>"000000010",
  5098=>"111000000",
  5099=>"111111111",
  5100=>"110100000",
  5101=>"000100100",
  5102=>"000101101",
  5103=>"111111111",
  5104=>"100100100",
  5105=>"000000111",
  5106=>"100111000",
  5107=>"100000000",
  5108=>"100110111",
  5109=>"000111000",
  5110=>"000000110",
  5111=>"000000100",
  5112=>"110100100",
  5113=>"100111101",
  5114=>"000000101",
  5115=>"111111111",
  5116=>"111111111",
  5117=>"000000000",
  5118=>"100000001",
  5119=>"000000000",
  5120=>"111111100",
  5121=>"111111111",
  5122=>"111011001",
  5123=>"111111111",
  5124=>"000110100",
  5125=>"111111110",
  5126=>"111111111",
  5127=>"000000000",
  5128=>"011011011",
  5129=>"000000000",
  5130=>"000000001",
  5131=>"111011111",
  5132=>"011011011",
  5133=>"111111111",
  5134=>"000000100",
  5135=>"111110111",
  5136=>"001000001",
  5137=>"111111000",
  5138=>"111111111",
  5139=>"110111111",
  5140=>"000111111",
  5141=>"000000000",
  5142=>"111111011",
  5143=>"111111111",
  5144=>"111111111",
  5145=>"001011111",
  5146=>"000000100",
  5147=>"111111110",
  5148=>"001011000",
  5149=>"011000100",
  5150=>"000000000",
  5151=>"011000000",
  5152=>"000111011",
  5153=>"111111111",
  5154=>"110111111",
  5155=>"110000011",
  5156=>"000001011",
  5157=>"111111110",
  5158=>"001101101",
  5159=>"000000000",
  5160=>"110110111",
  5161=>"000111111",
  5162=>"000000000",
  5163=>"000110111",
  5164=>"000000111",
  5165=>"000000000",
  5166=>"111111111",
  5167=>"000000000",
  5168=>"111111111",
  5169=>"000000000",
  5170=>"000000100",
  5171=>"000000111",
  5172=>"111111110",
  5173=>"111001000",
  5174=>"011111100",
  5175=>"110110110",
  5176=>"000000000",
  5177=>"110000000",
  5178=>"000100111",
  5179=>"000111111",
  5180=>"111011011",
  5181=>"000110000",
  5182=>"011001001",
  5183=>"111111111",
  5184=>"000000000",
  5185=>"111011010",
  5186=>"111111101",
  5187=>"111111111",
  5188=>"000000000",
  5189=>"000000000",
  5190=>"000000111",
  5191=>"111111111",
  5192=>"001001000",
  5193=>"111001101",
  5194=>"001000001",
  5195=>"101111101",
  5196=>"111011011",
  5197=>"000000001",
  5198=>"000000000",
  5199=>"100101101",
  5200=>"000000000",
  5201=>"000100000",
  5202=>"000000000",
  5203=>"000110001",
  5204=>"001111111",
  5205=>"000000000",
  5206=>"001101111",
  5207=>"001001011",
  5208=>"000000100",
  5209=>"100000000",
  5210=>"000010111",
  5211=>"011001001",
  5212=>"111111111",
  5213=>"010111011",
  5214=>"000000000",
  5215=>"011011000",
  5216=>"000000101",
  5217=>"110110110",
  5218=>"111111111",
  5219=>"111111111",
  5220=>"000000111",
  5221=>"110110110",
  5222=>"000001001",
  5223=>"110100000",
  5224=>"111111111",
  5225=>"000000000",
  5226=>"000000000",
  5227=>"111111111",
  5228=>"111111111",
  5229=>"111111111",
  5230=>"001001000",
  5231=>"111111000",
  5232=>"000000111",
  5233=>"110111100",
  5234=>"000000000",
  5235=>"001100110",
  5236=>"000000100",
  5237=>"000000000",
  5238=>"000110111",
  5239=>"111111111",
  5240=>"111111111",
  5241=>"111011000",
  5242=>"111111100",
  5243=>"011111111",
  5244=>"100000100",
  5245=>"111011011",
  5246=>"111111111",
  5247=>"000001001",
  5248=>"111111001",
  5249=>"011111111",
  5250=>"111111111",
  5251=>"000000000",
  5252=>"011111111",
  5253=>"101000000",
  5254=>"111011111",
  5255=>"000000000",
  5256=>"000110111",
  5257=>"111110111",
  5258=>"101101111",
  5259=>"000110110",
  5260=>"000000000",
  5261=>"000000000",
  5262=>"000000000",
  5263=>"000000110",
  5264=>"000000001",
  5265=>"000000111",
  5266=>"000010011",
  5267=>"000000001",
  5268=>"110100110",
  5269=>"001001011",
  5270=>"000000000",
  5271=>"111110110",
  5272=>"011111111",
  5273=>"000001111",
  5274=>"111100100",
  5275=>"001000000",
  5276=>"000111111",
  5277=>"111100000",
  5278=>"111111111",
  5279=>"001001000",
  5280=>"111110111",
  5281=>"110110111",
  5282=>"000111101",
  5283=>"000110111",
  5284=>"001010011",
  5285=>"000111111",
  5286=>"000100100",
  5287=>"001011011",
  5288=>"000100001",
  5289=>"001000000",
  5290=>"100000000",
  5291=>"110011110",
  5292=>"111111000",
  5293=>"111111111",
  5294=>"000100110",
  5295=>"000000010",
  5296=>"000000000",
  5297=>"111111011",
  5298=>"000101100",
  5299=>"100111111",
  5300=>"001001000",
  5301=>"111111111",
  5302=>"011011011",
  5303=>"110010111",
  5304=>"000001000",
  5305=>"000000000",
  5306=>"000000000",
  5307=>"011111011",
  5308=>"000001000",
  5309=>"000000000",
  5310=>"000000010",
  5311=>"111111111",
  5312=>"100000000",
  5313=>"101101111",
  5314=>"111111111",
  5315=>"010111000",
  5316=>"110100000",
  5317=>"000111011",
  5318=>"111011000",
  5319=>"111111111",
  5320=>"000011000",
  5321=>"111111111",
  5322=>"100000100",
  5323=>"111111111",
  5324=>"000000000",
  5325=>"111000000",
  5326=>"011001101",
  5327=>"111001001",
  5328=>"110010000",
  5329=>"011100110",
  5330=>"000011101",
  5331=>"101000000",
  5332=>"110111111",
  5333=>"111111111",
  5334=>"000000001",
  5335=>"000000000",
  5336=>"010011011",
  5337=>"000000110",
  5338=>"111111010",
  5339=>"000000010",
  5340=>"001000001",
  5341=>"000111111",
  5342=>"000110100",
  5343=>"000000000",
  5344=>"110111111",
  5345=>"000001001",
  5346=>"111111000",
  5347=>"100111111",
  5348=>"111111111",
  5349=>"110100000",
  5350=>"001001001",
  5351=>"111111111",
  5352=>"110111110",
  5353=>"111111111",
  5354=>"111111111",
  5355=>"001101111",
  5356=>"111111111",
  5357=>"000010010",
  5358=>"100111111",
  5359=>"000000000",
  5360=>"111111000",
  5361=>"000101111",
  5362=>"000111110",
  5363=>"000000000",
  5364=>"111010111",
  5365=>"000000000",
  5366=>"111111111",
  5367=>"111111111",
  5368=>"111111111",
  5369=>"000000000",
  5370=>"000000001",
  5371=>"000000000",
  5372=>"001001010",
  5373=>"001001111",
  5374=>"011111111",
  5375=>"001111011",
  5376=>"100111000",
  5377=>"011011000",
  5378=>"000000000",
  5379=>"000010011",
  5380=>"000000000",
  5381=>"000000000",
  5382=>"000000111",
  5383=>"000000100",
  5384=>"111111000",
  5385=>"000000111",
  5386=>"111111111",
  5387=>"110000110",
  5388=>"000000000",
  5389=>"011111010",
  5390=>"000101111",
  5391=>"111111000",
  5392=>"000000110",
  5393=>"000001000",
  5394=>"111011001",
  5395=>"111111011",
  5396=>"000000100",
  5397=>"000000110",
  5398=>"010110110",
  5399=>"111111011",
  5400=>"010000100",
  5401=>"001111111",
  5402=>"111111101",
  5403=>"110110000",
  5404=>"000010000",
  5405=>"000111110",
  5406=>"000000000",
  5407=>"011111111",
  5408=>"010110111",
  5409=>"000100000",
  5410=>"000100111",
  5411=>"111111110",
  5412=>"110111111",
  5413=>"000000000",
  5414=>"111010000",
  5415=>"111111110",
  5416=>"111000000",
  5417=>"000000001",
  5418=>"000001111",
  5419=>"000111111",
  5420=>"011011000",
  5421=>"000110110",
  5422=>"111111111",
  5423=>"111111001",
  5424=>"110110110",
  5425=>"000000000",
  5426=>"010000011",
  5427=>"101111111",
  5428=>"000000000",
  5429=>"111111111",
  5430=>"110110111",
  5431=>"000110111",
  5432=>"111111100",
  5433=>"000000101",
  5434=>"001101111",
  5435=>"100000000",
  5436=>"000110111",
  5437=>"011011011",
  5438=>"000010011",
  5439=>"001111111",
  5440=>"000000000",
  5441=>"010011011",
  5442=>"111111111",
  5443=>"011110110",
  5444=>"010000000",
  5445=>"000000000",
  5446=>"011000000",
  5447=>"011011111",
  5448=>"000010111",
  5449=>"111111111",
  5450=>"000000000",
  5451=>"110000000",
  5452=>"000000000",
  5453=>"101111110",
  5454=>"110111111",
  5455=>"000110110",
  5456=>"011011000",
  5457=>"000000000",
  5458=>"100000000",
  5459=>"001111111",
  5460=>"001000000",
  5461=>"011001011",
  5462=>"000000000",
  5463=>"111111100",
  5464=>"000000000",
  5465=>"111111111",
  5466=>"110111000",
  5467=>"110100100",
  5468=>"000000000",
  5469=>"001000100",
  5470=>"111000011",
  5471=>"110110110",
  5472=>"111111101",
  5473=>"000000000",
  5474=>"011000000",
  5475=>"000000000",
  5476=>"001001011",
  5477=>"000000000",
  5478=>"000000010",
  5479=>"011111011",
  5480=>"011000000",
  5481=>"110111111",
  5482=>"000000000",
  5483=>"011011110",
  5484=>"001111001",
  5485=>"000000000",
  5486=>"000000000",
  5487=>"000000000",
  5488=>"000000101",
  5489=>"000000000",
  5490=>"111111111",
  5491=>"111111111",
  5492=>"000100111",
  5493=>"001000110",
  5494=>"011001000",
  5495=>"111111111",
  5496=>"111111111",
  5497=>"000000100",
  5498=>"111110111",
  5499=>"111101000",
  5500=>"111110111",
  5501=>"111000000",
  5502=>"100000000",
  5503=>"000000000",
  5504=>"000000000",
  5505=>"111101101",
  5506=>"000001001",
  5507=>"000100111",
  5508=>"111111111",
  5509=>"000000000",
  5510=>"010011000",
  5511=>"111111111",
  5512=>"000000100",
  5513=>"000000000",
  5514=>"100100100",
  5515=>"111111111",
  5516=>"111111111",
  5517=>"010011010",
  5518=>"011010000",
  5519=>"000010111",
  5520=>"111000000",
  5521=>"111111111",
  5522=>"010000000",
  5523=>"000011111",
  5524=>"111111111",
  5525=>"000101011",
  5526=>"101001101",
  5527=>"000001001",
  5528=>"000000000",
  5529=>"110110111",
  5530=>"100111111",
  5531=>"000100111",
  5532=>"100101001",
  5533=>"000110110",
  5534=>"000000000",
  5535=>"111111000",
  5536=>"111111011",
  5537=>"011010000",
  5538=>"000010001",
  5539=>"111111111",
  5540=>"011011110",
  5541=>"011111000",
  5542=>"111000000",
  5543=>"111111111",
  5544=>"100110110",
  5545=>"101100110",
  5546=>"000110111",
  5547=>"111011110",
  5548=>"000000000",
  5549=>"111100100",
  5550=>"000111111",
  5551=>"000100000",
  5552=>"000111111",
  5553=>"000001111",
  5554=>"000000000",
  5555=>"111110110",
  5556=>"000000000",
  5557=>"000000010",
  5558=>"001111010",
  5559=>"110111111",
  5560=>"100101111",
  5561=>"000111111",
  5562=>"111111111",
  5563=>"001001011",
  5564=>"101000000",
  5565=>"011001101",
  5566=>"111100100",
  5567=>"001000000",
  5568=>"110110111",
  5569=>"101101100",
  5570=>"000000000",
  5571=>"000100000",
  5572=>"110110111",
  5573=>"000000000",
  5574=>"110111111",
  5575=>"111110000",
  5576=>"000111110",
  5577=>"111111111",
  5578=>"111111111",
  5579=>"111100000",
  5580=>"000000000",
  5581=>"000000000",
  5582=>"000000000",
  5583=>"000000001",
  5584=>"000000000",
  5585=>"011111111",
  5586=>"000000001",
  5587=>"111111111",
  5588=>"111111110",
  5589=>"100110111",
  5590=>"100110111",
  5591=>"110111111",
  5592=>"000000000",
  5593=>"111111011",
  5594=>"010000100",
  5595=>"010111110",
  5596=>"111111111",
  5597=>"001100101",
  5598=>"100000000",
  5599=>"111011000",
  5600=>"000000100",
  5601=>"111111111",
  5602=>"100100000",
  5603=>"111111111",
  5604=>"000000010",
  5605=>"000001111",
  5606=>"000000110",
  5607=>"000000011",
  5608=>"000000100",
  5609=>"001000001",
  5610=>"111111110",
  5611=>"000000000",
  5612=>"001001111",
  5613=>"101001101",
  5614=>"000000000",
  5615=>"010010000",
  5616=>"111000000",
  5617=>"110111111",
  5618=>"000110110",
  5619=>"000000000",
  5620=>"111111111",
  5621=>"000000000",
  5622=>"000000011",
  5623=>"000000000",
  5624=>"000010111",
  5625=>"000000100",
  5626=>"011011111",
  5627=>"100000000",
  5628=>"111111111",
  5629=>"000000000",
  5630=>"000110000",
  5631=>"000001011",
  5632=>"010010110",
  5633=>"011000000",
  5634=>"101000000",
  5635=>"111111000",
  5636=>"100111111",
  5637=>"000000000",
  5638=>"000000000",
  5639=>"000101111",
  5640=>"111110000",
  5641=>"000111111",
  5642=>"111000000",
  5643=>"111111001",
  5644=>"110110000",
  5645=>"001000000",
  5646=>"111111011",
  5647=>"000000111",
  5648=>"111111111",
  5649=>"000010011",
  5650=>"001001001",
  5651=>"000100111",
  5652=>"111111000",
  5653=>"001111111",
  5654=>"000000000",
  5655=>"110111000",
  5656=>"001001001",
  5657=>"000000110",
  5658=>"111001000",
  5659=>"111111111",
  5660=>"000000111",
  5661=>"000000111",
  5662=>"100111111",
  5663=>"110000000",
  5664=>"000110010",
  5665=>"111111111",
  5666=>"111111111",
  5667=>"100100101",
  5668=>"111000000",
  5669=>"000000111",
  5670=>"000111111",
  5671=>"000000010",
  5672=>"110000000",
  5673=>"010111011",
  5674=>"111111111",
  5675=>"001111111",
  5676=>"000000111",
  5677=>"100110110",
  5678=>"111000100",
  5679=>"100111111",
  5680=>"000000111",
  5681=>"000000100",
  5682=>"000110111",
  5683=>"101100000",
  5684=>"010111110",
  5685=>"000111011",
  5686=>"001000000",
  5687=>"000110000",
  5688=>"000001011",
  5689=>"000000001",
  5690=>"111111000",
  5691=>"000000000",
  5692=>"100100111",
  5693=>"011011011",
  5694=>"011101111",
  5695=>"000111111",
  5696=>"110100100",
  5697=>"010010000",
  5698=>"111000000",
  5699=>"000100110",
  5700=>"110110000",
  5701=>"111111000",
  5702=>"111111000",
  5703=>"101111111",
  5704=>"100111111",
  5705=>"111000111",
  5706=>"000111111",
  5707=>"000101111",
  5708=>"111111100",
  5709=>"111001000",
  5710=>"111011111",
  5711=>"101111111",
  5712=>"000111111",
  5713=>"111110110",
  5714=>"000000000",
  5715=>"110110001",
  5716=>"000000110",
  5717=>"111000000",
  5718=>"000000000",
  5719=>"111111100",
  5720=>"000000101",
  5721=>"000000000",
  5722=>"111111111",
  5723=>"111001000",
  5724=>"011111000",
  5725=>"000010111",
  5726=>"000000000",
  5727=>"000000000",
  5728=>"000000000",
  5729=>"111000000",
  5730=>"000100000",
  5731=>"000000000",
  5732=>"001110000",
  5733=>"000000100",
  5734=>"000001111",
  5735=>"111111111",
  5736=>"111000111",
  5737=>"000110111",
  5738=>"000000111",
  5739=>"000000001",
  5740=>"111001100",
  5741=>"111100000",
  5742=>"111011000",
  5743=>"111110111",
  5744=>"110111111",
  5745=>"111111111",
  5746=>"110010010",
  5747=>"011010000",
  5748=>"000000101",
  5749=>"100111111",
  5750=>"010000000",
  5751=>"000000000",
  5752=>"111111000",
  5753=>"000111111",
  5754=>"000000100",
  5755=>"111000000",
  5756=>"000111111",
  5757=>"001000000",
  5758=>"111111111",
  5759=>"000000000",
  5760=>"000000000",
  5761=>"111111000",
  5762=>"011000001",
  5763=>"011001000",
  5764=>"100111111",
  5765=>"000000111",
  5766=>"111111100",
  5767=>"111111000",
  5768=>"000000111",
  5769=>"000000000",
  5770=>"000000000",
  5771=>"000001111",
  5772=>"111111111",
  5773=>"100000000",
  5774=>"011000111",
  5775=>"000111000",
  5776=>"111111110",
  5777=>"000000000",
  5778=>"011000000",
  5779=>"111000000",
  5780=>"111111111",
  5781=>"111111000",
  5782=>"111111000",
  5783=>"100000000",
  5784=>"111111000",
  5785=>"111101111",
  5786=>"111001000",
  5787=>"010000000",
  5788=>"111111000",
  5789=>"111111111",
  5790=>"000000111",
  5791=>"111111000",
  5792=>"111111010",
  5793=>"000011000",
  5794=>"000000001",
  5795=>"011111110",
  5796=>"100000000",
  5797=>"100111000",
  5798=>"010001111",
  5799=>"111010111",
  5800=>"000000111",
  5801=>"000000000",
  5802=>"000111000",
  5803=>"000000111",
  5804=>"000000101",
  5805=>"100100000",
  5806=>"111000000",
  5807=>"000010111",
  5808=>"000111111",
  5809=>"100000000",
  5810=>"110111111",
  5811=>"010001000",
  5812=>"000111111",
  5813=>"000000111",
  5814=>"100000111",
  5815=>"000000000",
  5816=>"111111111",
  5817=>"100101001",
  5818=>"110000000",
  5819=>"011000000",
  5820=>"100010000",
  5821=>"111111111",
  5822=>"111111000",
  5823=>"000011111",
  5824=>"000000000",
  5825=>"001000100",
  5826=>"000000111",
  5827=>"000000111",
  5828=>"000000000",
  5829=>"111111110",
  5830=>"111111111",
  5831=>"000000000",
  5832=>"111101111",
  5833=>"000000001",
  5834=>"000111110",
  5835=>"000000000",
  5836=>"000000011",
  5837=>"000100111",
  5838=>"110111011",
  5839=>"000000000",
  5840=>"000000111",
  5841=>"000000000",
  5842=>"111111000",
  5843=>"000000000",
  5844=>"100111011",
  5845=>"001001001",
  5846=>"111111111",
  5847=>"000000000",
  5848=>"111111000",
  5849=>"000000110",
  5850=>"111011000",
  5851=>"011000000",
  5852=>"000000000",
  5853=>"001000000",
  5854=>"110111111",
  5855=>"110110100",
  5856=>"111111000",
  5857=>"011111111",
  5858=>"110111111",
  5859=>"000011000",
  5860=>"111111111",
  5861=>"100100100",
  5862=>"000000100",
  5863=>"001000000",
  5864=>"111111000",
  5865=>"000000111",
  5866=>"111000001",
  5867=>"000000000",
  5868=>"000010111",
  5869=>"010000111",
  5870=>"010011111",
  5871=>"111111100",
  5872=>"000100111",
  5873=>"000010101",
  5874=>"111111100",
  5875=>"010000000",
  5876=>"111000000",
  5877=>"000000001",
  5878=>"000000011",
  5879=>"111000000",
  5880=>"000000011",
  5881=>"000100111",
  5882=>"111011000",
  5883=>"110100000",
  5884=>"001001001",
  5885=>"100100111",
  5886=>"000000101",
  5887=>"000000000",
  5888=>"010000100",
  5889=>"111111110",
  5890=>"111010111",
  5891=>"000000000",
  5892=>"100100100",
  5893=>"000000000",
  5894=>"100000000",
  5895=>"000000110",
  5896=>"000000000",
  5897=>"000111111",
  5898=>"111000000",
  5899=>"111100111",
  5900=>"111111111",
  5901=>"000111111",
  5902=>"101000100",
  5903=>"110110100",
  5904=>"000000111",
  5905=>"000000000",
  5906=>"011000000",
  5907=>"000001000",
  5908=>"000000000",
  5909=>"000111111",
  5910=>"111000011",
  5911=>"111111000",
  5912=>"000000111",
  5913=>"111010001",
  5914=>"000111000",
  5915=>"111111000",
  5916=>"110111100",
  5917=>"111111111",
  5918=>"111000000",
  5919=>"111011000",
  5920=>"000100100",
  5921=>"011001011",
  5922=>"000110111",
  5923=>"100000000",
  5924=>"111111101",
  5925=>"111111000",
  5926=>"100111110",
  5927=>"000000000",
  5928=>"000000000",
  5929=>"111111110",
  5930=>"111000111",
  5931=>"000000110",
  5932=>"111001000",
  5933=>"000001011",
  5934=>"101111000",
  5935=>"000000000",
  5936=>"001011000",
  5937=>"111111110",
  5938=>"000110110",
  5939=>"000000111",
  5940=>"111000000",
  5941=>"100111111",
  5942=>"111000000",
  5943=>"000111111",
  5944=>"111111111",
  5945=>"101111001",
  5946=>"000000101",
  5947=>"000000000",
  5948=>"000000000",
  5949=>"111000000",
  5950=>"000000000",
  5951=>"111000000",
  5952=>"000000111",
  5953=>"111111000",
  5954=>"111111000",
  5955=>"011001000",
  5956=>"000000110",
  5957=>"111111111",
  5958=>"100111111",
  5959=>"111001000",
  5960=>"000000100",
  5961=>"111111000",
  5962=>"010001000",
  5963=>"010100110",
  5964=>"010000100",
  5965=>"000000011",
  5966=>"101110111",
  5967=>"011111111",
  5968=>"111110100",
  5969=>"000111111",
  5970=>"111111111",
  5971=>"110111000",
  5972=>"000000011",
  5973=>"111111001",
  5974=>"110000100",
  5975=>"110000000",
  5976=>"111111111",
  5977=>"111001111",
  5978=>"000000000",
  5979=>"001000000",
  5980=>"100000101",
  5981=>"100000000",
  5982=>"011011001",
  5983=>"111111111",
  5984=>"010011011",
  5985=>"111000000",
  5986=>"011111111",
  5987=>"111000010",
  5988=>"110000000",
  5989=>"000000110",
  5990=>"111111111",
  5991=>"111111111",
  5992=>"011001110",
  5993=>"011010101",
  5994=>"000000000",
  5995=>"000000111",
  5996=>"100000001",
  5997=>"000001111",
  5998=>"000000000",
  5999=>"111111110",
  6000=>"000000000",
  6001=>"000000000",
  6002=>"111110111",
  6003=>"011001000",
  6004=>"000000101",
  6005=>"001101100",
  6006=>"000000000",
  6007=>"000000000",
  6008=>"111000000",
  6009=>"111111111",
  6010=>"000000000",
  6011=>"111111111",
  6012=>"111011000",
  6013=>"110111111",
  6014=>"000000111",
  6015=>"110000101",
  6016=>"111001000",
  6017=>"111111101",
  6018=>"111111110",
  6019=>"010010000",
  6020=>"011111001",
  6021=>"101101111",
  6022=>"111110111",
  6023=>"111111111",
  6024=>"111010000",
  6025=>"000000000",
  6026=>"000011000",
  6027=>"011101111",
  6028=>"111110111",
  6029=>"011011011",
  6030=>"111111000",
  6031=>"000000000",
  6032=>"111110111",
  6033=>"000000000",
  6034=>"000001001",
  6035=>"000000000",
  6036=>"111010110",
  6037=>"000000000",
  6038=>"111110000",
  6039=>"110000100",
  6040=>"000000000",
  6041=>"000011000",
  6042=>"111111111",
  6043=>"111000100",
  6044=>"111010000",
  6045=>"111111110",
  6046=>"100100111",
  6047=>"000000000",
  6048=>"100100000",
  6049=>"000100100",
  6050=>"011000000",
  6051=>"000000000",
  6052=>"011100111",
  6053=>"111111110",
  6054=>"010101000",
  6055=>"111000000",
  6056=>"001000000",
  6057=>"000110000",
  6058=>"111001001",
  6059=>"100110110",
  6060=>"100111001",
  6061=>"000000000",
  6062=>"000000000",
  6063=>"000011011",
  6064=>"000111000",
  6065=>"000000110",
  6066=>"110000000",
  6067=>"000111111",
  6068=>"101000000",
  6069=>"110000000",
  6070=>"000001000",
  6071=>"000000111",
  6072=>"000000000",
  6073=>"011111111",
  6074=>"111001000",
  6075=>"000000000",
  6076=>"001001111",
  6077=>"111001000",
  6078=>"000001111",
  6079=>"111110110",
  6080=>"111000000",
  6081=>"111100000",
  6082=>"110000111",
  6083=>"111100000",
  6084=>"111110010",
  6085=>"011000001",
  6086=>"000000111",
  6087=>"000000111",
  6088=>"000000000",
  6089=>"111111000",
  6090=>"111100000",
  6091=>"000000000",
  6092=>"111110100",
  6093=>"000000111",
  6094=>"110110000",
  6095=>"111111111",
  6096=>"000010000",
  6097=>"111111111",
  6098=>"000111111",
  6099=>"000000000",
  6100=>"010111111",
  6101=>"111111000",
  6102=>"000010001",
  6103=>"111011001",
  6104=>"111110000",
  6105=>"000000110",
  6106=>"000000111",
  6107=>"000000111",
  6108=>"000000000",
  6109=>"000000111",
  6110=>"111111000",
  6111=>"111101000",
  6112=>"010010011",
  6113=>"111111111",
  6114=>"110000000",
  6115=>"111111110",
  6116=>"110000111",
  6117=>"001111111",
  6118=>"000110110",
  6119=>"000011001",
  6120=>"111111111",
  6121=>"000000000",
  6122=>"000000111",
  6123=>"000000000",
  6124=>"111111000",
  6125=>"000000100",
  6126=>"101111111",
  6127=>"111111111",
  6128=>"101000000",
  6129=>"101001101",
  6130=>"000000000",
  6131=>"011111010",
  6132=>"111000000",
  6133=>"000000000",
  6134=>"111111111",
  6135=>"111001000",
  6136=>"000110111",
  6137=>"100111100",
  6138=>"000000001",
  6139=>"111111000",
  6140=>"011010000",
  6141=>"111111001",
  6142=>"100000000",
  6143=>"111110110",
  6144=>"111111000",
  6145=>"000000000",
  6146=>"111111111",
  6147=>"100111011",
  6148=>"000000000",
  6149=>"011111001",
  6150=>"001000101",
  6151=>"001001111",
  6152=>"111101111",
  6153=>"000000000",
  6154=>"000000100",
  6155=>"111111110",
  6156=>"000000100",
  6157=>"111111111",
  6158=>"000000000",
  6159=>"001001001",
  6160=>"111111111",
  6161=>"111111111",
  6162=>"000000110",
  6163=>"111111111",
  6164=>"100000000",
  6165=>"111101000",
  6166=>"111010010",
  6167=>"111000000",
  6168=>"011111011",
  6169=>"000001000",
  6170=>"000111111",
  6171=>"001001000",
  6172=>"000001000",
  6173=>"110110110",
  6174=>"001001010",
  6175=>"101100111",
  6176=>"001000111",
  6177=>"010010011",
  6178=>"111110110",
  6179=>"000000110",
  6180=>"111111111",
  6181=>"000000100",
  6182=>"000000000",
  6183=>"000000000",
  6184=>"000101001",
  6185=>"000000000",
  6186=>"001000000",
  6187=>"000010111",
  6188=>"000000000",
  6189=>"111111110",
  6190=>"000000111",
  6191=>"010010000",
  6192=>"100000110",
  6193=>"001001111",
  6194=>"111111111",
  6195=>"111111000",
  6196=>"000011110",
  6197=>"001001001",
  6198=>"100100111",
  6199=>"000000000",
  6200=>"111111000",
  6201=>"000001000",
  6202=>"000000000",
  6203=>"110000000",
  6204=>"000000111",
  6205=>"000110100",
  6206=>"000000000",
  6207=>"011001001",
  6208=>"000010001",
  6209=>"000000111",
  6210=>"001000001",
  6211=>"000000110",
  6212=>"111111110",
  6213=>"111111111",
  6214=>"110111111",
  6215=>"000011100",
  6216=>"000001011",
  6217=>"000000101",
  6218=>"000000000",
  6219=>"111111000",
  6220=>"011111111",
  6221=>"001000000",
  6222=>"100000000",
  6223=>"000000000",
  6224=>"000011000",
  6225=>"000110100",
  6226=>"011111011",
  6227=>"000001011",
  6228=>"111111111",
  6229=>"111111110",
  6230=>"100000000",
  6231=>"011100000",
  6232=>"100100000",
  6233=>"000000000",
  6234=>"110010110",
  6235=>"010001011",
  6236=>"111111000",
  6237=>"001111110",
  6238=>"000000000",
  6239=>"111100111",
  6240=>"000000001",
  6241=>"001000000",
  6242=>"000000111",
  6243=>"111110110",
  6244=>"000000000",
  6245=>"111111111",
  6246=>"111110011",
  6247=>"111111100",
  6248=>"111111111",
  6249=>"111111100",
  6250=>"010000111",
  6251=>"001011111",
  6252=>"000001011",
  6253=>"000000000",
  6254=>"100000000",
  6255=>"111111101",
  6256=>"000000000",
  6257=>"001001111",
  6258=>"000000001",
  6259=>"110111111",
  6260=>"001101101",
  6261=>"111111111",
  6262=>"110110110",
  6263=>"000010011",
  6264=>"000001011",
  6265=>"111111111",
  6266=>"110100100",
  6267=>"100001111",
  6268=>"011011011",
  6269=>"111110111",
  6270=>"000000000",
  6271=>"000000001",
  6272=>"000000000",
  6273=>"000000010",
  6274=>"000000001",
  6275=>"110111101",
  6276=>"000000000",
  6277=>"000000000",
  6278=>"110100110",
  6279=>"000000000",
  6280=>"100111111",
  6281=>"111100100",
  6282=>"000000001",
  6283=>"111111000",
  6284=>"000001111",
  6285=>"011110000",
  6286=>"011000000",
  6287=>"001001001",
  6288=>"110000000",
  6289=>"101111111",
  6290=>"100110000",
  6291=>"010111011",
  6292=>"000000100",
  6293=>"111111011",
  6294=>"111111000",
  6295=>"000110110",
  6296=>"110111111",
  6297=>"111111111",
  6298=>"000000011",
  6299=>"111111111",
  6300=>"000000000",
  6301=>"111111011",
  6302=>"001000110",
  6303=>"111111111",
  6304=>"000000000",
  6305=>"111111111",
  6306=>"111111111",
  6307=>"111111011",
  6308=>"101000000",
  6309=>"111000001",
  6310=>"000111111",
  6311=>"001000000",
  6312=>"000110000",
  6313=>"000000000",
  6314=>"111111111",
  6315=>"111111111",
  6316=>"110010111",
  6317=>"111111011",
  6318=>"000000011",
  6319=>"000011000",
  6320=>"000111111",
  6321=>"011000001",
  6322=>"001011001",
  6323=>"010111111",
  6324=>"100110100",
  6325=>"000000000",
  6326=>"001000111",
  6327=>"000000011",
  6328=>"011111111",
  6329=>"111100000",
  6330=>"111011001",
  6331=>"011000000",
  6332=>"000000000",
  6333=>"011000011",
  6334=>"000000000",
  6335=>"111111110",
  6336=>"111110111",
  6337=>"111001001",
  6338=>"111100111",
  6339=>"000111111",
  6340=>"000000000",
  6341=>"000000110",
  6342=>"000111111",
  6343=>"111111100",
  6344=>"111111110",
  6345=>"000010111",
  6346=>"000000000",
  6347=>"011111111",
  6348=>"110110100",
  6349=>"000111110",
  6350=>"000000001",
  6351=>"111111111",
  6352=>"100111011",
  6353=>"000000000",
  6354=>"111010011",
  6355=>"011001101",
  6356=>"111010000",
  6357=>"001001111",
  6358=>"000010010",
  6359=>"000000111",
  6360=>"000000000",
  6361=>"111111110",
  6362=>"000110111",
  6363=>"111111111",
  6364=>"111001001",
  6365=>"000100100",
  6366=>"000000000",
  6367=>"011000001",
  6368=>"000000000",
  6369=>"000000000",
  6370=>"111100000",
  6371=>"111111111",
  6372=>"111001100",
  6373=>"000000100",
  6374=>"111111111",
  6375=>"111111101",
  6376=>"111110111",
  6377=>"000000111",
  6378=>"111111001",
  6379=>"111111111",
  6380=>"001001001",
  6381=>"010010000",
  6382=>"000110000",
  6383=>"001111111",
  6384=>"111111111",
  6385=>"001011011",
  6386=>"111111111",
  6387=>"111111111",
  6388=>"000001111",
  6389=>"000000001",
  6390=>"110110111",
  6391=>"100100110",
  6392=>"111111111",
  6393=>"011111111",
  6394=>"110110001",
  6395=>"000110111",
  6396=>"101101101",
  6397=>"000000000",
  6398=>"100000010",
  6399=>"111111111",
  6400=>"111110111",
  6401=>"000010000",
  6402=>"111111111",
  6403=>"000000000",
  6404=>"111111011",
  6405=>"110011011",
  6406=>"111110000",
  6407=>"000111001",
  6408=>"110000000",
  6409=>"111111100",
  6410=>"110010011",
  6411=>"110111111",
  6412=>"110000000",
  6413=>"111111111",
  6414=>"000000000",
  6415=>"110110000",
  6416=>"101001001",
  6417=>"000000011",
  6418=>"000000111",
  6419=>"000100000",
  6420=>"111011100",
  6421=>"000111111",
  6422=>"011011010",
  6423=>"100000000",
  6424=>"000000000",
  6425=>"000000000",
  6426=>"000000011",
  6427=>"111011001",
  6428=>"000110110",
  6429=>"000100111",
  6430=>"111111111",
  6431=>"111000001",
  6432=>"100000000",
  6433=>"110000000",
  6434=>"111110000",
  6435=>"110111111",
  6436=>"000000000",
  6437=>"011000000",
  6438=>"000001011",
  6439=>"000011110",
  6440=>"011001011",
  6441=>"000001001",
  6442=>"110000111",
  6443=>"011011111",
  6444=>"100101001",
  6445=>"000000000",
  6446=>"111111111",
  6447=>"000000100",
  6448=>"001001001",
  6449=>"011011111",
  6450=>"000000000",
  6451=>"111111111",
  6452=>"111100000",
  6453=>"100111111",
  6454=>"111100100",
  6455=>"000000110",
  6456=>"111111111",
  6457=>"111110100",
  6458=>"101111101",
  6459=>"111111010",
  6460=>"000110010",
  6461=>"110111000",
  6462=>"000000110",
  6463=>"000000101",
  6464=>"000000000",
  6465=>"011110100",
  6466=>"000001111",
  6467=>"110110000",
  6468=>"111111111",
  6469=>"111000100",
  6470=>"101000110",
  6471=>"011011010",
  6472=>"111111111",
  6473=>"111111111",
  6474=>"000000011",
  6475=>"000000110",
  6476=>"011011100",
  6477=>"000111110",
  6478=>"000000111",
  6479=>"000010000",
  6480=>"101100100",
  6481=>"011111110",
  6482=>"000001111",
  6483=>"111111111",
  6484=>"111111111",
  6485=>"111111101",
  6486=>"111010000",
  6487=>"000000111",
  6488=>"001000000",
  6489=>"101001011",
  6490=>"001011111",
  6491=>"111111111",
  6492=>"000000000",
  6493=>"000000000",
  6494=>"000001001",
  6495=>"001110110",
  6496=>"000001000",
  6497=>"111111010",
  6498=>"100100100",
  6499=>"001001000",
  6500=>"001100111",
  6501=>"000000011",
  6502=>"001111011",
  6503=>"010000110",
  6504=>"000000011",
  6505=>"111111111",
  6506=>"001001101",
  6507=>"000011111",
  6508=>"001001001",
  6509=>"100000011",
  6510=>"000000000",
  6511=>"001001011",
  6512=>"000001111",
  6513=>"000000000",
  6514=>"011000000",
  6515=>"001000000",
  6516=>"101111111",
  6517=>"000001011",
  6518=>"111111110",
  6519=>"100000000",
  6520=>"000000000",
  6521=>"000000000",
  6522=>"111001001",
  6523=>"001001011",
  6524=>"110010111",
  6525=>"000000111",
  6526=>"001000100",
  6527=>"001000000",
  6528=>"000000000",
  6529=>"111001111",
  6530=>"110111111",
  6531=>"000001000",
  6532=>"110111101",
  6533=>"000000000",
  6534=>"110000000",
  6535=>"000000000",
  6536=>"001001001",
  6537=>"011111111",
  6538=>"001001001",
  6539=>"000100111",
  6540=>"000000000",
  6541=>"001000001",
  6542=>"111111001",
  6543=>"011111011",
  6544=>"110111111",
  6545=>"010110111",
  6546=>"000000001",
  6547=>"110011001",
  6548=>"000000000",
  6549=>"111110111",
  6550=>"111110110",
  6551=>"111011000",
  6552=>"111111111",
  6553=>"111111001",
  6554=>"000000111",
  6555=>"111111111",
  6556=>"100100111",
  6557=>"011011111",
  6558=>"001001001",
  6559=>"110111110",
  6560=>"111111111",
  6561=>"000000010",
  6562=>"110110011",
  6563=>"110110100",
  6564=>"000100111",
  6565=>"111111111",
  6566=>"110111010",
  6567=>"110000001",
  6568=>"000000000",
  6569=>"000000100",
  6570=>"010000000",
  6571=>"111011011",
  6572=>"111111101",
  6573=>"101111111",
  6574=>"011110110",
  6575=>"000000111",
  6576=>"111000000",
  6577=>"100100000",
  6578=>"001011011",
  6579=>"111111110",
  6580=>"000000000",
  6581=>"000000111",
  6582=>"000000111",
  6583=>"111001000",
  6584=>"111111111",
  6585=>"111111111",
  6586=>"000001001",
  6587=>"110111111",
  6588=>"111000000",
  6589=>"111111111",
  6590=>"000000000",
  6591=>"010010010",
  6592=>"000000000",
  6593=>"110000001",
  6594=>"000000000",
  6595=>"000100000",
  6596=>"000000000",
  6597=>"000010010",
  6598=>"001000100",
  6599=>"000000000",
  6600=>"111100111",
  6601=>"111111111",
  6602=>"000001111",
  6603=>"000000111",
  6604=>"111111111",
  6605=>"011011011",
  6606=>"110111101",
  6607=>"100000001",
  6608=>"111111000",
  6609=>"000100110",
  6610=>"011010000",
  6611=>"000111111",
  6612=>"100100111",
  6613=>"000011011",
  6614=>"001101100",
  6615=>"111111011",
  6616=>"000101001",
  6617=>"111111111",
  6618=>"000111101",
  6619=>"000111111",
  6620=>"011000000",
  6621=>"011000000",
  6622=>"110110110",
  6623=>"000010000",
  6624=>"000000000",
  6625=>"111001111",
  6626=>"011001001",
  6627=>"011001111",
  6628=>"000000111",
  6629=>"110110111",
  6630=>"000111110",
  6631=>"000100111",
  6632=>"000000001",
  6633=>"100100000",
  6634=>"100111111",
  6635=>"111000000",
  6636=>"111000011",
  6637=>"111111100",
  6638=>"001001001",
  6639=>"110110000",
  6640=>"111111111",
  6641=>"111000100",
  6642=>"111011011",
  6643=>"000000100",
  6644=>"110111111",
  6645=>"101111111",
  6646=>"000010110",
  6647=>"011111111",
  6648=>"000111111",
  6649=>"001100111",
  6650=>"011111111",
  6651=>"000110100",
  6652=>"011011011",
  6653=>"001000000",
  6654=>"000111111",
  6655=>"000000001",
  6656=>"000000000",
  6657=>"111001111",
  6658=>"000000001",
  6659=>"111011111",
  6660=>"000111111",
  6661=>"000000110",
  6662=>"111000000",
  6663=>"111100111",
  6664=>"000000000",
  6665=>"111000000",
  6666=>"110000000",
  6667=>"111111111",
  6668=>"000000110",
  6669=>"111011000",
  6670=>"001111111",
  6671=>"100111111",
  6672=>"111100000",
  6673=>"000000101",
  6674=>"110110110",
  6675=>"000000001",
  6676=>"100000000",
  6677=>"110110111",
  6678=>"100110111",
  6679=>"111111111",
  6680=>"110110111",
  6681=>"001000100",
  6682=>"100000000",
  6683=>"101111100",
  6684=>"000100111",
  6685=>"000110000",
  6686=>"000111111",
  6687=>"111111111",
  6688=>"101111101",
  6689=>"100100000",
  6690=>"010110100",
  6691=>"100100000",
  6692=>"111111111",
  6693=>"111000000",
  6694=>"000000100",
  6695=>"001000000",
  6696=>"000000000",
  6697=>"000000111",
  6698=>"000000000",
  6699=>"000001100",
  6700=>"000000100",
  6701=>"111011000",
  6702=>"110000000",
  6703=>"100000100",
  6704=>"111111000",
  6705=>"011011000",
  6706=>"111111111",
  6707=>"101101100",
  6708=>"001010111",
  6709=>"111111110",
  6710=>"111111111",
  6711=>"111000000",
  6712=>"011011111",
  6713=>"101001000",
  6714=>"000000000",
  6715=>"000000000",
  6716=>"111111111",
  6717=>"100111001",
  6718=>"011101100",
  6719=>"000000000",
  6720=>"110111111",
  6721=>"000100111",
  6722=>"111111111",
  6723=>"000000110",
  6724=>"111111111",
  6725=>"111111000",
  6726=>"111111011",
  6727=>"000000000",
  6728=>"001000000",
  6729=>"111100000",
  6730=>"001000100",
  6731=>"111010010",
  6732=>"001101111",
  6733=>"111111111",
  6734=>"111111111",
  6735=>"000000000",
  6736=>"000000000",
  6737=>"100100110",
  6738=>"111111110",
  6739=>"011110000",
  6740=>"000000000",
  6741=>"100000000",
  6742=>"000000100",
  6743=>"100000000",
  6744=>"111111111",
  6745=>"000110111",
  6746=>"111100000",
  6747=>"111111110",
  6748=>"000111111",
  6749=>"000000111",
  6750=>"000111111",
  6751=>"100000000",
  6752=>"110111111",
  6753=>"111101000",
  6754=>"110100111",
  6755=>"111001000",
  6756=>"000110000",
  6757=>"100000110",
  6758=>"100110110",
  6759=>"000111111",
  6760=>"000000000",
  6761=>"000000001",
  6762=>"101001111",
  6763=>"111111110",
  6764=>"111001000",
  6765=>"000000000",
  6766=>"000000111",
  6767=>"111111111",
  6768=>"111111111",
  6769=>"110001000",
  6770=>"000100110",
  6771=>"111100000",
  6772=>"111000000",
  6773=>"111110000",
  6774=>"000000111",
  6775=>"000001111",
  6776=>"001111100",
  6777=>"000000100",
  6778=>"000111000",
  6779=>"111111000",
  6780=>"110100000",
  6781=>"111001001",
  6782=>"000000000",
  6783=>"111111111",
  6784=>"110100000",
  6785=>"000100011",
  6786=>"010000010",
  6787=>"001111111",
  6788=>"100110111",
  6789=>"100000000",
  6790=>"100110111",
  6791=>"111111000",
  6792=>"111111011",
  6793=>"100000111",
  6794=>"111001000",
  6795=>"111100000",
  6796=>"010000110",
  6797=>"001000000",
  6798=>"111111000",
  6799=>"000000000",
  6800=>"000000100",
  6801=>"001101000",
  6802=>"000000000",
  6803=>"111111111",
  6804=>"000110110",
  6805=>"000000110",
  6806=>"111000000",
  6807=>"000000000",
  6808=>"001000100",
  6809=>"100010010",
  6810=>"111111111",
  6811=>"111111000",
  6812=>"111111110",
  6813=>"111111000",
  6814=>"001001000",
  6815=>"000000111",
  6816=>"111111100",
  6817=>"011000000",
  6818=>"111010110",
  6819=>"111111111",
  6820=>"000111111",
  6821=>"111010100",
  6822=>"000000000",
  6823=>"100100011",
  6824=>"000000111",
  6825=>"000101111",
  6826=>"111111010",
  6827=>"000000000",
  6828=>"111001011",
  6829=>"111110100",
  6830=>"000111111",
  6831=>"011100110",
  6832=>"000000000",
  6833=>"111111011",
  6834=>"011101001",
  6835=>"000000001",
  6836=>"110100100",
  6837=>"001111111",
  6838=>"111111001",
  6839=>"011111111",
  6840=>"000000000",
  6841=>"000001111",
  6842=>"011001001",
  6843=>"101000100",
  6844=>"101100100",
  6845=>"111100111",
  6846=>"000000000",
  6847=>"101100110",
  6848=>"111111000",
  6849=>"100110000",
  6850=>"100110001",
  6851=>"000111111",
  6852=>"111111111",
  6853=>"101001111",
  6854=>"011000000",
  6855=>"111111000",
  6856=>"000110010",
  6857=>"000000001",
  6858=>"100100000",
  6859=>"110101101",
  6860=>"111000000",
  6861=>"010000000",
  6862=>"000000111",
  6863=>"000000000",
  6864=>"000000000",
  6865=>"000111111",
  6866=>"001000000",
  6867=>"000000000",
  6868=>"000000001",
  6869=>"001001000",
  6870=>"111111111",
  6871=>"000000100",
  6872=>"000111111",
  6873=>"000111000",
  6874=>"000000000",
  6875=>"111000000",
  6876=>"000000000",
  6877=>"000000000",
  6878=>"000111111",
  6879=>"000000100",
  6880=>"110110000",
  6881=>"000110000",
  6882=>"110000111",
  6883=>"111111100",
  6884=>"101111111",
  6885=>"110100100",
  6886=>"000000000",
  6887=>"101101011",
  6888=>"111111111",
  6889=>"100100001",
  6890=>"011111000",
  6891=>"100000011",
  6892=>"001001111",
  6893=>"000000000",
  6894=>"111001111",
  6895=>"101000000",
  6896=>"010000101",
  6897=>"000000000",
  6898=>"100111111",
  6899=>"000100100",
  6900=>"111000000",
  6901=>"111111000",
  6902=>"011000111",
  6903=>"111111111",
  6904=>"011010000",
  6905=>"111111111",
  6906=>"111100000",
  6907=>"111111011",
  6908=>"001111101",
  6909=>"110100111",
  6910=>"000001001",
  6911=>"000000101",
  6912=>"000000000",
  6913=>"011111111",
  6914=>"111000000",
  6915=>"000111100",
  6916=>"100000000",
  6917=>"111111111",
  6918=>"000000000",
  6919=>"000000000",
  6920=>"000000000",
  6921=>"011000000",
  6922=>"111110110",
  6923=>"111111110",
  6924=>"101000000",
  6925=>"101101000",
  6926=>"100001000",
  6927=>"000011111",
  6928=>"000111001",
  6929=>"000000000",
  6930=>"000000000",
  6931=>"010000011",
  6932=>"010110011",
  6933=>"100000000",
  6934=>"110110110",
  6935=>"000101111",
  6936=>"000000000",
  6937=>"111001001",
  6938=>"000000000",
  6939=>"000000111",
  6940=>"111111011",
  6941=>"000111100",
  6942=>"000000000",
  6943=>"000000001",
  6944=>"011001000",
  6945=>"101111111",
  6946=>"111111111",
  6947=>"001011111",
  6948=>"010000000",
  6949=>"111111110",
  6950=>"100101000",
  6951=>"011011111",
  6952=>"000000000",
  6953=>"111011111",
  6954=>"011000000",
  6955=>"000111100",
  6956=>"000000110",
  6957=>"111000000",
  6958=>"001000010",
  6959=>"000000111",
  6960=>"111111000",
  6961=>"111000000",
  6962=>"000000111",
  6963=>"111110100",
  6964=>"000000100",
  6965=>"000111001",
  6966=>"111111000",
  6967=>"111111100",
  6968=>"111111100",
  6969=>"111000011",
  6970=>"000000000",
  6971=>"111111001",
  6972=>"000100101",
  6973=>"111111110",
  6974=>"000000101",
  6975=>"000000000",
  6976=>"011001000",
  6977=>"000000100",
  6978=>"111100000",
  6979=>"000000111",
  6980=>"100000000",
  6981=>"101111000",
  6982=>"000000000",
  6983=>"111111100",
  6984=>"100000111",
  6985=>"001000011",
  6986=>"011001000",
  6987=>"100101100",
  6988=>"000000000",
  6989=>"111000000",
  6990=>"111111000",
  6991=>"000000000",
  6992=>"001101101",
  6993=>"000000000",
  6994=>"111100110",
  6995=>"001101111",
  6996=>"001111111",
  6997=>"111111111",
  6998=>"000000000",
  6999=>"100000100",
  7000=>"000111110",
  7001=>"011001001",
  7002=>"000011000",
  7003=>"111111100",
  7004=>"100100000",
  7005=>"001000000",
  7006=>"001111111",
  7007=>"000001111",
  7008=>"000000000",
  7009=>"000000000",
  7010=>"001001101",
  7011=>"000000000",
  7012=>"000000111",
  7013=>"111010000",
  7014=>"111010100",
  7015=>"111110111",
  7016=>"000100111",
  7017=>"000110111",
  7018=>"111111111",
  7019=>"110000100",
  7020=>"010010111",
  7021=>"000000100",
  7022=>"000011011",
  7023=>"011011000",
  7024=>"111000100",
  7025=>"111111000",
  7026=>"000000111",
  7027=>"001011011",
  7028=>"000111111",
  7029=>"000000000",
  7030=>"110000111",
  7031=>"001010000",
  7032=>"111000000",
  7033=>"111101001",
  7034=>"101000000",
  7035=>"001101011",
  7036=>"000001111",
  7037=>"000000001",
  7038=>"000111111",
  7039=>"111111111",
  7040=>"110110000",
  7041=>"000000100",
  7042=>"111111000",
  7043=>"000000110",
  7044=>"111111000",
  7045=>"100110001",
  7046=>"111111011",
  7047=>"111111111",
  7048=>"000000000",
  7049=>"100000010",
  7050=>"101000100",
  7051=>"000011000",
  7052=>"111111010",
  7053=>"111100100",
  7054=>"000000000",
  7055=>"001000000",
  7056=>"000101101",
  7057=>"000000011",
  7058=>"000000000",
  7059=>"000000111",
  7060=>"011111111",
  7061=>"010010000",
  7062=>"110110110",
  7063=>"111111000",
  7064=>"111111111",
  7065=>"111111000",
  7066=>"111001000",
  7067=>"111011000",
  7068=>"000000111",
  7069=>"111101111",
  7070=>"011000000",
  7071=>"111111111",
  7072=>"100111111",
  7073=>"111110100",
  7074=>"100100000",
  7075=>"000000000",
  7076=>"010111100",
  7077=>"111111000",
  7078=>"110111111",
  7079=>"000000111",
  7080=>"110000110",
  7081=>"001000000",
  7082=>"100000111",
  7083=>"000000000",
  7084=>"000000101",
  7085=>"111111000",
  7086=>"111111010",
  7087=>"000000000",
  7088=>"111111110",
  7089=>"000000001",
  7090=>"000011000",
  7091=>"100100100",
  7092=>"000100111",
  7093=>"111111111",
  7094=>"010011000",
  7095=>"111111111",
  7096=>"111111110",
  7097=>"000000100",
  7098=>"111111000",
  7099=>"000000000",
  7100=>"111100100",
  7101=>"111111100",
  7102=>"000001001",
  7103=>"101100111",
  7104=>"000000000",
  7105=>"111100111",
  7106=>"111000000",
  7107=>"111111111",
  7108=>"100100000",
  7109=>"001001011",
  7110=>"100011011",
  7111=>"111111111",
  7112=>"001001100",
  7113=>"111111100",
  7114=>"101100110",
  7115=>"111111010",
  7116=>"111111000",
  7117=>"111111111",
  7118=>"111011000",
  7119=>"000000001",
  7120=>"000111111",
  7121=>"000000110",
  7122=>"000111111",
  7123=>"111000010",
  7124=>"111111111",
  7125=>"000001000",
  7126=>"101111100",
  7127=>"000110111",
  7128=>"111111100",
  7129=>"111111111",
  7130=>"111110110",
  7131=>"111101111",
  7132=>"110000000",
  7133=>"111111011",
  7134=>"111011000",
  7135=>"111101111",
  7136=>"000000000",
  7137=>"000000000",
  7138=>"001000100",
  7139=>"000000011",
  7140=>"000000000",
  7141=>"111110111",
  7142=>"111100000",
  7143=>"111000000",
  7144=>"011111111",
  7145=>"100111111",
  7146=>"111110101",
  7147=>"001000000",
  7148=>"000111001",
  7149=>"110110111",
  7150=>"000000111",
  7151=>"111111100",
  7152=>"011000000",
  7153=>"100111111",
  7154=>"001011001",
  7155=>"000111111",
  7156=>"000100000",
  7157=>"111111111",
  7158=>"000001001",
  7159=>"111001111",
  7160=>"110111111",
  7161=>"110110000",
  7162=>"000000110",
  7163=>"111000000",
  7164=>"111001001",
  7165=>"110111111",
  7166=>"111111111",
  7167=>"111100000",
  7168=>"011000000",
  7169=>"000000000",
  7170=>"111111111",
  7171=>"000000000",
  7172=>"110111001",
  7173=>"000000001",
  7174=>"111010010",
  7175=>"000111111",
  7176=>"111100000",
  7177=>"110111110",
  7178=>"100101101",
  7179=>"000000001",
  7180=>"111111111",
  7181=>"111111111",
  7182=>"100111111",
  7183=>"110000000",
  7184=>"111111111",
  7185=>"001000000",
  7186=>"011000100",
  7187=>"000111111",
  7188=>"100000000",
  7189=>"111101001",
  7190=>"111110111",
  7191=>"111111111",
  7192=>"011010110",
  7193=>"000000110",
  7194=>"111000000",
  7195=>"110110100",
  7196=>"000001000",
  7197=>"111111000",
  7198=>"111011111",
  7199=>"100000000",
  7200=>"000001001",
  7201=>"000011011",
  7202=>"100001011",
  7203=>"110100000",
  7204=>"100000000",
  7205=>"111000000",
  7206=>"100100111",
  7207=>"000110110",
  7208=>"010111110",
  7209=>"010000000",
  7210=>"000000000",
  7211=>"000000000",
  7212=>"000000000",
  7213=>"000000000",
  7214=>"000000000",
  7215=>"111000000",
  7216=>"010111000",
  7217=>"000000000",
  7218=>"110110110",
  7219=>"100111111",
  7220=>"101101111",
  7221=>"110011111",
  7222=>"011010111",
  7223=>"110111111",
  7224=>"000000011",
  7225=>"000001000",
  7226=>"001001111",
  7227=>"111000000",
  7228=>"000000000",
  7229=>"110110110",
  7230=>"010010000",
  7231=>"000100111",
  7232=>"111111100",
  7233=>"000000100",
  7234=>"000001111",
  7235=>"000001011",
  7236=>"100000000",
  7237=>"011000000",
  7238=>"111010000",
  7239=>"111111111",
  7240=>"100110010",
  7241=>"000000000",
  7242=>"001001111",
  7243=>"000110011",
  7244=>"000000111",
  7245=>"111001111",
  7246=>"011001000",
  7247=>"111000000",
  7248=>"000000001",
  7249=>"111000111",
  7250=>"110010011",
  7251=>"011000000",
  7252=>"111111111",
  7253=>"110110110",
  7254=>"000110000",
  7255=>"000000111",
  7256=>"000010000",
  7257=>"000000101",
  7258=>"111110111",
  7259=>"111101111",
  7260=>"110110110",
  7261=>"000100000",
  7262=>"000111100",
  7263=>"000000000",
  7264=>"111111100",
  7265=>"011010000",
  7266=>"110110010",
  7267=>"111111110",
  7268=>"000100110",
  7269=>"000111111",
  7270=>"100100111",
  7271=>"000000000",
  7272=>"001001000",
  7273=>"111111111",
  7274=>"000000000",
  7275=>"111000000",
  7276=>"000011000",
  7277=>"110100000",
  7278=>"111110110",
  7279=>"100000000",
  7280=>"000101000",
  7281=>"001111111",
  7282=>"101001111",
  7283=>"000000111",
  7284=>"000111111",
  7285=>"111111001",
  7286=>"111111100",
  7287=>"111110111",
  7288=>"000000110",
  7289=>"000000000",
  7290=>"000000100",
  7291=>"000000110",
  7292=>"100100100",
  7293=>"110011111",
  7294=>"110111000",
  7295=>"100100100",
  7296=>"000000001",
  7297=>"110111111",
  7298=>"111111111",
  7299=>"100111010",
  7300=>"110110000",
  7301=>"000000000",
  7302=>"000000100",
  7303=>"000000011",
  7304=>"011111111",
  7305=>"000000001",
  7306=>"000010000",
  7307=>"111111111",
  7308=>"110111111",
  7309=>"111111000",
  7310=>"100111111",
  7311=>"111100000",
  7312=>"010000111",
  7313=>"111101101",
  7314=>"000000000",
  7315=>"011011111",
  7316=>"111110000",
  7317=>"111111111",
  7318=>"000000000",
  7319=>"101000000",
  7320=>"001101111",
  7321=>"010110001",
  7322=>"000000111",
  7323=>"000000000",
  7324=>"111111100",
  7325=>"000000001",
  7326=>"000110111",
  7327=>"000001011",
  7328=>"100000000",
  7329=>"000101111",
  7330=>"111111111",
  7331=>"001001000",
  7332=>"110100001",
  7333=>"110011000",
  7334=>"111111111",
  7335=>"111101111",
  7336=>"000000000",
  7337=>"000000110",
  7338=>"000000000",
  7339=>"011001000",
  7340=>"000111110",
  7341=>"110111111",
  7342=>"000000111",
  7343=>"000000001",
  7344=>"000000111",
  7345=>"000000000",
  7346=>"111111111",
  7347=>"000000000",
  7348=>"000110000",
  7349=>"110111101",
  7350=>"100000111",
  7351=>"111000010",
  7352=>"111000001",
  7353=>"000100111",
  7354=>"110011010",
  7355=>"100001001",
  7356=>"000111000",
  7357=>"000100110",
  7358=>"111110110",
  7359=>"101011000",
  7360=>"111000000",
  7361=>"110110000",
  7362=>"011011011",
  7363=>"111000111",
  7364=>"000000000",
  7365=>"111000001",
  7366=>"001000000",
  7367=>"000001011",
  7368=>"110001111",
  7369=>"111111011",
  7370=>"111011011",
  7371=>"111111111",
  7372=>"101111011",
  7373=>"110111111",
  7374=>"000000000",
  7375=>"110000000",
  7376=>"111110101",
  7377=>"111111000",
  7378=>"111000000",
  7379=>"110110011",
  7380=>"111111111",
  7381=>"111111111",
  7382=>"000111111",
  7383=>"000010110",
  7384=>"000000010",
  7385=>"000111111",
  7386=>"111000000",
  7387=>"011110100",
  7388=>"000001111",
  7389=>"011000000",
  7390=>"000000000",
  7391=>"111011000",
  7392=>"000111111",
  7393=>"101000000",
  7394=>"000111111",
  7395=>"000000000",
  7396=>"100110110",
  7397=>"011011011",
  7398=>"110000000",
  7399=>"110111011",
  7400=>"000000000",
  7401=>"000111111",
  7402=>"110100000",
  7403=>"010111111",
  7404=>"000011011",
  7405=>"000110111",
  7406=>"000011111",
  7407=>"000001000",
  7408=>"110110000",
  7409=>"111100111",
  7410=>"000000000",
  7411=>"000001110",
  7412=>"110001000",
  7413=>"001000000",
  7414=>"111000100",
  7415=>"010000000",
  7416=>"011011111",
  7417=>"111000000",
  7418=>"000100101",
  7419=>"100100000",
  7420=>"110010110",
  7421=>"001011111",
  7422=>"010110110",
  7423=>"111111111",
  7424=>"111111111",
  7425=>"100111110",
  7426=>"000011111",
  7427=>"110111001",
  7428=>"100100000",
  7429=>"101100110",
  7430=>"110110000",
  7431=>"000011011",
  7432=>"111111000",
  7433=>"110111001",
  7434=>"111111111",
  7435=>"010111000",
  7436=>"111000111",
  7437=>"000110010",
  7438=>"111111111",
  7439=>"000100000",
  7440=>"110110110",
  7441=>"011111111",
  7442=>"000000001",
  7443=>"000000000",
  7444=>"110110110",
  7445=>"001000000",
  7446=>"100001111",
  7447=>"001111111",
  7448=>"100100111",
  7449=>"111111111",
  7450=>"001111111",
  7451=>"111110111",
  7452=>"100111111",
  7453=>"000000000",
  7454=>"000000111",
  7455=>"111100001",
  7456=>"100000111",
  7457=>"101111111",
  7458=>"000000011",
  7459=>"111111111",
  7460=>"000011111",
  7461=>"111100111",
  7462=>"001000000",
  7463=>"110100000",
  7464=>"000001111",
  7465=>"011111111",
  7466=>"000000001",
  7467=>"001000001",
  7468=>"100000111",
  7469=>"000000110",
  7470=>"111111000",
  7471=>"010011011",
  7472=>"000000000",
  7473=>"000000001",
  7474=>"000001010",
  7475=>"010000000",
  7476=>"000110111",
  7477=>"001000000",
  7478=>"000000000",
  7479=>"000001011",
  7480=>"001101101",
  7481=>"101111111",
  7482=>"111000000",
  7483=>"111111111",
  7484=>"000100100",
  7485=>"001111111",
  7486=>"110011000",
  7487=>"110111110",
  7488=>"011111011",
  7489=>"111110110",
  7490=>"000001000",
  7491=>"101101000",
  7492=>"110100111",
  7493=>"000000000",
  7494=>"000000000",
  7495=>"111111110",
  7496=>"000111111",
  7497=>"011000000",
  7498=>"111111101",
  7499=>"110100000",
  7500=>"100000101",
  7501=>"000000000",
  7502=>"000000000",
  7503=>"001010111",
  7504=>"011011110",
  7505=>"110110110",
  7506=>"000010111",
  7507=>"110010000",
  7508=>"111101001",
  7509=>"000000100",
  7510=>"111000110",
  7511=>"000000000",
  7512=>"000000100",
  7513=>"111111110",
  7514=>"001110110",
  7515=>"001111011",
  7516=>"000000000",
  7517=>"101111111",
  7518=>"011011011",
  7519=>"000001111",
  7520=>"110000010",
  7521=>"111110110",
  7522=>"111110110",
  7523=>"000000000",
  7524=>"110110110",
  7525=>"100000001",
  7526=>"011111111",
  7527=>"000001001",
  7528=>"111001111",
  7529=>"000000000",
  7530=>"111111000",
  7531=>"000000001",
  7532=>"000000001",
  7533=>"000100100",
  7534=>"111011011",
  7535=>"000000000",
  7536=>"000000100",
  7537=>"000111111",
  7538=>"111111111",
  7539=>"011111011",
  7540=>"111111000",
  7541=>"100000001",
  7542=>"000010000",
  7543=>"100101111",
  7544=>"000000100",
  7545=>"000111100",
  7546=>"111111110",
  7547=>"110001011",
  7548=>"100000000",
  7549=>"100100000",
  7550=>"110111111",
  7551=>"000000000",
  7552=>"111111111",
  7553=>"110110000",
  7554=>"110110110",
  7555=>"000000000",
  7556=>"110111111",
  7557=>"111111100",
  7558=>"000000111",
  7559=>"111110000",
  7560=>"000000111",
  7561=>"000000000",
  7562=>"000000000",
  7563=>"100111111",
  7564=>"111111111",
  7565=>"111111111",
  7566=>"100100100",
  7567=>"111111111",
  7568=>"000100111",
  7569=>"111111111",
  7570=>"111000100",
  7571=>"110110000",
  7572=>"000111111",
  7573=>"110000000",
  7574=>"110000000",
  7575=>"000001110",
  7576=>"010000001",
  7577=>"010111111",
  7578=>"000000000",
  7579=>"111111011",
  7580=>"111111010",
  7581=>"000000001",
  7582=>"111111111",
  7583=>"000000000",
  7584=>"110000010",
  7585=>"000010110",
  7586=>"011100110",
  7587=>"000111111",
  7588=>"000110000",
  7589=>"101100001",
  7590=>"000100000",
  7591=>"000000000",
  7592=>"101111001",
  7593=>"000000001",
  7594=>"000000111",
  7595=>"111001011",
  7596=>"000000111",
  7597=>"110110000",
  7598=>"000000110",
  7599=>"111111111",
  7600=>"110000000",
  7601=>"111101000",
  7602=>"111100001",
  7603=>"000001000",
  7604=>"111111001",
  7605=>"111111111",
  7606=>"000000100",
  7607=>"111011000",
  7608=>"100011011",
  7609=>"110110111",
  7610=>"011001001",
  7611=>"111000000",
  7612=>"000000001",
  7613=>"000000111",
  7614=>"010111111",
  7615=>"100101100",
  7616=>"000111111",
  7617=>"011001001",
  7618=>"000000000",
  7619=>"000000000",
  7620=>"110111111",
  7621=>"000111111",
  7622=>"001000011",
  7623=>"001100111",
  7624=>"000000100",
  7625=>"111111100",
  7626=>"000000000",
  7627=>"001111111",
  7628=>"001111111",
  7629=>"111111111",
  7630=>"111111111",
  7631=>"111000000",
  7632=>"000000111",
  7633=>"111001111",
  7634=>"100000000",
  7635=>"100111111",
  7636=>"110111111",
  7637=>"000110100",
  7638=>"000100111",
  7639=>"111110111",
  7640=>"000111000",
  7641=>"101101111",
  7642=>"110000000",
  7643=>"000000100",
  7644=>"111011111",
  7645=>"001001001",
  7646=>"000000000",
  7647=>"110111111",
  7648=>"111000000",
  7649=>"111111111",
  7650=>"110100000",
  7651=>"000000100",
  7652=>"000000000",
  7653=>"000011001",
  7654=>"001100111",
  7655=>"000000000",
  7656=>"001101111",
  7657=>"111111100",
  7658=>"000000000",
  7659=>"111111111",
  7660=>"111111111",
  7661=>"011100111",
  7662=>"111111111",
  7663=>"011111001",
  7664=>"011000000",
  7665=>"111000000",
  7666=>"000000110",
  7667=>"000000101",
  7668=>"100111111",
  7669=>"100000100",
  7670=>"000000010",
  7671=>"111100000",
  7672=>"111000000",
  7673=>"011000100",
  7674=>"111111111",
  7675=>"011111111",
  7676=>"000001000",
  7677=>"010000000",
  7678=>"000100000",
  7679=>"000011001",
  7680=>"000001110",
  7681=>"000000000",
  7682=>"000000000",
  7683=>"111111100",
  7684=>"011001011",
  7685=>"110100100",
  7686=>"000000001",
  7687=>"000000100",
  7688=>"011011001",
  7689=>"000000000",
  7690=>"111100001",
  7691=>"000000000",
  7692=>"000100111",
  7693=>"111000000",
  7694=>"100000100",
  7695=>"000000000",
  7696=>"001000001",
  7697=>"000010000",
  7698=>"111111111",
  7699=>"001001011",
  7700=>"111111111",
  7701=>"001001111",
  7702=>"101110111",
  7703=>"111111101",
  7704=>"110110101",
  7705=>"000000100",
  7706=>"000000000",
  7707=>"111111001",
  7708=>"001001111",
  7709=>"001000000",
  7710=>"000000000",
  7711=>"110110000",
  7712=>"101111011",
  7713=>"111111111",
  7714=>"111111111",
  7715=>"111111111",
  7716=>"101000000",
  7717=>"111111111",
  7718=>"000000000",
  7719=>"000001000",
  7720=>"111100001",
  7721=>"000000000",
  7722=>"111111011",
  7723=>"000000000",
  7724=>"000100111",
  7725=>"000000000",
  7726=>"000000000",
  7727=>"000010100",
  7728=>"101101111",
  7729=>"111111111",
  7730=>"001011001",
  7731=>"010110110",
  7732=>"000000000",
  7733=>"111000001",
  7734=>"001000000",
  7735=>"101101100",
  7736=>"000000000",
  7737=>"000000111",
  7738=>"111110110",
  7739=>"000110000",
  7740=>"000000000",
  7741=>"111111001",
  7742=>"000001001",
  7743=>"001000001",
  7744=>"010100100",
  7745=>"000110110",
  7746=>"110110111",
  7747=>"110110010",
  7748=>"110110010",
  7749=>"000100100",
  7750=>"000000000",
  7751=>"111111111",
  7752=>"001011001",
  7753=>"000000001",
  7754=>"111111111",
  7755=>"111111000",
  7756=>"110000000",
  7757=>"111110010",
  7758=>"000000000",
  7759=>"110000000",
  7760=>"101000000",
  7761=>"100100111",
  7762=>"000000000",
  7763=>"110111111",
  7764=>"000000000",
  7765=>"111111111",
  7766=>"111110011",
  7767=>"111111001",
  7768=>"011101100",
  7769=>"001000101",
  7770=>"110110000",
  7771=>"111111010",
  7772=>"111001000",
  7773=>"110111011",
  7774=>"000010000",
  7775=>"111111111",
  7776=>"010111100",
  7777=>"100001100",
  7778=>"111111111",
  7779=>"011000000",
  7780=>"111111000",
  7781=>"100000001",
  7782=>"000000010",
  7783=>"001000101",
  7784=>"000000000",
  7785=>"111111111",
  7786=>"100000000",
  7787=>"110010000",
  7788=>"000000001",
  7789=>"000000101",
  7790=>"110111010",
  7791=>"111111111",
  7792=>"000001101",
  7793=>"101001001",
  7794=>"100000011",
  7795=>"000000100",
  7796=>"000000000",
  7797=>"000000000",
  7798=>"000001110",
  7799=>"000000000",
  7800=>"110001001",
  7801=>"000000001",
  7802=>"111111111",
  7803=>"100100111",
  7804=>"110100000",
  7805=>"111001001",
  7806=>"111111111",
  7807=>"111111111",
  7808=>"000101111",
  7809=>"111111111",
  7810=>"000010010",
  7811=>"001001101",
  7812=>"000000101",
  7813=>"111111111",
  7814=>"100100000",
  7815=>"111111000",
  7816=>"111111000",
  7817=>"000000000",
  7818=>"100000000",
  7819=>"111111011",
  7820=>"000000001",
  7821=>"111100111",
  7822=>"101000000",
  7823=>"111111111",
  7824=>"110111111",
  7825=>"111111111",
  7826=>"000110101",
  7827=>"010001011",
  7828=>"111111000",
  7829=>"101111111",
  7830=>"110111011",
  7831=>"001001000",
  7832=>"001000101",
  7833=>"000100111",
  7834=>"100101101",
  7835=>"010010000",
  7836=>"110000000",
  7837=>"100111001",
  7838=>"001111010",
  7839=>"010111000",
  7840=>"000000101",
  7841=>"000000000",
  7842=>"000100101",
  7843=>"111111111",
  7844=>"001001001",
  7845=>"000000110",
  7846=>"000000000",
  7847=>"100100000",
  7848=>"111111111",
  7849=>"001101101",
  7850=>"111000111",
  7851=>"111111011",
  7852=>"111111111",
  7853=>"100100001",
  7854=>"000000001",
  7855=>"000000000",
  7856=>"111111111",
  7857=>"000001011",
  7858=>"111111111",
  7859=>"010011010",
  7860=>"110111111",
  7861=>"000100111",
  7862=>"111001001",
  7863=>"000000111",
  7864=>"000000001",
  7865=>"000000000",
  7866=>"001011111",
  7867=>"111111010",
  7868=>"101101111",
  7869=>"001000000",
  7870=>"111111111",
  7871=>"110111010",
  7872=>"111100111",
  7873=>"000000001",
  7874=>"000000100",
  7875=>"111101101",
  7876=>"111111111",
  7877=>"111111111",
  7878=>"110100000",
  7879=>"000000001",
  7880=>"000011000",
  7881=>"000000111",
  7882=>"101001001",
  7883=>"111011001",
  7884=>"110111111",
  7885=>"000010000",
  7886=>"010111101",
  7887=>"100000011",
  7888=>"000000000",
  7889=>"110000000",
  7890=>"100100100",
  7891=>"010000000",
  7892=>"000101111",
  7893=>"111111111",
  7894=>"000000111",
  7895=>"110000000",
  7896=>"000000001",
  7897=>"100111011",
  7898=>"000000000",
  7899=>"000000000",
  7900=>"111110000",
  7901=>"111001001",
  7902=>"000010101",
  7903=>"000000000",
  7904=>"111000111",
  7905=>"000000000",
  7906=>"011111111",
  7907=>"111111111",
  7908=>"000000000",
  7909=>"111111101",
  7910=>"111111010",
  7911=>"100111111",
  7912=>"000000010",
  7913=>"000000000",
  7914=>"000001010",
  7915=>"111111111",
  7916=>"111111111",
  7917=>"000000000",
  7918=>"000000000",
  7919=>"111111100",
  7920=>"011011000",
  7921=>"011111011",
  7922=>"001111011",
  7923=>"111000100",
  7924=>"000000000",
  7925=>"110111111",
  7926=>"000000100",
  7927=>"111110111",
  7928=>"000001001",
  7929=>"000000001",
  7930=>"100111111",
  7931=>"110111000",
  7932=>"001001111",
  7933=>"000101111",
  7934=>"111111011",
  7935=>"000000000",
  7936=>"111001001",
  7937=>"100101001",
  7938=>"000000000",
  7939=>"000000101",
  7940=>"000000000",
  7941=>"111001000",
  7942=>"001111111",
  7943=>"010011000",
  7944=>"001001001",
  7945=>"000000000",
  7946=>"111111000",
  7947=>"000000000",
  7948=>"111111101",
  7949=>"000000000",
  7950=>"111111111",
  7951=>"000100110",
  7952=>"111111111",
  7953=>"101101100",
  7954=>"101001001",
  7955=>"000010000",
  7956=>"001000111",
  7957=>"000000001",
  7958=>"111111100",
  7959=>"000000111",
  7960=>"001011001",
  7961=>"000010011",
  7962=>"000000000",
  7963=>"111111000",
  7964=>"100100100",
  7965=>"100000000",
  7966=>"111100000",
  7967=>"000111001",
  7968=>"101100101",
  7969=>"010111111",
  7970=>"111100100",
  7971=>"100000101",
  7972=>"100000000",
  7973=>"111111111",
  7974=>"100001101",
  7975=>"000000000",
  7976=>"111101111",
  7977=>"010111011",
  7978=>"111101101",
  7979=>"100000111",
  7980=>"111111000",
  7981=>"001001001",
  7982=>"111111110",
  7983=>"000000000",
  7984=>"000000000",
  7985=>"000000001",
  7986=>"111010000",
  7987=>"000000010",
  7988=>"110100000",
  7989=>"000000000",
  7990=>"000000000",
  7991=>"111011001",
  7992=>"000000000",
  7993=>"000001101",
  7994=>"111001000",
  7995=>"000000100",
  7996=>"000001011",
  7997=>"111111011",
  7998=>"000000000",
  7999=>"100001000",
  8000=>"000101101",
  8001=>"000111111",
  8002=>"101001001",
  8003=>"111111111",
  8004=>"001101111",
  8005=>"010111111",
  8006=>"111111101",
  8007=>"001001111",
  8008=>"011000000",
  8009=>"010010000",
  8010=>"100110001",
  8011=>"001001011",
  8012=>"101000000",
  8013=>"111111000",
  8014=>"000000000",
  8015=>"001001001",
  8016=>"111111011",
  8017=>"000110110",
  8018=>"111111011",
  8019=>"000000001",
  8020=>"010110000",
  8021=>"001001001",
  8022=>"010010010",
  8023=>"111111111",
  8024=>"111100111",
  8025=>"010011010",
  8026=>"000000000",
  8027=>"000111111",
  8028=>"000000000",
  8029=>"010110010",
  8030=>"000000000",
  8031=>"000000001",
  8032=>"111111111",
  8033=>"101101101",
  8034=>"000000100",
  8035=>"111011000",
  8036=>"110110001",
  8037=>"111100111",
  8038=>"000000100",
  8039=>"100100110",
  8040=>"000000110",
  8041=>"010111111",
  8042=>"100100000",
  8043=>"110111111",
  8044=>"000000000",
  8045=>"011000000",
  8046=>"001000101",
  8047=>"000000000",
  8048=>"111101000",
  8049=>"111110111",
  8050=>"000000000",
  8051=>"111110111",
  8052=>"010110110",
  8053=>"110000000",
  8054=>"000000001",
  8055=>"000110000",
  8056=>"111111010",
  8057=>"110111111",
  8058=>"111111111",
  8059=>"110111010",
  8060=>"100000100",
  8061=>"110111111",
  8062=>"101111111",
  8063=>"111000101",
  8064=>"011010001",
  8065=>"011001101",
  8066=>"011011001",
  8067=>"111111110",
  8068=>"011011111",
  8069=>"000000000",
  8070=>"100000000",
  8071=>"111110111",
  8072=>"000000000",
  8073=>"011111000",
  8074=>"000000000",
  8075=>"110000000",
  8076=>"111111111",
  8077=>"100101110",
  8078=>"100001001",
  8079=>"010101011",
  8080=>"000000000",
  8081=>"100000000",
  8082=>"111111001",
  8083=>"001000111",
  8084=>"000110111",
  8085=>"010110000",
  8086=>"011001111",
  8087=>"000000011",
  8088=>"111111111",
  8089=>"111111111",
  8090=>"101000111",
  8091=>"011000001",
  8092=>"111111111",
  8093=>"111111101",
  8094=>"000000000",
  8095=>"000000000",
  8096=>"110110110",
  8097=>"100100000",
  8098=>"111101000",
  8099=>"010000000",
  8100=>"001001111",
  8101=>"010010110",
  8102=>"001001111",
  8103=>"000111111",
  8104=>"000000000",
  8105=>"000000000",
  8106=>"000000111",
  8107=>"111001101",
  8108=>"000000000",
  8109=>"000000001",
  8110=>"000000101",
  8111=>"111111011",
  8112=>"000000000",
  8113=>"000000101",
  8114=>"000001001",
  8115=>"111111111",
  8116=>"001000000",
  8117=>"111101111",
  8118=>"000000001",
  8119=>"001001001",
  8120=>"110110111",
  8121=>"111111111",
  8122=>"000000101",
  8123=>"101101101",
  8124=>"110111111",
  8125=>"100101111",
  8126=>"111100101",
  8127=>"110111000",
  8128=>"111111111",
  8129=>"000000001",
  8130=>"111111110",
  8131=>"101001111",
  8132=>"110011001",
  8133=>"101001001",
  8134=>"000000111",
  8135=>"100000000",
  8136=>"111100000",
  8137=>"111111100",
  8138=>"100000000",
  8139=>"110110111",
  8140=>"000000000",
  8141=>"110111111",
  8142=>"110000000",
  8143=>"000110110",
  8144=>"110100100",
  8145=>"111111111",
  8146=>"111001000",
  8147=>"111111111",
  8148=>"100100110",
  8149=>"111111000",
  8150=>"100111110",
  8151=>"110000000",
  8152=>"000001100",
  8153=>"111000000",
  8154=>"111111111",
  8155=>"000000111",
  8156=>"001001001",
  8157=>"110111001",
  8158=>"111111000",
  8159=>"100000000",
  8160=>"000000000",
  8161=>"111111111",
  8162=>"111001001",
  8163=>"000000000",
  8164=>"111011111",
  8165=>"001001000",
  8166=>"111101111",
  8167=>"000010110",
  8168=>"010011011",
  8169=>"000000101",
  8170=>"001001011",
  8171=>"110111111",
  8172=>"001111011",
  8173=>"100110110",
  8174=>"000001111",
  8175=>"110000000",
  8176=>"101101111",
  8177=>"000110111",
  8178=>"111111111",
  8179=>"011010000",
  8180=>"000001111",
  8181=>"111001100",
  8182=>"111111110",
  8183=>"100100001",
  8184=>"011111111",
  8185=>"101100001",
  8186=>"000000000",
  8187=>"000000000",
  8188=>"111011000",
  8189=>"111111110",
  8190=>"000000101",
  8191=>"000111111",
  8192=>"111111111",
  8193=>"000000000",
  8194=>"001001111",
  8195=>"000000000",
  8196=>"000000001",
  8197=>"001000011",
  8198=>"111100100",
  8199=>"000000000",
  8200=>"000000000",
  8201=>"111111111",
  8202=>"000000000",
  8203=>"111111111",
  8204=>"000000100",
  8205=>"001001000",
  8206=>"000000000",
  8207=>"111111111",
  8208=>"000000000",
  8209=>"111111111",
  8210=>"011000000",
  8211=>"111101111",
  8212=>"000110000",
  8213=>"000000111",
  8214=>"011000000",
  8215=>"001000010",
  8216=>"111111111",
  8217=>"001000000",
  8218=>"000000111",
  8219=>"100110000",
  8220=>"111110000",
  8221=>"000000100",
  8222=>"000000100",
  8223=>"100111111",
  8224=>"000000001",
  8225=>"110111111",
  8226=>"000000000",
  8227=>"100101001",
  8228=>"111111111",
  8229=>"111111000",
  8230=>"111111111",
  8231=>"111111111",
  8232=>"001111111",
  8233=>"000000011",
  8234=>"000000000",
  8235=>"000000000",
  8236=>"111111111",
  8237=>"000000100",
  8238=>"100100111",
  8239=>"110111110",
  8240=>"000000001",
  8241=>"111111111",
  8242=>"000000000",
  8243=>"000110001",
  8244=>"000000000",
  8245=>"001000000",
  8246=>"100100111",
  8247=>"111100000",
  8248=>"000000000",
  8249=>"000000000",
  8250=>"000000000",
  8251=>"101000000",
  8252=>"111111111",
  8253=>"110110110",
  8254=>"111111011",
  8255=>"011011000",
  8256=>"100110111",
  8257=>"100000000",
  8258=>"000011110",
  8259=>"100100111",
  8260=>"110111111",
  8261=>"010100000",
  8262=>"001001011",
  8263=>"111111111",
  8264=>"101111111",
  8265=>"101001110",
  8266=>"111111111",
  8267=>"111111111",
  8268=>"111111111",
  8269=>"011011010",
  8270=>"011011011",
  8271=>"010110111",
  8272=>"111111000",
  8273=>"000000000",
  8274=>"110111111",
  8275=>"010010000",
  8276=>"111111110",
  8277=>"000000000",
  8278=>"000000101",
  8279=>"111111100",
  8280=>"000000000",
  8281=>"111111111",
  8282=>"110111100",
  8283=>"111101111",
  8284=>"000010000",
  8285=>"111111111",
  8286=>"000000100",
  8287=>"111111111",
  8288=>"000000000",
  8289=>"011000000",
  8290=>"000000111",
  8291=>"011010111",
  8292=>"110110111",
  8293=>"111111111",
  8294=>"000000000",
  8295=>"000000000",
  8296=>"100111111",
  8297=>"000011011",
  8298=>"111110000",
  8299=>"000000000",
  8300=>"111110110",
  8301=>"111100111",
  8302=>"111111100",
  8303=>"110111111",
  8304=>"011011110",
  8305=>"000000000",
  8306=>"000000101",
  8307=>"000000110",
  8308=>"101001000",
  8309=>"111111111",
  8310=>"000000000",
  8311=>"001000000",
  8312=>"111111111",
  8313=>"111110100",
  8314=>"000000000",
  8315=>"000000000",
  8316=>"111110111",
  8317=>"000000000",
  8318=>"111100000",
  8319=>"111111111",
  8320=>"000000000",
  8321=>"100101100",
  8322=>"111111111",
  8323=>"000110110",
  8324=>"000000000",
  8325=>"000000000",
  8326=>"000000000",
  8327=>"000000000",
  8328=>"000010110",
  8329=>"000000000",
  8330=>"010000111",
  8331=>"000111111",
  8332=>"111111111",
  8333=>"000000111",
  8334=>"110110110",
  8335=>"011101111",
  8336=>"011111000",
  8337=>"111111111",
  8338=>"011111111",
  8339=>"111111111",
  8340=>"001010111",
  8341=>"000000000",
  8342=>"000000000",
  8343=>"000110000",
  8344=>"000000110",
  8345=>"111111111",
  8346=>"000011011",
  8347=>"100100100",
  8348=>"111111111",
  8349=>"000111011",
  8350=>"111111110",
  8351=>"111111111",
  8352=>"000000000",
  8353=>"011111111",
  8354=>"000001100",
  8355=>"111111111",
  8356=>"000000000",
  8357=>"010111110",
  8358=>"011111111",
  8359=>"000000001",
  8360=>"111111111",
  8361=>"001111011",
  8362=>"000000010",
  8363=>"000000000",
  8364=>"000000000",
  8365=>"000000111",
  8366=>"000000000",
  8367=>"111111000",
  8368=>"111111111",
  8369=>"011011111",
  8370=>"111111111",
  8371=>"000000000",
  8372=>"111111111",
  8373=>"100111111",
  8374=>"000000000",
  8375=>"000000000",
  8376=>"101111111",
  8377=>"000000000",
  8378=>"000100100",
  8379=>"110000000",
  8380=>"000000001",
  8381=>"111111111",
  8382=>"110011111",
  8383=>"101111111",
  8384=>"111110100",
  8385=>"111111011",
  8386=>"000000001",
  8387=>"000000000",
  8388=>"111111100",
  8389=>"111111011",
  8390=>"111111101",
  8391=>"000001111",
  8392=>"111111111",
  8393=>"111101111",
  8394=>"111111011",
  8395=>"111111111",
  8396=>"111111111",
  8397=>"111101001",
  8398=>"111111111",
  8399=>"000000000",
  8400=>"111111111",
  8401=>"000000000",
  8402=>"000111111",
  8403=>"111101111",
  8404=>"000000000",
  8405=>"000001001",
  8406=>"110110010",
  8407=>"110000000",
  8408=>"111111111",
  8409=>"100100001",
  8410=>"110110110",
  8411=>"000000111",
  8412=>"111111111",
  8413=>"110100100",
  8414=>"111111000",
  8415=>"000100000",
  8416=>"111111111",
  8417=>"111000111",
  8418=>"111111011",
  8419=>"100101111",
  8420=>"111111100",
  8421=>"111111111",
  8422=>"111100000",
  8423=>"110111111",
  8424=>"000100111",
  8425=>"001001000",
  8426=>"000000111",
  8427=>"000000000",
  8428=>"111111111",
  8429=>"000010010",
  8430=>"101000000",
  8431=>"000000111",
  8432=>"011001000",
  8433=>"111111110",
  8434=>"111010111",
  8435=>"000000000",
  8436=>"110110111",
  8437=>"111000000",
  8438=>"110110111",
  8439=>"110111111",
  8440=>"000000100",
  8441=>"000001111",
  8442=>"111111111",
  8443=>"110100111",
  8444=>"111011000",
  8445=>"000000000",
  8446=>"011001000",
  8447=>"100000100",
  8448=>"000000010",
  8449=>"000100110",
  8450=>"100110111",
  8451=>"000000000",
  8452=>"111111111",
  8453=>"000000000",
  8454=>"111111000",
  8455=>"100111000",
  8456=>"001111011",
  8457=>"000000000",
  8458=>"111111100",
  8459=>"000001001",
  8460=>"000000000",
  8461=>"000000100",
  8462=>"110001011",
  8463=>"111101000",
  8464=>"010000010",
  8465=>"000000000",
  8466=>"000011001",
  8467=>"010110100",
  8468=>"000000000",
  8469=>"011000000",
  8470=>"000000110",
  8471=>"111111111",
  8472=>"111111111",
  8473=>"100110111",
  8474=>"101111111",
  8475=>"111000000",
  8476=>"101101111",
  8477=>"011111000",
  8478=>"011111110",
  8479=>"111111111",
  8480=>"111011011",
  8481=>"000000100",
  8482=>"110110000",
  8483=>"111111111",
  8484=>"000000000",
  8485=>"111111111",
  8486=>"000000000",
  8487=>"000000000",
  8488=>"111111111",
  8489=>"000000000",
  8490=>"110110110",
  8491=>"000001000",
  8492=>"000000000",
  8493=>"000100000",
  8494=>"111100111",
  8495=>"111111011",
  8496=>"111111111",
  8497=>"101111111",
  8498=>"000000000",
  8499=>"010000000",
  8500=>"000010010",
  8501=>"001101111",
  8502=>"111111111",
  8503=>"011010000",
  8504=>"000000000",
  8505=>"111111111",
  8506=>"000100000",
  8507=>"000001000",
  8508=>"010010000",
  8509=>"100100000",
  8510=>"001011000",
  8511=>"000000000",
  8512=>"000000000",
  8513=>"111100111",
  8514=>"111111000",
  8515=>"111111111",
  8516=>"111111111",
  8517=>"000000000",
  8518=>"000000000",
  8519=>"000000100",
  8520=>"100000110",
  8521=>"111111111",
  8522=>"001001000",
  8523=>"101111111",
  8524=>"111011000",
  8525=>"000110111",
  8526=>"110110000",
  8527=>"111111011",
  8528=>"111101100",
  8529=>"000000000",
  8530=>"111111111",
  8531=>"111010000",
  8532=>"000000000",
  8533=>"111111111",
  8534=>"000000000",
  8535=>"111111111",
  8536=>"111111111",
  8537=>"111111111",
  8538=>"111111111",
  8539=>"000000111",
  8540=>"000000101",
  8541=>"111110000",
  8542=>"001000011",
  8543=>"111110111",
  8544=>"010010010",
  8545=>"000010010",
  8546=>"000001011",
  8547=>"000100111",
  8548=>"000000000",
  8549=>"000000000",
  8550=>"000000000",
  8551=>"111111000",
  8552=>"110111111",
  8553=>"111100000",
  8554=>"111111111",
  8555=>"000000000",
  8556=>"111111111",
  8557=>"000101111",
  8558=>"110110000",
  8559=>"001001100",
  8560=>"000000111",
  8561=>"000000111",
  8562=>"111111111",
  8563=>"010111110",
  8564=>"101000000",
  8565=>"001001001",
  8566=>"100000000",
  8567=>"000010110",
  8568=>"100111111",
  8569=>"111011011",
  8570=>"000000000",
  8571=>"111111111",
  8572=>"000110110",
  8573=>"111011011",
  8574=>"000000000",
  8575=>"111111111",
  8576=>"110110110",
  8577=>"001111111",
  8578=>"111111111",
  8579=>"001000000",
  8580=>"111011001",
  8581=>"111111111",
  8582=>"111111111",
  8583=>"000000010",
  8584=>"000010010",
  8585=>"100000000",
  8586=>"111111110",
  8587=>"011000000",
  8588=>"111111111",
  8589=>"100100000",
  8590=>"000000000",
  8591=>"100100000",
  8592=>"000000000",
  8593=>"100110111",
  8594=>"000010010",
  8595=>"011011011",
  8596=>"000000000",
  8597=>"000000000",
  8598=>"000001000",
  8599=>"001001001",
  8600=>"000000111",
  8601=>"111111111",
  8602=>"111111111",
  8603=>"000001001",
  8604=>"000000000",
  8605=>"111000001",
  8606=>"011000000",
  8607=>"000000111",
  8608=>"111111111",
  8609=>"111111111",
  8610=>"110100100",
  8611=>"111010111",
  8612=>"000000000",
  8613=>"000010000",
  8614=>"000000100",
  8615=>"000111111",
  8616=>"000000000",
  8617=>"100011111",
  8618=>"000110010",
  8619=>"011001010",
  8620=>"000000000",
  8621=>"000000000",
  8622=>"000001101",
  8623=>"011111111",
  8624=>"011111111",
  8625=>"000111111",
  8626=>"000000001",
  8627=>"111111110",
  8628=>"000000000",
  8629=>"000000000",
  8630=>"001101101",
  8631=>"001000000",
  8632=>"011100001",
  8633=>"111111111",
  8634=>"000000010",
  8635=>"111101101",
  8636=>"001011000",
  8637=>"111111111",
  8638=>"010000111",
  8639=>"111101100",
  8640=>"010011010",
  8641=>"111111111",
  8642=>"000000000",
  8643=>"000011000",
  8644=>"100001000",
  8645=>"111110111",
  8646=>"000100100",
  8647=>"001000000",
  8648=>"110110010",
  8649=>"000000000",
  8650=>"000000001",
  8651=>"111111010",
  8652=>"110110111",
  8653=>"111111111",
  8654=>"001110111",
  8655=>"000000101",
  8656=>"000000000",
  8657=>"111111111",
  8658=>"010000000",
  8659=>"000000000",
  8660=>"000111111",
  8661=>"000000100",
  8662=>"000000000",
  8663=>"011011000",
  8664=>"111111111",
  8665=>"111111000",
  8666=>"000000000",
  8667=>"100000000",
  8668=>"000000000",
  8669=>"000010111",
  8670=>"111111111",
  8671=>"000000000",
  8672=>"101100110",
  8673=>"111111111",
  8674=>"111010000",
  8675=>"111001000",
  8676=>"111111101",
  8677=>"010000000",
  8678=>"011011000",
  8679=>"111111111",
  8680=>"001111111",
  8681=>"000000000",
  8682=>"111111111",
  8683=>"000111111",
  8684=>"111000000",
  8685=>"000100100",
  8686=>"001001111",
  8687=>"111111111",
  8688=>"000000000",
  8689=>"111111111",
  8690=>"000000000",
  8691=>"111111111",
  8692=>"000000000",
  8693=>"010000000",
  8694=>"000000000",
  8695=>"111111001",
  8696=>"111111111",
  8697=>"001001001",
  8698=>"111111011",
  8699=>"111111111",
  8700=>"110000000",
  8701=>"000000000",
  8702=>"011000000",
  8703=>"111111110",
  8704=>"100000111",
  8705=>"111110110",
  8706=>"111100111",
  8707=>"000000000",
  8708=>"000011001",
  8709=>"011000001",
  8710=>"000000000",
  8711=>"000000011",
  8712=>"111111100",
  8713=>"111000000",
  8714=>"111000100",
  8715=>"111000000",
  8716=>"110110110",
  8717=>"111000000",
  8718=>"010110111",
  8719=>"111001000",
  8720=>"001001000",
  8721=>"000010111",
  8722=>"000000001",
  8723=>"000111111",
  8724=>"110000000",
  8725=>"000000000",
  8726=>"111000001",
  8727=>"111010000",
  8728=>"100110000",
  8729=>"001100100",
  8730=>"111111000",
  8731=>"111111011",
  8732=>"000000000",
  8733=>"000000111",
  8734=>"111111111",
  8735=>"000011001",
  8736=>"010010011",
  8737=>"111111111",
  8738=>"110110100",
  8739=>"000111111",
  8740=>"111111111",
  8741=>"000000000",
  8742=>"000000111",
  8743=>"000111111",
  8744=>"000011101",
  8745=>"111111111",
  8746=>"111110000",
  8747=>"000010000",
  8748=>"111111000",
  8749=>"101100111",
  8750=>"110000100",
  8751=>"000001111",
  8752=>"101111111",
  8753=>"000000011",
  8754=>"110110000",
  8755=>"111110111",
  8756=>"101101100",
  8757=>"111111110",
  8758=>"111001111",
  8759=>"111111111",
  8760=>"111010000",
  8761=>"110010011",
  8762=>"111111000",
  8763=>"000000111",
  8764=>"111111111",
  8765=>"110111110",
  8766=>"100100001",
  8767=>"110000000",
  8768=>"010000000",
  8769=>"110000000",
  8770=>"011111111",
  8771=>"010111101",
  8772=>"110110000",
  8773=>"111111000",
  8774=>"111100100",
  8775=>"111111110",
  8776=>"001111111",
  8777=>"000000000",
  8778=>"101111011",
  8779=>"100111000",
  8780=>"111010110",
  8781=>"111100000",
  8782=>"111111111",
  8783=>"011000000",
  8784=>"000000000",
  8785=>"100000000",
  8786=>"001011111",
  8787=>"000001111",
  8788=>"000110110",
  8789=>"011010111",
  8790=>"111011111",
  8791=>"000000000",
  8792=>"000100000",
  8793=>"000101001",
  8794=>"111001011",
  8795=>"101000000",
  8796=>"001000111",
  8797=>"111111111",
  8798=>"110111111",
  8799=>"111010000",
  8800=>"111000111",
  8801=>"111010010",
  8802=>"000000000",
  8803=>"000111111",
  8804=>"111111111",
  8805=>"000000000",
  8806=>"111111000",
  8807=>"000000000",
  8808=>"111000000",
  8809=>"111001111",
  8810=>"111100111",
  8811=>"000001001",
  8812=>"000110110",
  8813=>"010000000",
  8814=>"000000111",
  8815=>"000111111",
  8816=>"000000100",
  8817=>"111000000",
  8818=>"111101111",
  8819=>"111011010",
  8820=>"010000110",
  8821=>"000000111",
  8822=>"111011010",
  8823=>"011000000",
  8824=>"011001000",
  8825=>"111011111",
  8826=>"110111110",
  8827=>"000000000",
  8828=>"111111110",
  8829=>"111111111",
  8830=>"000000000",
  8831=>"011111111",
  8832=>"000000101",
  8833=>"000000000",
  8834=>"111000000",
  8835=>"111111110",
  8836=>"000010111",
  8837=>"111111000",
  8838=>"101000000",
  8839=>"000000111",
  8840=>"000101111",
  8841=>"001101101",
  8842=>"000110000",
  8843=>"000000000",
  8844=>"000111101",
  8845=>"111111111",
  8846=>"111011000",
  8847=>"000010000",
  8848=>"111111111",
  8849=>"000000000",
  8850=>"110000000",
  8851=>"111100000",
  8852=>"010000000",
  8853=>"000000111",
  8854=>"000000111",
  8855=>"100000101",
  8856=>"000000111",
  8857=>"000110111",
  8858=>"000000111",
  8859=>"000000000",
  8860=>"111000000",
  8861=>"110100111",
  8862=>"100000000",
  8863=>"111110000",
  8864=>"111111001",
  8865=>"000111111",
  8866=>"000111111",
  8867=>"111111001",
  8868=>"000011111",
  8869=>"100110111",
  8870=>"000111010",
  8871=>"111011011",
  8872=>"111001000",
  8873=>"101001101",
  8874=>"111111011",
  8875=>"000110110",
  8876=>"111000000",
  8877=>"100100100",
  8878=>"111111111",
  8879=>"111000000",
  8880=>"000111111",
  8881=>"001010100",
  8882=>"010011011",
  8883=>"111111111",
  8884=>"111011001",
  8885=>"111111001",
  8886=>"111000000",
  8887=>"111111111",
  8888=>"111111111",
  8889=>"111111111",
  8890=>"000001111",
  8891=>"110110111",
  8892=>"000000001",
  8893=>"111111111",
  8894=>"101000000",
  8895=>"000100110",
  8896=>"101111111",
  8897=>"000010110",
  8898=>"000000111",
  8899=>"111111111",
  8900=>"000000111",
  8901=>"100000100",
  8902=>"010111010",
  8903=>"000010000",
  8904=>"000000000",
  8905=>"001000000",
  8906=>"111011011",
  8907=>"000000100",
  8908=>"111100100",
  8909=>"000101111",
  8910=>"001001011",
  8911=>"111111000",
  8912=>"001000100",
  8913=>"010000000",
  8914=>"101111111",
  8915=>"001000000",
  8916=>"100000000",
  8917=>"111001000",
  8918=>"000100111",
  8919=>"111111000",
  8920=>"110111011",
  8921=>"111111101",
  8922=>"011000000",
  8923=>"001101101",
  8924=>"001001101",
  8925=>"100111101",
  8926=>"111111111",
  8927=>"011000000",
  8928=>"000000111",
  8929=>"000101000",
  8930=>"000000111",
  8931=>"111011011",
  8932=>"000111101",
  8933=>"111111001",
  8934=>"000000000",
  8935=>"000000111",
  8936=>"010000000",
  8937=>"001001000",
  8938=>"001000000",
  8939=>"101111111",
  8940=>"111000001",
  8941=>"000000101",
  8942=>"111011000",
  8943=>"000111111",
  8944=>"111111111",
  8945=>"110100100",
  8946=>"111101000",
  8947=>"000000001",
  8948=>"000000000",
  8949=>"111111011",
  8950=>"010010110",
  8951=>"111111111",
  8952=>"010111011",
  8953=>"111000000",
  8954=>"111010101",
  8955=>"101000010",
  8956=>"110000100",
  8957=>"010000000",
  8958=>"111000001",
  8959=>"000010110",
  8960=>"000000000",
  8961=>"111010000",
  8962=>"000000000",
  8963=>"010010001",
  8964=>"000000000",
  8965=>"110111111",
  8966=>"111111111",
  8967=>"111100000",
  8968=>"011000111",
  8969=>"000100111",
  8970=>"000100111",
  8971=>"001111111",
  8972=>"111001000",
  8973=>"111011000",
  8974=>"111111111",
  8975=>"000000000",
  8976=>"111000000",
  8977=>"111101101",
  8978=>"000001000",
  8979=>"100110111",
  8980=>"000000111",
  8981=>"111111000",
  8982=>"100110100",
  8983=>"000000110",
  8984=>"000111111",
  8985=>"000000111",
  8986=>"111111100",
  8987=>"110110111",
  8988=>"110100100",
  8989=>"111111111",
  8990=>"111000000",
  8991=>"000000000",
  8992=>"000100111",
  8993=>"000000111",
  8994=>"000011110",
  8995=>"000101111",
  8996=>"111010111",
  8997=>"111000110",
  8998=>"011000000",
  8999=>"000111111",
  9000=>"000011111",
  9001=>"011011000",
  9002=>"111111111",
  9003=>"110000010",
  9004=>"000100110",
  9005=>"001000001",
  9006=>"111111111",
  9007=>"000111111",
  9008=>"110110000",
  9009=>"010000000",
  9010=>"111111111",
  9011=>"000111111",
  9012=>"111111111",
  9013=>"011010000",
  9014=>"111111011",
  9015=>"111111000",
  9016=>"011001000",
  9017=>"000000000",
  9018=>"000000000",
  9019=>"111111111",
  9020=>"110110010",
  9021=>"111111111",
  9022=>"111011000",
  9023=>"111000000",
  9024=>"111111100",
  9025=>"110110110",
  9026=>"110111111",
  9027=>"000000000",
  9028=>"111111111",
  9029=>"111000111",
  9030=>"000110111",
  9031=>"101101100",
  9032=>"110011111",
  9033=>"111111000",
  9034=>"110111111",
  9035=>"011011000",
  9036=>"000101111",
  9037=>"001001111",
  9038=>"001111111",
  9039=>"111000100",
  9040=>"110011001",
  9041=>"000000000",
  9042=>"111001111",
  9043=>"111000000",
  9044=>"101111010",
  9045=>"001100111",
  9046=>"010010001",
  9047=>"111111111",
  9048=>"110110111",
  9049=>"111111110",
  9050=>"110000000",
  9051=>"011111111",
  9052=>"000001101",
  9053=>"000110100",
  9054=>"101001001",
  9055=>"001011011",
  9056=>"001001001",
  9057=>"111111111",
  9058=>"110111111",
  9059=>"101101000",
  9060=>"100000000",
  9061=>"000000111",
  9062=>"000000000",
  9063=>"000000111",
  9064=>"110111011",
  9065=>"000111111",
  9066=>"010111111",
  9067=>"111000000",
  9068=>"001001111",
  9069=>"010111111",
  9070=>"111111001",
  9071=>"011000000",
  9072=>"111111011",
  9073=>"100000000",
  9074=>"000001000",
  9075=>"011111100",
  9076=>"000010011",
  9077=>"111100101",
  9078=>"100000001",
  9079=>"111111000",
  9080=>"111111000",
  9081=>"000000000",
  9082=>"111000000",
  9083=>"111111000",
  9084=>"101000000",
  9085=>"000000000",
  9086=>"111011000",
  9087=>"111000000",
  9088=>"111111111",
  9089=>"000110110",
  9090=>"111110000",
  9091=>"100100000",
  9092=>"011000000",
  9093=>"001001101",
  9094=>"100111111",
  9095=>"100000111",
  9096=>"111111000",
  9097=>"011000000",
  9098=>"000000011",
  9099=>"000000000",
  9100=>"101000101",
  9101=>"000110110",
  9102=>"111001101",
  9103=>"000000010",
  9104=>"111011000",
  9105=>"000000111",
  9106=>"000111101",
  9107=>"111111111",
  9108=>"000101111",
  9109=>"001011000",
  9110=>"101111111",
  9111=>"000000000",
  9112=>"000000100",
  9113=>"100000110",
  9114=>"111111110",
  9115=>"111000100",
  9116=>"111111000",
  9117=>"000111111",
  9118=>"000001000",
  9119=>"111100110",
  9120=>"111111000",
  9121=>"100100100",
  9122=>"101000000",
  9123=>"111001101",
  9124=>"111111111",
  9125=>"111101000",
  9126=>"111111111",
  9127=>"000000110",
  9128=>"011000000",
  9129=>"000111111",
  9130=>"000000101",
  9131=>"000000000",
  9132=>"000111001",
  9133=>"010110000",
  9134=>"110111000",
  9135=>"111001000",
  9136=>"000100111",
  9137=>"001000000",
  9138=>"110011111",
  9139=>"010111011",
  9140=>"000000111",
  9141=>"001001111",
  9142=>"110111111",
  9143=>"000000000",
  9144=>"000111111",
  9145=>"000000000",
  9146=>"111111111",
  9147=>"111111111",
  9148=>"000000111",
  9149=>"000000000",
  9150=>"101100111",
  9151=>"100100100",
  9152=>"100111111",
  9153=>"001100000",
  9154=>"111000000",
  9155=>"111111000",
  9156=>"111111110",
  9157=>"111110000",
  9158=>"111110111",
  9159=>"111101101",
  9160=>"111111000",
  9161=>"000000000",
  9162=>"111101000",
  9163=>"111111111",
  9164=>"111001111",
  9165=>"111110111",
  9166=>"110111111",
  9167=>"111011111",
  9168=>"101111111",
  9169=>"000001111",
  9170=>"001111111",
  9171=>"010110111",
  9172=>"111111110",
  9173=>"111111100",
  9174=>"010010000",
  9175=>"011011011",
  9176=>"100100100",
  9177=>"101000000",
  9178=>"110010010",
  9179=>"110010001",
  9180=>"000011010",
  9181=>"100001101",
  9182=>"001111111",
  9183=>"001111011",
  9184=>"111001000",
  9185=>"000000111",
  9186=>"111111111",
  9187=>"001000011",
  9188=>"111111111",
  9189=>"110110000",
  9190=>"101000000",
  9191=>"111001001",
  9192=>"011000000",
  9193=>"110111101",
  9194=>"010111110",
  9195=>"001001111",
  9196=>"100110000",
  9197=>"010000000",
  9198=>"000000000",
  9199=>"101111111",
  9200=>"000000000",
  9201=>"111111101",
  9202=>"001011111",
  9203=>"000000000",
  9204=>"100000000",
  9205=>"001101111",
  9206=>"111111111",
  9207=>"111111000",
  9208=>"001111000",
  9209=>"001001001",
  9210=>"111011000",
  9211=>"111111101",
  9212=>"000001000",
  9213=>"110110111",
  9214=>"000000110",
  9215=>"100000100",
  9216=>"111111111",
  9217=>"011111111",
  9218=>"011000000",
  9219=>"000000110",
  9220=>"000100100",
  9221=>"010011000",
  9222=>"000111111",
  9223=>"111000000",
  9224=>"111100000",
  9225=>"111111111",
  9226=>"000000000",
  9227=>"111111111",
  9228=>"000000111",
  9229=>"111111111",
  9230=>"111111000",
  9231=>"110110000",
  9232=>"110111111",
  9233=>"000111111",
  9234=>"000111111",
  9235=>"000000000",
  9236=>"111111011",
  9237=>"000000000",
  9238=>"001001000",
  9239=>"110111111",
  9240=>"000100110",
  9241=>"011001000",
  9242=>"101000111",
  9243=>"000000000",
  9244=>"111110100",
  9245=>"111000100",
  9246=>"111111101",
  9247=>"111111111",
  9248=>"000000000",
  9249=>"111111101",
  9250=>"111001000",
  9251=>"100000001",
  9252=>"111111111",
  9253=>"000000000",
  9254=>"011001000",
  9255=>"001001000",
  9256=>"111111001",
  9257=>"111111000",
  9258=>"111111111",
  9259=>"111111111",
  9260=>"111000011",
  9261=>"101100001",
  9262=>"000011011",
  9263=>"001111111",
  9264=>"110000000",
  9265=>"111111111",
  9266=>"000000000",
  9267=>"000000000",
  9268=>"000000000",
  9269=>"000011001",
  9270=>"000000010",
  9271=>"011000110",
  9272=>"111111000",
  9273=>"111111011",
  9274=>"111111111",
  9275=>"000000000",
  9276=>"000000000",
  9277=>"001000000",
  9278=>"000111111",
  9279=>"000000000",
  9280=>"011000000",
  9281=>"100111111",
  9282=>"111110111",
  9283=>"001000111",
  9284=>"001101001",
  9285=>"001011111",
  9286=>"000000000",
  9287=>"111111011",
  9288=>"000110100",
  9289=>"010010001",
  9290=>"000001011",
  9291=>"000000111",
  9292=>"000000000",
  9293=>"110111111",
  9294=>"000000001",
  9295=>"000000110",
  9296=>"010000000",
  9297=>"000000100",
  9298=>"000000000",
  9299=>"111111100",
  9300=>"000000000",
  9301=>"001010010",
  9302=>"111111100",
  9303=>"011111111",
  9304=>"011101100",
  9305=>"111000000",
  9306=>"000000000",
  9307=>"011111001",
  9308=>"111111111",
  9309=>"000000000",
  9310=>"111110000",
  9311=>"000010110",
  9312=>"000000010",
  9313=>"000000000",
  9314=>"111011010",
  9315=>"011011111",
  9316=>"001101111",
  9317=>"000000000",
  9318=>"001000000",
  9319=>"000000000",
  9320=>"111111111",
  9321=>"111111111",
  9322=>"111111111",
  9323=>"001011011",
  9324=>"000101001",
  9325=>"111111111",
  9326=>"111111111",
  9327=>"111101001",
  9328=>"011011000",
  9329=>"001111110",
  9330=>"110100000",
  9331=>"111111101",
  9332=>"000000000",
  9333=>"111000000",
  9334=>"111111111",
  9335=>"000000011",
  9336=>"111111110",
  9337=>"100000111",
  9338=>"000000011",
  9339=>"111111010",
  9340=>"100000001",
  9341=>"110110000",
  9342=>"000000000",
  9343=>"000000000",
  9344=>"111111111",
  9345=>"011011000",
  9346=>"100100110",
  9347=>"111111001",
  9348=>"000000000",
  9349=>"000000000",
  9350=>"111111110",
  9351=>"111111111",
  9352=>"011111000",
  9353=>"011111110",
  9354=>"111111111",
  9355=>"000000110",
  9356=>"111110010",
  9357=>"111111111",
  9358=>"001001000",
  9359=>"111111111",
  9360=>"111111111",
  9361=>"000000000",
  9362=>"000000101",
  9363=>"001001111",
  9364=>"001000000",
  9365=>"110110000",
  9366=>"100111100",
  9367=>"011011000",
  9368=>"111111000",
  9369=>"111101011",
  9370=>"000110110",
  9371=>"100000000",
  9372=>"000000000",
  9373=>"010000000",
  9374=>"111000111",
  9375=>"111111010",
  9376=>"000110111",
  9377=>"110110110",
  9378=>"111111111",
  9379=>"000000000",
  9380=>"000111111",
  9381=>"111000000",
  9382=>"111111111",
  9383=>"000111111",
  9384=>"000000000",
  9385=>"000000000",
  9386=>"000000000",
  9387=>"000000000",
  9388=>"001101000",
  9389=>"000000011",
  9390=>"011111000",
  9391=>"111111111",
  9392=>"011111111",
  9393=>"000000000",
  9394=>"010111111",
  9395=>"000000000",
  9396=>"111001000",
  9397=>"111110111",
  9398=>"111111111",
  9399=>"000000000",
  9400=>"111101111",
  9401=>"111111000",
  9402=>"000000000",
  9403=>"000000000",
  9404=>"000110100",
  9405=>"000000000",
  9406=>"111111111",
  9407=>"010000000",
  9408=>"010101101",
  9409=>"000000000",
  9410=>"110110100",
  9411=>"000010111",
  9412=>"000000000",
  9413=>"001011010",
  9414=>"000001001",
  9415=>"000000000",
  9416=>"111111110",
  9417=>"111110000",
  9418=>"010110100",
  9419=>"000000000",
  9420=>"111111011",
  9421=>"000100000",
  9422=>"001001011",
  9423=>"000001011",
  9424=>"111001000",
  9425=>"111111111",
  9426=>"111111111",
  9427=>"011111011",
  9428=>"111001000",
  9429=>"011110110",
  9430=>"111000000",
  9431=>"111111111",
  9432=>"011111111",
  9433=>"111111000",
  9434=>"111111100",
  9435=>"000000000",
  9436=>"000000000",
  9437=>"111111111",
  9438=>"010000000",
  9439=>"011010000",
  9440=>"000000000",
  9441=>"000000000",
  9442=>"110000000",
  9443=>"100000000",
  9444=>"000000110",
  9445=>"100101100",
  9446=>"000001111",
  9447=>"000011111",
  9448=>"111110111",
  9449=>"000000000",
  9450=>"111111100",
  9451=>"000000000",
  9452=>"110111110",
  9453=>"000000011",
  9454=>"111111110",
  9455=>"000111111",
  9456=>"111011111",
  9457=>"111111111",
  9458=>"111111111",
  9459=>"111111000",
  9460=>"000000000",
  9461=>"000010000",
  9462=>"111111111",
  9463=>"111111000",
  9464=>"111111111",
  9465=>"000000000",
  9466=>"111000000",
  9467=>"000000000",
  9468=>"000011001",
  9469=>"001100000",
  9470=>"000010000",
  9471=>"000110000",
  9472=>"001000000",
  9473=>"000110001",
  9474=>"011111111",
  9475=>"011111111",
  9476=>"110100000",
  9477=>"000000000",
  9478=>"111100000",
  9479=>"001111111",
  9480=>"111110000",
  9481=>"000000000",
  9482=>"000000000",
  9483=>"000000001",
  9484=>"111111111",
  9485=>"000001111",
  9486=>"000000000",
  9487=>"100101000",
  9488=>"000100000",
  9489=>"100100100",
  9490=>"000000000",
  9491=>"110000001",
  9492=>"000111011",
  9493=>"111111111",
  9494=>"001001011",
  9495=>"101111111",
  9496=>"000000001",
  9497=>"111110111",
  9498=>"010000000",
  9499=>"011111110",
  9500=>"000000011",
  9501=>"111000000",
  9502=>"000000111",
  9503=>"010111010",
  9504=>"100111111",
  9505=>"000011111",
  9506=>"110111000",
  9507=>"010111111",
  9508=>"000000000",
  9509=>"111111111",
  9510=>"000111111",
  9511=>"011110000",
  9512=>"000000000",
  9513=>"000000010",
  9514=>"111111111",
  9515=>"000000000",
  9516=>"000000000",
  9517=>"111111111",
  9518=>"111111000",
  9519=>"000111011",
  9520=>"000000000",
  9521=>"000000000",
  9522=>"000011011",
  9523=>"111000111",
  9524=>"000000111",
  9525=>"111111011",
  9526=>"000010011",
  9527=>"000000000",
  9528=>"000001000",
  9529=>"110000100",
  9530=>"111111111",
  9531=>"100011011",
  9532=>"111111111",
  9533=>"111110111",
  9534=>"101101111",
  9535=>"001001001",
  9536=>"111111100",
  9537=>"111011111",
  9538=>"011111001",
  9539=>"000000000",
  9540=>"111111111",
  9541=>"111110000",
  9542=>"100111111",
  9543=>"000000000",
  9544=>"011000000",
  9545=>"111111111",
  9546=>"111111111",
  9547=>"000000000",
  9548=>"000000000",
  9549=>"010000111",
  9550=>"111111111",
  9551=>"001001001",
  9552=>"001011011",
  9553=>"001000000",
  9554=>"000110111",
  9555=>"000000000",
  9556=>"000000000",
  9557=>"011001111",
  9558=>"000100111",
  9559=>"000000100",
  9560=>"001001001",
  9561=>"111111111",
  9562=>"111001011",
  9563=>"000010000",
  9564=>"000000111",
  9565=>"111100111",
  9566=>"001000000",
  9567=>"100100001",
  9568=>"111111011",
  9569=>"000000000",
  9570=>"111111011",
  9571=>"001000000",
  9572=>"000001111",
  9573=>"111111111",
  9574=>"111111111",
  9575=>"111100100",
  9576=>"100110001",
  9577=>"001001000",
  9578=>"111111111",
  9579=>"000100100",
  9580=>"110110110",
  9581=>"000111111",
  9582=>"000000000",
  9583=>"111111111",
  9584=>"010010000",
  9585=>"110110111",
  9586=>"111111110",
  9587=>"111100100",
  9588=>"000000000",
  9589=>"010110010",
  9590=>"110110000",
  9591=>"000000111",
  9592=>"000000111",
  9593=>"111000000",
  9594=>"001001011",
  9595=>"000000000",
  9596=>"001111111",
  9597=>"000111111",
  9598=>"111111111",
  9599=>"111111111",
  9600=>"110000001",
  9601=>"010010000",
  9602=>"000110111",
  9603=>"111000000",
  9604=>"000111111",
  9605=>"000000000",
  9606=>"010010000",
  9607=>"010111111",
  9608=>"010011001",
  9609=>"111111110",
  9610=>"111000000",
  9611=>"010111011",
  9612=>"111111111",
  9613=>"111111110",
  9614=>"000001000",
  9615=>"000000100",
  9616=>"000000000",
  9617=>"000111111",
  9618=>"111011110",
  9619=>"111111111",
  9620=>"000000000",
  9621=>"001001011",
  9622=>"001011111",
  9623=>"011011011",
  9624=>"000001111",
  9625=>"011000000",
  9626=>"100000010",
  9627=>"000111111",
  9628=>"111111111",
  9629=>"000100111",
  9630=>"000000100",
  9631=>"111111111",
  9632=>"000000000",
  9633=>"100100110",
  9634=>"000001011",
  9635=>"110000011",
  9636=>"100110110",
  9637=>"011011000",
  9638=>"001001001",
  9639=>"111000000",
  9640=>"111111111",
  9641=>"000000000",
  9642=>"010111111",
  9643=>"111101101",
  9644=>"111000000",
  9645=>"000100000",
  9646=>"111111000",
  9647=>"101111111",
  9648=>"111111111",
  9649=>"100101111",
  9650=>"111101111",
  9651=>"100111111",
  9652=>"111111111",
  9653=>"111111111",
  9654=>"000111111",
  9655=>"111100001",
  9656=>"111111111",
  9657=>"000000101",
  9658=>"000000000",
  9659=>"000010000",
  9660=>"000000000",
  9661=>"000000111",
  9662=>"000000000",
  9663=>"010110001",
  9664=>"111111000",
  9665=>"100111111",
  9666=>"000000000",
  9667=>"111001000",
  9668=>"001001001",
  9669=>"001001111",
  9670=>"101111111",
  9671=>"000000001",
  9672=>"001011000",
  9673=>"001111111",
  9674=>"000000110",
  9675=>"110110000",
  9676=>"000000000",
  9677=>"011011001",
  9678=>"111011111",
  9679=>"000000000",
  9680=>"000011111",
  9681=>"111110000",
  9682=>"010111111",
  9683=>"111111000",
  9684=>"001101101",
  9685=>"000000000",
  9686=>"111010000",
  9687=>"011001001",
  9688=>"101000000",
  9689=>"111000000",
  9690=>"000100111",
  9691=>"111111111",
  9692=>"000000111",
  9693=>"011000000",
  9694=>"000000001",
  9695=>"110110000",
  9696=>"101101000",
  9697=>"000000000",
  9698=>"111111111",
  9699=>"011011111",
  9700=>"001001000",
  9701=>"000000110",
  9702=>"011000000",
  9703=>"010010000",
  9704=>"011011001",
  9705=>"000000000",
  9706=>"110111111",
  9707=>"111100000",
  9708=>"000000000",
  9709=>"000100111",
  9710=>"100111001",
  9711=>"011111111",
  9712=>"101111111",
  9713=>"011111010",
  9714=>"000101011",
  9715=>"100000000",
  9716=>"111100000",
  9717=>"111111000",
  9718=>"111111111",
  9719=>"001010010",
  9720=>"111111011",
  9721=>"000001100",
  9722=>"000000000",
  9723=>"010111110",
  9724=>"101101101",
  9725=>"000000000",
  9726=>"000000000",
  9727=>"111100111",
  9728=>"000000000",
  9729=>"000000000",
  9730=>"101001000",
  9731=>"100000001",
  9732=>"110110101",
  9733=>"011001111",
  9734=>"000001011",
  9735=>"111111111",
  9736=>"000000111",
  9737=>"000000000",
  9738=>"110111111",
  9739=>"000000000",
  9740=>"100110100",
  9741=>"110110111",
  9742=>"111110100",
  9743=>"011000000",
  9744=>"110110111",
  9745=>"000000000",
  9746=>"000111111",
  9747=>"000001111",
  9748=>"011010111",
  9749=>"000000000",
  9750=>"000000000",
  9751=>"111111111",
  9752=>"000100100",
  9753=>"011111111",
  9754=>"111111010",
  9755=>"111000000",
  9756=>"011111111",
  9757=>"101111010",
  9758=>"001000000",
  9759=>"111111111",
  9760=>"000000111",
  9761=>"111111111",
  9762=>"111110110",
  9763=>"111101111",
  9764=>"000000000",
  9765=>"111111111",
  9766=>"101000111",
  9767=>"000100111",
  9768=>"110100000",
  9769=>"000000000",
  9770=>"001111111",
  9771=>"100100000",
  9772=>"111111111",
  9773=>"000111111",
  9774=>"110111111",
  9775=>"111111111",
  9776=>"111111011",
  9777=>"111000000",
  9778=>"001001001",
  9779=>"001000111",
  9780=>"000111111",
  9781=>"110100111",
  9782=>"111111111",
  9783=>"000000001",
  9784=>"111111111",
  9785=>"000000010",
  9786=>"011001001",
  9787=>"000101101",
  9788=>"100111111",
  9789=>"011010000",
  9790=>"001101100",
  9791=>"001000111",
  9792=>"111111000",
  9793=>"000000000",
  9794=>"000000111",
  9795=>"111011111",
  9796=>"000000111",
  9797=>"000100110",
  9798=>"011000111",
  9799=>"000000000",
  9800=>"000000000",
  9801=>"101000111",
  9802=>"100111011",
  9803=>"000111111",
  9804=>"111001000",
  9805=>"000010000",
  9806=>"001000111",
  9807=>"111111111",
  9808=>"000000010",
  9809=>"111111001",
  9810=>"000000000",
  9811=>"100100110",
  9812=>"000111111",
  9813=>"000000000",
  9814=>"111111111",
  9815=>"111111111",
  9816=>"111110000",
  9817=>"111000000",
  9818=>"000000000",
  9819=>"000000010",
  9820=>"011111111",
  9821=>"000000011",
  9822=>"111001001",
  9823=>"111000001",
  9824=>"000001000",
  9825=>"010010011",
  9826=>"111111111",
  9827=>"001001111",
  9828=>"100010111",
  9829=>"111111000",
  9830=>"010110000",
  9831=>"111000000",
  9832=>"101000111",
  9833=>"111111111",
  9834=>"000110000",
  9835=>"000000000",
  9836=>"110010000",
  9837=>"110000000",
  9838=>"010000111",
  9839=>"111111010",
  9840=>"111110111",
  9841=>"111110100",
  9842=>"000000000",
  9843=>"000111111",
  9844=>"011111111",
  9845=>"000000000",
  9846=>"001000000",
  9847=>"000000010",
  9848=>"000000111",
  9849=>"011000100",
  9850=>"000000000",
  9851=>"000100100",
  9852=>"110111011",
  9853=>"001100100",
  9854=>"000000000",
  9855=>"111000000",
  9856=>"100000011",
  9857=>"000000001",
  9858=>"111110111",
  9859=>"011011001",
  9860=>"001001000",
  9861=>"101111111",
  9862=>"110000010",
  9863=>"000010111",
  9864=>"111110000",
  9865=>"010000111",
  9866=>"010000000",
  9867=>"011111111",
  9868=>"100000111",
  9869=>"000000000",
  9870=>"111111001",
  9871=>"111111111",
  9872=>"000000000",
  9873=>"010010010",
  9874=>"000000111",
  9875=>"000000000",
  9876=>"000010000",
  9877=>"000000000",
  9878=>"000111110",
  9879=>"100000000",
  9880=>"000000000",
  9881=>"100100111",
  9882=>"000000000",
  9883=>"011011111",
  9884=>"000000110",
  9885=>"000000000",
  9886=>"011000000",
  9887=>"000000111",
  9888=>"100000101",
  9889=>"011010000",
  9890=>"011000111",
  9891=>"000000000",
  9892=>"001000000",
  9893=>"000010001",
  9894=>"111111000",
  9895=>"001011111",
  9896=>"001000111",
  9897=>"000000000",
  9898=>"010010000",
  9899=>"000011110",
  9900=>"111111111",
  9901=>"111110000",
  9902=>"011000011",
  9903=>"111111111",
  9904=>"000000111",
  9905=>"010111111",
  9906=>"111111000",
  9907=>"000101110",
  9908=>"111111000",
  9909=>"111110000",
  9910=>"011011000",
  9911=>"100111111",
  9912=>"100100111",
  9913=>"110110110",
  9914=>"000000101",
  9915=>"001000000",
  9916=>"110111111",
  9917=>"010111111",
  9918=>"111111111",
  9919=>"000000000",
  9920=>"000000000",
  9921=>"000000000",
  9922=>"111111111",
  9923=>"111111011",
  9924=>"000000010",
  9925=>"000101111",
  9926=>"001100000",
  9927=>"101111110",
  9928=>"000011111",
  9929=>"111111111",
  9930=>"111111111",
  9931=>"000100111",
  9932=>"011011000",
  9933=>"000010011",
  9934=>"110111111",
  9935=>"011111000",
  9936=>"001000000",
  9937=>"111000000",
  9938=>"000000001",
  9939=>"111101111",
  9940=>"111111111",
  9941=>"000000111",
  9942=>"000000000",
  9943=>"000000111",
  9944=>"110110010",
  9945=>"000000000",
  9946=>"000000011",
  9947=>"000011111",
  9948=>"111100100",
  9949=>"000000000",
  9950=>"010000000",
  9951=>"100000000",
  9952=>"111111000",
  9953=>"111111000",
  9954=>"111001001",
  9955=>"000000011",
  9956=>"000100100",
  9957=>"000000111",
  9958=>"000000111",
  9959=>"000000011",
  9960=>"111111111",
  9961=>"111000000",
  9962=>"111110100",
  9963=>"011000000",
  9964=>"011111111",
  9965=>"000000000",
  9966=>"111111111",
  9967=>"010110111",
  9968=>"000000000",
  9969=>"000000000",
  9970=>"011111111",
  9971=>"011000000",
  9972=>"000011111",
  9973=>"111000000",
  9974=>"011111111",
  9975=>"000000000",
  9976=>"100000111",
  9977=>"111111000",
  9978=>"111111111",
  9979=>"111111001",
  9980=>"100110100",
  9981=>"101000000",
  9982=>"010110010",
  9983=>"100000000",
  9984=>"000100111",
  9985=>"110100011",
  9986=>"110110110",
  9987=>"001011111",
  9988=>"111111101",
  9989=>"111010000",
  9990=>"000000101",
  9991=>"010111101",
  9992=>"000000101",
  9993=>"100000111",
  9994=>"100111101",
  9995=>"111111111",
  9996=>"001001111",
  9997=>"000000000",
  9998=>"000000001",
  9999=>"111111010",
  10000=>"111111101",
  10001=>"000000000",
  10002=>"110100001",
  10003=>"000000000",
  10004=>"110100000",
  10005=>"000011011",
  10006=>"100110110",
  10007=>"000000000",
  10008=>"000010000",
  10009=>"111100000",
  10010=>"000000000",
  10011=>"110111111",
  10012=>"110011011",
  10013=>"111000000",
  10014=>"111100100",
  10015=>"010000000",
  10016=>"000100000",
  10017=>"111000000",
  10018=>"000000010",
  10019=>"111001001",
  10020=>"111111111",
  10021=>"000000100",
  10022=>"000000110",
  10023=>"010100000",
  10024=>"111111000",
  10025=>"000001111",
  10026=>"010010110",
  10027=>"111111000",
  10028=>"000000111",
  10029=>"000110110",
  10030=>"111110010",
  10031=>"000000000",
  10032=>"011011110",
  10033=>"100000000",
  10034=>"101000000",
  10035=>"000000000",
  10036=>"111101011",
  10037=>"000111111",
  10038=>"000100111",
  10039=>"111000000",
  10040=>"111111001",
  10041=>"111101111",
  10042=>"101000000",
  10043=>"111111001",
  10044=>"000000000",
  10045=>"111111001",
  10046=>"110111100",
  10047=>"111110110",
  10048=>"000000000",
  10049=>"111111111",
  10050=>"110111110",
  10051=>"000000100",
  10052=>"000000111",
  10053=>"000011011",
  10054=>"000000111",
  10055=>"000100100",
  10056=>"111111011",
  10057=>"000000000",
  10058=>"011000101",
  10059=>"000111111",
  10060=>"000111111",
  10061=>"111111011",
  10062=>"000000111",
  10063=>"111110100",
  10064=>"111111111",
  10065=>"111111000",
  10066=>"110100000",
  10067=>"111010000",
  10068=>"000000000",
  10069=>"000011011",
  10070=>"111110000",
  10071=>"111111111",
  10072=>"111111110",
  10073=>"000000000",
  10074=>"110110000",
  10075=>"111111101",
  10076=>"000000000",
  10077=>"111111101",
  10078=>"010010000",
  10079=>"000010110",
  10080=>"100100000",
  10081=>"000110111",
  10082=>"110000000",
  10083=>"000000000",
  10084=>"110110100",
  10085=>"000000000",
  10086=>"000111111",
  10087=>"000000000",
  10088=>"000110111",
  10089=>"111111110",
  10090=>"000000000",
  10091=>"111000001",
  10092=>"100000000",
  10093=>"111111111",
  10094=>"000000111",
  10095=>"101111001",
  10096=>"100111111",
  10097=>"111010011",
  10098=>"010010111",
  10099=>"111110100",
  10100=>"000000110",
  10101=>"101000000",
  10102=>"111111111",
  10103=>"000000000",
  10104=>"000000110",
  10105=>"111101000",
  10106=>"100111111",
  10107=>"000010011",
  10108=>"111011001",
  10109=>"111111100",
  10110=>"000000000",
  10111=>"000000000",
  10112=>"111111101",
  10113=>"000000000",
  10114=>"001001011",
  10115=>"000000000",
  10116=>"000100111",
  10117=>"000100111",
  10118=>"101000111",
  10119=>"111111111",
  10120=>"000000011",
  10121=>"110110000",
  10122=>"111111111",
  10123=>"000000000",
  10124=>"111101111",
  10125=>"001111110",
  10126=>"110000000",
  10127=>"111010010",
  10128=>"000000000",
  10129=>"110111111",
  10130=>"011011011",
  10131=>"000000001",
  10132=>"111000000",
  10133=>"000011010",
  10134=>"111111111",
  10135=>"000000001",
  10136=>"111111111",
  10137=>"111000010",
  10138=>"100111111",
  10139=>"000000000",
  10140=>"111111111",
  10141=>"111100000",
  10142=>"000101101",
  10143=>"111000111",
  10144=>"010110000",
  10145=>"000000000",
  10146=>"001100101",
  10147=>"000000101",
  10148=>"111100100",
  10149=>"000000000",
  10150=>"111111000",
  10151=>"000110111",
  10152=>"111111111",
  10153=>"000000000",
  10154=>"100110110",
  10155=>"010010001",
  10156=>"000000000",
  10157=>"010110111",
  10158=>"111111000",
  10159=>"000111011",
  10160=>"111111110",
  10161=>"111111111",
  10162=>"111110111",
  10163=>"010111000",
  10164=>"000000000",
  10165=>"001000000",
  10166=>"000100101",
  10167=>"000000001",
  10168=>"000001000",
  10169=>"000000011",
  10170=>"110000000",
  10171=>"111111101",
  10172=>"111101000",
  10173=>"100000111",
  10174=>"111000000",
  10175=>"001001000",
  10176=>"000000000",
  10177=>"000000000",
  10178=>"111111111",
  10179=>"111111111",
  10180=>"111100000",
  10181=>"000000111",
  10182=>"010110110",
  10183=>"000000111",
  10184=>"010000000",
  10185=>"010011001",
  10186=>"001001011",
  10187=>"000001001",
  10188=>"111111000",
  10189=>"011111010",
  10190=>"111111111",
  10191=>"001111111",
  10192=>"000000111",
  10193=>"000000000",
  10194=>"000000000",
  10195=>"111111111",
  10196=>"000000111",
  10197=>"111111111",
  10198=>"000000111",
  10199=>"011011011",
  10200=>"000001111",
  10201=>"011000000",
  10202=>"011111111",
  10203=>"000101111",
  10204=>"111100100",
  10205=>"011100000",
  10206=>"000000000",
  10207=>"001000111",
  10208=>"000111111",
  10209=>"000000000",
  10210=>"111111111",
  10211=>"000000111",
  10212=>"111000111",
  10213=>"011111111",
  10214=>"111111111",
  10215=>"011000010",
  10216=>"000000001",
  10217=>"000010011",
  10218=>"000000000",
  10219=>"101101100",
  10220=>"000000111",
  10221=>"000000000",
  10222=>"001111111",
  10223=>"000011111",
  10224=>"001000000",
  10225=>"111011011",
  10226=>"111000000",
  10227=>"000000110",
  10228=>"110110000",
  10229=>"111111111",
  10230=>"000000110",
  10231=>"111111100",
  10232=>"011111000",
  10233=>"000000001",
  10234=>"100111111",
  10235=>"111111000",
  10236=>"011111000",
  10237=>"000000000",
  10238=>"010011000",
  10239=>"001001111",
  10240=>"111111111",
  10241=>"000001000",
  10242=>"111000000",
  10243=>"000000000",
  10244=>"110100110",
  10245=>"000000100",
  10246=>"000011111",
  10247=>"100000000",
  10248=>"100000000",
  10249=>"111110110",
  10250=>"111111000",
  10251=>"111101001",
  10252=>"100100101",
  10253=>"100101111",
  10254=>"111111111",
  10255=>"111111000",
  10256=>"111100100",
  10257=>"011111111",
  10258=>"000000000",
  10259=>"000000000",
  10260=>"000000000",
  10261=>"111111110",
  10262=>"011111111",
  10263=>"100110111",
  10264=>"111100111",
  10265=>"000011011",
  10266=>"110111011",
  10267=>"001000000",
  10268=>"000000000",
  10269=>"000011110",
  10270=>"001011111",
  10271=>"000011111",
  10272=>"000000000",
  10273=>"111001000",
  10274=>"111111111",
  10275=>"011011011",
  10276=>"000000000",
  10277=>"111001000",
  10278=>"000000000",
  10279=>"111101011",
  10280=>"001101111",
  10281=>"110111111",
  10282=>"000000000",
  10283=>"111111111",
  10284=>"100000001",
  10285=>"000000000",
  10286=>"111110110",
  10287=>"101001001",
  10288=>"100000000",
  10289=>"000000000",
  10290=>"001000011",
  10291=>"100100111",
  10292=>"000000000",
  10293=>"100000000",
  10294=>"010111111",
  10295=>"111001001",
  10296=>"001000111",
  10297=>"001111111",
  10298=>"111111111",
  10299=>"111000000",
  10300=>"111111101",
  10301=>"111111111",
  10302=>"001000110",
  10303=>"000000000",
  10304=>"001000000",
  10305=>"001111111",
  10306=>"111111111",
  10307=>"001101111",
  10308=>"110110100",
  10309=>"001001111",
  10310=>"011010111",
  10311=>"000000000",
  10312=>"111110111",
  10313=>"111111111",
  10314=>"000000110",
  10315=>"010000111",
  10316=>"000000111",
  10317=>"111111100",
  10318=>"100100100",
  10319=>"000000000",
  10320=>"000001111",
  10321=>"111111111",
  10322=>"000000000",
  10323=>"111100001",
  10324=>"110111000",
  10325=>"110011001",
  10326=>"110110111",
  10327=>"000000001",
  10328=>"100000000",
  10329=>"000000100",
  10330=>"111101111",
  10331=>"001001001",
  10332=>"111111111",
  10333=>"011011000",
  10334=>"001001011",
  10335=>"000000000",
  10336=>"111111111",
  10337=>"000001011",
  10338=>"011000000",
  10339=>"000111111",
  10340=>"000000010",
  10341=>"010011110",
  10342=>"110110110",
  10343=>"111000000",
  10344=>"111111111",
  10345=>"111000000",
  10346=>"001000000",
  10347=>"111111111",
  10348=>"110101111",
  10349=>"111010010",
  10350=>"111111111",
  10351=>"011011011",
  10352=>"001000000",
  10353=>"000000000",
  10354=>"000010010",
  10355=>"000000001",
  10356=>"000000000",
  10357=>"011010010",
  10358=>"001001111",
  10359=>"000000000",
  10360=>"000000000",
  10361=>"001001000",
  10362=>"000000000",
  10363=>"000000000",
  10364=>"111111001",
  10365=>"000110110",
  10366=>"000000000",
  10367=>"101111111",
  10368=>"111101000",
  10369=>"111100000",
  10370=>"100110000",
  10371=>"110110111",
  10372=>"011111011",
  10373=>"110000000",
  10374=>"011101000",
  10375=>"001010000",
  10376=>"000000101",
  10377=>"011111111",
  10378=>"111100111",
  10379=>"000100000",
  10380=>"111001001",
  10381=>"100000000",
  10382=>"001000000",
  10383=>"110010010",
  10384=>"111000000",
  10385=>"011000010",
  10386=>"110110111",
  10387=>"111111111",
  10388=>"011000000",
  10389=>"110010000",
  10390=>"111000001",
  10391=>"000000000",
  10392=>"110111110",
  10393=>"000001001",
  10394=>"111111111",
  10395=>"000000000",
  10396=>"111111111",
  10397=>"000100000",
  10398=>"111101000",
  10399=>"111111111",
  10400=>"001000000",
  10401=>"000001111",
  10402=>"111101111",
  10403=>"000000000",
  10404=>"000110111",
  10405=>"111111111",
  10406=>"111111111",
  10407=>"000111110",
  10408=>"111111111",
  10409=>"000111111",
  10410=>"111110111",
  10411=>"111111001",
  10412=>"001111111",
  10413=>"111111111",
  10414=>"111111111",
  10415=>"000000000",
  10416=>"100100100",
  10417=>"111110110",
  10418=>"111111111",
  10419=>"110000111",
  10420=>"101000000",
  10421=>"010000000",
  10422=>"000000000",
  10423=>"111111111",
  10424=>"111011001",
  10425=>"111111111",
  10426=>"000000000",
  10427=>"101111111",
  10428=>"101000111",
  10429=>"011011001",
  10430=>"000000000",
  10431=>"111111010",
  10432=>"000110111",
  10433=>"000000000",
  10434=>"000000000",
  10435=>"111011011",
  10436=>"111111111",
  10437=>"111111111",
  10438=>"011011011",
  10439=>"000000110",
  10440=>"000011000",
  10441=>"111111111",
  10442=>"101111101",
  10443=>"000000001",
  10444=>"001000000",
  10445=>"000001000",
  10446=>"010000000",
  10447=>"000100010",
  10448=>"001011011",
  10449=>"011011011",
  10450=>"111001111",
  10451=>"010010000",
  10452=>"000000000",
  10453=>"111111111",
  10454=>"000000000",
  10455=>"111111111",
  10456=>"000000000",
  10457=>"111111000",
  10458=>"000000111",
  10459=>"111001000",
  10460=>"000000000",
  10461=>"000000111",
  10462=>"001111111",
  10463=>"001011000",
  10464=>"111001111",
  10465=>"000000000",
  10466=>"000000000",
  10467=>"000100000",
  10468=>"110110000",
  10469=>"110100100",
  10470=>"011011000",
  10471=>"111111111",
  10472=>"000000000",
  10473=>"000000010",
  10474=>"000000000",
  10475=>"011000100",
  10476=>"000000000",
  10477=>"110111111",
  10478=>"000111111",
  10479=>"000000000",
  10480=>"111000000",
  10481=>"011111111",
  10482=>"111100100",
  10483=>"000100100",
  10484=>"001111111",
  10485=>"110010000",
  10486=>"110110100",
  10487=>"000000000",
  10488=>"000000101",
  10489=>"111111111",
  10490=>"111001000",
  10491=>"111111111",
  10492=>"000101111",
  10493=>"011011001",
  10494=>"000001000",
  10495=>"010000000",
  10496=>"011111111",
  10497=>"100111110",
  10498=>"000000000",
  10499=>"100111111",
  10500=>"111111101",
  10501=>"111101100",
  10502=>"111111111",
  10503=>"000000000",
  10504=>"000000000",
  10505=>"111111111",
  10506=>"011000000",
  10507=>"111110111",
  10508=>"111111011",
  10509=>"111101101",
  10510=>"011011001",
  10511=>"000000000",
  10512=>"000010110",
  10513=>"100000100",
  10514=>"000000000",
  10515=>"111111111",
  10516=>"000001001",
  10517=>"111111000",
  10518=>"011111111",
  10519=>"111000000",
  10520=>"100100100",
  10521=>"000000100",
  10522=>"000000000",
  10523=>"111111111",
  10524=>"101100101",
  10525=>"111111111",
  10526=>"000111111",
  10527=>"000000000",
  10528=>"111111111",
  10529=>"111100111",
  10530=>"100000111",
  10531=>"111111111",
  10532=>"000000011",
  10533=>"000000100",
  10534=>"111111111",
  10535=>"101110000",
  10536=>"000000000",
  10537=>"110110000",
  10538=>"101101111",
  10539=>"000000000",
  10540=>"000000000",
  10541=>"001111110",
  10542=>"011111111",
  10543=>"000000000",
  10544=>"001000001",
  10545=>"111111111",
  10546=>"000000000",
  10547=>"100000001",
  10548=>"000000000",
  10549=>"001101000",
  10550=>"000000000",
  10551=>"111100010",
  10552=>"000000000",
  10553=>"000000000",
  10554=>"110010000",
  10555=>"000000000",
  10556=>"000000100",
  10557=>"101111111",
  10558=>"111101111",
  10559=>"111111111",
  10560=>"100111101",
  10561=>"111111111",
  10562=>"100111111",
  10563=>"100100101",
  10564=>"100011000",
  10565=>"111111111",
  10566=>"110111101",
  10567=>"011111011",
  10568=>"000000000",
  10569=>"000000000",
  10570=>"111111111",
  10571=>"100100110",
  10572=>"000000000",
  10573=>"111111111",
  10574=>"001000000",
  10575=>"000100100",
  10576=>"111111101",
  10577=>"000000000",
  10578=>"111110110",
  10579=>"100111111",
  10580=>"111111110",
  10581=>"011011011",
  10582=>"000000100",
  10583=>"111111111",
  10584=>"001111111",
  10585=>"000000100",
  10586=>"001000000",
  10587=>"000000001",
  10588=>"000000000",
  10589=>"111111111",
  10590=>"000000000",
  10591=>"111101111",
  10592=>"001010010",
  10593=>"111001001",
  10594=>"111111111",
  10595=>"000000100",
  10596=>"000111111",
  10597=>"000000000",
  10598=>"000000000",
  10599=>"000000000",
  10600=>"101111111",
  10601=>"000000000",
  10602=>"100100100",
  10603=>"111011111",
  10604=>"100111111",
  10605=>"000100100",
  10606=>"000000001",
  10607=>"100100111",
  10608=>"001111111",
  10609=>"111111111",
  10610=>"000000000",
  10611=>"110100100",
  10612=>"111111110",
  10613=>"000000011",
  10614=>"000000000",
  10615=>"010000001",
  10616=>"000000000",
  10617=>"111111111",
  10618=>"111111111",
  10619=>"000000101",
  10620=>"110100000",
  10621=>"100000111",
  10622=>"000011111",
  10623=>"111111111",
  10624=>"111111111",
  10625=>"011000000",
  10626=>"000011011",
  10627=>"111000101",
  10628=>"000010100",
  10629=>"000000000",
  10630=>"000000011",
  10631=>"100000000",
  10632=>"000000001",
  10633=>"111111111",
  10634=>"101000000",
  10635=>"110111111",
  10636=>"111111111",
  10637=>"011111111",
  10638=>"111101011",
  10639=>"011111111",
  10640=>"000000000",
  10641=>"000000000",
  10642=>"111101000",
  10643=>"100001111",
  10644=>"111111111",
  10645=>"000000010",
  10646=>"111001111",
  10647=>"000001011",
  10648=>"111111111",
  10649=>"111111000",
  10650=>"111101000",
  10651=>"111101111",
  10652=>"011000000",
  10653=>"101001101",
  10654=>"100000000",
  10655=>"111111111",
  10656=>"000000000",
  10657=>"111000000",
  10658=>"101001111",
  10659=>"111111111",
  10660=>"000100111",
  10661=>"000000000",
  10662=>"000000000",
  10663=>"000001000",
  10664=>"110000111",
  10665=>"110000000",
  10666=>"000000111",
  10667=>"100100000",
  10668=>"000010110",
  10669=>"111111111",
  10670=>"011111110",
  10671=>"000000000",
  10672=>"111111000",
  10673=>"100000000",
  10674=>"000011001",
  10675=>"000000011",
  10676=>"110101001",
  10677=>"000110010",
  10678=>"111000000",
  10679=>"000000000",
  10680=>"111111111",
  10681=>"110100100",
  10682=>"000111110",
  10683=>"111111111",
  10684=>"000000000",
  10685=>"111010000",
  10686=>"100000100",
  10687=>"001001000",
  10688=>"100111111",
  10689=>"001001011",
  10690=>"000000100",
  10691=>"111111111",
  10692=>"101101111",
  10693=>"010111111",
  10694=>"111111011",
  10695=>"000000011",
  10696=>"000000111",
  10697=>"000100100",
  10698=>"000110010",
  10699=>"000000000",
  10700=>"000000010",
  10701=>"000000000",
  10702=>"111111111",
  10703=>"101111111",
  10704=>"111111111",
  10705=>"100101101",
  10706=>"000000000",
  10707=>"000010000",
  10708=>"000000000",
  10709=>"000000000",
  10710=>"111111000",
  10711=>"011011011",
  10712=>"100100000",
  10713=>"110111111",
  10714=>"000000000",
  10715=>"100000110",
  10716=>"000000011",
  10717=>"001001100",
  10718=>"000000011",
  10719=>"000000000",
  10720=>"001011011",
  10721=>"111111011",
  10722=>"000011011",
  10723=>"000000000",
  10724=>"100111111",
  10725=>"000000111",
  10726=>"000000000",
  10727=>"000000011",
  10728=>"111101001",
  10729=>"111111111",
  10730=>"100110110",
  10731=>"111111111",
  10732=>"111000000",
  10733=>"001110110",
  10734=>"100001001",
  10735=>"000000000",
  10736=>"000100000",
  10737=>"000000000",
  10738=>"111111111",
  10739=>"000000000",
  10740=>"000011111",
  10741=>"100000001",
  10742=>"000000111",
  10743=>"010010110",
  10744=>"000001000",
  10745=>"001001110",
  10746=>"000000000",
  10747=>"000110111",
  10748=>"000100001",
  10749=>"011001000",
  10750=>"000110000",
  10751=>"000000000",
  10752=>"000011000",
  10753=>"111001111",
  10754=>"111101111",
  10755=>"111111001",
  10756=>"000110000",
  10757=>"111111111",
  10758=>"111111000",
  10759=>"111111111",
  10760=>"000111101",
  10761=>"111101000",
  10762=>"111111010",
  10763=>"000000000",
  10764=>"000000000",
  10765=>"110111111",
  10766=>"100000111",
  10767=>"111011000",
  10768=>"000000111",
  10769=>"000100111",
  10770=>"000000010",
  10771=>"000000000",
  10772=>"000111111",
  10773=>"000000000",
  10774=>"000000111",
  10775=>"101110100",
  10776=>"110010000",
  10777=>"011011000",
  10778=>"000110111",
  10779=>"111101001",
  10780=>"111111000",
  10781=>"111000111",
  10782=>"110100100",
  10783=>"000000000",
  10784=>"000000000",
  10785=>"110110110",
  10786=>"000000111",
  10787=>"001000000",
  10788=>"001000001",
  10789=>"110110000",
  10790=>"111111111",
  10791=>"110111100",
  10792=>"111111001",
  10793=>"000000010",
  10794=>"000101111",
  10795=>"111111111",
  10796=>"000000111",
  10797=>"000000111",
  10798=>"101111111",
  10799=>"111011010",
  10800=>"000000000",
  10801=>"110110000",
  10802=>"000100000",
  10803=>"100111111",
  10804=>"111111111",
  10805=>"000000100",
  10806=>"111100100",
  10807=>"001000000",
  10808=>"000000111",
  10809=>"110000000",
  10810=>"000000000",
  10811=>"101101111",
  10812=>"111111111",
  10813=>"000111111",
  10814=>"110111101",
  10815=>"000000100",
  10816=>"000100111",
  10817=>"011111100",
  10818=>"000000000",
  10819=>"000000000",
  10820=>"000000000",
  10821=>"100110111",
  10822=>"111111111",
  10823=>"111111111",
  10824=>"011010000",
  10825=>"110111000",
  10826=>"111111111",
  10827=>"001000000",
  10828=>"001001000",
  10829=>"000000110",
  10830=>"110110111",
  10831=>"100000000",
  10832=>"000000110",
  10833=>"011000000",
  10834=>"000000000",
  10835=>"001100101",
  10836=>"000000000",
  10837=>"111111110",
  10838=>"111001001",
  10839=>"000000111",
  10840=>"111111011",
  10841=>"111000001",
  10842=>"000000000",
  10843=>"110110100",
  10844=>"000101000",
  10845=>"000000000",
  10846=>"111110111",
  10847=>"100111111",
  10848=>"000000000",
  10849=>"111111011",
  10850=>"111111111",
  10851=>"000000000",
  10852=>"010010010",
  10853=>"000000111",
  10854=>"111111000",
  10855=>"111111000",
  10856=>"011111001",
  10857=>"111111111",
  10858=>"000000010",
  10859=>"111000000",
  10860=>"011010000",
  10861=>"111111000",
  10862=>"111111111",
  10863=>"110111000",
  10864=>"010111111",
  10865=>"000001111",
  10866=>"111111111",
  10867=>"111011011",
  10868=>"000000000",
  10869=>"101001100",
  10870=>"111001111",
  10871=>"111111000",
  10872=>"000000000",
  10873=>"000000000",
  10874=>"111111111",
  10875=>"010011011",
  10876=>"111111110",
  10877=>"101111011",
  10878=>"101000000",
  10879=>"011111111",
  10880=>"000000010",
  10881=>"111000000",
  10882=>"111111111",
  10883=>"000011111",
  10884=>"000000000",
  10885=>"000111111",
  10886=>"001110100",
  10887=>"000000010",
  10888=>"011001011",
  10889=>"011111111",
  10890=>"000000000",
  10891=>"111101000",
  10892=>"101000000",
  10893=>"000011000",
  10894=>"110111111",
  10895=>"111001000",
  10896=>"111111111",
  10897=>"110010010",
  10898=>"000000110",
  10899=>"000000011",
  10900=>"000000111",
  10901=>"000111001",
  10902=>"111111000",
  10903=>"111111100",
  10904=>"111101111",
  10905=>"111111001",
  10906=>"100111111",
  10907=>"111000111",
  10908=>"111111000",
  10909=>"000000000",
  10910=>"111111001",
  10911=>"111000000",
  10912=>"111101111",
  10913=>"001101111",
  10914=>"001111111",
  10915=>"000000100",
  10916=>"111001000",
  10917=>"000000100",
  10918=>"111111000",
  10919=>"111111011",
  10920=>"010000000",
  10921=>"110000000",
  10922=>"111101000",
  10923=>"111000000",
  10924=>"111111111",
  10925=>"000000000",
  10926=>"001000100",
  10927=>"000000010",
  10928=>"001011000",
  10929=>"001011011",
  10930=>"110110110",
  10931=>"111111101",
  10932=>"111111111",
  10933=>"111111111",
  10934=>"000000010",
  10935=>"000000001",
  10936=>"111000110",
  10937=>"000000111",
  10938=>"011001001",
  10939=>"000000111",
  10940=>"000000111",
  10941=>"000111111",
  10942=>"100100100",
  10943=>"000000000",
  10944=>"000000100",
  10945=>"111111111",
  10946=>"000001111",
  10947=>"010000111",
  10948=>"110000000",
  10949=>"000000000",
  10950=>"011011101",
  10951=>"111000000",
  10952=>"111111111",
  10953=>"111000000",
  10954=>"111000110",
  10955=>"111111110",
  10956=>"101101111",
  10957=>"000001111",
  10958=>"110111100",
  10959=>"100000000",
  10960=>"111111010",
  10961=>"011010110",
  10962=>"111111111",
  10963=>"000000110",
  10964=>"111011010",
  10965=>"000000111",
  10966=>"011111111",
  10967=>"111010000",
  10968=>"111111111",
  10969=>"101111111",
  10970=>"111110000",
  10971=>"111100111",
  10972=>"001000001",
  10973=>"111101001",
  10974=>"011110111",
  10975=>"001000100",
  10976=>"000000000",
  10977=>"011110111",
  10978=>"001111111",
  10979=>"111011000",
  10980=>"000000111",
  10981=>"011011001",
  10982=>"000000101",
  10983=>"000000101",
  10984=>"000000000",
  10985=>"001111111",
  10986=>"011000000",
  10987=>"111111111",
  10988=>"000011000",
  10989=>"000110111",
  10990=>"000010000",
  10991=>"000000000",
  10992=>"000111001",
  10993=>"100000000",
  10994=>"000000000",
  10995=>"001111111",
  10996=>"111111000",
  10997=>"101111111",
  10998=>"001101100",
  10999=>"000000101",
  11000=>"000000000",
  11001=>"000000000",
  11002=>"000000111",
  11003=>"000000011",
  11004=>"111111000",
  11005=>"101001111",
  11006=>"000000000",
  11007=>"111001000",
  11008=>"000000000",
  11009=>"011011001",
  11010=>"000000110",
  11011=>"111000000",
  11012=>"000000111",
  11013=>"000000000",
  11014=>"000000001",
  11015=>"110111111",
  11016=>"110100101",
  11017=>"010010010",
  11018=>"000000000",
  11019=>"101111111",
  11020=>"110110110",
  11021=>"111111011",
  11022=>"100000000",
  11023=>"000000111",
  11024=>"100110111",
  11025=>"100100000",
  11026=>"111111000",
  11027=>"000001101",
  11028=>"000000000",
  11029=>"111111111",
  11030=>"100100000",
  11031=>"110111111",
  11032=>"101111111",
  11033=>"000000000",
  11034=>"111111110",
  11035=>"111001011",
  11036=>"000111000",
  11037=>"000111100",
  11038=>"000000010",
  11039=>"100111000",
  11040=>"100111111",
  11041=>"001001001",
  11042=>"101111111",
  11043=>"000000100",
  11044=>"011011111",
  11045=>"000000111",
  11046=>"101011000",
  11047=>"111111000",
  11048=>"111111111",
  11049=>"000000000",
  11050=>"000101110",
  11051=>"100111111",
  11052=>"000000000",
  11053=>"000001011",
  11054=>"010111111",
  11055=>"111011000",
  11056=>"001010111",
  11057=>"000110110",
  11058=>"111000100",
  11059=>"000010000",
  11060=>"000000000",
  11061=>"100100111",
  11062=>"111110111",
  11063=>"111111000",
  11064=>"111111001",
  11065=>"111001111",
  11066=>"111110000",
  11067=>"000111111",
  11068=>"000000000",
  11069=>"000000000",
  11070=>"000000111",
  11071=>"000011000",
  11072=>"011000000",
  11073=>"111111111",
  11074=>"000000111",
  11075=>"001100000",
  11076=>"101010010",
  11077=>"111010000",
  11078=>"000001000",
  11079=>"011001111",
  11080=>"011100000",
  11081=>"001000000",
  11082=>"101110110",
  11083=>"001001111",
  11084=>"000000111",
  11085=>"000000110",
  11086=>"000100110",
  11087=>"100000000",
  11088=>"100000100",
  11089=>"111111100",
  11090=>"110010111",
  11091=>"111000000",
  11092=>"000000000",
  11093=>"001000000",
  11094=>"111110111",
  11095=>"111111101",
  11096=>"111111111",
  11097=>"000000000",
  11098=>"000000111",
  11099=>"000100110",
  11100=>"000000000",
  11101=>"111111111",
  11102=>"001111111",
  11103=>"111110111",
  11104=>"101001011",
  11105=>"111000000",
  11106=>"111011001",
  11107=>"010000000",
  11108=>"100110110",
  11109=>"111111011",
  11110=>"000000000",
  11111=>"000100111",
  11112=>"100110110",
  11113=>"000010000",
  11114=>"000100000",
  11115=>"000000000",
  11116=>"101101001",
  11117=>"111000001",
  11118=>"000000000",
  11119=>"111111010",
  11120=>"011011111",
  11121=>"111011001",
  11122=>"100000000",
  11123=>"001000001",
  11124=>"000100100",
  11125=>"111000000",
  11126=>"111000000",
  11127=>"110100110",
  11128=>"111111011",
  11129=>"111111111",
  11130=>"100000000",
  11131=>"111111111",
  11132=>"011000111",
  11133=>"000000000",
  11134=>"111111111",
  11135=>"111000000",
  11136=>"110100110",
  11137=>"111101000",
  11138=>"001011111",
  11139=>"000000110",
  11140=>"010111111",
  11141=>"111110011",
  11142=>"010111110",
  11143=>"111100111",
  11144=>"000011111",
  11145=>"011011011",
  11146=>"000011101",
  11147=>"111111111",
  11148=>"111001001",
  11149=>"000000000",
  11150=>"110111111",
  11151=>"110111111",
  11152=>"011111111",
  11153=>"011110110",
  11154=>"001111011",
  11155=>"100011000",
  11156=>"111111111",
  11157=>"000010110",
  11158=>"011000000",
  11159=>"001011010",
  11160=>"000000000",
  11161=>"111111011",
  11162=>"001000000",
  11163=>"101111011",
  11164=>"000000011",
  11165=>"000000111",
  11166=>"000111111",
  11167=>"000110010",
  11168=>"000000000",
  11169=>"111111100",
  11170=>"000000111",
  11171=>"011101000",
  11172=>"001000011",
  11173=>"111000000",
  11174=>"000000000",
  11175=>"000000110",
  11176=>"000000000",
  11177=>"111111111",
  11178=>"000100100",
  11179=>"100100111",
  11180=>"000000000",
  11181=>"000000000",
  11182=>"000001101",
  11183=>"100000001",
  11184=>"111111110",
  11185=>"000000000",
  11186=>"000000111",
  11187=>"100100111",
  11188=>"000011111",
  11189=>"111001111",
  11190=>"001111111",
  11191=>"111111111",
  11192=>"100111111",
  11193=>"000111111",
  11194=>"111111100",
  11195=>"000001111",
  11196=>"111111111",
  11197=>"111011001",
  11198=>"111111111",
  11199=>"011001001",
  11200=>"100110110",
  11201=>"000000000",
  11202=>"111111111",
  11203=>"000010100",
  11204=>"001000101",
  11205=>"111111000",
  11206=>"110000111",
  11207=>"010011111",
  11208=>"111111111",
  11209=>"000000000",
  11210=>"000000100",
  11211=>"000111111",
  11212=>"111111111",
  11213=>"111111111",
  11214=>"111011011",
  11215=>"111111111",
  11216=>"000000011",
  11217=>"100111111",
  11218=>"000000001",
  11219=>"000000000",
  11220=>"001001000",
  11221=>"001000000",
  11222=>"000000000",
  11223=>"000001100",
  11224=>"111111100",
  11225=>"100001001",
  11226=>"111111000",
  11227=>"000000000",
  11228=>"001001001",
  11229=>"101111111",
  11230=>"101000111",
  11231=>"000001011",
  11232=>"000000000",
  11233=>"011111111",
  11234=>"000011001",
  11235=>"111001000",
  11236=>"110110110",
  11237=>"111111111",
  11238=>"110000011",
  11239=>"000111111",
  11240=>"000000001",
  11241=>"101111111",
  11242=>"110110000",
  11243=>"000000000",
  11244=>"111001110",
  11245=>"000000000",
  11246=>"000001111",
  11247=>"000000000",
  11248=>"001000010",
  11249=>"100111111",
  11250=>"100000000",
  11251=>"111111111",
  11252=>"101111111",
  11253=>"111111111",
  11254=>"111111011",
  11255=>"111111001",
  11256=>"000000110",
  11257=>"011001001",
  11258=>"111101000",
  11259=>"111111111",
  11260=>"001000000",
  11261=>"100100100",
  11262=>"000100111",
  11263=>"111111100",
  11264=>"111111011",
  11265=>"000000000",
  11266=>"111111111",
  11267=>"111111011",
  11268=>"111111111",
  11269=>"000000000",
  11270=>"000000000",
  11271=>"111111111",
  11272=>"000000011",
  11273=>"011010000",
  11274=>"100101111",
  11275=>"001011111",
  11276=>"000000100",
  11277=>"111111111",
  11278=>"000000001",
  11279=>"011010000",
  11280=>"001110111",
  11281=>"111001000",
  11282=>"000000000",
  11283=>"111111111",
  11284=>"000000000",
  11285=>"111000001",
  11286=>"111111000",
  11287=>"000000111",
  11288=>"001101111",
  11289=>"001001101",
  11290=>"000000000",
  11291=>"111111101",
  11292=>"000000000",
  11293=>"111111111",
  11294=>"000100100",
  11295=>"111001000",
  11296=>"000000110",
  11297=>"111111111",
  11298=>"111101111",
  11299=>"111110110",
  11300=>"000100111",
  11301=>"000111110",
  11302=>"000100111",
  11303=>"000010000",
  11304=>"101111111",
  11305=>"000000000",
  11306=>"000111111",
  11307=>"001001100",
  11308=>"110000000",
  11309=>"010111000",
  11310=>"100000000",
  11311=>"000000000",
  11312=>"111101001",
  11313=>"000000000",
  11314=>"000011011",
  11315=>"000000000",
  11316=>"001001111",
  11317=>"000000001",
  11318=>"000000111",
  11319=>"111111011",
  11320=>"000000010",
  11321=>"101001100",
  11322=>"000000000",
  11323=>"111111111",
  11324=>"000001111",
  11325=>"110100000",
  11326=>"100110110",
  11327=>"111011000",
  11328=>"000000000",
  11329=>"000000000",
  11330=>"001001000",
  11331=>"000000000",
  11332=>"000000000",
  11333=>"111110111",
  11334=>"000000000",
  11335=>"101100111",
  11336=>"110111111",
  11337=>"000000000",
  11338=>"111111111",
  11339=>"111111001",
  11340=>"000011011",
  11341=>"100100101",
  11342=>"101100111",
  11343=>"000000000",
  11344=>"010000000",
  11345=>"001011000",
  11346=>"000011010",
  11347=>"000000111",
  11348=>"111101001",
  11349=>"111010111",
  11350=>"100111100",
  11351=>"000000100",
  11352=>"000000010",
  11353=>"000000000",
  11354=>"010010000",
  11355=>"001011011",
  11356=>"110000000",
  11357=>"000110111",
  11358=>"111111111",
  11359=>"111111001",
  11360=>"111111101",
  11361=>"111001000",
  11362=>"000000000",
  11363=>"000000000",
  11364=>"111101111",
  11365=>"111111111",
  11366=>"111000111",
  11367=>"000111111",
  11368=>"111000111",
  11369=>"000100000",
  11370=>"001001000",
  11371=>"000000110",
  11372=>"011011111",
  11373=>"000000111",
  11374=>"110111111",
  11375=>"000000000",
  11376=>"000100001",
  11377=>"001011000",
  11378=>"111111111",
  11379=>"000101111",
  11380=>"101100000",
  11381=>"000000111",
  11382=>"000000101",
  11383=>"000000001",
  11384=>"110111111",
  11385=>"111111111",
  11386=>"111011111",
  11387=>"111111101",
  11388=>"001001001",
  11389=>"000110111",
  11390=>"000010111",
  11391=>"111111101",
  11392=>"001000000",
  11393=>"000000000",
  11394=>"000000000",
  11395=>"100110111",
  11396=>"111111111",
  11397=>"000000000",
  11398=>"110111111",
  11399=>"111111111",
  11400=>"111111000",
  11401=>"010010000",
  11402=>"011000000",
  11403=>"000000010",
  11404=>"111111111",
  11405=>"101000000",
  11406=>"001000000",
  11407=>"011001111",
  11408=>"000000000",
  11409=>"111111111",
  11410=>"000010000",
  11411=>"000110000",
  11412=>"000000001",
  11413=>"111111111",
  11414=>"000011111",
  11415=>"011111000",
  11416=>"111000000",
  11417=>"000000111",
  11418=>"000111111",
  11419=>"111111000",
  11420=>"111011000",
  11421=>"000000111",
  11422=>"011110110",
  11423=>"011001001",
  11424=>"000000000",
  11425=>"011000001",
  11426=>"111000000",
  11427=>"101101111",
  11428=>"000000100",
  11429=>"111000000",
  11430=>"011111111",
  11431=>"111100100",
  11432=>"000000000",
  11433=>"000000000",
  11434=>"111111111",
  11435=>"111111001",
  11436=>"011001111",
  11437=>"011111001",
  11438=>"000011001",
  11439=>"111111001",
  11440=>"000000000",
  11441=>"111111111",
  11442=>"111111111",
  11443=>"000110111",
  11444=>"000000000",
  11445=>"000000000",
  11446=>"000000000",
  11447=>"111000000",
  11448=>"011011111",
  11449=>"111111100",
  11450=>"110000000",
  11451=>"000010000",
  11452=>"000000000",
  11453=>"010110110",
  11454=>"000000000",
  11455=>"100000000",
  11456=>"110110110",
  11457=>"000000011",
  11458=>"001111111",
  11459=>"000001001",
  11460=>"001001000",
  11461=>"101100000",
  11462=>"000000000",
  11463=>"111111111",
  11464=>"111111011",
  11465=>"000000000",
  11466=>"001001001",
  11467=>"111011010",
  11468=>"011001000",
  11469=>"001001001",
  11470=>"001000010",
  11471=>"110000111",
  11472=>"000110111",
  11473=>"000000000",
  11474=>"000011101",
  11475=>"000000000",
  11476=>"111001001",
  11477=>"001111101",
  11478=>"111111000",
  11479=>"000111111",
  11480=>"001111111",
  11481=>"111111111",
  11482=>"111111100",
  11483=>"111111001",
  11484=>"110110111",
  11485=>"000101111",
  11486=>"000000111",
  11487=>"011000110",
  11488=>"000000000",
  11489=>"000000000",
  11490=>"111111111",
  11491=>"011011000",
  11492=>"101000101",
  11493=>"011110100",
  11494=>"111111111",
  11495=>"111111111",
  11496=>"111000111",
  11497=>"001001011",
  11498=>"111000000",
  11499=>"111111111",
  11500=>"000000000",
  11501=>"000000111",
  11502=>"001001001",
  11503=>"001000000",
  11504=>"111111111",
  11505=>"111011000",
  11506=>"000011000",
  11507=>"000000110",
  11508=>"000010110",
  11509=>"100000100",
  11510=>"111110110",
  11511=>"000000000",
  11512=>"000001001",
  11513=>"011001011",
  11514=>"111111111",
  11515=>"111111111",
  11516=>"101001011",
  11517=>"011011111",
  11518=>"110000110",
  11519=>"110000100",
  11520=>"010111010",
  11521=>"001010000",
  11522=>"111111100",
  11523=>"000110110",
  11524=>"010011011",
  11525=>"111111000",
  11526=>"100111001",
  11527=>"001001011",
  11528=>"111111111",
  11529=>"000001011",
  11530=>"111111011",
  11531=>"101110111",
  11532=>"100100100",
  11533=>"111111100",
  11534=>"000000011",
  11535=>"110111111",
  11536=>"101000000",
  11537=>"000111111",
  11538=>"100100110",
  11539=>"000001000",
  11540=>"111111000",
  11541=>"100101111",
  11542=>"111111000",
  11543=>"110111111",
  11544=>"110111111",
  11545=>"000000000",
  11546=>"000001111",
  11547=>"000000000",
  11548=>"100100100",
  11549=>"110011000",
  11550=>"000000000",
  11551=>"010111101",
  11552=>"100100111",
  11553=>"111010100",
  11554=>"000100111",
  11555=>"000100011",
  11556=>"000000000",
  11557=>"110110000",
  11558=>"100000000",
  11559=>"000000000",
  11560=>"111101000",
  11561=>"111011001",
  11562=>"111001000",
  11563=>"000111010",
  11564=>"100000111",
  11565=>"001011111",
  11566=>"000111000",
  11567=>"011111111",
  11568=>"011011011",
  11569=>"111001101",
  11570=>"110000000",
  11571=>"011000000",
  11572=>"110001111",
  11573=>"001001000",
  11574=>"000000000",
  11575=>"000110111",
  11576=>"000000000",
  11577=>"111111101",
  11578=>"011000101",
  11579=>"000111000",
  11580=>"000000000",
  11581=>"010010011",
  11582=>"000000000",
  11583=>"111101111",
  11584=>"000000000",
  11585=>"010100111",
  11586=>"111111111",
  11587=>"000000000",
  11588=>"110110001",
  11589=>"001001000",
  11590=>"111000010",
  11591=>"111000000",
  11592=>"011111111",
  11593=>"100000000",
  11594=>"000000000",
  11595=>"010111111",
  11596=>"000110111",
  11597=>"000001111",
  11598=>"000111111",
  11599=>"000001000",
  11600=>"011000000",
  11601=>"000000000",
  11602=>"000000000",
  11603=>"111111111",
  11604=>"000000101",
  11605=>"100100100",
  11606=>"010000110",
  11607=>"000000001",
  11608=>"001000000",
  11609=>"111111111",
  11610=>"001000001",
  11611=>"111111000",
  11612=>"000000000",
  11613=>"111101100",
  11614=>"000000000",
  11615=>"111111110",
  11616=>"111001111",
  11617=>"110000000",
  11618=>"000001001",
  11619=>"001000000",
  11620=>"000100110",
  11621=>"111111000",
  11622=>"000000000",
  11623=>"100011111",
  11624=>"000110110",
  11625=>"000100000",
  11626=>"101000101",
  11627=>"000111111",
  11628=>"011001011",
  11629=>"000000111",
  11630=>"000000000",
  11631=>"011111010",
  11632=>"000001101",
  11633=>"111110111",
  11634=>"111111111",
  11635=>"001000101",
  11636=>"110111110",
  11637=>"000000001",
  11638=>"000000110",
  11639=>"000000101",
  11640=>"111110000",
  11641=>"000000000",
  11642=>"111111111",
  11643=>"000000000",
  11644=>"100100111",
  11645=>"110111111",
  11646=>"100000000",
  11647=>"010000000",
  11648=>"011000000",
  11649=>"111000010",
  11650=>"000000111",
  11651=>"000100111",
  11652=>"101100000",
  11653=>"111111111",
  11654=>"000000100",
  11655=>"000000000",
  11656=>"000000000",
  11657=>"000000000",
  11658=>"000001001",
  11659=>"000000000",
  11660=>"000001001",
  11661=>"111111111",
  11662=>"000100000",
  11663=>"011001011",
  11664=>"111110100",
  11665=>"111110100",
  11666=>"111111111",
  11667=>"110000000",
  11668=>"111111111",
  11669=>"100000000",
  11670=>"100100000",
  11671=>"000011000",
  11672=>"111111111",
  11673=>"111100000",
  11674=>"100110100",
  11675=>"000110111",
  11676=>"111011111",
  11677=>"111111111",
  11678=>"111101111",
  11679=>"000010000",
  11680=>"000111111",
  11681=>"011011001",
  11682=>"001110000",
  11683=>"000011011",
  11684=>"000000100",
  11685=>"111111111",
  11686=>"100100100",
  11687=>"111110111",
  11688=>"000000011",
  11689=>"111100110",
  11690=>"000010100",
  11691=>"110111111",
  11692=>"000000000",
  11693=>"111101001",
  11694=>"001000110",
  11695=>"000000101",
  11696=>"110000000",
  11697=>"000000000",
  11698=>"001000000",
  11699=>"000000000",
  11700=>"111111100",
  11701=>"111001111",
  11702=>"000010011",
  11703=>"010000000",
  11704=>"000000000",
  11705=>"000000000",
  11706=>"111101000",
  11707=>"011011110",
  11708=>"000000101",
  11709=>"000000000",
  11710=>"000000000",
  11711=>"111111000",
  11712=>"011000000",
  11713=>"100000000",
  11714=>"111010000",
  11715=>"110000000",
  11716=>"001011001",
  11717=>"000111110",
  11718=>"000000000",
  11719=>"011000000",
  11720=>"000000010",
  11721=>"111111000",
  11722=>"000000000",
  11723=>"000001000",
  11724=>"000111111",
  11725=>"111111111",
  11726=>"000000000",
  11727=>"111111110",
  11728=>"011000000",
  11729=>"000000000",
  11730=>"111111111",
  11731=>"111111111",
  11732=>"111001011",
  11733=>"101110111",
  11734=>"101101111",
  11735=>"000000001",
  11736=>"001111111",
  11737=>"111101111",
  11738=>"110100000",
  11739=>"011111111",
  11740=>"111000000",
  11741=>"001011000",
  11742=>"100111111",
  11743=>"110000000",
  11744=>"000000000",
  11745=>"000000000",
  11746=>"100100000",
  11747=>"000000001",
  11748=>"000101101",
  11749=>"111000111",
  11750=>"000101111",
  11751=>"000111100",
  11752=>"011010000",
  11753=>"111111000",
  11754=>"000111111",
  11755=>"111111001",
  11756=>"111001001",
  11757=>"001111011",
  11758=>"001111011",
  11759=>"111111010",
  11760=>"111111111",
  11761=>"000000000",
  11762=>"111000000",
  11763=>"001000000",
  11764=>"111111101",
  11765=>"111111111",
  11766=>"110110100",
  11767=>"000000100",
  11768=>"000000000",
  11769=>"011011111",
  11770=>"000000000",
  11771=>"111111111",
  11772=>"001000000",
  11773=>"000101000",
  11774=>"000000000",
  11775=>"000000000",
  11776=>"001111111",
  11777=>"000011111",
  11778=>"111101111",
  11779=>"000000000",
  11780=>"001011011",
  11781=>"000000000",
  11782=>"110111110",
  11783=>"111101001",
  11784=>"110110111",
  11785=>"000111011",
  11786=>"111110000",
  11787=>"000001000",
  11788=>"100100000",
  11789=>"011011011",
  11790=>"111111111",
  11791=>"000000000",
  11792=>"001001011",
  11793=>"110110111",
  11794=>"111111111",
  11795=>"000000000",
  11796=>"000110110",
  11797=>"011000001",
  11798=>"111000000",
  11799=>"111111001",
  11800=>"110000000",
  11801=>"000000101",
  11802=>"101000000",
  11803=>"110100000",
  11804=>"111111100",
  11805=>"100110110",
  11806=>"111000000",
  11807=>"100100110",
  11808=>"000110111",
  11809=>"111001000",
  11810=>"111111110",
  11811=>"000000000",
  11812=>"111111111",
  11813=>"011001111",
  11814=>"111111111",
  11815=>"000000000",
  11816=>"011111111",
  11817=>"110100000",
  11818=>"110111111",
  11819=>"111111111",
  11820=>"001000000",
  11821=>"111111111",
  11822=>"011111111",
  11823=>"110100100",
  11824=>"000000111",
  11825=>"111111111",
  11826=>"111111011",
  11827=>"010110100",
  11828=>"001111111",
  11829=>"010001001",
  11830=>"001000001",
  11831=>"000000000",
  11832=>"100110000",
  11833=>"010000000",
  11834=>"010111111",
  11835=>"000000000",
  11836=>"000000111",
  11837=>"000000000",
  11838=>"000000000",
  11839=>"000011111",
  11840=>"010100100",
  11841=>"011011111",
  11842=>"000001000",
  11843=>"111000000",
  11844=>"000000111",
  11845=>"111000010",
  11846=>"110110100",
  11847=>"111111000",
  11848=>"000100110",
  11849=>"000110111",
  11850=>"000111111",
  11851=>"111111111",
  11852=>"001001011",
  11853=>"000000000",
  11854=>"101111011",
  11855=>"000000000",
  11856=>"000110110",
  11857=>"111111111",
  11858=>"111000000",
  11859=>"000000000",
  11860=>"000000000",
  11861=>"110110100",
  11862=>"111101001",
  11863=>"111111111",
  11864=>"111111011",
  11865=>"000000000",
  11866=>"000000000",
  11867=>"010000000",
  11868=>"111111111",
  11869=>"000000111",
  11870=>"100000000",
  11871=>"111001111",
  11872=>"000101111",
  11873=>"000000000",
  11874=>"000000100",
  11875=>"000000000",
  11876=>"101000000",
  11877=>"111100100",
  11878=>"110110111",
  11879=>"111111111",
  11880=>"000010000",
  11881=>"100000111",
  11882=>"110110000",
  11883=>"000000110",
  11884=>"000000000",
  11885=>"000000111",
  11886=>"111100000",
  11887=>"010110110",
  11888=>"000000000",
  11889=>"011111111",
  11890=>"111100111",
  11891=>"000000000",
  11892=>"000000011",
  11893=>"000111111",
  11894=>"000010000",
  11895=>"000000000",
  11896=>"000000000",
  11897=>"111111000",
  11898=>"100000000",
  11899=>"111001000",
  11900=>"111011011",
  11901=>"111111000",
  11902=>"000000000",
  11903=>"000000000",
  11904=>"000000000",
  11905=>"111011011",
  11906=>"001111100",
  11907=>"000000000",
  11908=>"110111111",
  11909=>"000000000",
  11910=>"110110111",
  11911=>"111111111",
  11912=>"111111111",
  11913=>"110000000",
  11914=>"110111000",
  11915=>"011111000",
  11916=>"111101111",
  11917=>"111111010",
  11918=>"011000000",
  11919=>"111111111",
  11920=>"000000001",
  11921=>"000000001",
  11922=>"000000000",
  11923=>"111000000",
  11924=>"000100100",
  11925=>"110110110",
  11926=>"011011010",
  11927=>"000000000",
  11928=>"100000100",
  11929=>"111111111",
  11930=>"111011111",
  11931=>"000000001",
  11932=>"000000101",
  11933=>"111000000",
  11934=>"000000000",
  11935=>"000000000",
  11936=>"000100100",
  11937=>"001111111",
  11938=>"111111111",
  11939=>"110000110",
  11940=>"001001001",
  11941=>"100110111",
  11942=>"101000000",
  11943=>"000000000",
  11944=>"110111010",
  11945=>"000000000",
  11946=>"111110100",
  11947=>"101000001",
  11948=>"011001000",
  11949=>"000000000",
  11950=>"000000111",
  11951=>"000000000",
  11952=>"111110111",
  11953=>"111111001",
  11954=>"111111111",
  11955=>"001101111",
  11956=>"000010110",
  11957=>"001000000",
  11958=>"000100110",
  11959=>"110010000",
  11960=>"111110111",
  11961=>"110000110",
  11962=>"101001101",
  11963=>"000000000",
  11964=>"100000000",
  11965=>"000000000",
  11966=>"011111111",
  11967=>"111111000",
  11968=>"011001011",
  11969=>"100111111",
  11970=>"000001111",
  11971=>"111111111",
  11972=>"000000000",
  11973=>"110111110",
  11974=>"111111111",
  11975=>"111111111",
  11976=>"000000100",
  11977=>"111111111",
  11978=>"101000001",
  11979=>"011011111",
  11980=>"000000000",
  11981=>"001111011",
  11982=>"001111111",
  11983=>"000000100",
  11984=>"111001011",
  11985=>"111111111",
  11986=>"000011111",
  11987=>"111111100",
  11988=>"111111100",
  11989=>"001000000",
  11990=>"000000110",
  11991=>"111001000",
  11992=>"000000000",
  11993=>"000000000",
  11994=>"111111111",
  11995=>"000000110",
  11996=>"111011000",
  11997=>"100000000",
  11998=>"000000111",
  11999=>"010000000",
  12000=>"011000000",
  12001=>"000000000",
  12002=>"000000000",
  12003=>"110110000",
  12004=>"111111001",
  12005=>"011000011",
  12006=>"111111101",
  12007=>"111111111",
  12008=>"000001111",
  12009=>"111000000",
  12010=>"000000101",
  12011=>"000000000",
  12012=>"011001001",
  12013=>"100100110",
  12014=>"011000000",
  12015=>"000000111",
  12016=>"000000000",
  12017=>"000000000",
  12018=>"000010000",
  12019=>"000000000",
  12020=>"111111111",
  12021=>"100110000",
  12022=>"110111111",
  12023=>"000111100",
  12024=>"000001111",
  12025=>"001001101",
  12026=>"000000100",
  12027=>"111000000",
  12028=>"001000000",
  12029=>"110100000",
  12030=>"111110100",
  12031=>"000000000",
  12032=>"111111000",
  12033=>"110110000",
  12034=>"100110111",
  12035=>"111110000",
  12036=>"000111000",
  12037=>"111111111",
  12038=>"000111011",
  12039=>"111000111",
  12040=>"111111111",
  12041=>"000000000",
  12042=>"000000000",
  12043=>"111111010",
  12044=>"001001000",
  12045=>"000100001",
  12046=>"001111111",
  12047=>"111001000",
  12048=>"111111111",
  12049=>"000000000",
  12050=>"111100100",
  12051=>"000000000",
  12052=>"110010011",
  12053=>"000100111",
  12054=>"111111011",
  12055=>"111111011",
  12056=>"001011111",
  12057=>"111111011",
  12058=>"000000000",
  12059=>"010001001",
  12060=>"111000000",
  12061=>"000000111",
  12062=>"111111111",
  12063=>"000001111",
  12064=>"001000000",
  12065=>"111111111",
  12066=>"000000000",
  12067=>"000000000",
  12068=>"111001000",
  12069=>"010000000",
  12070=>"111111111",
  12071=>"000100100",
  12072=>"000000000",
  12073=>"110100100",
  12074=>"000100000",
  12075=>"000000110",
  12076=>"110111111",
  12077=>"111111011",
  12078=>"111111111",
  12079=>"000000000",
  12080=>"100100111",
  12081=>"111110000",
  12082=>"111111111",
  12083=>"001000000",
  12084=>"000000100",
  12085=>"101100100",
  12086=>"001111111",
  12087=>"101101111",
  12088=>"000000000",
  12089=>"110000111",
  12090=>"111110100",
  12091=>"010010000",
  12092=>"010000100",
  12093=>"000111111",
  12094=>"111011001",
  12095=>"111000001",
  12096=>"011001001",
  12097=>"110100000",
  12098=>"000000000",
  12099=>"101111111",
  12100=>"111111110",
  12101=>"011111111",
  12102=>"000000010",
  12103=>"000000000",
  12104=>"000000001",
  12105=>"000000100",
  12106=>"110010000",
  12107=>"101100101",
  12108=>"010011011",
  12109=>"001001111",
  12110=>"111111111",
  12111=>"001001011",
  12112=>"000000110",
  12113=>"100110000",
  12114=>"111111111",
  12115=>"101111101",
  12116=>"111111111",
  12117=>"001011010",
  12118=>"111111111",
  12119=>"111111001",
  12120=>"110111111",
  12121=>"000000000",
  12122=>"000000011",
  12123=>"000000000",
  12124=>"111000000",
  12125=>"000000000",
  12126=>"000000000",
  12127=>"111111000",
  12128=>"111111000",
  12129=>"111111101",
  12130=>"000000000",
  12131=>"000000101",
  12132=>"100000000",
  12133=>"000011000",
  12134=>"000000111",
  12135=>"000000000",
  12136=>"100100100",
  12137=>"000001111",
  12138=>"000000000",
  12139=>"010010110",
  12140=>"000001011",
  12141=>"000111011",
  12142=>"111111011",
  12143=>"011001000",
  12144=>"110111111",
  12145=>"000110100",
  12146=>"000000011",
  12147=>"111111011",
  12148=>"001000000",
  12149=>"011101111",
  12150=>"000000000",
  12151=>"111010001",
  12152=>"000000000",
  12153=>"111111011",
  12154=>"111111011",
  12155=>"000000001",
  12156=>"111111111",
  12157=>"111101101",
  12158=>"000000101",
  12159=>"000000000",
  12160=>"100111000",
  12161=>"001111111",
  12162=>"000000000",
  12163=>"100110100",
  12164=>"000000000",
  12165=>"111000000",
  12166=>"001001000",
  12167=>"111001000",
  12168=>"000000001",
  12169=>"000100111",
  12170=>"111110101",
  12171=>"000100100",
  12172=>"111111111",
  12173=>"001001000",
  12174=>"000000001",
  12175=>"000000001",
  12176=>"111111111",
  12177=>"010001110",
  12178=>"001001001",
  12179=>"111011011",
  12180=>"111111111",
  12181=>"000000000",
  12182=>"111110000",
  12183=>"001011010",
  12184=>"110100000",
  12185=>"110101110",
  12186=>"000000000",
  12187=>"111111000",
  12188=>"111111000",
  12189=>"001000000",
  12190=>"111111111",
  12191=>"110010000",
  12192=>"000000000",
  12193=>"100000000",
  12194=>"010010000",
  12195=>"011011000",
  12196=>"000001000",
  12197=>"000011111",
  12198=>"100000000",
  12199=>"111011011",
  12200=>"100000000",
  12201=>"100111111",
  12202=>"111000000",
  12203=>"001001111",
  12204=>"111111111",
  12205=>"000100110",
  12206=>"101101000",
  12207=>"111011111",
  12208=>"101101001",
  12209=>"111000000",
  12210=>"000001111",
  12211=>"110111111",
  12212=>"111111111",
  12213=>"000000000",
  12214=>"000000000",
  12215=>"111111000",
  12216=>"000000000",
  12217=>"100111111",
  12218=>"011000000",
  12219=>"001001001",
  12220=>"000000000",
  12221=>"000000000",
  12222=>"000101000",
  12223=>"101101101",
  12224=>"011111000",
  12225=>"111111111",
  12226=>"000000111",
  12227=>"000011011",
  12228=>"000000000",
  12229=>"111001001",
  12230=>"000000000",
  12231=>"110110010",
  12232=>"000000000",
  12233=>"001000000",
  12234=>"000000001",
  12235=>"000001000",
  12236=>"111000010",
  12237=>"001000111",
  12238=>"001101111",
  12239=>"110111011",
  12240=>"011000000",
  12241=>"000000001",
  12242=>"011111111",
  12243=>"000000000",
  12244=>"000000111",
  12245=>"000000000",
  12246=>"111111001",
  12247=>"010110000",
  12248=>"111111111",
  12249=>"000000000",
  12250=>"100000110",
  12251=>"111111111",
  12252=>"110101111",
  12253=>"010000111",
  12254=>"111101111",
  12255=>"000000000",
  12256=>"110110110",
  12257=>"000000000",
  12258=>"011111111",
  12259=>"001111111",
  12260=>"000000000",
  12261=>"111000100",
  12262=>"001000001",
  12263=>"000000110",
  12264=>"110101100",
  12265=>"011111111",
  12266=>"100101011",
  12267=>"000000000",
  12268=>"111011111",
  12269=>"111110110",
  12270=>"111101110",
  12271=>"010010011",
  12272=>"111111111",
  12273=>"000000011",
  12274=>"000100000",
  12275=>"000000111",
  12276=>"000000000",
  12277=>"000000001",
  12278=>"111100000",
  12279=>"001111110",
  12280=>"111001000",
  12281=>"011011011",
  12282=>"000000000",
  12283=>"000000000",
  12284=>"100111111",
  12285=>"100111110",
  12286=>"010111111",
  12287=>"001001111",
  12288=>"000010010",
  12289=>"000000111",
  12290=>"111111111",
  12291=>"101001000",
  12292=>"010011000",
  12293=>"111001000",
  12294=>"000000111",
  12295=>"000111011",
  12296=>"011111111",
  12297=>"000011110",
  12298=>"000000000",
  12299=>"000100100",
  12300=>"111111011",
  12301=>"001000000",
  12302=>"111100101",
  12303=>"111111111",
  12304=>"000001000",
  12305=>"111111000",
  12306=>"000000000",
  12307=>"011000101",
  12308=>"111010000",
  12309=>"000111011",
  12310=>"000111111",
  12311=>"001111111",
  12312=>"100110111",
  12313=>"001000001",
  12314=>"101100100",
  12315=>"111111111",
  12316=>"000000000",
  12317=>"111111110",
  12318=>"110111100",
  12319=>"000011000",
  12320=>"011110111",
  12321=>"000000000",
  12322=>"001111001",
  12323=>"111111000",
  12324=>"111111111",
  12325=>"111111001",
  12326=>"000000000",
  12327=>"000000000",
  12328=>"000000000",
  12329=>"000000110",
  12330=>"111111111",
  12331=>"110110110",
  12332=>"000000110",
  12333=>"111111100",
  12334=>"111000000",
  12335=>"111100111",
  12336=>"011000000",
  12337=>"000111111",
  12338=>"001011011",
  12339=>"100000000",
  12340=>"111111111",
  12341=>"000001001",
  12342=>"000000010",
  12343=>"010010000",
  12344=>"011001000",
  12345=>"000010000",
  12346=>"111000011",
  12347=>"011000000",
  12348=>"111011110",
  12349=>"110000000",
  12350=>"000000000",
  12351=>"000000000",
  12352=>"011100110",
  12353=>"101100100",
  12354=>"000111111",
  12355=>"000000000",
  12356=>"111111111",
  12357=>"000000011",
  12358=>"000111111",
  12359=>"011011000",
  12360=>"111000000",
  12361=>"111000111",
  12362=>"000001111",
  12363=>"010110111",
  12364=>"000000000",
  12365=>"000110110",
  12366=>"000001101",
  12367=>"101111111",
  12368=>"000000000",
  12369=>"000000000",
  12370=>"111111110",
  12371=>"111110111",
  12372=>"000000000",
  12373=>"100110110",
  12374=>"000000000",
  12375=>"000000000",
  12376=>"000000110",
  12377=>"111001000",
  12378=>"011011111",
  12379=>"011000010",
  12380=>"111111000",
  12381=>"111000000",
  12382=>"011011001",
  12383=>"110110100",
  12384=>"111110100",
  12385=>"000100111",
  12386=>"111000100",
  12387=>"111111111",
  12388=>"001001000",
  12389=>"000111111",
  12390=>"111111011",
  12391=>"110111110",
  12392=>"111000101",
  12393=>"111111111",
  12394=>"000000000",
  12395=>"100000000",
  12396=>"011011111",
  12397=>"111111110",
  12398=>"110000111",
  12399=>"000000000",
  12400=>"010000000",
  12401=>"000001001",
  12402=>"101101101",
  12403=>"010000111",
  12404=>"111110000",
  12405=>"111000100",
  12406=>"111111111",
  12407=>"111111111",
  12408=>"000110111",
  12409=>"100000110",
  12410=>"110100000",
  12411=>"110111000",
  12412=>"011011011",
  12413=>"111111111",
  12414=>"000000111",
  12415=>"000110111",
  12416=>"111000000",
  12417=>"110111011",
  12418=>"111110111",
  12419=>"100100000",
  12420=>"000000001",
  12421=>"111110111",
  12422=>"000001011",
  12423=>"111111110",
  12424=>"001000000",
  12425=>"000000000",
  12426=>"111111111",
  12427=>"000001111",
  12428=>"000000000",
  12429=>"000110000",
  12430=>"010000000",
  12431=>"000101000",
  12432=>"100101111",
  12433=>"111100000",
  12434=>"000000000",
  12435=>"010110110",
  12436=>"110110000",
  12437=>"011000110",
  12438=>"000000011",
  12439=>"111000001",
  12440=>"000000000",
  12441=>"000110100",
  12442=>"111111000",
  12443=>"111111101",
  12444=>"000000001",
  12445=>"000000111",
  12446=>"001000001",
  12447=>"111110111",
  12448=>"000000000",
  12449=>"001001001",
  12450=>"110000001",
  12451=>"000010110",
  12452=>"111001001",
  12453=>"111111111",
  12454=>"101111111",
  12455=>"000111110",
  12456=>"111111001",
  12457=>"000111110",
  12458=>"111111101",
  12459=>"100100101",
  12460=>"000000000",
  12461=>"110110000",
  12462=>"111111000",
  12463=>"111001111",
  12464=>"111111111",
  12465=>"000000111",
  12466=>"111111001",
  12467=>"111111111",
  12468=>"000000010",
  12469=>"000000111",
  12470=>"111111111",
  12471=>"000111001",
  12472=>"010010111",
  12473=>"110110111",
  12474=>"100000000",
  12475=>"111110110",
  12476=>"111000000",
  12477=>"000000000",
  12478=>"010111111",
  12479=>"011111111",
  12480=>"100101111",
  12481=>"000000000",
  12482=>"000000000",
  12483=>"111111111",
  12484=>"110000000",
  12485=>"111111111",
  12486=>"000000011",
  12487=>"000000100",
  12488=>"000000001",
  12489=>"111001001",
  12490=>"110101111",
  12491=>"000000100",
  12492=>"111110110",
  12493=>"100001001",
  12494=>"111111111",
  12495=>"111000000",
  12496=>"100000111",
  12497=>"001000100",
  12498=>"010011111",
  12499=>"000000000",
  12500=>"111100000",
  12501=>"000110110",
  12502=>"111000000",
  12503=>"000001000",
  12504=>"110110000",
  12505=>"011110110",
  12506=>"000111111",
  12507=>"110111111",
  12508=>"010111110",
  12509=>"111111111",
  12510=>"111111111",
  12511=>"000010011",
  12512=>"100000000",
  12513=>"001111000",
  12514=>"111001000",
  12515=>"001001101",
  12516=>"001010111",
  12517=>"100000111",
  12518=>"000000111",
  12519=>"000000110",
  12520=>"111111111",
  12521=>"000000111",
  12522=>"000000110",
  12523=>"001110010",
  12524=>"000001111",
  12525=>"101000110",
  12526=>"111111111",
  12527=>"000000000",
  12528=>"000000111",
  12529=>"111111111",
  12530=>"000000000",
  12531=>"100000000",
  12532=>"000111111",
  12533=>"011011010",
  12534=>"000011111",
  12535=>"000000000",
  12536=>"111111111",
  12537=>"000000011",
  12538=>"011000000",
  12539=>"000000000",
  12540=>"110110000",
  12541=>"111011010",
  12542=>"000000000",
  12543=>"110000000",
  12544=>"000000011",
  12545=>"100100100",
  12546=>"110111110",
  12547=>"000110100",
  12548=>"000000000",
  12549=>"000011111",
  12550=>"111000100",
  12551=>"000000000",
  12552=>"111111000",
  12553=>"000000000",
  12554=>"111000000",
  12555=>"000000111",
  12556=>"001001111",
  12557=>"110110110",
  12558=>"000001111",
  12559=>"111111111",
  12560=>"000110111",
  12561=>"111000011",
  12562=>"111011111",
  12563=>"110000000",
  12564=>"000000011",
  12565=>"111111111",
  12566=>"001001001",
  12567=>"111111111",
  12568=>"111011011",
  12569=>"111111000",
  12570=>"111000000",
  12571=>"011110111",
  12572=>"000000110",
  12573=>"111111111",
  12574=>"000000111",
  12575=>"111000001",
  12576=>"000000001",
  12577=>"000000000",
  12578=>"111111000",
  12579=>"011100111",
  12580=>"100000010",
  12581=>"000101001",
  12582=>"111111111",
  12583=>"101101111",
  12584=>"111111111",
  12585=>"001000000",
  12586=>"110000001",
  12587=>"010000000",
  12588=>"100000111",
  12589=>"000010000",
  12590=>"000000111",
  12591=>"000000101",
  12592=>"000100000",
  12593=>"100110000",
  12594=>"000111111",
  12595=>"111011000",
  12596=>"000000000",
  12597=>"000101101",
  12598=>"000010010",
  12599=>"000000001",
  12600=>"111111111",
  12601=>"011111111",
  12602=>"001000111",
  12603=>"001000000",
  12604=>"011000100",
  12605=>"000000000",
  12606=>"111110110",
  12607=>"000000111",
  12608=>"111111000",
  12609=>"111111100",
  12610=>"111111111",
  12611=>"000000000",
  12612=>"000111111",
  12613=>"000000000",
  12614=>"110111000",
  12615=>"111111111",
  12616=>"000100111",
  12617=>"011000011",
  12618=>"111000111",
  12619=>"010011000",
  12620=>"001110111",
  12621=>"000110000",
  12622=>"001111001",
  12623=>"000011001",
  12624=>"000001011",
  12625=>"000001111",
  12626=>"001000010",
  12627=>"000110111",
  12628=>"000101000",
  12629=>"111111110",
  12630=>"111010111",
  12631=>"011000110",
  12632=>"001000011",
  12633=>"100111111",
  12634=>"000010111",
  12635=>"110000111",
  12636=>"000001001",
  12637=>"101000000",
  12638=>"111001001",
  12639=>"111111111",
  12640=>"000000011",
  12641=>"000111111",
  12642=>"111111111",
  12643=>"101111110",
  12644=>"000000000",
  12645=>"101001111",
  12646=>"111111100",
  12647=>"011110111",
  12648=>"001101011",
  12649=>"110000010",
  12650=>"111111111",
  12651=>"000001001",
  12652=>"001001011",
  12653=>"110110110",
  12654=>"000000000",
  12655=>"000000110",
  12656=>"111111011",
  12657=>"000000111",
  12658=>"110111111",
  12659=>"110100111",
  12660=>"000000000",
  12661=>"000000111",
  12662=>"000000000",
  12663=>"111111111",
  12664=>"000000110",
  12665=>"000000000",
  12666=>"000000110",
  12667=>"000100100",
  12668=>"000000000",
  12669=>"011111101",
  12670=>"000000000",
  12671=>"010011111",
  12672=>"111111111",
  12673=>"110000000",
  12674=>"000000100",
  12675=>"111111111",
  12676=>"100111111",
  12677=>"111000000",
  12678=>"000111111",
  12679=>"111100000",
  12680=>"111111010",
  12681=>"111111100",
  12682=>"000000000",
  12683=>"000011011",
  12684=>"110010000",
  12685=>"111111111",
  12686=>"000000000",
  12687=>"000000000",
  12688=>"000000001",
  12689=>"011001100",
  12690=>"111111011",
  12691=>"110111111",
  12692=>"010111111",
  12693=>"000010000",
  12694=>"000000111",
  12695=>"000000011",
  12696=>"111111111",
  12697=>"000010010",
  12698=>"111000000",
  12699=>"111101000",
  12700=>"111111111",
  12701=>"110010111",
  12702=>"000001000",
  12703=>"111110111",
  12704=>"111001000",
  12705=>"000100110",
  12706=>"100100100",
  12707=>"000111111",
  12708=>"110000111",
  12709=>"111001001",
  12710=>"111101111",
  12711=>"111111110",
  12712=>"101001111",
  12713=>"111110110",
  12714=>"111000000",
  12715=>"001001111",
  12716=>"000001001",
  12717=>"000111110",
  12718=>"000111111",
  12719=>"011000000",
  12720=>"111011010",
  12721=>"111111111",
  12722=>"000000111",
  12723=>"000001111",
  12724=>"111111111",
  12725=>"111111000",
  12726=>"111010001",
  12727=>"111000000",
  12728=>"111101110",
  12729=>"111111111",
  12730=>"000000000",
  12731=>"111011011",
  12732=>"000000001",
  12733=>"110000000",
  12734=>"001000001",
  12735=>"111000000",
  12736=>"111111111",
  12737=>"001001111",
  12738=>"000000000",
  12739=>"111111001",
  12740=>"011001001",
  12741=>"000001111",
  12742=>"100110111",
  12743=>"110000000",
  12744=>"111111111",
  12745=>"000000100",
  12746=>"000000001",
  12747=>"110000000",
  12748=>"100111000",
  12749=>"000000111",
  12750=>"000100111",
  12751=>"111111111",
  12752=>"000111111",
  12753=>"000000011",
  12754=>"000000110",
  12755=>"111111111",
  12756=>"100111111",
  12757=>"000000000",
  12758=>"000000100",
  12759=>"111000000",
  12760=>"000100100",
  12761=>"000000000",
  12762=>"000000010",
  12763=>"000000000",
  12764=>"000000001",
  12765=>"000000000",
  12766=>"111111111",
  12767=>"001001111",
  12768=>"000111111",
  12769=>"111111111",
  12770=>"000100100",
  12771=>"000001001",
  12772=>"111000000",
  12773=>"000000000",
  12774=>"011100111",
  12775=>"111111000",
  12776=>"011000000",
  12777=>"111111111",
  12778=>"111111110",
  12779=>"000001001",
  12780=>"000111111",
  12781=>"100111011",
  12782=>"011001000",
  12783=>"111100000",
  12784=>"000000111",
  12785=>"000011011",
  12786=>"111111000",
  12787=>"111111001",
  12788=>"110110000",
  12789=>"110100100",
  12790=>"000110111",
  12791=>"000010110",
  12792=>"111111000",
  12793=>"000011001",
  12794=>"111111111",
  12795=>"100110111",
  12796=>"101000100",
  12797=>"111110111",
  12798=>"000001000",
  12799=>"011001111",
  12800=>"110111111",
  12801=>"111001001",
  12802=>"111101111",
  12803=>"111111111",
  12804=>"000100000",
  12805=>"101101111",
  12806=>"101101100",
  12807=>"111111111",
  12808=>"111111111",
  12809=>"110110110",
  12810=>"000000000",
  12811=>"111111000",
  12812=>"001001001",
  12813=>"000110000",
  12814=>"010011100",
  12815=>"101101111",
  12816=>"000110110",
  12817=>"001000111",
  12818=>"000000111",
  12819=>"000000000",
  12820=>"011001001",
  12821=>"111111111",
  12822=>"000000010",
  12823=>"001001000",
  12824=>"101111111",
  12825=>"001001101",
  12826=>"001101001",
  12827=>"111111111",
  12828=>"010000000",
  12829=>"111111001",
  12830=>"000000001",
  12831=>"000000000",
  12832=>"111111111",
  12833=>"000000000",
  12834=>"001001011",
  12835=>"111111100",
  12836=>"000000111",
  12837=>"000000110",
  12838=>"000000000",
  12839=>"001000000",
  12840=>"001000000",
  12841=>"101001101",
  12842=>"111000111",
  12843=>"000000111",
  12844=>"001001111",
  12845=>"001000000",
  12846=>"000000100",
  12847=>"111111000",
  12848=>"111110111",
  12849=>"000001000",
  12850=>"001100100",
  12851=>"000000110",
  12852=>"000001101",
  12853=>"110110000",
  12854=>"110111001",
  12855=>"001001110",
  12856=>"110000000",
  12857=>"001000111",
  12858=>"101101101",
  12859=>"111101000",
  12860=>"111111111",
  12861=>"011001001",
  12862=>"001001111",
  12863=>"100100100",
  12864=>"011111100",
  12865=>"001101111",
  12866=>"001000100",
  12867=>"001101111",
  12868=>"110110100",
  12869=>"110111011",
  12870=>"101000001",
  12871=>"110111100",
  12872=>"000111101",
  12873=>"000001101",
  12874=>"111111011",
  12875=>"110000000",
  12876=>"000001010",
  12877=>"011001001",
  12878=>"010010000",
  12879=>"000000101",
  12880=>"010111111",
  12881=>"111110000",
  12882=>"111111111",
  12883=>"110100001",
  12884=>"001000001",
  12885=>"010111111",
  12886=>"000001001",
  12887=>"110010010",
  12888=>"111110000",
  12889=>"111111111",
  12890=>"000000111",
  12891=>"000100001",
  12892=>"001000010",
  12893=>"000011001",
  12894=>"001001001",
  12895=>"000010011",
  12896=>"000011000",
  12897=>"000000101",
  12898=>"000000000",
  12899=>"100101000",
  12900=>"000000110",
  12901=>"111011001",
  12902=>"110110000",
  12903=>"111111111",
  12904=>"000000001",
  12905=>"111111111",
  12906=>"001000111",
  12907=>"101101000",
  12908=>"000001001",
  12909=>"000000001",
  12910=>"101001001",
  12911=>"000000100",
  12912=>"110111000",
  12913=>"111110001",
  12914=>"110111000",
  12915=>"000110111",
  12916=>"000000101",
  12917=>"001001000",
  12918=>"111101101",
  12919=>"110100000",
  12920=>"110110110",
  12921=>"000110110",
  12922=>"001001001",
  12923=>"001001000",
  12924=>"110110110",
  12925=>"000000111",
  12926=>"111001000",
  12927=>"011111111",
  12928=>"010111100",
  12929=>"000000001",
  12930=>"000000000",
  12931=>"000100100",
  12932=>"111001001",
  12933=>"111101111",
  12934=>"111111111",
  12935=>"001001111",
  12936=>"000100000",
  12937=>"111110010",
  12938=>"000000100",
  12939=>"101100000",
  12940=>"010110100",
  12941=>"110110111",
  12942=>"001001001",
  12943=>"100111110",
  12944=>"000000110",
  12945=>"000010111",
  12946=>"000101111",
  12947=>"011001100",
  12948=>"000000001",
  12949=>"100111111",
  12950=>"101001001",
  12951=>"111001111",
  12952=>"111111001",
  12953=>"111010000",
  12954=>"010110001",
  12955=>"101100001",
  12956=>"111111111",
  12957=>"110110110",
  12958=>"110110111",
  12959=>"111111111",
  12960=>"111101111",
  12961=>"000000100",
  12962=>"100101000",
  12963=>"110111000",
  12964=>"110111000",
  12965=>"101000000",
  12966=>"110111000",
  12967=>"111111000",
  12968=>"111000001",
  12969=>"001001000",
  12970=>"101000101",
  12971=>"001001001",
  12972=>"110110110",
  12973=>"000000111",
  12974=>"111101110",
  12975=>"000001100",
  12976=>"111000111",
  12977=>"000000110",
  12978=>"110111010",
  12979=>"011111000",
  12980=>"000000101",
  12981=>"000000101",
  12982=>"010000110",
  12983=>"111100100",
  12984=>"000000000",
  12985=>"111101111",
  12986=>"111000001",
  12987=>"110001001",
  12988=>"011000000",
  12989=>"010010111",
  12990=>"000000000",
  12991=>"111111111",
  12992=>"110000010",
  12993=>"110111110",
  12994=>"000000101",
  12995=>"111011101",
  12996=>"000111111",
  12997=>"011001111",
  12998=>"111001101",
  12999=>"010110101",
  13000=>"101101000",
  13001=>"001001111",
  13002=>"000000111",
  13003=>"101101100",
  13004=>"111111111",
  13005=>"111111110",
  13006=>"001001111",
  13007=>"000000111",
  13008=>"100100010",
  13009=>"101101101",
  13010=>"110110111",
  13011=>"000001101",
  13012=>"110111011",
  13013=>"010000111",
  13014=>"010111001",
  13015=>"111101111",
  13016=>"111111111",
  13017=>"001000100",
  13018=>"000001011",
  13019=>"010010111",
  13020=>"110110110",
  13021=>"000111111",
  13022=>"000000000",
  13023=>"010011010",
  13024=>"001000001",
  13025=>"111101111",
  13026=>"111111111",
  13027=>"000000001",
  13028=>"001000000",
  13029=>"001001001",
  13030=>"001000111",
  13031=>"000000000",
  13032=>"101111001",
  13033=>"010001001",
  13034=>"100110110",
  13035=>"101001101",
  13036=>"000000000",
  13037=>"111111010",
  13038=>"100001001",
  13039=>"001111000",
  13040=>"000001011",
  13041=>"110111000",
  13042=>"100000000",
  13043=>"110001000",
  13044=>"001000000",
  13045=>"000100110",
  13046=>"011111100",
  13047=>"000111111",
  13048=>"001101100",
  13049=>"101101101",
  13050=>"110000111",
  13051=>"001100000",
  13052=>"000010000",
  13053=>"000011011",
  13054=>"001000000",
  13055=>"111000000",
  13056=>"001000100",
  13057=>"011001001",
  13058=>"111111111",
  13059=>"001001000",
  13060=>"111111100",
  13061=>"111101000",
  13062=>"110100100",
  13063=>"111111001",
  13064=>"111110000",
  13065=>"101001001",
  13066=>"011111101",
  13067=>"011000000",
  13068=>"111101111",
  13069=>"110110110",
  13070=>"111111100",
  13071=>"100100100",
  13072=>"111110110",
  13073=>"100110111",
  13074=>"010010010",
  13075=>"001000100",
  13076=>"000000000",
  13077=>"100110010",
  13078=>"001000001",
  13079=>"111110000",
  13080=>"001000110",
  13081=>"000001001",
  13082=>"100111011",
  13083=>"001001111",
  13084=>"011001001",
  13085=>"111111101",
  13086=>"001101111",
  13087=>"000001111",
  13088=>"010111111",
  13089=>"010010010",
  13090=>"111111111",
  13091=>"001111001",
  13092=>"000000010",
  13093=>"000000100",
  13094=>"000000000",
  13095=>"011000110",
  13096=>"000000111",
  13097=>"111111000",
  13098=>"000000000",
  13099=>"001001000",
  13100=>"001001100",
  13101=>"110110110",
  13102=>"001000000",
  13103=>"111110000",
  13104=>"110110111",
  13105=>"000001001",
  13106=>"000000000",
  13107=>"000100100",
  13108=>"010111000",
  13109=>"111100111",
  13110=>"111111101",
  13111=>"111011000",
  13112=>"000111000",
  13113=>"101101111",
  13114=>"000001001",
  13115=>"110111011",
  13116=>"000000000",
  13117=>"000000000",
  13118=>"110100110",
  13119=>"010010000",
  13120=>"000001000",
  13121=>"000100111",
  13122=>"000000111",
  13123=>"101000110",
  13124=>"100110000",
  13125=>"000000101",
  13126=>"000000111",
  13127=>"001000000",
  13128=>"101101101",
  13129=>"000000000",
  13130=>"001010110",
  13131=>"000001001",
  13132=>"000000111",
  13133=>"000000100",
  13134=>"001000111",
  13135=>"110110110",
  13136=>"011010000",
  13137=>"011110111",
  13138=>"110110000",
  13139=>"111111110",
  13140=>"000001000",
  13141=>"001001001",
  13142=>"010000110",
  13143=>"101001111",
  13144=>"001001001",
  13145=>"111010000",
  13146=>"000110110",
  13147=>"111111101",
  13148=>"111111111",
  13149=>"000010011",
  13150=>"110110110",
  13151=>"111111111",
  13152=>"111111000",
  13153=>"000110011",
  13154=>"001000000",
  13155=>"111111011",
  13156=>"110110010",
  13157=>"000011111",
  13158=>"111110000",
  13159=>"000010000",
  13160=>"001001101",
  13161=>"000111111",
  13162=>"000000111",
  13163=>"001111110",
  13164=>"000000001",
  13165=>"111001111",
  13166=>"000000111",
  13167=>"000000100",
  13168=>"000000010",
  13169=>"000110111",
  13170=>"111111101",
  13171=>"001001110",
  13172=>"111111111",
  13173=>"111111110",
  13174=>"000000000",
  13175=>"110010000",
  13176=>"000000000",
  13177=>"000100111",
  13178=>"000000001",
  13179=>"110111111",
  13180=>"110110000",
  13181=>"000010000",
  13182=>"010111010",
  13183=>"101101101",
  13184=>"000110111",
  13185=>"111000000",
  13186=>"111110100",
  13187=>"101001101",
  13188=>"010000000",
  13189=>"110111010",
  13190=>"001000000",
  13191=>"000000000",
  13192=>"000000000",
  13193=>"010000011",
  13194=>"001101111",
  13195=>"000000001",
  13196=>"000000111",
  13197=>"000000000",
  13198=>"000100101",
  13199=>"111010000",
  13200=>"001111000",
  13201=>"000001001",
  13202=>"111110000",
  13203=>"000000001",
  13204=>"111000000",
  13205=>"000000111",
  13206=>"001000000",
  13207=>"110111000",
  13208=>"000101100",
  13209=>"000110110",
  13210=>"111111001",
  13211=>"111000100",
  13212=>"111111011",
  13213=>"000000000",
  13214=>"000111111",
  13215=>"001011000",
  13216=>"111111111",
  13217=>"001011011",
  13218=>"111011001",
  13219=>"110111001",
  13220=>"110111101",
  13221=>"000110110",
  13222=>"111001000",
  13223=>"011111111",
  13224=>"001101101",
  13225=>"000010111",
  13226=>"000000000",
  13227=>"101001101",
  13228=>"000011001",
  13229=>"000000000",
  13230=>"100000110",
  13231=>"011100110",
  13232=>"101101111",
  13233=>"000000111",
  13234=>"001001000",
  13235=>"011001111",
  13236=>"010110101",
  13237=>"011001011",
  13238=>"111111111",
  13239=>"000111001",
  13240=>"000111001",
  13241=>"111010100",
  13242=>"000001111",
  13243=>"110110111",
  13244=>"001001001",
  13245=>"111111000",
  13246=>"001001111",
  13247=>"011000011",
  13248=>"010000000",
  13249=>"101111111",
  13250=>"111111111",
  13251=>"000001000",
  13252=>"001000001",
  13253=>"110010111",
  13254=>"001000101",
  13255=>"000101111",
  13256=>"001000000",
  13257=>"010000000",
  13258=>"001000101",
  13259=>"101111111",
  13260=>"111101000",
  13261=>"111111000",
  13262=>"110111101",
  13263=>"110111011",
  13264=>"000100110",
  13265=>"111001111",
  13266=>"111000111",
  13267=>"111101111",
  13268=>"000000000",
  13269=>"110110100",
  13270=>"001101111",
  13271=>"100000000",
  13272=>"111110110",
  13273=>"111111110",
  13274=>"111111000",
  13275=>"000000000",
  13276=>"000000000",
  13277=>"111111111",
  13278=>"111011001",
  13279=>"000110010",
  13280=>"101001111",
  13281=>"000000110",
  13282=>"000000000",
  13283=>"111111000",
  13284=>"110111101",
  13285=>"110111101",
  13286=>"110110111",
  13287=>"111111000",
  13288=>"000010110",
  13289=>"000000000",
  13290=>"000011111",
  13291=>"000110110",
  13292=>"011111111",
  13293=>"000001000",
  13294=>"000000010",
  13295=>"000001001",
  13296=>"001000000",
  13297=>"101111111",
  13298=>"100111111",
  13299=>"111111001",
  13300=>"000000110",
  13301=>"110110010",
  13302=>"111101110",
  13303=>"000000011",
  13304=>"111111111",
  13305=>"101001101",
  13306=>"000000110",
  13307=>"000111000",
  13308=>"101000001",
  13309=>"001100111",
  13310=>"110110111",
  13311=>"100101111",
  13312=>"011001001",
  13313=>"000000111",
  13314=>"111111111",
  13315=>"111011001",
  13316=>"111101111",
  13317=>"001000000",
  13318=>"000000100",
  13319=>"111111111",
  13320=>"110000100",
  13321=>"000000111",
  13322=>"000100100",
  13323=>"111111110",
  13324=>"000100100",
  13325=>"000000011",
  13326=>"110110110",
  13327=>"000000111",
  13328=>"000000000",
  13329=>"111111011",
  13330=>"111110101",
  13331=>"000000000",
  13332=>"111111101",
  13333=>"000000101",
  13334=>"100000000",
  13335=>"100101111",
  13336=>"000000000",
  13337=>"000100111",
  13338=>"000000000",
  13339=>"011111111",
  13340=>"111111000",
  13341=>"000000011",
  13342=>"110100000",
  13343=>"110111111",
  13344=>"000110000",
  13345=>"001001000",
  13346=>"111111111",
  13347=>"111111111",
  13348=>"000000110",
  13349=>"000000001",
  13350=>"111111000",
  13351=>"000000100",
  13352=>"111001000",
  13353=>"000000000",
  13354=>"100000000",
  13355=>"000001111",
  13356=>"000000000",
  13357=>"000000000",
  13358=>"000000000",
  13359=>"110111011",
  13360=>"000000001",
  13361=>"111111111",
  13362=>"110101111",
  13363=>"111111000",
  13364=>"111111100",
  13365=>"000000000",
  13366=>"100100111",
  13367=>"011011000",
  13368=>"011000000",
  13369=>"000000100",
  13370=>"000000000",
  13371=>"100000000",
  13372=>"000000111",
  13373=>"111111100",
  13374=>"000111111",
  13375=>"000001000",
  13376=>"001110000",
  13377=>"110111111",
  13378=>"000000000",
  13379=>"000000000",
  13380=>"100110111",
  13381=>"000000100",
  13382=>"101000000",
  13383=>"111001001",
  13384=>"010111111",
  13385=>"000000000",
  13386=>"000000000",
  13387=>"111111100",
  13388=>"000000000",
  13389=>"000000111",
  13390=>"000000110",
  13391=>"111111111",
  13392=>"000000000",
  13393=>"011011111",
  13394=>"100100100",
  13395=>"111111111",
  13396=>"000000111",
  13397=>"110111111",
  13398=>"101101101",
  13399=>"111011011",
  13400=>"111111110",
  13401=>"101100110",
  13402=>"011111111",
  13403=>"011111110",
  13404=>"111000000",
  13405=>"111111111",
  13406=>"001000000",
  13407=>"110110100",
  13408=>"000000000",
  13409=>"000000000",
  13410=>"111111101",
  13411=>"111111000",
  13412=>"001001001",
  13413=>"001010010",
  13414=>"000000000",
  13415=>"000000100",
  13416=>"111111111",
  13417=>"000000000",
  13418=>"000000000",
  13419=>"110000000",
  13420=>"111111111",
  13421=>"000000100",
  13422=>"001000000",
  13423=>"111111011",
  13424=>"000000000",
  13425=>"000000000",
  13426=>"000000000",
  13427=>"000001001",
  13428=>"101111111",
  13429=>"000000000",
  13430=>"000000000",
  13431=>"100100000",
  13432=>"000000000",
  13433=>"111001001",
  13434=>"111111111",
  13435=>"000000000",
  13436=>"111111111",
  13437=>"010000000",
  13438=>"101001101",
  13439=>"000000000",
  13440=>"000000000",
  13441=>"111111000",
  13442=>"000111111",
  13443=>"110110000",
  13444=>"000100111",
  13445=>"000000011",
  13446=>"100110010",
  13447=>"000111100",
  13448=>"000000000",
  13449=>"000000000",
  13450=>"100100111",
  13451=>"100100110",
  13452=>"001101001",
  13453=>"111111111",
  13454=>"000000000",
  13455=>"110111111",
  13456=>"111111111",
  13457=>"000001011",
  13458=>"000000000",
  13459=>"111111001",
  13460=>"011111001",
  13461=>"110110110",
  13462=>"000000000",
  13463=>"000001011",
  13464=>"111011000",
  13465=>"111111111",
  13466=>"111111111",
  13467=>"011011000",
  13468=>"011010000",
  13469=>"000100110",
  13470=>"101000000",
  13471=>"111000110",
  13472=>"000010000",
  13473=>"111110110",
  13474=>"000010110",
  13475=>"001011111",
  13476=>"111001001",
  13477=>"100000111",
  13478=>"110010000",
  13479=>"000000000",
  13480=>"110111011",
  13481=>"100111111",
  13482=>"000000000",
  13483=>"001100110",
  13484=>"110101011",
  13485=>"011011111",
  13486=>"000000000",
  13487=>"110110100",
  13488=>"010111111",
  13489=>"000110100",
  13490=>"111001000",
  13491=>"111111111",
  13492=>"010000111",
  13493=>"000000000",
  13494=>"111001011",
  13495=>"111111111",
  13496=>"000100000",
  13497=>"111000000",
  13498=>"111001001",
  13499=>"101101101",
  13500=>"100000000",
  13501=>"000000000",
  13502=>"000000000",
  13503=>"111111111",
  13504=>"100100111",
  13505=>"000000101",
  13506=>"000110111",
  13507=>"111111110",
  13508=>"000000000",
  13509=>"011000000",
  13510=>"111010000",
  13511=>"000000100",
  13512=>"001111000",
  13513=>"000000000",
  13514=>"111011001",
  13515=>"000000001",
  13516=>"110111010",
  13517=>"110111111",
  13518=>"010110100",
  13519=>"001111111",
  13520=>"111111111",
  13521=>"000001001",
  13522=>"010010010",
  13523=>"000000001",
  13524=>"100100000",
  13525=>"111111111",
  13526=>"000111111",
  13527=>"111111111",
  13528=>"000000000",
  13529=>"111111111",
  13530=>"000000000",
  13531=>"110110010",
  13532=>"111111111",
  13533=>"000000010",
  13534=>"111000000",
  13535=>"000000000",
  13536=>"000000100",
  13537=>"111111111",
  13538=>"100000000",
  13539=>"111111101",
  13540=>"010110100",
  13541=>"110010000",
  13542=>"000000000",
  13543=>"001000000",
  13544=>"110010010",
  13545=>"101101101",
  13546=>"000000001",
  13547=>"000000000",
  13548=>"000000000",
  13549=>"000000000",
  13550=>"111111110",
  13551=>"011011011",
  13552=>"000100111",
  13553=>"111101101",
  13554=>"110111110",
  13555=>"100000000",
  13556=>"111111111",
  13557=>"011011011",
  13558=>"011111011",
  13559=>"111111111",
  13560=>"101111111",
  13561=>"001000000",
  13562=>"000001101",
  13563=>"000000000",
  13564=>"000000100",
  13565=>"001001111",
  13566=>"111111011",
  13567=>"110110100",
  13568=>"011111111",
  13569=>"011001011",
  13570=>"011011001",
  13571=>"000000110",
  13572=>"010100100",
  13573=>"000000000",
  13574=>"000000000",
  13575=>"101111111",
  13576=>"111111111",
  13577=>"111111100",
  13578=>"000000000",
  13579=>"000000111",
  13580=>"000000000",
  13581=>"000000111",
  13582=>"000000111",
  13583=>"000101000",
  13584=>"111101001",
  13585=>"100000000",
  13586=>"000011111",
  13587=>"111110110",
  13588=>"000000000",
  13589=>"110110111",
  13590=>"011011010",
  13591=>"011111111",
  13592=>"000001001",
  13593=>"011111000",
  13594=>"000000000",
  13595=>"111111111",
  13596=>"000000100",
  13597=>"111111111",
  13598=>"111111111",
  13599=>"010111110",
  13600=>"011111011",
  13601=>"000000000",
  13602=>"000000000",
  13603=>"111111111",
  13604=>"001000000",
  13605=>"111111111",
  13606=>"111111111",
  13607=>"111111111",
  13608=>"001000110",
  13609=>"011111010",
  13610=>"000000000",
  13611=>"000000000",
  13612=>"111111011",
  13613=>"110110110",
  13614=>"110010111",
  13615=>"000000000",
  13616=>"111111000",
  13617=>"000111111",
  13618=>"111100000",
  13619=>"100000111",
  13620=>"000000000",
  13621=>"111110010",
  13622=>"001001010",
  13623=>"000000000",
  13624=>"000000000",
  13625=>"000000000",
  13626=>"101111111",
  13627=>"100000001",
  13628=>"111111001",
  13629=>"010110110",
  13630=>"001001111",
  13631=>"101111111",
  13632=>"000000000",
  13633=>"111111111",
  13634=>"000000100",
  13635=>"101001111",
  13636=>"011000000",
  13637=>"110010110",
  13638=>"110111110",
  13639=>"000000000",
  13640=>"000001001",
  13641=>"010010000",
  13642=>"110000111",
  13643=>"000000000",
  13644=>"110111000",
  13645=>"000000000",
  13646=>"100101111",
  13647=>"110111111",
  13648=>"100000000",
  13649=>"100000111",
  13650=>"111111111",
  13651=>"000000111",
  13652=>"000000000",
  13653=>"111111111",
  13654=>"001110111",
  13655=>"111111000",
  13656=>"000000000",
  13657=>"111111011",
  13658=>"111111111",
  13659=>"000100111",
  13660=>"000111000",
  13661=>"111110111",
  13662=>"000100111",
  13663=>"111111111",
  13664=>"000001001",
  13665=>"000000000",
  13666=>"011001001",
  13667=>"110111111",
  13668=>"111111100",
  13669=>"000000111",
  13670=>"110110111",
  13671=>"110111000",
  13672=>"100110000",
  13673=>"000111111",
  13674=>"111111111",
  13675=>"000111111",
  13676=>"000011000",
  13677=>"001001111",
  13678=>"000000000",
  13679=>"000000001",
  13680=>"001000000",
  13681=>"111111000",
  13682=>"111111111",
  13683=>"111111110",
  13684=>"111111111",
  13685=>"000000000",
  13686=>"001000000",
  13687=>"110111111",
  13688=>"000000001",
  13689=>"000000100",
  13690=>"000000000",
  13691=>"010111111",
  13692=>"111101100",
  13693=>"001001001",
  13694=>"111100111",
  13695=>"111111111",
  13696=>"010010000",
  13697=>"000001000",
  13698=>"011011011",
  13699=>"000000001",
  13700=>"000000110",
  13701=>"000000000",
  13702=>"110100000",
  13703=>"000000111",
  13704=>"000000000",
  13705=>"111111110",
  13706=>"100111111",
  13707=>"111111110",
  13708=>"111111111",
  13709=>"001011011",
  13710=>"000000111",
  13711=>"111111000",
  13712=>"111110000",
  13713=>"111111000",
  13714=>"000000010",
  13715=>"011001111",
  13716=>"101111000",
  13717=>"000010000",
  13718=>"111111111",
  13719=>"101001001",
  13720=>"000000111",
  13721=>"101001111",
  13722=>"000000110",
  13723=>"101111111",
  13724=>"011111111",
  13725=>"010000111",
  13726=>"100000000",
  13727=>"111011001",
  13728=>"000000000",
  13729=>"001001111",
  13730=>"110110111",
  13731=>"000000000",
  13732=>"110111001",
  13733=>"010010000",
  13734=>"000000001",
  13735=>"111011101",
  13736=>"100000000",
  13737=>"100000000",
  13738=>"000000000",
  13739=>"100100100",
  13740=>"111111010",
  13741=>"111110010",
  13742=>"111111111",
  13743=>"111111111",
  13744=>"000000000",
  13745=>"000111111",
  13746=>"100110111",
  13747=>"111111010",
  13748=>"111111111",
  13749=>"000000011",
  13750=>"111110111",
  13751=>"100000110",
  13752=>"000111111",
  13753=>"000000111",
  13754=>"000111111",
  13755=>"000010111",
  13756=>"010010000",
  13757=>"100011111",
  13758=>"000000000",
  13759=>"011011011",
  13760=>"111111111",
  13761=>"111110000",
  13762=>"000000000",
  13763=>"111111111",
  13764=>"110110110",
  13765=>"111110111",
  13766=>"110111011",
  13767=>"111111010",
  13768=>"000000000",
  13769=>"000001111",
  13770=>"000000000",
  13771=>"000000111",
  13772=>"000000000",
  13773=>"000101111",
  13774=>"000000000",
  13775=>"001000001",
  13776=>"111111111",
  13777=>"011001111",
  13778=>"111111110",
  13779=>"010111011",
  13780=>"000111011",
  13781=>"000000000",
  13782=>"000111111",
  13783=>"000000000",
  13784=>"000111011",
  13785=>"000000000",
  13786=>"000000000",
  13787=>"111110111",
  13788=>"111010010",
  13789=>"000100000",
  13790=>"000000000",
  13791=>"001000110",
  13792=>"000000000",
  13793=>"111111111",
  13794=>"000000001",
  13795=>"000000000",
  13796=>"000001111",
  13797=>"110110111",
  13798=>"001001011",
  13799=>"000000000",
  13800=>"010111111",
  13801=>"111111110",
  13802=>"000000000",
  13803=>"111010111",
  13804=>"000110111",
  13805=>"111110111",
  13806=>"000000000",
  13807=>"000000110",
  13808=>"000000101",
  13809=>"000000000",
  13810=>"010110110",
  13811=>"110010000",
  13812=>"000000000",
  13813=>"000000000",
  13814=>"111111111",
  13815=>"000000100",
  13816=>"010111111",
  13817=>"100100100",
  13818=>"000000000",
  13819=>"111111110",
  13820=>"000000000",
  13821=>"000001001",
  13822=>"000000000",
  13823=>"000001101",
  13824=>"011111111",
  13825=>"000000000",
  13826=>"000000000",
  13827=>"111100000",
  13828=>"000000000",
  13829=>"111101001",
  13830=>"010010011",
  13831=>"101000000",
  13832=>"001011000",
  13833=>"110111111",
  13834=>"101000000",
  13835=>"000001100",
  13836=>"011000000",
  13837=>"000000000",
  13838=>"001001111",
  13839=>"111111111",
  13840=>"000000001",
  13841=>"111011001",
  13842=>"111111111",
  13843=>"000000000",
  13844=>"100000100",
  13845=>"111111111",
  13846=>"101111011",
  13847=>"100100001",
  13848=>"001110100",
  13849=>"001011000",
  13850=>"001111111",
  13851=>"011000010",
  13852=>"011000000",
  13853=>"111101001",
  13854=>"111101000",
  13855=>"000101111",
  13856=>"111111100",
  13857=>"110000000",
  13858=>"011011011",
  13859=>"000000000",
  13860=>"000110110",
  13861=>"000111111",
  13862=>"111111000",
  13863=>"111111111",
  13864=>"000111111",
  13865=>"111111111",
  13866=>"000000000",
  13867=>"000000000",
  13868=>"000000011",
  13869=>"111101001",
  13870=>"011001011",
  13871=>"111111111",
  13872=>"000000000",
  13873=>"111111111",
  13874=>"000110010",
  13875=>"000111101",
  13876=>"010111111",
  13877=>"001011011",
  13878=>"000000000",
  13879=>"000000111",
  13880=>"011111110",
  13881=>"000011000",
  13882=>"000000010",
  13883=>"000000110",
  13884=>"000000110",
  13885=>"000000000",
  13886=>"111111001",
  13887=>"111000000",
  13888=>"110000000",
  13889=>"010010000",
  13890=>"010111111",
  13891=>"100100000",
  13892=>"111001001",
  13893=>"111111101",
  13894=>"000000000",
  13895=>"111111111",
  13896=>"110000000",
  13897=>"111111111",
  13898=>"111111100",
  13899=>"001011000",
  13900=>"101101100",
  13901=>"111111111",
  13902=>"101111101",
  13903=>"000000111",
  13904=>"111111111",
  13905=>"111110000",
  13906=>"000000000",
  13907=>"010110111",
  13908=>"000000111",
  13909=>"000001111",
  13910=>"111000001",
  13911=>"111111000",
  13912=>"111111110",
  13913=>"111101111",
  13914=>"111111111",
  13915=>"110110001",
  13916=>"111111111",
  13917=>"110110111",
  13918=>"000000101",
  13919=>"100001000",
  13920=>"111111011",
  13921=>"110100101",
  13922=>"000000000",
  13923=>"000111011",
  13924=>"000000000",
  13925=>"011000001",
  13926=>"111111111",
  13927=>"111100000",
  13928=>"111110000",
  13929=>"100000000",
  13930=>"111111111",
  13931=>"000000110",
  13932=>"001001000",
  13933=>"111111111",
  13934=>"100100000",
  13935=>"100100100",
  13936=>"100000110",
  13937=>"011011111",
  13938=>"000010000",
  13939=>"100110110",
  13940=>"001000000",
  13941=>"111111111",
  13942=>"000000000",
  13943=>"001111111",
  13944=>"111111011",
  13945=>"111001000",
  13946=>"001000101",
  13947=>"111100000",
  13948=>"110111111",
  13949=>"000110111",
  13950=>"000000000",
  13951=>"011111111",
  13952=>"000000000",
  13953=>"100000000",
  13954=>"111000000",
  13955=>"001001000",
  13956=>"000000000",
  13957=>"111111111",
  13958=>"110100000",
  13959=>"111000000",
  13960=>"000000000",
  13961=>"110100000",
  13962=>"000010001",
  13963=>"000000111",
  13964=>"000000000",
  13965=>"111110000",
  13966=>"011000011",
  13967=>"000000111",
  13968=>"000000000",
  13969=>"111111111",
  13970=>"000000000",
  13971=>"000011111",
  13972=>"000110111",
  13973=>"111111111",
  13974=>"111000000",
  13975=>"100100000",
  13976=>"000000001",
  13977=>"111111100",
  13978=>"000000000",
  13979=>"000000000",
  13980=>"000000101",
  13981=>"111111010",
  13982=>"111111111",
  13983=>"000001011",
  13984=>"100111111",
  13985=>"111111110",
  13986=>"000000011",
  13987=>"000000000",
  13988=>"011111111",
  13989=>"111111111",
  13990=>"000000000",
  13991=>"111100111",
  13992=>"111111111",
  13993=>"100101111",
  13994=>"111111111",
  13995=>"111100110",
  13996=>"111010111",
  13997=>"001111111",
  13998=>"111010000",
  13999=>"000000000",
  14000=>"000000000",
  14001=>"111111111",
  14002=>"100110110",
  14003=>"000000000",
  14004=>"000000000",
  14005=>"111111111",
  14006=>"111111000",
  14007=>"000110111",
  14008=>"100100001",
  14009=>"111111111",
  14010=>"000000100",
  14011=>"000000001",
  14012=>"111110110",
  14013=>"001001001",
  14014=>"000001111",
  14015=>"001001001",
  14016=>"001001011",
  14017=>"110111111",
  14018=>"000001111",
  14019=>"010000000",
  14020=>"011011111",
  14021=>"011111011",
  14022=>"111101111",
  14023=>"100111000",
  14024=>"110110110",
  14025=>"011111000",
  14026=>"000100110",
  14027=>"111111111",
  14028=>"000000000",
  14029=>"000000111",
  14030=>"111000001",
  14031=>"000011111",
  14032=>"111100000",
  14033=>"000000010",
  14034=>"000000010",
  14035=>"111011000",
  14036=>"000000000",
  14037=>"111111111",
  14038=>"111111111",
  14039=>"000000000",
  14040=>"011000100",
  14041=>"011011011",
  14042=>"000010010",
  14043=>"000001000",
  14044=>"110000111",
  14045=>"100000000",
  14046=>"000000111",
  14047=>"000110110",
  14048=>"000000000",
  14049=>"100101100",
  14050=>"111010000",
  14051=>"000000000",
  14052=>"000000000",
  14053=>"100110110",
  14054=>"101101100",
  14055=>"101111111",
  14056=>"011111111",
  14057=>"101000110",
  14058=>"000000001",
  14059=>"000000000",
  14060=>"111111111",
  14061=>"100110111",
  14062=>"111111000",
  14063=>"111100111",
  14064=>"111110100",
  14065=>"000000000",
  14066=>"000000000",
  14067=>"011010000",
  14068=>"000000010",
  14069=>"111011000",
  14070=>"000000001",
  14071=>"111010111",
  14072=>"111111111",
  14073=>"000000000",
  14074=>"111111111",
  14075=>"100101101",
  14076=>"101111011",
  14077=>"000100110",
  14078=>"000000000",
  14079=>"111111111",
  14080=>"000000100",
  14081=>"001011110",
  14082=>"000000000",
  14083=>"110111101",
  14084=>"000000000",
  14085=>"011011001",
  14086=>"000001111",
  14087=>"011011100",
  14088=>"111111111",
  14089=>"111111111",
  14090=>"110100100",
  14091=>"001111111",
  14092=>"110100110",
  14093=>"111011011",
  14094=>"111110101",
  14095=>"111111110",
  14096=>"111111101",
  14097=>"000000000",
  14098=>"100000111",
  14099=>"111000000",
  14100=>"011010000",
  14101=>"111111111",
  14102=>"111110110",
  14103=>"111111111",
  14104=>"111111111",
  14105=>"111111111",
  14106=>"100000100",
  14107=>"111100111",
  14108=>"011011001",
  14109=>"111111111",
  14110=>"000000000",
  14111=>"001111111",
  14112=>"101000111",
  14113=>"110000000",
  14114=>"000000100",
  14115=>"111111111",
  14116=>"101111000",
  14117=>"000000001",
  14118=>"111000111",
  14119=>"011011000",
  14120=>"000000000",
  14121=>"111111111",
  14122=>"111111100",
  14123=>"111111000",
  14124=>"000000000",
  14125=>"011011000",
  14126=>"000010000",
  14127=>"111111111",
  14128=>"001001011",
  14129=>"000000100",
  14130=>"000000011",
  14131=>"000000110",
  14132=>"000000000",
  14133=>"000101111",
  14134=>"000000111",
  14135=>"001000000",
  14136=>"110111110",
  14137=>"000000011",
  14138=>"000000000",
  14139=>"110110100",
  14140=>"000000001",
  14141=>"001001100",
  14142=>"000000000",
  14143=>"000000000",
  14144=>"001001001",
  14145=>"111011011",
  14146=>"001100000",
  14147=>"111111111",
  14148=>"011110000",
  14149=>"000000000",
  14150=>"111111111",
  14151=>"111111001",
  14152=>"000110111",
  14153=>"000000000",
  14154=>"000000000",
  14155=>"010011010",
  14156=>"111111111",
  14157=>"010000111",
  14158=>"101110111",
  14159=>"110110110",
  14160=>"000100110",
  14161=>"101101100",
  14162=>"111111111",
  14163=>"000000001",
  14164=>"101001001",
  14165=>"001010011",
  14166=>"000000000",
  14167=>"100001001",
  14168=>"001011000",
  14169=>"111001000",
  14170=>"110001000",
  14171=>"000000000",
  14172=>"101101001",
  14173=>"111111111",
  14174=>"011010110",
  14175=>"111111111",
  14176=>"111111111",
  14177=>"111000000",
  14178=>"111011011",
  14179=>"000000011",
  14180=>"001000000",
  14181=>"000000000",
  14182=>"111111111",
  14183=>"111111111",
  14184=>"101000000",
  14185=>"011010111",
  14186=>"010000111",
  14187=>"110110111",
  14188=>"111111111",
  14189=>"000000000",
  14190=>"111111111",
  14191=>"000011011",
  14192=>"111100010",
  14193=>"111111111",
  14194=>"110110111",
  14195=>"111111010",
  14196=>"000000000",
  14197=>"010000000",
  14198=>"111111000",
  14199=>"000010000",
  14200=>"000000000",
  14201=>"101110110",
  14202=>"111111111",
  14203=>"000001111",
  14204=>"111111111",
  14205=>"111111101",
  14206=>"100100100",
  14207=>"111111000",
  14208=>"100000000",
  14209=>"111001101",
  14210=>"111111111",
  14211=>"000000000",
  14212=>"111010000",
  14213=>"001000101",
  14214=>"001101111",
  14215=>"011111011",
  14216=>"000000110",
  14217=>"000000000",
  14218=>"110111111",
  14219=>"110010000",
  14220=>"000000000",
  14221=>"001011000",
  14222=>"101111100",
  14223=>"110110110",
  14224=>"000000000",
  14225=>"111111111",
  14226=>"100000000",
  14227=>"000000100",
  14228=>"000000100",
  14229=>"000100000",
  14230=>"000000000",
  14231=>"111110111",
  14232=>"001000000",
  14233=>"110000000",
  14234=>"000111111",
  14235=>"000111111",
  14236=>"000000011",
  14237=>"001011011",
  14238=>"101000000",
  14239=>"000000100",
  14240=>"111101111",
  14241=>"100101111",
  14242=>"010000000",
  14243=>"111111111",
  14244=>"011111111",
  14245=>"111111111",
  14246=>"111111111",
  14247=>"011111111",
  14248=>"111010001",
  14249=>"010100111",
  14250=>"101111111",
  14251=>"000011000",
  14252=>"000000000",
  14253=>"101001111",
  14254=>"100011011",
  14255=>"111111011",
  14256=>"111111111",
  14257=>"011010000",
  14258=>"000000110",
  14259=>"000000000",
  14260=>"111000000",
  14261=>"111111111",
  14262=>"010000000",
  14263=>"000000000",
  14264=>"000000111",
  14265=>"000000000",
  14266=>"110000000",
  14267=>"000000000",
  14268=>"100000000",
  14269=>"111111101",
  14270=>"111111111",
  14271=>"001001011",
  14272=>"001001000",
  14273=>"000000000",
  14274=>"111000101",
  14275=>"000000000",
  14276=>"111011000",
  14277=>"001111000",
  14278=>"111011111",
  14279=>"000000000",
  14280=>"000000111",
  14281=>"111111000",
  14282=>"011110000",
  14283=>"111111111",
  14284=>"000000111",
  14285=>"101000110",
  14286=>"000000000",
  14287=>"111111001",
  14288=>"000000100",
  14289=>"000000010",
  14290=>"000100000",
  14291=>"111010000",
  14292=>"000000000",
  14293=>"111000101",
  14294=>"111111100",
  14295=>"000000000",
  14296=>"001000001",
  14297=>"111111001",
  14298=>"000111110",
  14299=>"000000000",
  14300=>"011011010",
  14301=>"001000000",
  14302=>"000000000",
  14303=>"001000000",
  14304=>"111111000",
  14305=>"011111111",
  14306=>"111111000",
  14307=>"000001111",
  14308=>"010010010",
  14309=>"111111111",
  14310=>"000010111",
  14311=>"111111111",
  14312=>"111111111",
  14313=>"100100111",
  14314=>"110000111",
  14315=>"000000011",
  14316=>"000110110",
  14317=>"011111111",
  14318=>"100111111",
  14319=>"110110100",
  14320=>"000000111",
  14321=>"110111000",
  14322=>"111111111",
  14323=>"000000000",
  14324=>"011111010",
  14325=>"000000111",
  14326=>"111111111",
  14327=>"011101111",
  14328=>"000000111",
  14329=>"000000110",
  14330=>"000010010",
  14331=>"000000000",
  14332=>"000000000",
  14333=>"111111111",
  14334=>"000000000",
  14335=>"111111111",
  14336=>"100000011",
  14337=>"111111111",
  14338=>"101000000",
  14339=>"000000110",
  14340=>"000000000",
  14341=>"100000000",
  14342=>"010000000",
  14343=>"111111111",
  14344=>"111111011",
  14345=>"111110110",
  14346=>"111110000",
  14347=>"100100000",
  14348=>"111111100",
  14349=>"000011000",
  14350=>"100111011",
  14351=>"000000111",
  14352=>"111100101",
  14353=>"011001111",
  14354=>"111001001",
  14355=>"000000000",
  14356=>"111111111",
  14357=>"111011000",
  14358=>"111111111",
  14359=>"001000000",
  14360=>"110111111",
  14361=>"010000000",
  14362=>"000110110",
  14363=>"100100100",
  14364=>"000000111",
  14365=>"000000000",
  14366=>"111111111",
  14367=>"000000000",
  14368=>"000111111",
  14369=>"111111000",
  14370=>"111111110",
  14371=>"000000000",
  14372=>"111110111",
  14373=>"000000000",
  14374=>"111111111",
  14375=>"111111000",
  14376=>"000000000",
  14377=>"111111101",
  14378=>"100000100",
  14379=>"000000000",
  14380=>"111101000",
  14381=>"100000010",
  14382=>"000110110",
  14383=>"100010000",
  14384=>"000010000",
  14385=>"000000000",
  14386=>"000000000",
  14387=>"111111011",
  14388=>"000000000",
  14389=>"110000100",
  14390=>"111111111",
  14391=>"011011111",
  14392=>"111011001",
  14393=>"001001111",
  14394=>"000000000",
  14395=>"111110000",
  14396=>"000110110",
  14397=>"000100111",
  14398=>"100111111",
  14399=>"011001011",
  14400=>"001000001",
  14401=>"001011011",
  14402=>"110000000",
  14403=>"110100000",
  14404=>"110100100",
  14405=>"110110111",
  14406=>"111000000",
  14407=>"111111111",
  14408=>"001011011",
  14409=>"000000000",
  14410=>"011111111",
  14411=>"000000000",
  14412=>"000000000",
  14413=>"100000000",
  14414=>"111000000",
  14415=>"100110000",
  14416=>"011111111",
  14417=>"111011000",
  14418=>"111001111",
  14419=>"000000100",
  14420=>"000000000",
  14421=>"111101110",
  14422=>"000101001",
  14423=>"111101001",
  14424=>"111110000",
  14425=>"000000000",
  14426=>"000000000",
  14427=>"000000000",
  14428=>"000111111",
  14429=>"000000000",
  14430=>"000001101",
  14431=>"101101101",
  14432=>"000001000",
  14433=>"110111111",
  14434=>"000111111",
  14435=>"001111111",
  14436=>"111111000",
  14437=>"001011001",
  14438=>"111111000",
  14439=>"000000111",
  14440=>"101001010",
  14441=>"000000000",
  14442=>"000000000",
  14443=>"000000000",
  14444=>"110110110",
  14445=>"000111111",
  14446=>"100100000",
  14447=>"000100111",
  14448=>"001000000",
  14449=>"011000100",
  14450=>"011011110",
  14451=>"011110001",
  14452=>"000000010",
  14453=>"000000011",
  14454=>"111100111",
  14455=>"000000111",
  14456=>"000000000",
  14457=>"000010000",
  14458=>"000000000",
  14459=>"000000000",
  14460=>"100110110",
  14461=>"000000000",
  14462=>"000000000",
  14463=>"111011001",
  14464=>"000000001",
  14465=>"111111100",
  14466=>"111111111",
  14467=>"000000000",
  14468=>"011000000",
  14469=>"000000000",
  14470=>"110100111",
  14471=>"000111111",
  14472=>"111111111",
  14473=>"100100000",
  14474=>"111011000",
  14475=>"001000011",
  14476=>"000000000",
  14477=>"111111110",
  14478=>"000000010",
  14479=>"000000000",
  14480=>"000111111",
  14481=>"111111000",
  14482=>"111111111",
  14483=>"111111111",
  14484=>"000100111",
  14485=>"110000000",
  14486=>"101000000",
  14487=>"111110010",
  14488=>"000000001",
  14489=>"111111010",
  14490=>"011111111",
  14491=>"111000000",
  14492=>"111011111",
  14493=>"000000000",
  14494=>"111111000",
  14495=>"000000001",
  14496=>"000000000",
  14497=>"000000000",
  14498=>"110100111",
  14499=>"000000001",
  14500=>"100100010",
  14501=>"000001001",
  14502=>"111001000",
  14503=>"011010000",
  14504=>"111111111",
  14505=>"000000111",
  14506=>"111111111",
  14507=>"101110111",
  14508=>"000000111",
  14509=>"000000000",
  14510=>"111111111",
  14511=>"000000110",
  14512=>"110111111",
  14513=>"000000100",
  14514=>"001001111",
  14515=>"111101000",
  14516=>"000111000",
  14517=>"000000000",
  14518=>"000000001",
  14519=>"001000000",
  14520=>"111111110",
  14521=>"111111111",
  14522=>"110110000",
  14523=>"111111110",
  14524=>"000000100",
  14525=>"110011000",
  14526=>"000000100",
  14527=>"111000001",
  14528=>"001111111",
  14529=>"010011111",
  14530=>"000010010",
  14531=>"000000000",
  14532=>"000000111",
  14533=>"000000000",
  14534=>"000001000",
  14535=>"111111111",
  14536=>"111111111",
  14537=>"000000111",
  14538=>"111111111",
  14539=>"100101111",
  14540=>"011110110",
  14541=>"000111111",
  14542=>"000011000",
  14543=>"011111000",
  14544=>"000000000",
  14545=>"001111111",
  14546=>"100100000",
  14547=>"110100111",
  14548=>"000000111",
  14549=>"001011000",
  14550=>"000000000",
  14551=>"111100010",
  14552=>"111111111",
  14553=>"111111110",
  14554=>"111111111",
  14555=>"011111110",
  14556=>"000000000",
  14557=>"000100110",
  14558=>"000000111",
  14559=>"111111111",
  14560=>"001000000",
  14561=>"111111111",
  14562=>"111000000",
  14563=>"000000011",
  14564=>"000010111",
  14565=>"010000000",
  14566=>"111111001",
  14567=>"111101000",
  14568=>"000010000",
  14569=>"001110111",
  14570=>"111111111",
  14571=>"111111101",
  14572=>"111111001",
  14573=>"100010000",
  14574=>"111111111",
  14575=>"000011000",
  14576=>"111111000",
  14577=>"011011011",
  14578=>"100000010",
  14579=>"111011000",
  14580=>"110000111",
  14581=>"111111100",
  14582=>"011111000",
  14583=>"111111111",
  14584=>"000000000",
  14585=>"111100110",
  14586=>"001011111",
  14587=>"101101111",
  14588=>"000111111",
  14589=>"111010000",
  14590=>"011000000",
  14591=>"111110000",
  14592=>"000000111",
  14593=>"111110110",
  14594=>"100100100",
  14595=>"111110110",
  14596=>"000110011",
  14597=>"001000000",
  14598=>"110000000",
  14599=>"111111111",
  14600=>"000000011",
  14601=>"111010110",
  14602=>"000001011",
  14603=>"000000000",
  14604=>"111001000",
  14605=>"000000000",
  14606=>"110000001",
  14607=>"000100100",
  14608=>"100100100",
  14609=>"000001000",
  14610=>"111111111",
  14611=>"000111111",
  14612=>"110001011",
  14613=>"111110111",
  14614=>"000000110",
  14615=>"011011010",
  14616=>"111111111",
  14617=>"110111111",
  14618=>"000000000",
  14619=>"000000000",
  14620=>"110111110",
  14621=>"011111111",
  14622=>"011111111",
  14623=>"101101111",
  14624=>"000001011",
  14625=>"101001001",
  14626=>"000000000",
  14627=>"111011111",
  14628=>"111111111",
  14629=>"111101000",
  14630=>"000111000",
  14631=>"111111000",
  14632=>"111111100",
  14633=>"011011111",
  14634=>"100000000",
  14635=>"101011000",
  14636=>"111111111",
  14637=>"000000100",
  14638=>"110000000",
  14639=>"000000001",
  14640=>"001111111",
  14641=>"111111111",
  14642=>"000000000",
  14643=>"000000000",
  14644=>"001000000",
  14645=>"011111111",
  14646=>"000000000",
  14647=>"111111111",
  14648=>"101000000",
  14649=>"100001000",
  14650=>"111111111",
  14651=>"000001000",
  14652=>"000000011",
  14653=>"001000000",
  14654=>"000000101",
  14655=>"111111110",
  14656=>"111100111",
  14657=>"001001001",
  14658=>"001000001",
  14659=>"111011111",
  14660=>"000000000",
  14661=>"111110000",
  14662=>"111011000",
  14663=>"000000000",
  14664=>"000111111",
  14665=>"000000000",
  14666=>"111110000",
  14667=>"111100101",
  14668=>"110100000",
  14669=>"000000000",
  14670=>"111111111",
  14671=>"110111111",
  14672=>"000000011",
  14673=>"111111110",
  14674=>"111110111",
  14675=>"111101001",
  14676=>"100000000",
  14677=>"011111011",
  14678=>"101110111",
  14679=>"000001000",
  14680=>"000000000",
  14681=>"111001000",
  14682=>"011000000",
  14683=>"011010000",
  14684=>"011000000",
  14685=>"101111111",
  14686=>"100010000",
  14687=>"110111111",
  14688=>"000100111",
  14689=>"000000000",
  14690=>"100110111",
  14691=>"011111011",
  14692=>"000000111",
  14693=>"111011001",
  14694=>"101101100",
  14695=>"111111111",
  14696=>"110011001",
  14697=>"000111111",
  14698=>"111001000",
  14699=>"111100000",
  14700=>"011000000",
  14701=>"110110010",
  14702=>"110111011",
  14703=>"000000000",
  14704=>"111111111",
  14705=>"001111111",
  14706=>"111111000",
  14707=>"000011001",
  14708=>"000000001",
  14709=>"111111000",
  14710=>"010011111",
  14711=>"101111111",
  14712=>"111111111",
  14713=>"000100100",
  14714=>"111111111",
  14715=>"010000000",
  14716=>"111111111",
  14717=>"000000111",
  14718=>"000100000",
  14719=>"100000010",
  14720=>"000111111",
  14721=>"111101111",
  14722=>"011011011",
  14723=>"000000110",
  14724=>"111010110",
  14725=>"011111011",
  14726=>"111111001",
  14727=>"001101101",
  14728=>"010000000",
  14729=>"110110100",
  14730=>"000000001",
  14731=>"000010110",
  14732=>"101111111",
  14733=>"000000001",
  14734=>"111111111",
  14735=>"000001111",
  14736=>"000100111",
  14737=>"111111111",
  14738=>"100000000",
  14739=>"000000011",
  14740=>"111111111",
  14741=>"000000000",
  14742=>"110100110",
  14743=>"101100000",
  14744=>"111111001",
  14745=>"111111111",
  14746=>"000000011",
  14747=>"100000000",
  14748=>"111111001",
  14749=>"111000000",
  14750=>"000000000",
  14751=>"000000000",
  14752=>"110110111",
  14753=>"000000000",
  14754=>"001000000",
  14755=>"000000010",
  14756=>"001001001",
  14757=>"101101000",
  14758=>"011000000",
  14759=>"111100100",
  14760=>"000000000",
  14761=>"111111111",
  14762=>"000000000",
  14763=>"000000000",
  14764=>"011011111",
  14765=>"000000000",
  14766=>"000000101",
  14767=>"111011000",
  14768=>"000000000",
  14769=>"001000000",
  14770=>"011011000",
  14771=>"000000000",
  14772=>"111111111",
  14773=>"111111111",
  14774=>"000000000",
  14775=>"110100110",
  14776=>"011000000",
  14777=>"111111000",
  14778=>"101100111",
  14779=>"111111011",
  14780=>"111111111",
  14781=>"000000100",
  14782=>"111001000",
  14783=>"000011011",
  14784=>"000000000",
  14785=>"001101001",
  14786=>"111111011",
  14787=>"000001000",
  14788=>"000000000",
  14789=>"010010010",
  14790=>"001000000",
  14791=>"000000110",
  14792=>"000000000",
  14793=>"111111111",
  14794=>"000001000",
  14795=>"101111110",
  14796=>"111100000",
  14797=>"111111111",
  14798=>"111001000",
  14799=>"000000000",
  14800=>"110000000",
  14801=>"011111111",
  14802=>"111111010",
  14803=>"101100111",
  14804=>"111111110",
  14805=>"000000000",
  14806=>"111111111",
  14807=>"111110000",
  14808=>"000000000",
  14809=>"111011110",
  14810=>"111101111",
  14811=>"111111000",
  14812=>"111100000",
  14813=>"000000111",
  14814=>"100110011",
  14815=>"000000110",
  14816=>"101110110",
  14817=>"111000000",
  14818=>"000000000",
  14819=>"001000011",
  14820=>"000000000",
  14821=>"000000000",
  14822=>"000000000",
  14823=>"111001000",
  14824=>"111111111",
  14825=>"000011011",
  14826=>"110000000",
  14827=>"111011011",
  14828=>"000110111",
  14829=>"000000000",
  14830=>"000111111",
  14831=>"000000000",
  14832=>"010110000",
  14833=>"000000111",
  14834=>"111111111",
  14835=>"000000111",
  14836=>"100110111",
  14837=>"000000000",
  14838=>"111111111",
  14839=>"111011000",
  14840=>"111000000",
  14841=>"010010010",
  14842=>"111111111",
  14843=>"001000000",
  14844=>"000100000",
  14845=>"011011110",
  14846=>"000000111",
  14847=>"000000000",
  14848=>"110001011",
  14849=>"000000000",
  14850=>"101000000",
  14851=>"000000000",
  14852=>"001000000",
  14853=>"011110100",
  14854=>"111111111",
  14855=>"111111111",
  14856=>"111110110",
  14857=>"111101000",
  14858=>"011000000",
  14859=>"000111111",
  14860=>"011000000",
  14861=>"000000000",
  14862=>"000000111",
  14863=>"111111111",
  14864=>"111000000",
  14865=>"111111111",
  14866=>"111111010",
  14867=>"000000000",
  14868=>"111000000",
  14869=>"011000110",
  14870=>"000000000",
  14871=>"110100100",
  14872=>"111111111",
  14873=>"011011000",
  14874=>"111111111",
  14875=>"111111110",
  14876=>"001001000",
  14877=>"011000000",
  14878=>"001111110",
  14879=>"101111001",
  14880=>"100000000",
  14881=>"000000000",
  14882=>"010010010",
  14883=>"000000000",
  14884=>"100111111",
  14885=>"100111111",
  14886=>"111110010",
  14887=>"000101001",
  14888=>"000000000",
  14889=>"111111111",
  14890=>"001111000",
  14891=>"100100001",
  14892=>"010000000",
  14893=>"011101000",
  14894=>"000000000",
  14895=>"111111100",
  14896=>"111011000",
  14897=>"000000000",
  14898=>"110110110",
  14899=>"000000101",
  14900=>"000000101",
  14901=>"011111110",
  14902=>"000000000",
  14903=>"111111111",
  14904=>"111111111",
  14905=>"010011000",
  14906=>"000000011",
  14907=>"000000000",
  14908=>"000000000",
  14909=>"000000010",
  14910=>"110110110",
  14911=>"000000000",
  14912=>"111000000",
  14913=>"000101111",
  14914=>"000111000",
  14915=>"111111100",
  14916=>"001001011",
  14917=>"011011011",
  14918=>"000000111",
  14919=>"000011111",
  14920=>"110110111",
  14921=>"000111111",
  14922=>"011111100",
  14923=>"011011111",
  14924=>"000100111",
  14925=>"000000000",
  14926=>"000000000",
  14927=>"000000000",
  14928=>"111111111",
  14929=>"110111011",
  14930=>"000000000",
  14931=>"100110000",
  14932=>"111000001",
  14933=>"001000000",
  14934=>"100000001",
  14935=>"111111111",
  14936=>"101001111",
  14937=>"100100000",
  14938=>"000000010",
  14939=>"110110000",
  14940=>"111111111",
  14941=>"000000110",
  14942=>"111111111",
  14943=>"000000000",
  14944=>"000001111",
  14945=>"110110000",
  14946=>"000000000",
  14947=>"110110000",
  14948=>"000000001",
  14949=>"010010000",
  14950=>"110111111",
  14951=>"000111011",
  14952=>"111111111",
  14953=>"000101111",
  14954=>"111110100",
  14955=>"111000000",
  14956=>"110111111",
  14957=>"101101111",
  14958=>"000000000",
  14959=>"001000000",
  14960=>"111000000",
  14961=>"000000110",
  14962=>"001011001",
  14963=>"000001001",
  14964=>"011011010",
  14965=>"011000111",
  14966=>"000000000",
  14967=>"011111111",
  14968=>"111100001",
  14969=>"111011010",
  14970=>"111001001",
  14971=>"000000000",
  14972=>"000000000",
  14973=>"100111111",
  14974=>"001000000",
  14975=>"000000011",
  14976=>"001001001",
  14977=>"000000000",
  14978=>"010010111",
  14979=>"000000100",
  14980=>"000000001",
  14981=>"111100111",
  14982=>"000111111",
  14983=>"000000010",
  14984=>"000000100",
  14985=>"111000000",
  14986=>"000111111",
  14987=>"111111111",
  14988=>"111110010",
  14989=>"000000000",
  14990=>"111000011",
  14991=>"111111111",
  14992=>"000000000",
  14993=>"011001001",
  14994=>"000010010",
  14995=>"000000000",
  14996=>"111111101",
  14997=>"111111001",
  14998=>"010111011",
  14999=>"000000000",
  15000=>"000000000",
  15001=>"000000000",
  15002=>"000000000",
  15003=>"000000000",
  15004=>"111111111",
  15005=>"000001001",
  15006=>"111111111",
  15007=>"111110110",
  15008=>"111111111",
  15009=>"100111111",
  15010=>"000000000",
  15011=>"000111111",
  15012=>"001001001",
  15013=>"111101101",
  15014=>"111111111",
  15015=>"111000000",
  15016=>"000000000",
  15017=>"000111111",
  15018=>"011111111",
  15019=>"111111111",
  15020=>"000000000",
  15021=>"000000111",
  15022=>"000000000",
  15023=>"000000111",
  15024=>"001001000",
  15025=>"111100111",
  15026=>"111111100",
  15027=>"111000001",
  15028=>"111111111",
  15029=>"000010000",
  15030=>"010010010",
  15031=>"111111111",
  15032=>"111110111",
  15033=>"010010110",
  15034=>"001001001",
  15035=>"000010010",
  15036=>"000000000",
  15037=>"010010011",
  15038=>"110111111",
  15039=>"000000000",
  15040=>"111111111",
  15041=>"001000000",
  15042=>"010110111",
  15043=>"000000111",
  15044=>"111111111",
  15045=>"010000000",
  15046=>"010010111",
  15047=>"100000000",
  15048=>"101110111",
  15049=>"000000000",
  15050=>"100100100",
  15051=>"111111111",
  15052=>"110111111",
  15053=>"001001001",
  15054=>"000000101",
  15055=>"000000001",
  15056=>"011000000",
  15057=>"000000000",
  15058=>"000010001",
  15059=>"101101101",
  15060=>"000000001",
  15061=>"110000000",
  15062=>"100100000",
  15063=>"111110110",
  15064=>"010010001",
  15065=>"110110110",
  15066=>"111111111",
  15067=>"100100111",
  15068=>"111110110",
  15069=>"000000000",
  15070=>"010000110",
  15071=>"111111111",
  15072=>"110000000",
  15073=>"111111010",
  15074=>"000011011",
  15075=>"000000000",
  15076=>"001101101",
  15077=>"011010000",
  15078=>"111101111",
  15079=>"111110000",
  15080=>"000000010",
  15081=>"111111001",
  15082=>"111111000",
  15083=>"001000000",
  15084=>"000000000",
  15085=>"111111111",
  15086=>"100111101",
  15087=>"000101110",
  15088=>"111101111",
  15089=>"000000000",
  15090=>"000010110",
  15091=>"000000111",
  15092=>"111101111",
  15093=>"010000000",
  15094=>"000000000",
  15095=>"000001111",
  15096=>"000101111",
  15097=>"100111101",
  15098=>"111111001",
  15099=>"000000000",
  15100=>"111101101",
  15101=>"000000000",
  15102=>"000000111",
  15103=>"111111011",
  15104=>"111111111",
  15105=>"011010000",
  15106=>"000000000",
  15107=>"111010000",
  15108=>"111111111",
  15109=>"110100110",
  15110=>"110111000",
  15111=>"011000000",
  15112=>"100000100",
  15113=>"111111010",
  15114=>"111111100",
  15115=>"111111100",
  15116=>"110111111",
  15117=>"111111111",
  15118=>"010010000",
  15119=>"000000000",
  15120=>"101000000",
  15121=>"000001000",
  15122=>"110111111",
  15123=>"101001001",
  15124=>"001101011",
  15125=>"110100011",
  15126=>"001111110",
  15127=>"000000001",
  15128=>"001111111",
  15129=>"111111111",
  15130=>"111111111",
  15131=>"111111111",
  15132=>"111011111",
  15133=>"111111011",
  15134=>"000000001",
  15135=>"000111111",
  15136=>"000011011",
  15137=>"111110000",
  15138=>"111111111",
  15139=>"101111111",
  15140=>"111110000",
  15141=>"110110001",
  15142=>"000110000",
  15143=>"010111111",
  15144=>"000010000",
  15145=>"000000000",
  15146=>"011111111",
  15147=>"001011111",
  15148=>"000000000",
  15149=>"100110110",
  15150=>"000111000",
  15151=>"000000000",
  15152=>"111111111",
  15153=>"000000000",
  15154=>"001000100",
  15155=>"111111101",
  15156=>"111000000",
  15157=>"011011111",
  15158=>"000111111",
  15159=>"000000001",
  15160=>"000000010",
  15161=>"000000000",
  15162=>"000000111",
  15163=>"111110111",
  15164=>"111111011",
  15165=>"000000010",
  15166=>"000000000",
  15167=>"111100101",
  15168=>"111111111",
  15169=>"100000000",
  15170=>"011011111",
  15171=>"000010111",
  15172=>"110110000",
  15173=>"011111011",
  15174=>"111110000",
  15175=>"000001001",
  15176=>"000000000",
  15177=>"000011011",
  15178=>"000000111",
  15179=>"100110000",
  15180=>"011111111",
  15181=>"000111111",
  15182=>"111100101",
  15183=>"000010000",
  15184=>"011001000",
  15185=>"000101101",
  15186=>"000010000",
  15187=>"011001001",
  15188=>"001111111",
  15189=>"111110011",
  15190=>"000000111",
  15191=>"100101100",
  15192=>"111111111",
  15193=>"101000000",
  15194=>"111000011",
  15195=>"111100100",
  15196=>"111100100",
  15197=>"111111111",
  15198=>"000111111",
  15199=>"110110010",
  15200=>"110000100",
  15201=>"111111011",
  15202=>"110110011",
  15203=>"000000000",
  15204=>"001001001",
  15205=>"000011011",
  15206=>"100000000",
  15207=>"000000010",
  15208=>"001001000",
  15209=>"101000001",
  15210=>"111111111",
  15211=>"011111111",
  15212=>"111111111",
  15213=>"000000111",
  15214=>"111000101",
  15215=>"000000000",
  15216=>"000000000",
  15217=>"111111111",
  15218=>"000100000",
  15219=>"110111111",
  15220=>"000000000",
  15221=>"000000111",
  15222=>"110100000",
  15223=>"110110100",
  15224=>"111100000",
  15225=>"000000000",
  15226=>"000000000",
  15227=>"101101000",
  15228=>"111001000",
  15229=>"000001001",
  15230=>"111001000",
  15231=>"111111111",
  15232=>"110110111",
  15233=>"110111111",
  15234=>"100100100",
  15235=>"000000000",
  15236=>"110000000",
  15237=>"000111111",
  15238=>"000000110",
  15239=>"001001001",
  15240=>"111011000",
  15241=>"111000000",
  15242=>"111100100",
  15243=>"000000000",
  15244=>"000000000",
  15245=>"110111110",
  15246=>"111110111",
  15247=>"111000100",
  15248=>"111000000",
  15249=>"000000000",
  15250=>"100111111",
  15251=>"111111111",
  15252=>"110110000",
  15253=>"001111111",
  15254=>"111100110",
  15255=>"010000101",
  15256=>"111111110",
  15257=>"000000010",
  15258=>"111111111",
  15259=>"000000111",
  15260=>"111110000",
  15261=>"010000000",
  15262=>"101101101",
  15263=>"001000000",
  15264=>"000000000",
  15265=>"011001011",
  15266=>"111110100",
  15267=>"000000111",
  15268=>"111111110",
  15269=>"000111101",
  15270=>"000111011",
  15271=>"001011111",
  15272=>"111111111",
  15273=>"011010110",
  15274=>"000000000",
  15275=>"001001101",
  15276=>"111111000",
  15277=>"001000111",
  15278=>"000000011",
  15279=>"011011000",
  15280=>"111100111",
  15281=>"000000000",
  15282=>"000000000",
  15283=>"000000000",
  15284=>"110100100",
  15285=>"110110010",
  15286=>"101000000",
  15287=>"111111111",
  15288=>"000000000",
  15289=>"001010000",
  15290=>"111000000",
  15291=>"000000000",
  15292=>"000100100",
  15293=>"111111010",
  15294=>"111111111",
  15295=>"000010010",
  15296=>"000000000",
  15297=>"111101111",
  15298=>"110111111",
  15299=>"111111000",
  15300=>"000000001",
  15301=>"100000010",
  15302=>"111111111",
  15303=>"000010011",
  15304=>"000001001",
  15305=>"111111111",
  15306=>"111001000",
  15307=>"010000000",
  15308=>"000000110",
  15309=>"110100000",
  15310=>"001000000",
  15311=>"000000111",
  15312=>"111111111",
  15313=>"000100000",
  15314=>"111111111",
  15315=>"010000000",
  15316=>"000000000",
  15317=>"110010000",
  15318=>"111100100",
  15319=>"111111000",
  15320=>"111111111",
  15321=>"111100100",
  15322=>"001101000",
  15323=>"111111111",
  15324=>"100100000",
  15325=>"100000000",
  15326=>"111111001",
  15327=>"111110100",
  15328=>"000110110",
  15329=>"111111000",
  15330=>"111011010",
  15331=>"111111011",
  15332=>"011010000",
  15333=>"111111111",
  15334=>"000010010",
  15335=>"111110000",
  15336=>"000000000",
  15337=>"111101000",
  15338=>"001011011",
  15339=>"000100100",
  15340=>"000010110",
  15341=>"011111111",
  15342=>"111111111",
  15343=>"000111111",
  15344=>"000000000",
  15345=>"110000000",
  15346=>"100111100",
  15347=>"111001000",
  15348=>"000000000",
  15349=>"001000000",
  15350=>"001001111",
  15351=>"000000000",
  15352=>"110000000",
  15353=>"000000010",
  15354=>"000000000",
  15355=>"000000000",
  15356=>"100111100",
  15357=>"111010100",
  15358=>"001111111",
  15359=>"001001111",
  15360=>"110110110",
  15361=>"001111111",
  15362=>"111111111",
  15363=>"001000000",
  15364=>"000000000",
  15365=>"001000000",
  15366=>"000000000",
  15367=>"100001001",
  15368=>"111111111",
  15369=>"111111000",
  15370=>"111000000",
  15371=>"111010011",
  15372=>"111100110",
  15373=>"111000001",
  15374=>"100000000",
  15375=>"111111111",
  15376=>"000000000",
  15377=>"000000000",
  15378=>"010111111",
  15379=>"101000000",
  15380=>"111000000",
  15381=>"111111101",
  15382=>"111111111",
  15383=>"001011111",
  15384=>"111111111",
  15385=>"100100000",
  15386=>"111100100",
  15387=>"000000001",
  15388=>"001001111",
  15389=>"011001011",
  15390=>"100100100",
  15391=>"000000000",
  15392=>"110111111",
  15393=>"100010010",
  15394=>"001111111",
  15395=>"000000100",
  15396=>"001001000",
  15397=>"110110110",
  15398=>"000000111",
  15399=>"000110000",
  15400=>"111111011",
  15401=>"000000000",
  15402=>"111010111",
  15403=>"011011011",
  15404=>"000100001",
  15405=>"111111011",
  15406=>"001001001",
  15407=>"111000000",
  15408=>"000011111",
  15409=>"111101001",
  15410=>"011001001",
  15411=>"111111111",
  15412=>"010110010",
  15413=>"001001000",
  15414=>"000000000",
  15415=>"000000000",
  15416=>"111011000",
  15417=>"000110110",
  15418=>"111100111",
  15419=>"001001111",
  15420=>"110100110",
  15421=>"110010000",
  15422=>"010011111",
  15423=>"101101101",
  15424=>"000011111",
  15425=>"000000100",
  15426=>"000101111",
  15427=>"110110010",
  15428=>"001001111",
  15429=>"110111110",
  15430=>"000000000",
  15431=>"101001101",
  15432=>"001101111",
  15433=>"101001001",
  15434=>"111111111",
  15435=>"111111001",
  15436=>"001011001",
  15437=>"000000100",
  15438=>"011000000",
  15439=>"000110111",
  15440=>"100000000",
  15441=>"000001101",
  15442=>"000001000",
  15443=>"100110110",
  15444=>"111111000",
  15445=>"101100000",
  15446=>"100011111",
  15447=>"000000000",
  15448=>"111011011",
  15449=>"111101111",
  15450=>"111111000",
  15451=>"000000000",
  15452=>"010110011",
  15453=>"000000000",
  15454=>"101111111",
  15455=>"111111000",
  15456=>"110100000",
  15457=>"111101001",
  15458=>"011011100",
  15459=>"111001000",
  15460=>"000001011",
  15461=>"000011111",
  15462=>"111110000",
  15463=>"000111011",
  15464=>"011011111",
  15465=>"010000010",
  15466=>"100110010",
  15467=>"111110000",
  15468=>"000000000",
  15469=>"111111111",
  15470=>"000000000",
  15471=>"111011000",
  15472=>"111111111",
  15473=>"111010000",
  15474=>"111010010",
  15475=>"111111111",
  15476=>"000000000",
  15477=>"111000000",
  15478=>"001000101",
  15479=>"100100111",
  15480=>"111111111",
  15481=>"000110110",
  15482=>"001000000",
  15483=>"111101000",
  15484=>"100110110",
  15485=>"000000000",
  15486=>"000000000",
  15487=>"001110011",
  15488=>"101101000",
  15489=>"100010000",
  15490=>"011000000",
  15491=>"000111011",
  15492=>"101001101",
  15493=>"000000000",
  15494=>"001001001",
  15495=>"011111111",
  15496=>"001000000",
  15497=>"000000111",
  15498=>"000110111",
  15499=>"000000000",
  15500=>"110110111",
  15501=>"000000000",
  15502=>"111111111",
  15503=>"111111111",
  15504=>"110111111",
  15505=>"000010001",
  15506=>"000000110",
  15507=>"000000000",
  15508=>"000000111",
  15509=>"001000000",
  15510=>"001001101",
  15511=>"001000000",
  15512=>"000000101",
  15513=>"000000000",
  15514=>"111111111",
  15515=>"000011011",
  15516=>"111111111",
  15517=>"000000000",
  15518=>"111111000",
  15519=>"111111111",
  15520=>"000100100",
  15521=>"000111111",
  15522=>"111111011",
  15523=>"111111111",
  15524=>"011000000",
  15525=>"111001000",
  15526=>"000010111",
  15527=>"111111000",
  15528=>"000000000",
  15529=>"001001000",
  15530=>"001000000",
  15531=>"111111111",
  15532=>"111001000",
  15533=>"001111111",
  15534=>"000000000",
  15535=>"001011001",
  15536=>"111111000",
  15537=>"100100100",
  15538=>"011111111",
  15539=>"111111111",
  15540=>"111111111",
  15541=>"111100000",
  15542=>"000000000",
  15543=>"010000100",
  15544=>"011011111",
  15545=>"000000100",
  15546=>"000001000",
  15547=>"100010110",
  15548=>"111000000",
  15549=>"100110111",
  15550=>"111111010",
  15551=>"100100110",
  15552=>"101011001",
  15553=>"010000000",
  15554=>"101101011",
  15555=>"001011000",
  15556=>"111111111",
  15557=>"000000110",
  15558=>"111111000",
  15559=>"000000011",
  15560=>"111111111",
  15561=>"000000000",
  15562=>"001001100",
  15563=>"001110111",
  15564=>"111111010",
  15565=>"000000000",
  15566=>"000000101",
  15567=>"000000000",
  15568=>"101100111",
  15569=>"001001000",
  15570=>"001011110",
  15571=>"111111111",
  15572=>"011111111",
  15573=>"111000001",
  15574=>"000011111",
  15575=>"110100000",
  15576=>"111000000",
  15577=>"000010110",
  15578=>"101000000",
  15579=>"000000000",
  15580=>"110110111",
  15581=>"111110010",
  15582=>"110000000",
  15583=>"001000000",
  15584=>"011000000",
  15585=>"011000010",
  15586=>"000000000",
  15587=>"111110000",
  15588=>"000000000",
  15589=>"000011011",
  15590=>"001011001",
  15591=>"110111110",
  15592=>"000110111",
  15593=>"000000000",
  15594=>"111111111",
  15595=>"001001010",
  15596=>"010110110",
  15597=>"110000000",
  15598=>"111111101",
  15599=>"000000111",
  15600=>"000000100",
  15601=>"000000111",
  15602=>"111000100",
  15603=>"011011001",
  15604=>"011001100",
  15605=>"111110001",
  15606=>"111111110",
  15607=>"101001000",
  15608=>"011111101",
  15609=>"111011000",
  15610=>"000000000",
  15611=>"111111111",
  15612=>"111111110",
  15613=>"000000000",
  15614=>"110000000",
  15615=>"101111111",
  15616=>"100100100",
  15617=>"100100000",
  15618=>"111111001",
  15619=>"111111001",
  15620=>"111011111",
  15621=>"111000000",
  15622=>"111110100",
  15623=>"100110011",
  15624=>"110000000",
  15625=>"011011000",
  15626=>"001000101",
  15627=>"111111111",
  15628=>"000001111",
  15629=>"000000000",
  15630=>"001111111",
  15631=>"000000000",
  15632=>"000000000",
  15633=>"110000000",
  15634=>"101101101",
  15635=>"111111000",
  15636=>"111111111",
  15637=>"111100000",
  15638=>"111011001",
  15639=>"000000001",
  15640=>"110110010",
  15641=>"000000000",
  15642=>"001001001",
  15643=>"111111111",
  15644=>"000000010",
  15645=>"010011010",
  15646=>"110110000",
  15647=>"000111011",
  15648=>"010011001",
  15649=>"110110011",
  15650=>"000000010",
  15651=>"000000001",
  15652=>"000000011",
  15653=>"001001001",
  15654=>"001001001",
  15655=>"110110110",
  15656=>"000000000",
  15657=>"000100010",
  15658=>"001011001",
  15659=>"001001000",
  15660=>"000011010",
  15661=>"000000000",
  15662=>"111011111",
  15663=>"101000001",
  15664=>"101111001",
  15665=>"111001000",
  15666=>"011011011",
  15667=>"001000000",
  15668=>"100000000",
  15669=>"110111111",
  15670=>"010000000",
  15671=>"110110011",
  15672=>"111011001",
  15673=>"111111101",
  15674=>"000000000",
  15675=>"111111111",
  15676=>"000011010",
  15677=>"110110010",
  15678=>"000001011",
  15679=>"100111111",
  15680=>"111111111",
  15681=>"111111111",
  15682=>"111111111",
  15683=>"000001001",
  15684=>"000001001",
  15685=>"111010000",
  15686=>"000011011",
  15687=>"111111011",
  15688=>"111101101",
  15689=>"111111111",
  15690=>"000000001",
  15691=>"000000000",
  15692=>"000000000",
  15693=>"000000000",
  15694=>"001111111",
  15695=>"001001000",
  15696=>"000000000",
  15697=>"011000100",
  15698=>"110110010",
  15699=>"111000011",
  15700=>"111010000",
  15701=>"011011011",
  15702=>"001001001",
  15703=>"001001001",
  15704=>"111111111",
  15705=>"011111011",
  15706=>"000010000",
  15707=>"010110010",
  15708=>"111000010",
  15709=>"000000000",
  15710=>"000000111",
  15711=>"111101011",
  15712=>"110110110",
  15713=>"111111111",
  15714=>"001001011",
  15715=>"111111111",
  15716=>"001001101",
  15717=>"100000000",
  15718=>"011111001",
  15719=>"000011011",
  15720=>"100100100",
  15721=>"011011111",
  15722=>"000000000",
  15723=>"111011011",
  15724=>"111111010",
  15725=>"100111111",
  15726=>"000111111",
  15727=>"111111111",
  15728=>"101001001",
  15729=>"000011000",
  15730=>"000000000",
  15731=>"100100000",
  15732=>"000000110",
  15733=>"111000000",
  15734=>"001001001",
  15735=>"001001000",
  15736=>"001101111",
  15737=>"011000000",
  15738=>"111111111",
  15739=>"111111111",
  15740=>"110111011",
  15741=>"111111111",
  15742=>"100111111",
  15743=>"100111111",
  15744=>"000000000",
  15745=>"001111111",
  15746=>"001100110",
  15747=>"000001111",
  15748=>"010000000",
  15749=>"010011000",
  15750=>"001000001",
  15751=>"101110010",
  15752=>"001000100",
  15753=>"111111111",
  15754=>"000101111",
  15755=>"111111001",
  15756=>"001001111",
  15757=>"011001000",
  15758=>"111111010",
  15759=>"111111111",
  15760=>"001000000",
  15761=>"111111111",
  15762=>"101000000",
  15763=>"011011000",
  15764=>"001001001",
  15765=>"000011000",
  15766=>"001000010",
  15767=>"001000000",
  15768=>"110110010",
  15769=>"111111101",
  15770=>"010010100",
  15771=>"000000000",
  15772=>"000100110",
  15773=>"111111101",
  15774=>"000000000",
  15775=>"000000000",
  15776=>"111111111",
  15777=>"011011001",
  15778=>"111111111",
  15779=>"000001000",
  15780=>"001001000",
  15781=>"010011111",
  15782=>"111100100",
  15783=>"101001000",
  15784=>"000000000",
  15785=>"110000000",
  15786=>"111100000",
  15787=>"001001000",
  15788=>"001000000",
  15789=>"101001000",
  15790=>"110010110",
  15791=>"010000000",
  15792=>"111111011",
  15793=>"111111101",
  15794=>"000000000",
  15795=>"111000000",
  15796=>"000000000",
  15797=>"111111000",
  15798=>"000000001",
  15799=>"101001001",
  15800=>"000000000",
  15801=>"011100110",
  15802=>"110110100",
  15803=>"110111111",
  15804=>"001111111",
  15805=>"001011011",
  15806=>"000000000",
  15807=>"111111111",
  15808=>"111011001",
  15809=>"000000000",
  15810=>"011011111",
  15811=>"101001000",
  15812=>"000000000",
  15813=>"111000000",
  15814=>"111110010",
  15815=>"011001000",
  15816=>"111011000",
  15817=>"110010001",
  15818=>"000000000",
  15819=>"000000111",
  15820=>"111111000",
  15821=>"001001001",
  15822=>"011000000",
  15823=>"000000000",
  15824=>"111011010",
  15825=>"001001000",
  15826=>"101111110",
  15827=>"000000011",
  15828=>"111111111",
  15829=>"000000011",
  15830=>"100100100",
  15831=>"101111111",
  15832=>"000000000",
  15833=>"111111000",
  15834=>"000000010",
  15835=>"011011100",
  15836=>"000000000",
  15837=>"110110010",
  15838=>"111111001",
  15839=>"100000000",
  15840=>"001000000",
  15841=>"000000000",
  15842=>"000111111",
  15843=>"111111111",
  15844=>"000000000",
  15845=>"111110110",
  15846=>"100100010",
  15847=>"111111111",
  15848=>"000000000",
  15849=>"000000000",
  15850=>"000000000",
  15851=>"000000001",
  15852=>"000000000",
  15853=>"100100001",
  15854=>"110111110",
  15855=>"111111111",
  15856=>"000111111",
  15857=>"111011000",
  15858=>"100110111",
  15859=>"000011011",
  15860=>"101001001",
  15861=>"110101100",
  15862=>"000000100",
  15863=>"100100100",
  15864=>"111111000",
  15865=>"100000000",
  15866=>"111111111",
  15867=>"111101111",
  15868=>"001001000",
  15869=>"001000001",
  15870=>"000000110",
  15871=>"000111111",
  15872=>"000000010",
  15873=>"000011101",
  15874=>"111111111",
  15875=>"110100101",
  15876=>"100001001",
  15877=>"010110111",
  15878=>"100010000",
  15879=>"111111011",
  15880=>"101001101",
  15881=>"110110000",
  15882=>"101001111",
  15883=>"010001111",
  15884=>"011011111",
  15885=>"101101100",
  15886=>"100111111",
  15887=>"101101111",
  15888=>"000100100",
  15889=>"000000000",
  15890=>"111111110",
  15891=>"011001001",
  15892=>"001001001",
  15893=>"111010010",
  15894=>"000110110",
  15895=>"111111111",
  15896=>"111001100",
  15897=>"011110100",
  15898=>"000000111",
  15899=>"111100000",
  15900=>"101101001",
  15901=>"001001111",
  15902=>"111010010",
  15903=>"000100111",
  15904=>"101101000",
  15905=>"101001001",
  15906=>"001000110",
  15907=>"111111111",
  15908=>"001100111",
  15909=>"111111100",
  15910=>"000001001",
  15911=>"100110110",
  15912=>"100100100",
  15913=>"111000000",
  15914=>"101101101",
  15915=>"101101100",
  15916=>"010010011",
  15917=>"100100110",
  15918=>"010000000",
  15919=>"000110111",
  15920=>"100000110",
  15921=>"111111111",
  15922=>"110110110",
  15923=>"111111110",
  15924=>"111011010",
  15925=>"010010010",
  15926=>"000000101",
  15927=>"000101101",
  15928=>"001011001",
  15929=>"101101011",
  15930=>"000100101",
  15931=>"011000000",
  15932=>"010010010",
  15933=>"100100000",
  15934=>"100110111",
  15935=>"101001100",
  15936=>"101101111",
  15937=>"011001001",
  15938=>"000000111",
  15939=>"101100000",
  15940=>"100111111",
  15941=>"110000000",
  15942=>"101101100",
  15943=>"101101101",
  15944=>"000000000",
  15945=>"101001101",
  15946=>"001101111",
  15947=>"101001000",
  15948=>"111111010",
  15949=>"100100001",
  15950=>"000010110",
  15951=>"001011001",
  15952=>"111111000",
  15953=>"111111111",
  15954=>"100100100",
  15955=>"010010110",
  15956=>"100101101",
  15957=>"101101101",
  15958=>"100101101",
  15959=>"010010010",
  15960=>"000000000",
  15961=>"111101101",
  15962=>"001000000",
  15963=>"000101100",
  15964=>"000101101",
  15965=>"111111111",
  15966=>"001001001",
  15967=>"000100100",
  15968=>"101101110",
  15969=>"000001001",
  15970=>"111111101",
  15971=>"000010111",
  15972=>"010000000",
  15973=>"101100000",
  15974=>"101101000",
  15975=>"110110000",
  15976=>"100100001",
  15977=>"011001000",
  15978=>"111111000",
  15979=>"000000001",
  15980=>"011011101",
  15981=>"010010010",
  15982=>"000010110",
  15983=>"111111000",
  15984=>"011011111",
  15985=>"110010010",
  15986=>"011001001",
  15987=>"000000000",
  15988=>"100101101",
  15989=>"001111111",
  15990=>"011001101",
  15991=>"100101001",
  15992=>"000100111",
  15993=>"100001001",
  15994=>"101101000",
  15995=>"011111000",
  15996=>"010010010",
  15997=>"111111101",
  15998=>"111101111",
  15999=>"000010010",
  16000=>"010010010",
  16001=>"101101101",
  16002=>"100000100",
  16003=>"000110110",
  16004=>"101101100",
  16005=>"100000101",
  16006=>"000000010",
  16007=>"001101101",
  16008=>"000000000",
  16009=>"111111001",
  16010=>"100100101",
  16011=>"011111101",
  16012=>"010010010",
  16013=>"110110111",
  16014=>"101101001",
  16015=>"000001000",
  16016=>"011010010",
  16017=>"000110111",
  16018=>"110000001",
  16019=>"101101101",
  16020=>"000001101",
  16021=>"100110100",
  16022=>"011010000",
  16023=>"011010000",
  16024=>"111011110",
  16025=>"111111111",
  16026=>"111101101",
  16027=>"001001001",
  16028=>"101101001",
  16029=>"100101101",
  16030=>"101101001",
  16031=>"100100100",
  16032=>"100101001",
  16033=>"000100110",
  16034=>"000000000",
  16035=>"100100100",
  16036=>"001101001",
  16037=>"100111100",
  16038=>"011010110",
  16039=>"010110110",
  16040=>"000000000",
  16041=>"111001000",
  16042=>"101101101",
  16043=>"000001010",
  16044=>"101101111",
  16045=>"001011011",
  16046=>"000010011",
  16047=>"101001000",
  16048=>"000100111",
  16049=>"110111000",
  16050=>"000010000",
  16051=>"110110110",
  16052=>"111101101",
  16053=>"101101101",
  16054=>"000000010",
  16055=>"101111110",
  16056=>"001101101",
  16057=>"110110010",
  16058=>"101100100",
  16059=>"101101000",
  16060=>"111111011",
  16061=>"000000000",
  16062=>"100100101",
  16063=>"000010010",
  16064=>"111100000",
  16065=>"011101111",
  16066=>"000000000",
  16067=>"100110010",
  16068=>"011010011",
  16069=>"000001001",
  16070=>"001101001",
  16071=>"101111111",
  16072=>"010110110",
  16073=>"001001000",
  16074=>"101101101",
  16075=>"010110010",
  16076=>"111111111",
  16077=>"000100100",
  16078=>"100100101",
  16079=>"100100100",
  16080=>"100101101",
  16081=>"010010010",
  16082=>"000111100",
  16083=>"110110110",
  16084=>"000100100",
  16085=>"101111111",
  16086=>"011010010",
  16087=>"111111000",
  16088=>"100100000",
  16089=>"111101111",
  16090=>"000000000",
  16091=>"100101111",
  16092=>"000000000",
  16093=>"010010010",
  16094=>"000001001",
  16095=>"100101001",
  16096=>"000001011",
  16097=>"101101101",
  16098=>"111110111",
  16099=>"100000000",
  16100=>"101101101",
  16101=>"110000100",
  16102=>"100101001",
  16103=>"000101001",
  16104=>"111101100",
  16105=>"110010011",
  16106=>"000110000",
  16107=>"101000000",
  16108=>"000110110",
  16109=>"000101101",
  16110=>"110010000",
  16111=>"000000000",
  16112=>"001101100",
  16113=>"100101101",
  16114=>"101001000",
  16115=>"101101001",
  16116=>"111000000",
  16117=>"000011111",
  16118=>"011010000",
  16119=>"100100000",
  16120=>"110110111",
  16121=>"100100100",
  16122=>"010000000",
  16123=>"010010010",
  16124=>"111110110",
  16125=>"000001111",
  16126=>"100101000",
  16127=>"111110000",
  16128=>"101001000",
  16129=>"011011001",
  16130=>"101101101",
  16131=>"100100111",
  16132=>"000000100",
  16133=>"100100101",
  16134=>"101101111",
  16135=>"000011000",
  16136=>"101101100",
  16137=>"100110110",
  16138=>"000000000",
  16139=>"101101111",
  16140=>"110000111",
  16141=>"000101101",
  16142=>"000000000",
  16143=>"000000000",
  16144=>"000101100",
  16145=>"000100000",
  16146=>"011001001",
  16147=>"100101101",
  16148=>"100100100",
  16149=>"100101101",
  16150=>"011011011",
  16151=>"101111111",
  16152=>"010011110",
  16153=>"111101101",
  16154=>"110000000",
  16155=>"110110101",
  16156=>"110011010",
  16157=>"101111101",
  16158=>"100101111",
  16159=>"000101101",
  16160=>"001011001",
  16161=>"000001011",
  16162=>"111111110",
  16163=>"111111111",
  16164=>"101001001",
  16165=>"001001100",
  16166=>"110111001",
  16167=>"100110100",
  16168=>"110111100",
  16169=>"100101000",
  16170=>"001001001",
  16171=>"001001000",
  16172=>"001100000",
  16173=>"110010110",
  16174=>"100100000",
  16175=>"000010010",
  16176=>"010011010",
  16177=>"000000000",
  16178=>"000000000",
  16179=>"001101101",
  16180=>"000000111",
  16181=>"011111101",
  16182=>"100111111",
  16183=>"100010110",
  16184=>"001000000",
  16185=>"001101111",
  16186=>"100100101",
  16187=>"000000000",
  16188=>"000000100",
  16189=>"110100000",
  16190=>"101101101",
  16191=>"100110010",
  16192=>"111101111",
  16193=>"011011000",
  16194=>"001110110",
  16195=>"010010010",
  16196=>"010010010",
  16197=>"011000000",
  16198=>"000000000",
  16199=>"001111111",
  16200=>"100000000",
  16201=>"100101101",
  16202=>"101100101",
  16203=>"110110110",
  16204=>"100101101",
  16205=>"010110110",
  16206=>"101101000",
  16207=>"110111110",
  16208=>"110010010",
  16209=>"101100001",
  16210=>"110101100",
  16211=>"000000000",
  16212=>"010011011",
  16213=>"110110111",
  16214=>"101000000",
  16215=>"111000001",
  16216=>"111011010",
  16217=>"000000000",
  16218=>"001000110",
  16219=>"101101110",
  16220=>"110110000",
  16221=>"111111101",
  16222=>"000110110",
  16223=>"110110111",
  16224=>"000100100",
  16225=>"101001001",
  16226=>"110110110",
  16227=>"011010010",
  16228=>"100110000",
  16229=>"000100100",
  16230=>"101101111",
  16231=>"101101111",
  16232=>"001011011",
  16233=>"101101111",
  16234=>"100100001",
  16235=>"000000001",
  16236=>"100110110",
  16237=>"101111001",
  16238=>"100101111",
  16239=>"000001001",
  16240=>"000100101",
  16241=>"111100000",
  16242=>"000000000",
  16243=>"111111110",
  16244=>"100100000",
  16245=>"111110110",
  16246=>"100000111",
  16247=>"101101001",
  16248=>"010000000",
  16249=>"000000001",
  16250=>"000000000",
  16251=>"101101101",
  16252=>"100101101",
  16253=>"111111111",
  16254=>"010000000",
  16255=>"111111111",
  16256=>"111000000",
  16257=>"000000000",
  16258=>"000000000",
  16259=>"001100101",
  16260=>"000001101",
  16261=>"000000000",
  16262=>"101101001",
  16263=>"111111101",
  16264=>"110110001",
  16265=>"110110111",
  16266=>"001001001",
  16267=>"000100100",
  16268=>"111001111",
  16269=>"100011011",
  16270=>"100100110",
  16271=>"111111110",
  16272=>"100000000",
  16273=>"101111111",
  16274=>"010000110",
  16275=>"100111101",
  16276=>"000010110",
  16277=>"000110110",
  16278=>"111101101",
  16279=>"001011011",
  16280=>"001100001",
  16281=>"101101101",
  16282=>"000101100",
  16283=>"101101101",
  16284=>"100000100",
  16285=>"001001001",
  16286=>"001001111",
  16287=>"000001001",
  16288=>"100100100",
  16289=>"011011011",
  16290=>"000011011",
  16291=>"101101111",
  16292=>"101101101",
  16293=>"111111000",
  16294=>"110110010",
  16295=>"111111100",
  16296=>"011010100",
  16297=>"101111111",
  16298=>"010010011",
  16299=>"100101101",
  16300=>"000110110",
  16301=>"100101000",
  16302=>"100101001",
  16303=>"100100100",
  16304=>"100000100",
  16305=>"000111000",
  16306=>"000000000",
  16307=>"000100101",
  16308=>"101100100",
  16309=>"111000000",
  16310=>"011111001",
  16311=>"001001111",
  16312=>"101101100",
  16313=>"111111101",
  16314=>"100100100",
  16315=>"011110000",
  16316=>"111011111",
  16317=>"100100101",
  16318=>"010010011",
  16319=>"001001011",
  16320=>"101001001",
  16321=>"010010010",
  16322=>"010010110",
  16323=>"010110111",
  16324=>"001101101",
  16325=>"111111011",
  16326=>"001001000",
  16327=>"011000000",
  16328=>"101000011",
  16329=>"100000001",
  16330=>"101100100",
  16331=>"000000010",
  16332=>"101000000",
  16333=>"001111001",
  16334=>"100000000",
  16335=>"101101101",
  16336=>"010110110",
  16337=>"111110110",
  16338=>"101101100",
  16339=>"111010010",
  16340=>"011011011",
  16341=>"000101101",
  16342=>"101101101",
  16343=>"100011111",
  16344=>"110010110",
  16345=>"100101101",
  16346=>"100100101",
  16347=>"000001000",
  16348=>"100100111",
  16349=>"000110010",
  16350=>"111111011",
  16351=>"001111011",
  16352=>"011011011",
  16353=>"100110010",
  16354=>"000100111",
  16355=>"000110100",
  16356=>"001101101",
  16357=>"100100100",
  16358=>"001111111",
  16359=>"101101100",
  16360=>"000010011",
  16361=>"100101100",
  16362=>"100101101",
  16363=>"000111111",
  16364=>"000100101",
  16365=>"111101100",
  16366=>"010010010",
  16367=>"000000101",
  16368=>"110111010",
  16369=>"000110111",
  16370=>"100000111",
  16371=>"000101100",
  16372=>"000000110",
  16373=>"100111110",
  16374=>"111100110",
  16375=>"001001010",
  16376=>"111111111",
  16377=>"110110110",
  16378=>"001111111",
  16379=>"001000111",
  16380=>"001100000",
  16381=>"111111011",
  16382=>"100000000",
  16383=>"000000100",
  16384=>"100110111",
  16385=>"111111111",
  16386=>"111010010",
  16387=>"001001111",
  16388=>"111111111",
  16389=>"111001001",
  16390=>"111111101",
  16391=>"000000111",
  16392=>"010111111",
  16393=>"101101101",
  16394=>"010110111",
  16395=>"111111100",
  16396=>"010000000",
  16397=>"101101000",
  16398=>"111111111",
  16399=>"011101001",
  16400=>"010111111",
  16401=>"000100110",
  16402=>"100100000",
  16403=>"111111110",
  16404=>"110010000",
  16405=>"100000000",
  16406=>"001010010",
  16407=>"101001000",
  16408=>"000000011",
  16409=>"001001000",
  16410=>"111110100",
  16411=>"100110101",
  16412=>"101001101",
  16413=>"111011010",
  16414=>"110100100",
  16415=>"110110000",
  16416=>"001001001",
  16417=>"000000000",
  16418=>"001001001",
  16419=>"011010011",
  16420=>"100000110",
  16421=>"000000000",
  16422=>"001001001",
  16423=>"010110110",
  16424=>"011000111",
  16425=>"000010010",
  16426=>"101101101",
  16427=>"011011111",
  16428=>"101100000",
  16429=>"001001101",
  16430=>"110110010",
  16431=>"111111110",
  16432=>"111101100",
  16433=>"000101110",
  16434=>"011001001",
  16435=>"110000000",
  16436=>"000000000",
  16437=>"011011011",
  16438=>"001001011",
  16439=>"000110110",
  16440=>"101101001",
  16441=>"100100111",
  16442=>"111111111",
  16443=>"100011001",
  16444=>"111000000",
  16445=>"101101001",
  16446=>"110100000",
  16447=>"101101001",
  16448=>"001001100",
  16449=>"000000010",
  16450=>"100101101",
  16451=>"101111111",
  16452=>"010010111",
  16453=>"000000000",
  16454=>"111111100",
  16455=>"110010010",
  16456=>"011011111",
  16457=>"000000000",
  16458=>"010110111",
  16459=>"110110100",
  16460=>"101101001",
  16461=>"100111111",
  16462=>"110111111",
  16463=>"000000000",
  16464=>"000111111",
  16465=>"001000000",
  16466=>"100101111",
  16467=>"101101101",
  16468=>"111111101",
  16469=>"000000111",
  16470=>"111100010",
  16471=>"011111111",
  16472=>"111001111",
  16473=>"100000000",
  16474=>"000000000",
  16475=>"000101001",
  16476=>"101000000",
  16477=>"000000000",
  16478=>"101101000",
  16479=>"001001001",
  16480=>"000010011",
  16481=>"000000000",
  16482=>"111111111",
  16483=>"100100001",
  16484=>"000000111",
  16485=>"000000000",
  16486=>"111100100",
  16487=>"000100100",
  16488=>"110100000",
  16489=>"110110110",
  16490=>"101101100",
  16491=>"111110110",
  16492=>"001001001",
  16493=>"000000000",
  16494=>"100100111",
  16495=>"110111110",
  16496=>"000100000",
  16497=>"010000010",
  16498=>"000000000",
  16499=>"110110000",
  16500=>"001001000",
  16501=>"110111111",
  16502=>"101100111",
  16503=>"101111111",
  16504=>"001001101",
  16505=>"000000001",
  16506=>"011001001",
  16507=>"111110100",
  16508=>"001001011",
  16509=>"100111011",
  16510=>"110110110",
  16511=>"100101111",
  16512=>"000000100",
  16513=>"110111110",
  16514=>"110110110",
  16515=>"111011000",
  16516=>"001000100",
  16517=>"000000000",
  16518=>"001000111",
  16519=>"110110011",
  16520=>"010000000",
  16521=>"000000001",
  16522=>"000100100",
  16523=>"111001000",
  16524=>"101101001",
  16525=>"001001000",
  16526=>"001000010",
  16527=>"111111110",
  16528=>"110111001",
  16529=>"101101101",
  16530=>"001000000",
  16531=>"101001001",
  16532=>"001101100",
  16533=>"000100001",
  16534=>"110111011",
  16535=>"111010010",
  16536=>"111111111",
  16537=>"111110110",
  16538=>"001110100",
  16539=>"000000001",
  16540=>"111101001",
  16541=>"010000000",
  16542=>"010000100",
  16543=>"001101101",
  16544=>"000000000",
  16545=>"000001101",
  16546=>"001101100",
  16547=>"000001001",
  16548=>"111110000",
  16549=>"111101111",
  16550=>"111111111",
  16551=>"001101001",
  16552=>"110100100",
  16553=>"110110110",
  16554=>"000010010",
  16555=>"111101101",
  16556=>"001000000",
  16557=>"000000000",
  16558=>"001100100",
  16559=>"001011011",
  16560=>"000000001",
  16561=>"100100111",
  16562=>"001001001",
  16563=>"111111101",
  16564=>"000100100",
  16565=>"100100111",
  16566=>"010000000",
  16567=>"010000001",
  16568=>"000000000",
  16569=>"111010000",
  16570=>"111111000",
  16571=>"001001001",
  16572=>"000001001",
  16573=>"001001000",
  16574=>"000110010",
  16575=>"110110111",
  16576=>"000001011",
  16577=>"010110111",
  16578=>"000001011",
  16579=>"001111010",
  16580=>"100110100",
  16581=>"011110111",
  16582=>"000000000",
  16583=>"001001101",
  16584=>"110100000",
  16585=>"001000001",
  16586=>"101101111",
  16587=>"111111111",
  16588=>"001001001",
  16589=>"101101111",
  16590=>"101001001",
  16591=>"111100110",
  16592=>"110110111",
  16593=>"000000001",
  16594=>"111111111",
  16595=>"111111111",
  16596=>"001101111",
  16597=>"011000000",
  16598=>"010110110",
  16599=>"100000110",
  16600=>"111111110",
  16601=>"111111111",
  16602=>"111110110",
  16603=>"111111111",
  16604=>"000000000",
  16605=>"010110110",
  16606=>"101101101",
  16607=>"000000001",
  16608=>"001110111",
  16609=>"000000000",
  16610=>"111111111",
  16611=>"111000000",
  16612=>"101111111",
  16613=>"000000100",
  16614=>"111110111",
  16615=>"111010000",
  16616=>"111111101",
  16617=>"111110110",
  16618=>"000001111",
  16619=>"010010111",
  16620=>"100100000",
  16621=>"000010110",
  16622=>"111111111",
  16623=>"011001001",
  16624=>"000000000",
  16625=>"000100101",
  16626=>"111110000",
  16627=>"000000000",
  16628=>"101001001",
  16629=>"100100100",
  16630=>"110111110",
  16631=>"011001000",
  16632=>"010011111",
  16633=>"001101101",
  16634=>"111110000",
  16635=>"100101111",
  16636=>"000001001",
  16637=>"111111111",
  16638=>"101100100",
  16639=>"001011110",
  16640=>"011001000",
  16641=>"000000000",
  16642=>"000000100",
  16643=>"101001001",
  16644=>"100101101",
  16645=>"000101111",
  16646=>"110110000",
  16647=>"011111111",
  16648=>"010000111",
  16649=>"000000100",
  16650=>"111111111",
  16651=>"010010011",
  16652=>"001001000",
  16653=>"000000000",
  16654=>"000100100",
  16655=>"111100000",
  16656=>"011100100",
  16657=>"000100000",
  16658=>"001111111",
  16659=>"111111001",
  16660=>"100111111",
  16661=>"001001001",
  16662=>"000000000",
  16663=>"101101101",
  16664=>"001001001",
  16665=>"110110110",
  16666=>"101100000",
  16667=>"111111111",
  16668=>"001001011",
  16669=>"111111111",
  16670=>"110111110",
  16671=>"100101001",
  16672=>"000000000",
  16673=>"011011010",
  16674=>"000000000",
  16675=>"111111101",
  16676=>"010110110",
  16677=>"111000000",
  16678=>"101001111",
  16679=>"110010110",
  16680=>"000100101",
  16681=>"001101101",
  16682=>"111001000",
  16683=>"110110000",
  16684=>"000000000",
  16685=>"001001001",
  16686=>"111111111",
  16687=>"000000000",
  16688=>"011011011",
  16689=>"001001001",
  16690=>"110110010",
  16691=>"110110111",
  16692=>"000000001",
  16693=>"111110010",
  16694=>"111111111",
  16695=>"111111111",
  16696=>"000000000",
  16697=>"110110111",
  16698=>"000000000",
  16699=>"110110110",
  16700=>"110011011",
  16701=>"001001001",
  16702=>"010110110",
  16703=>"101001001",
  16704=>"101100101",
  16705=>"011101001",
  16706=>"000000110",
  16707=>"000000001",
  16708=>"000000001",
  16709=>"111111110",
  16710=>"100000000",
  16711=>"000000001",
  16712=>"100000000",
  16713=>"101100101",
  16714=>"000000001",
  16715=>"111101001",
  16716=>"110110100",
  16717=>"111101111",
  16718=>"001101101",
  16719=>"011111111",
  16720=>"001001001",
  16721=>"100100110",
  16722=>"000001001",
  16723=>"000000000",
  16724=>"001001001",
  16725=>"000000101",
  16726=>"111111111",
  16727=>"000000000",
  16728=>"110111111",
  16729=>"010011011",
  16730=>"101101101",
  16731=>"000010110",
  16732=>"000000100",
  16733=>"100110100",
  16734=>"110011111",
  16735=>"111111100",
  16736=>"000010110",
  16737=>"100101101",
  16738=>"011011011",
  16739=>"111111111",
  16740=>"001001011",
  16741=>"101001001",
  16742=>"010110110",
  16743=>"001001001",
  16744=>"000001001",
  16745=>"110100110",
  16746=>"101101101",
  16747=>"100100101",
  16748=>"001001111",
  16749=>"111101101",
  16750=>"000111111",
  16751=>"111110111",
  16752=>"100100100",
  16753=>"011111110",
  16754=>"000001111",
  16755=>"101101100",
  16756=>"110110100",
  16757=>"111111111",
  16758=>"000000001",
  16759=>"111111111",
  16760=>"010111111",
  16761=>"000000001",
  16762=>"111111111",
  16763=>"000000100",
  16764=>"110010000",
  16765=>"111111111",
  16766=>"000100101",
  16767=>"000011111",
  16768=>"000000001",
  16769=>"001101000",
  16770=>"100110110",
  16771=>"101101101",
  16772=>"111111111",
  16773=>"010000000",
  16774=>"000010110",
  16775=>"000010000",
  16776=>"110110111",
  16777=>"011011111",
  16778=>"101111111",
  16779=>"110111111",
  16780=>"111111101",
  16781=>"110100110",
  16782=>"001001000",
  16783=>"000000100",
  16784=>"011011011",
  16785=>"011011001",
  16786=>"000010110",
  16787=>"110110100",
  16788=>"111100000",
  16789=>"011111101",
  16790=>"011011110",
  16791=>"111011011",
  16792=>"000100000",
  16793=>"101101001",
  16794=>"001000000",
  16795=>"010010010",
  16796=>"111111101",
  16797=>"110010111",
  16798=>"000000100",
  16799=>"111001001",
  16800=>"001000000",
  16801=>"111100000",
  16802=>"001001010",
  16803=>"100000010",
  16804=>"111101100",
  16805=>"110110111",
  16806=>"000001011",
  16807=>"100100111",
  16808=>"101000001",
  16809=>"010111111",
  16810=>"111110110",
  16811=>"000110111",
  16812=>"000000100",
  16813=>"110110110",
  16814=>"110000000",
  16815=>"111101111",
  16816=>"001101001",
  16817=>"101000101",
  16818=>"000111111",
  16819=>"111111111",
  16820=>"000111111",
  16821=>"111110110",
  16822=>"001001101",
  16823=>"100101011",
  16824=>"101101101",
  16825=>"001101111",
  16826=>"111101101",
  16827=>"001011011",
  16828=>"001000110",
  16829=>"000000000",
  16830=>"000000000",
  16831=>"000001001",
  16832=>"101111011",
  16833=>"101101101",
  16834=>"111111111",
  16835=>"111111111",
  16836=>"001000011",
  16837=>"011001111",
  16838=>"101001011",
  16839=>"110110110",
  16840=>"001001101",
  16841=>"101100100",
  16842=>"010010010",
  16843=>"000000000",
  16844=>"111111110",
  16845=>"001001011",
  16846=>"001001001",
  16847=>"110110110",
  16848=>"001111111",
  16849=>"001101111",
  16850=>"001001101",
  16851=>"111111111",
  16852=>"111001001",
  16853=>"111000001",
  16854=>"101101000",
  16855=>"101101000",
  16856=>"101111000",
  16857=>"110000000",
  16858=>"111111111",
  16859=>"111101101",
  16860=>"011011111",
  16861=>"110110110",
  16862=>"111111111",
  16863=>"100100101",
  16864=>"000100100",
  16865=>"101111001",
  16866=>"111011000",
  16867=>"010010111",
  16868=>"111111111",
  16869=>"110110110",
  16870=>"010110110",
  16871=>"110110110",
  16872=>"101001001",
  16873=>"110110100",
  16874=>"010010011",
  16875=>"001001111",
  16876=>"110101111",
  16877=>"111001000",
  16878=>"001101101",
  16879=>"111101111",
  16880=>"101100101",
  16881=>"101111101",
  16882=>"101101101",
  16883=>"010000000",
  16884=>"001001111",
  16885=>"000000000",
  16886=>"100000010",
  16887=>"000000000",
  16888=>"011001000",
  16889=>"001001001",
  16890=>"110111111",
  16891=>"101001000",
  16892=>"101101111",
  16893=>"000000110",
  16894=>"000000011",
  16895=>"010011011",
  16896=>"111111110",
  16897=>"000000111",
  16898=>"100010111",
  16899=>"100000000",
  16900=>"001000000",
  16901=>"111111111",
  16902=>"000000001",
  16903=>"111111111",
  16904=>"111001000",
  16905=>"111111111",
  16906=>"000111111",
  16907=>"000111111",
  16908=>"011000000",
  16909=>"000000000",
  16910=>"011001000",
  16911=>"011000001",
  16912=>"100000000",
  16913=>"001011001",
  16914=>"111111000",
  16915=>"000110110",
  16916=>"111111111",
  16917=>"000100111",
  16918=>"101000000",
  16919=>"011011010",
  16920=>"100000000",
  16921=>"000001111",
  16922=>"001000000",
  16923=>"000110100",
  16924=>"111111111",
  16925=>"111011111",
  16926=>"001111000",
  16927=>"001111111",
  16928=>"001001000",
  16929=>"110110000",
  16930=>"100000001",
  16931=>"111100000",
  16932=>"000000100",
  16933=>"111110000",
  16934=>"000111111",
  16935=>"110000000",
  16936=>"001100100",
  16937=>"000000000",
  16938=>"111111000",
  16939=>"111000101",
  16940=>"111101000",
  16941=>"111000010",
  16942=>"001111111",
  16943=>"001000111",
  16944=>"000000000",
  16945=>"000000111",
  16946=>"100111011",
  16947=>"111001111",
  16948=>"111111000",
  16949=>"000000000",
  16950=>"000000000",
  16951=>"110111101",
  16952=>"000100111",
  16953=>"111000000",
  16954=>"111111111",
  16955=>"000000011",
  16956=>"001000000",
  16957=>"101000000",
  16958=>"111111001",
  16959=>"000000000",
  16960=>"111111110",
  16961=>"111000000",
  16962=>"111111111",
  16963=>"111111101",
  16964=>"100110010",
  16965=>"111100110",
  16966=>"000111100",
  16967=>"000001111",
  16968=>"011011001",
  16969=>"000111111",
  16970=>"110111111",
  16971=>"111111111",
  16972=>"000000111",
  16973=>"110110000",
  16974=>"000111111",
  16975=>"100111111",
  16976=>"111111001",
  16977=>"111111101",
  16978=>"000000111",
  16979=>"000000001",
  16980=>"111110110",
  16981=>"000110100",
  16982=>"110000000",
  16983=>"110000000",
  16984=>"011001001",
  16985=>"100100111",
  16986=>"000000100",
  16987=>"000001001",
  16988=>"000000000",
  16989=>"000000011",
  16990=>"111111111",
  16991=>"000100111",
  16992=>"000000111",
  16993=>"111111000",
  16994=>"000111111",
  16995=>"101111000",
  16996=>"101001111",
  16997=>"111011111",
  16998=>"000110111",
  16999=>"101111111",
  17000=>"101111111",
  17001=>"000000010",
  17002=>"110110111",
  17003=>"000110000",
  17004=>"110111110",
  17005=>"000000010",
  17006=>"111111111",
  17007=>"000111101",
  17008=>"000000001",
  17009=>"100111111",
  17010=>"000000000",
  17011=>"000000110",
  17012=>"110000000",
  17013=>"000100111",
  17014=>"000000110",
  17015=>"000111111",
  17016=>"111001000",
  17017=>"111101000",
  17018=>"001111100",
  17019=>"000111111",
  17020=>"110111000",
  17021=>"000000000",
  17022=>"000111111",
  17023=>"000000010",
  17024=>"101111111",
  17025=>"000001111",
  17026=>"000001111",
  17027=>"111000000",
  17028=>"001000001",
  17029=>"000000000",
  17030=>"100100000",
  17031=>"000000010",
  17032=>"000000010",
  17033=>"000000000",
  17034=>"111111111",
  17035=>"110111011",
  17036=>"000000000",
  17037=>"111111000",
  17038=>"111111111",
  17039=>"000000000",
  17040=>"000000000",
  17041=>"111000000",
  17042=>"000000110",
  17043=>"111111000",
  17044=>"100111111",
  17045=>"001110100",
  17046=>"111111111",
  17047=>"111111111",
  17048=>"101001001",
  17049=>"100000000",
  17050=>"101000001",
  17051=>"100000000",
  17052=>"111111101",
  17053=>"000111111",
  17054=>"111111100",
  17055=>"111111000",
  17056=>"000100110",
  17057=>"100111111",
  17058=>"111111111",
  17059=>"000101000",
  17060=>"011111000",
  17061=>"000000001",
  17062=>"111000000",
  17063=>"011001000",
  17064=>"100000011",
  17065=>"001001111",
  17066=>"111111110",
  17067=>"111111111",
  17068=>"111100000",
  17069=>"000001011",
  17070=>"000000000",
  17071=>"001000100",
  17072=>"000000000",
  17073=>"000100000",
  17074=>"110010110",
  17075=>"111000111",
  17076=>"000000001",
  17077=>"000000000",
  17078=>"000000011",
  17079=>"111111111",
  17080=>"011111111",
  17081=>"111111111",
  17082=>"000000100",
  17083=>"000000001",
  17084=>"111110000",
  17085=>"011111111",
  17086=>"100000111",
  17087=>"111111111",
  17088=>"111111111",
  17089=>"111100111",
  17090=>"111110000",
  17091=>"000111111",
  17092=>"001111111",
  17093=>"111001000",
  17094=>"111100000",
  17095=>"101001001",
  17096=>"000000101",
  17097=>"111000000",
  17098=>"000000000",
  17099=>"001111111",
  17100=>"111001000",
  17101=>"000111111",
  17102=>"111111110",
  17103=>"111111011",
  17104=>"000011011",
  17105=>"000000001",
  17106=>"010000000",
  17107=>"111101101",
  17108=>"111111000",
  17109=>"110110110",
  17110=>"000000000",
  17111=>"100101111",
  17112=>"000000000",
  17113=>"111111101",
  17114=>"000110000",
  17115=>"001100111",
  17116=>"110010000",
  17117=>"000000000",
  17118=>"111111111",
  17119=>"111111001",
  17120=>"111111111",
  17121=>"000000100",
  17122=>"000111110",
  17123=>"000000000",
  17124=>"000000000",
  17125=>"001101111",
  17126=>"111101000",
  17127=>"000000000",
  17128=>"000000000",
  17129=>"101111111",
  17130=>"110000101",
  17131=>"011111100",
  17132=>"011111111",
  17133=>"000000101",
  17134=>"100100000",
  17135=>"000111111",
  17136=>"101111111",
  17137=>"111111011",
  17138=>"111000000",
  17139=>"000000001",
  17140=>"111111111",
  17141=>"000000000",
  17142=>"001011011",
  17143=>"001100110",
  17144=>"111111000",
  17145=>"111111000",
  17146=>"111000111",
  17147=>"000000000",
  17148=>"110000000",
  17149=>"110110111",
  17150=>"111111111",
  17151=>"000000100",
  17152=>"111111101",
  17153=>"110110000",
  17154=>"101100000",
  17155=>"101111111",
  17156=>"000100111",
  17157=>"000111111",
  17158=>"111111111",
  17159=>"110000000",
  17160=>"001011011",
  17161=>"000000000",
  17162=>"111111111",
  17163=>"111000101",
  17164=>"111111000",
  17165=>"111110111",
  17166=>"110001111",
  17167=>"111000000",
  17168=>"000000111",
  17169=>"000011100",
  17170=>"111111111",
  17171=>"000100111",
  17172=>"111111111",
  17173=>"000000101",
  17174=>"000000000",
  17175=>"111111110",
  17176=>"110111111",
  17177=>"011111001",
  17178=>"001000100",
  17179=>"011111110",
  17180=>"001011011",
  17181=>"111101111",
  17182=>"000101100",
  17183=>"000010100",
  17184=>"111011011",
  17185=>"000000001",
  17186=>"000101111",
  17187=>"000100111",
  17188=>"111111011",
  17189=>"001111111",
  17190=>"001000011",
  17191=>"111111110",
  17192=>"000100000",
  17193=>"110110000",
  17194=>"011000000",
  17195=>"000001111",
  17196=>"010111001",
  17197=>"110100000",
  17198=>"000111000",
  17199=>"000000001",
  17200=>"000111111",
  17201=>"000000000",
  17202=>"111111111",
  17203=>"000111111",
  17204=>"000010111",
  17205=>"100111111",
  17206=>"000000000",
  17207=>"111111100",
  17208=>"000000111",
  17209=>"000000000",
  17210=>"111100101",
  17211=>"111101111",
  17212=>"110000000",
  17213=>"000000000",
  17214=>"001111000",
  17215=>"111111100",
  17216=>"101101100",
  17217=>"111111001",
  17218=>"000000000",
  17219=>"111111100",
  17220=>"000000110",
  17221=>"111101100",
  17222=>"000000111",
  17223=>"000000000",
  17224=>"111000000",
  17225=>"000000000",
  17226=>"111111111",
  17227=>"111111000",
  17228=>"111110001",
  17229=>"101111111",
  17230=>"010110000",
  17231=>"011011111",
  17232=>"111101111",
  17233=>"000111111",
  17234=>"111111010",
  17235=>"000000000",
  17236=>"000000000",
  17237=>"001001111",
  17238=>"000000000",
  17239=>"011011000",
  17240=>"011111000",
  17241=>"000000111",
  17242=>"000000101",
  17243=>"111000000",
  17244=>"111000000",
  17245=>"111010010",
  17246=>"000000111",
  17247=>"000000000",
  17248=>"101000000",
  17249=>"111010111",
  17250=>"111111010",
  17251=>"111111000",
  17252=>"110000000",
  17253=>"111000000",
  17254=>"001000111",
  17255=>"111001111",
  17256=>"111011000",
  17257=>"000111110",
  17258=>"110110000",
  17259=>"111111110",
  17260=>"111111111",
  17261=>"000001111",
  17262=>"101000111",
  17263=>"111011000",
  17264=>"100100111",
  17265=>"000000000",
  17266=>"000000000",
  17267=>"000000100",
  17268=>"000000000",
  17269=>"011111111",
  17270=>"000111111",
  17271=>"000111111",
  17272=>"011111011",
  17273=>"101111111",
  17274=>"000000000",
  17275=>"001111111",
  17276=>"000001000",
  17277=>"110100001",
  17278=>"000000000",
  17279=>"111001000",
  17280=>"000000000",
  17281=>"000000010",
  17282=>"001011011",
  17283=>"000000000",
  17284=>"000000000",
  17285=>"010010110",
  17286=>"000000100",
  17287=>"000000011",
  17288=>"000000100",
  17289=>"111111001",
  17290=>"001111111",
  17291=>"111111111",
  17292=>"111000111",
  17293=>"110100000",
  17294=>"111000011",
  17295=>"111111101",
  17296=>"000000111",
  17297=>"111111011",
  17298=>"111111111",
  17299=>"011001000",
  17300=>"000000000",
  17301=>"111000000",
  17302=>"000000111",
  17303=>"000000010",
  17304=>"001111111",
  17305=>"000000000",
  17306=>"111111000",
  17307=>"100101111",
  17308=>"111111110",
  17309=>"110000000",
  17310=>"111000100",
  17311=>"101101001",
  17312=>"000000000",
  17313=>"101111001",
  17314=>"111100000",
  17315=>"000100111",
  17316=>"111111000",
  17317=>"101001011",
  17318=>"000000000",
  17319=>"010111111",
  17320=>"111000000",
  17321=>"100000000",
  17322=>"111111000",
  17323=>"111000000",
  17324=>"000000111",
  17325=>"000000000",
  17326=>"111001001",
  17327=>"000000000",
  17328=>"110000000",
  17329=>"101111000",
  17330=>"000110100",
  17331=>"000000111",
  17332=>"100000000",
  17333=>"101001000",
  17334=>"111111111",
  17335=>"000010111",
  17336=>"111111111",
  17337=>"101001011",
  17338=>"111111111",
  17339=>"000000000",
  17340=>"000000111",
  17341=>"001000000",
  17342=>"101001010",
  17343=>"000011011",
  17344=>"010001101",
  17345=>"111000001",
  17346=>"110000000",
  17347=>"000001011",
  17348=>"101000001",
  17349=>"011001000",
  17350=>"110000111",
  17351=>"111001000",
  17352=>"111000000",
  17353=>"000000001",
  17354=>"011000000",
  17355=>"000111111",
  17356=>"000000100",
  17357=>"011000000",
  17358=>"001000000",
  17359=>"000000101",
  17360=>"111111111",
  17361=>"111111100",
  17362=>"110100000",
  17363=>"111000000",
  17364=>"000000000",
  17365=>"111111110",
  17366=>"011111000",
  17367=>"111101111",
  17368=>"101001111",
  17369=>"110110000",
  17370=>"011101000",
  17371=>"001000011",
  17372=>"111111110",
  17373=>"110000000",
  17374=>"001111111",
  17375=>"110100001",
  17376=>"000111000",
  17377=>"000000000",
  17378=>"100111111",
  17379=>"111101101",
  17380=>"000000100",
  17381=>"111000000",
  17382=>"110111111",
  17383=>"110000111",
  17384=>"000000111",
  17385=>"000111111",
  17386=>"011111111",
  17387=>"110110000",
  17388=>"101000000",
  17389=>"001000010",
  17390=>"000000000",
  17391=>"111111100",
  17392=>"011000000",
  17393=>"110100111",
  17394=>"000000011",
  17395=>"000000000",
  17396=>"111111001",
  17397=>"000000000",
  17398=>"111111000",
  17399=>"110111110",
  17400=>"000011111",
  17401=>"001000100",
  17402=>"100000111",
  17403=>"000111010",
  17404=>"110000000",
  17405=>"000000001",
  17406=>"000001000",
  17407=>"100000111",
  17408=>"111100111",
  17409=>"111111001",
  17410=>"111000000",
  17411=>"000100111",
  17412=>"111011000",
  17413=>"000000001",
  17414=>"111111100",
  17415=>"111111111",
  17416=>"111111111",
  17417=>"111110100",
  17418=>"000010011",
  17419=>"111011001",
  17420=>"110011111",
  17421=>"100101100",
  17422=>"000001001",
  17423=>"111111111",
  17424=>"001000001",
  17425=>"111111011",
  17426=>"110110000",
  17427=>"100100111",
  17428=>"000000000",
  17429=>"101000000",
  17430=>"011001100",
  17431=>"001011110",
  17432=>"001000000",
  17433=>"111111000",
  17434=>"111000000",
  17435=>"011100101",
  17436=>"000110111",
  17437=>"001000000",
  17438=>"010100110",
  17439=>"000111111",
  17440=>"000100100",
  17441=>"111111111",
  17442=>"100110110",
  17443=>"111011000",
  17444=>"000100110",
  17445=>"000000111",
  17446=>"011000100",
  17447=>"000100110",
  17448=>"000000000",
  17449=>"111100000",
  17450=>"111111111",
  17451=>"000000100",
  17452=>"011111111",
  17453=>"110000000",
  17454=>"011000000",
  17455=>"000000110",
  17456=>"000001011",
  17457=>"001000000",
  17458=>"000101111",
  17459=>"000000011",
  17460=>"000000000",
  17461=>"111111001",
  17462=>"000011000",
  17463=>"111111100",
  17464=>"101111111",
  17465=>"110111111",
  17466=>"000000000",
  17467=>"000000000",
  17468=>"111000000",
  17469=>"000000110",
  17470=>"111111111",
  17471=>"000000100",
  17472=>"000000111",
  17473=>"111001111",
  17474=>"000000111",
  17475=>"000001111",
  17476=>"000000011",
  17477=>"000001110",
  17478=>"111111010",
  17479=>"111111111",
  17480=>"001001000",
  17481=>"000001000",
  17482=>"111001001",
  17483=>"010001001",
  17484=>"000110000",
  17485=>"111000011",
  17486=>"000000000",
  17487=>"111111111",
  17488=>"000111111",
  17489=>"110111100",
  17490=>"000000001",
  17491=>"011011011",
  17492=>"111000000",
  17493=>"000011001",
  17494=>"010000000",
  17495=>"111011000",
  17496=>"000000000",
  17497=>"000000000",
  17498=>"000010111",
  17499=>"011011000",
  17500=>"101101100",
  17501=>"111111111",
  17502=>"111011010",
  17503=>"011001011",
  17504=>"000000000",
  17505=>"010111011",
  17506=>"111111111",
  17507=>"111111000",
  17508=>"001101001",
  17509=>"100100000",
  17510=>"000101111",
  17511=>"111011011",
  17512=>"011011000",
  17513=>"000101000",
  17514=>"000000000",
  17515=>"111111111",
  17516=>"010110111",
  17517=>"111111111",
  17518=>"011111110",
  17519=>"111000000",
  17520=>"000011111",
  17521=>"101101011",
  17522=>"110111100",
  17523=>"000010011",
  17524=>"111110100",
  17525=>"111111111",
  17526=>"000000000",
  17527=>"000000000",
  17528=>"111111001",
  17529=>"000000000",
  17530=>"111011001",
  17531=>"111110000",
  17532=>"100001001",
  17533=>"111001000",
  17534=>"111111111",
  17535=>"111110011",
  17536=>"111000000",
  17537=>"111111011",
  17538=>"001000111",
  17539=>"111111000",
  17540=>"111111111",
  17541=>"110000000",
  17542=>"111101111",
  17543=>"000000101",
  17544=>"000000000",
  17545=>"000000000",
  17546=>"100100111",
  17547=>"000010000",
  17548=>"001101111",
  17549=>"000110000",
  17550=>"100100000",
  17551=>"000000111",
  17552=>"000000111",
  17553=>"001000111",
  17554=>"100111111",
  17555=>"000000100",
  17556=>"100000000",
  17557=>"001111101",
  17558=>"001101111",
  17559=>"111000000",
  17560=>"111011011",
  17561=>"000000010",
  17562=>"111001000",
  17563=>"010010010",
  17564=>"000011110",
  17565=>"011001011",
  17566=>"100111111",
  17567=>"100000000",
  17568=>"001000000",
  17569=>"000000111",
  17570=>"000111000",
  17571=>"111110110",
  17572=>"101011001",
  17573=>"111011101",
  17574=>"111111110",
  17575=>"000111110",
  17576=>"111100000",
  17577=>"000000011",
  17578=>"000000000",
  17579=>"110111111",
  17580=>"111111111",
  17581=>"111111101",
  17582=>"000000000",
  17583=>"000000111",
  17584=>"000000001",
  17585=>"111011010",
  17586=>"100110100",
  17587=>"111111111",
  17588=>"111001001",
  17589=>"111111111",
  17590=>"000100111",
  17591=>"100111000",
  17592=>"111111000",
  17593=>"011000000",
  17594=>"111111000",
  17595=>"111111111",
  17596=>"000111011",
  17597=>"100000000",
  17598=>"000000111",
  17599=>"001111111",
  17600=>"111111011",
  17601=>"110111011",
  17602=>"010111111",
  17603=>"000111111",
  17604=>"110000000",
  17605=>"000111111",
  17606=>"000000000",
  17607=>"001000000",
  17608=>"011000000",
  17609=>"111111011",
  17610=>"000000010",
  17611=>"111011000",
  17612=>"000111111",
  17613=>"000110000",
  17614=>"000000111",
  17615=>"000000000",
  17616=>"111111111",
  17617=>"011001000",
  17618=>"000000100",
  17619=>"111111001",
  17620=>"101000000",
  17621=>"110111101",
  17622=>"111011011",
  17623=>"011010010",
  17624=>"000001000",
  17625=>"001000000",
  17626=>"011000000",
  17627=>"000000000",
  17628=>"001000100",
  17629=>"111111111",
  17630=>"110111111",
  17631=>"110000000",
  17632=>"100101111",
  17633=>"111111001",
  17634=>"000111111",
  17635=>"111000000",
  17636=>"010001000",
  17637=>"011000100",
  17638=>"111001111",
  17639=>"111111111",
  17640=>"101111111",
  17641=>"000101111",
  17642=>"101111100",
  17643=>"111111011",
  17644=>"110000000",
  17645=>"001111111",
  17646=>"000000101",
  17647=>"111101111",
  17648=>"001111101",
  17649=>"111001100",
  17650=>"000011111",
  17651=>"111101111",
  17652=>"111111111",
  17653=>"000100111",
  17654=>"000001001",
  17655=>"000000001",
  17656=>"111111111",
  17657=>"000100111",
  17658=>"000000100",
  17659=>"011000000",
  17660=>"111111011",
  17661=>"000110100",
  17662=>"010010000",
  17663=>"000000000",
  17664=>"111000000",
  17665=>"100100111",
  17666=>"111111101",
  17667=>"000000101",
  17668=>"000000000",
  17669=>"110000100",
  17670=>"001000001",
  17671=>"111111111",
  17672=>"111111000",
  17673=>"000000000",
  17674=>"111111110",
  17675=>"111111111",
  17676=>"110100100",
  17677=>"111111010",
  17678=>"000000100",
  17679=>"000111111",
  17680=>"100110111",
  17681=>"111111111",
  17682=>"000100000",
  17683=>"100000000",
  17684=>"000100101",
  17685=>"000000001",
  17686=>"001001101",
  17687=>"000000100",
  17688=>"000110000",
  17689=>"011011000",
  17690=>"001111100",
  17691=>"000100111",
  17692=>"011110100",
  17693=>"111111111",
  17694=>"100100111",
  17695=>"000001111",
  17696=>"110111101",
  17697=>"111111101",
  17698=>"100000000",
  17699=>"111011001",
  17700=>"111100111",
  17701=>"100100101",
  17702=>"111110110",
  17703=>"111111011",
  17704=>"111111000",
  17705=>"000000100",
  17706=>"001000111",
  17707=>"110110111",
  17708=>"111111000",
  17709=>"010110110",
  17710=>"111010111",
  17711=>"001000110",
  17712=>"111100100",
  17713=>"111111111",
  17714=>"111111001",
  17715=>"111111001",
  17716=>"001001000",
  17717=>"000010011",
  17718=>"000000100",
  17719=>"110011111",
  17720=>"001111000",
  17721=>"111101011",
  17722=>"001001000",
  17723=>"000000000",
  17724=>"110110111",
  17725=>"010000001",
  17726=>"001000100",
  17727=>"111101110",
  17728=>"111111000",
  17729=>"111001000",
  17730=>"000000111",
  17731=>"111000000",
  17732=>"000001111",
  17733=>"111111000",
  17734=>"001000001",
  17735=>"111001000",
  17736=>"000111111",
  17737=>"000111111",
  17738=>"100000001",
  17739=>"111000100",
  17740=>"001111111",
  17741=>"111011000",
  17742=>"111001001",
  17743=>"011111110",
  17744=>"000000000",
  17745=>"111111111",
  17746=>"100000000",
  17747=>"011000000",
  17748=>"100100000",
  17749=>"111111001",
  17750=>"111111111",
  17751=>"000111100",
  17752=>"111111000",
  17753=>"000011111",
  17754=>"111111000",
  17755=>"100100110",
  17756=>"111000000",
  17757=>"111111111",
  17758=>"000000111",
  17759=>"001111111",
  17760=>"000000111",
  17761=>"111111001",
  17762=>"111001001",
  17763=>"000000011",
  17764=>"000000010",
  17765=>"111111011",
  17766=>"000000111",
  17767=>"111000110",
  17768=>"001101111",
  17769=>"000001001",
  17770=>"000000000",
  17771=>"000000111",
  17772=>"111001000",
  17773=>"000001000",
  17774=>"000110111",
  17775=>"000100100",
  17776=>"111000000",
  17777=>"000000000",
  17778=>"111111110",
  17779=>"111111110",
  17780=>"011111111",
  17781=>"111000001",
  17782=>"000000001",
  17783=>"111111001",
  17784=>"111111101",
  17785=>"000000011",
  17786=>"111000000",
  17787=>"111000000",
  17788=>"000000011",
  17789=>"110110001",
  17790=>"111111111",
  17791=>"000000100",
  17792=>"110110110",
  17793=>"101001000",
  17794=>"011011001",
  17795=>"000000000",
  17796=>"111111000",
  17797=>"000000000",
  17798=>"000011111",
  17799=>"111100000",
  17800=>"011111100",
  17801=>"001000111",
  17802=>"111011000",
  17803=>"000011111",
  17804=>"111111111",
  17805=>"100110100",
  17806=>"011011010",
  17807=>"000000000",
  17808=>"111111110",
  17809=>"101000100",
  17810=>"110111111",
  17811=>"001001101",
  17812=>"000000111",
  17813=>"001000000",
  17814=>"111111111",
  17815=>"111111011",
  17816=>"000000111",
  17817=>"111011001",
  17818=>"111111110",
  17819=>"011100000",
  17820=>"001001100",
  17821=>"000000101",
  17822=>"000000000",
  17823=>"111110111",
  17824=>"011000000",
  17825=>"110111111",
  17826=>"000000000",
  17827=>"111000000",
  17828=>"100000000",
  17829=>"110111011",
  17830=>"111111100",
  17831=>"111111111",
  17832=>"000000010",
  17833=>"111111111",
  17834=>"000000100",
  17835=>"011000000",
  17836=>"000001111",
  17837=>"000001010",
  17838=>"000000000",
  17839=>"000000000",
  17840=>"011000000",
  17841=>"011111111",
  17842=>"101000000",
  17843=>"010011000",
  17844=>"000000011",
  17845=>"011111111",
  17846=>"011011000",
  17847=>"000000010",
  17848=>"011000100",
  17849=>"111100100",
  17850=>"111011000",
  17851=>"111001000",
  17852=>"000111111",
  17853=>"111111111",
  17854=>"000000000",
  17855=>"111100100",
  17856=>"111111100",
  17857=>"010011000",
  17858=>"000000000",
  17859=>"000111111",
  17860=>"010001111",
  17861=>"100110110",
  17862=>"000001000",
  17863=>"111011010",
  17864=>"111111111",
  17865=>"000000000",
  17866=>"110000000",
  17867=>"000000110",
  17868=>"000110001",
  17869=>"000000000",
  17870=>"000000100",
  17871=>"100111111",
  17872=>"000000000",
  17873=>"001011111",
  17874=>"000001111",
  17875=>"110011111",
  17876=>"111111111",
  17877=>"010011001",
  17878=>"011000000",
  17879=>"100000010",
  17880=>"000000000",
  17881=>"111110100",
  17882=>"101101111",
  17883=>"000111111",
  17884=>"100111111",
  17885=>"000111111",
  17886=>"000000111",
  17887=>"000111011",
  17888=>"111111110",
  17889=>"111111001",
  17890=>"000110110",
  17891=>"001001001",
  17892=>"011001000",
  17893=>"111101000",
  17894=>"000000000",
  17895=>"000001111",
  17896=>"111110000",
  17897=>"001111111",
  17898=>"111101000",
  17899=>"000000000",
  17900=>"111001000",
  17901=>"110110100",
  17902=>"111010000",
  17903=>"000000000",
  17904=>"001000000",
  17905=>"000111111",
  17906=>"111111000",
  17907=>"111000000",
  17908=>"000000010",
  17909=>"111111010",
  17910=>"000001111",
  17911=>"111111110",
  17912=>"000111111",
  17913=>"000000100",
  17914=>"111111111",
  17915=>"000111111",
  17916=>"010011000",
  17917=>"101001011",
  17918=>"000000000",
  17919=>"111011001",
  17920=>"110110110",
  17921=>"000010111",
  17922=>"111001000",
  17923=>"111100100",
  17924=>"001111000",
  17925=>"110000000",
  17926=>"000000000",
  17927=>"111111111",
  17928=>"101101111",
  17929=>"110000000",
  17930=>"000000000",
  17931=>"110001000",
  17932=>"000000000",
  17933=>"000001110",
  17934=>"111111010",
  17935=>"100000000",
  17936=>"100100100",
  17937=>"000000101",
  17938=>"000001111",
  17939=>"111110100",
  17940=>"000110000",
  17941=>"111111111",
  17942=>"000000000",
  17943=>"011000000",
  17944=>"000001001",
  17945=>"101000000",
  17946=>"100000000",
  17947=>"000111011",
  17948=>"001001000",
  17949=>"001111001",
  17950=>"001001001",
  17951=>"001101111",
  17952=>"111111000",
  17953=>"111001000",
  17954=>"001001111",
  17955=>"101111111",
  17956=>"111001111",
  17957=>"111111111",
  17958=>"000000000",
  17959=>"000000100",
  17960=>"010111111",
  17961=>"111000111",
  17962=>"001111111",
  17963=>"001001000",
  17964=>"111111111",
  17965=>"111111110",
  17966=>"001001011",
  17967=>"110111111",
  17968=>"111001011",
  17969=>"001000000",
  17970=>"001100100",
  17971=>"011010010",
  17972=>"000010000",
  17973=>"000000000",
  17974=>"001001011",
  17975=>"000111111",
  17976=>"000000011",
  17977=>"001000111",
  17978=>"000000000",
  17979=>"000000111",
  17980=>"111111111",
  17981=>"000000011",
  17982=>"000111111",
  17983=>"000001111",
  17984=>"001100100",
  17985=>"000111111",
  17986=>"000000000",
  17987=>"000110111",
  17988=>"011011011",
  17989=>"000000000",
  17990=>"000111111",
  17991=>"111111111",
  17992=>"000000000",
  17993=>"000111111",
  17994=>"111110010",
  17995=>"111001111",
  17996=>"111000000",
  17997=>"111111001",
  17998=>"010000000",
  17999=>"011000001",
  18000=>"000010000",
  18001=>"110111111",
  18002=>"000000000",
  18003=>"110111101",
  18004=>"000000000",
  18005=>"111110000",
  18006=>"000111111",
  18007=>"000000000",
  18008=>"001011010",
  18009=>"000000000",
  18010=>"110010000",
  18011=>"111111000",
  18012=>"011001000",
  18013=>"111111110",
  18014=>"000000111",
  18015=>"111001001",
  18016=>"000001000",
  18017=>"111000000",
  18018=>"000011010",
  18019=>"000111111",
  18020=>"000001000",
  18021=>"111111000",
  18022=>"111000111",
  18023=>"100100111",
  18024=>"101001000",
  18025=>"111111111",
  18026=>"110000010",
  18027=>"000000111",
  18028=>"100111111",
  18029=>"110010111",
  18030=>"100000111",
  18031=>"111111000",
  18032=>"000000111",
  18033=>"000000111",
  18034=>"111111111",
  18035=>"000000000",
  18036=>"000000000",
  18037=>"000000000",
  18038=>"001000111",
  18039=>"000000000",
  18040=>"111000000",
  18041=>"000000000",
  18042=>"000011111",
  18043=>"000000000",
  18044=>"110110110",
  18045=>"110000111",
  18046=>"001000000",
  18047=>"000000111",
  18048=>"000000000",
  18049=>"100010111",
  18050=>"110000000",
  18051=>"110111010",
  18052=>"111000000",
  18053=>"111111000",
  18054=>"110110110",
  18055=>"001001001",
  18056=>"000110010",
  18057=>"111111111",
  18058=>"000000000",
  18059=>"000000000",
  18060=>"000000000",
  18061=>"001000000",
  18062=>"111111001",
  18063=>"111111000",
  18064=>"111111000",
  18065=>"111111011",
  18066=>"000000001",
  18067=>"001011011",
  18068=>"111000111",
  18069=>"111111000",
  18070=>"000000010",
  18071=>"000000111",
  18072=>"000000100",
  18073=>"111111000",
  18074=>"111111111",
  18075=>"000001111",
  18076=>"000100110",
  18077=>"110110110",
  18078=>"011111001",
  18079=>"111111111",
  18080=>"111000111",
  18081=>"000111111",
  18082=>"111101101",
  18083=>"111000000",
  18084=>"001000010",
  18085=>"001000001",
  18086=>"000111111",
  18087=>"110000000",
  18088=>"011000001",
  18089=>"100001111",
  18090=>"111100101",
  18091=>"000000001",
  18092=>"101101101",
  18093=>"001001011",
  18094=>"000000000",
  18095=>"111111001",
  18096=>"111111111",
  18097=>"111001000",
  18098=>"111111111",
  18099=>"001000000",
  18100=>"111000000",
  18101=>"000000000",
  18102=>"111000000",
  18103=>"110000000",
  18104=>"111111111",
  18105=>"000000000",
  18106=>"000000000",
  18107=>"001101000",
  18108=>"000010110",
  18109=>"001001101",
  18110=>"111111000",
  18111=>"111111101",
  18112=>"111111111",
  18113=>"110111111",
  18114=>"001001101",
  18115=>"000000000",
  18116=>"000001000",
  18117=>"111111111",
  18118=>"111101101",
  18119=>"001111011",
  18120=>"000000000",
  18121=>"101111111",
  18122=>"101101110",
  18123=>"110110110",
  18124=>"000000111",
  18125=>"101001000",
  18126=>"000001001",
  18127=>"000001111",
  18128=>"000000000",
  18129=>"000111111",
  18130=>"100000000",
  18131=>"111100111",
  18132=>"101000000",
  18133=>"011011011",
  18134=>"000000111",
  18135=>"111000001",
  18136=>"001000101",
  18137=>"001111111",
  18138=>"000000000",
  18139=>"111111100",
  18140=>"111100000",
  18141=>"000000000",
  18142=>"101000101",
  18143=>"011000000",
  18144=>"101001001",
  18145=>"000000111",
  18146=>"111000000",
  18147=>"100111111",
  18148=>"010111000",
  18149=>"111110000",
  18150=>"000111111",
  18151=>"111111111",
  18152=>"111111111",
  18153=>"111110000",
  18154=>"001000110",
  18155=>"101001111",
  18156=>"111111111",
  18157=>"111111100",
  18158=>"111000000",
  18159=>"000110111",
  18160=>"100000000",
  18161=>"010111111",
  18162=>"111100110",
  18163=>"000000000",
  18164=>"000000000",
  18165=>"111111101",
  18166=>"101000000",
  18167=>"111111111",
  18168=>"000011011",
  18169=>"111000000",
  18170=>"001001000",
  18171=>"000001000",
  18172=>"000100110",
  18173=>"000111111",
  18174=>"000000000",
  18175=>"000100111",
  18176=>"000000001",
  18177=>"111001001",
  18178=>"000000111",
  18179=>"100101111",
  18180=>"111101111",
  18181=>"000000000",
  18182=>"101111111",
  18183=>"000000111",
  18184=>"000000101",
  18185=>"000000000",
  18186=>"110000100",
  18187=>"000100111",
  18188=>"111111111",
  18189=>"000001001",
  18190=>"000000000",
  18191=>"000110111",
  18192=>"111000000",
  18193=>"000001111",
  18194=>"000000000",
  18195=>"100111000",
  18196=>"101010011",
  18197=>"111100111",
  18198=>"011011000",
  18199=>"000111111",
  18200=>"111001001",
  18201=>"100111111",
  18202=>"010011011",
  18203=>"111111100",
  18204=>"111111011",
  18205=>"000000110",
  18206=>"111111111",
  18207=>"000101111",
  18208=>"000000111",
  18209=>"000111111",
  18210=>"110111111",
  18211=>"110000111",
  18212=>"110010010",
  18213=>"111111111",
  18214=>"100000000",
  18215=>"110000101",
  18216=>"111111111",
  18217=>"011011111",
  18218=>"000000000",
  18219=>"111111000",
  18220=>"000100100",
  18221=>"111000001",
  18222=>"111000111",
  18223=>"100000100",
  18224=>"111110110",
  18225=>"000000000",
  18226=>"111011111",
  18227=>"111111110",
  18228=>"000000000",
  18229=>"011111111",
  18230=>"110101111",
  18231=>"111101001",
  18232=>"111000000",
  18233=>"110111100",
  18234=>"000000000",
  18235=>"011100100",
  18236=>"011011011",
  18237=>"000111111",
  18238=>"011011111",
  18239=>"011000000",
  18240=>"000000110",
  18241=>"100110000",
  18242=>"000000101",
  18243=>"000111011",
  18244=>"001101111",
  18245=>"111111111",
  18246=>"000000000",
  18247=>"100110000",
  18248=>"111000000",
  18249=>"000000110",
  18250=>"001001000",
  18251=>"011111111",
  18252=>"111111000",
  18253=>"001000001",
  18254=>"000000110",
  18255=>"111101111",
  18256=>"011111111",
  18257=>"000000000",
  18258=>"111111111",
  18259=>"111111111",
  18260=>"111111111",
  18261=>"011011011",
  18262=>"000000100",
  18263=>"000101111",
  18264=>"101001111",
  18265=>"111111010",
  18266=>"000000000",
  18267=>"111000000",
  18268=>"111100111",
  18269=>"011011000",
  18270=>"000100000",
  18271=>"110001111",
  18272=>"000000101",
  18273=>"000100011",
  18274=>"100000000",
  18275=>"111111100",
  18276=>"111111111",
  18277=>"000101111",
  18278=>"000000000",
  18279=>"000000111",
  18280=>"110111111",
  18281=>"111111111",
  18282=>"001111011",
  18283=>"011000000",
  18284=>"000000000",
  18285=>"000000000",
  18286=>"110010000",
  18287=>"011001000",
  18288=>"001000000",
  18289=>"001000000",
  18290=>"110100000",
  18291=>"100000100",
  18292=>"111000111",
  18293=>"011111110",
  18294=>"111111111",
  18295=>"000111111",
  18296=>"111000000",
  18297=>"000000111",
  18298=>"000000000",
  18299=>"111011111",
  18300=>"101100100",
  18301=>"000010110",
  18302=>"111000000",
  18303=>"111111111",
  18304=>"111111111",
  18305=>"010010000",
  18306=>"001001001",
  18307=>"111100100",
  18308=>"111000000",
  18309=>"000111111",
  18310=>"000001000",
  18311=>"110010010",
  18312=>"000000000",
  18313=>"010110111",
  18314=>"000000000",
  18315=>"111111111",
  18316=>"101100000",
  18317=>"000001111",
  18318=>"111111100",
  18319=>"110100000",
  18320=>"000111111",
  18321=>"000000000",
  18322=>"000001000",
  18323=>"001110110",
  18324=>"111111111",
  18325=>"000010010",
  18326=>"111111000",
  18327=>"011011001",
  18328=>"000101000",
  18329=>"001001000",
  18330=>"000000001",
  18331=>"001000000",
  18332=>"000111111",
  18333=>"000111000",
  18334=>"000111000",
  18335=>"000111000",
  18336=>"111111111",
  18337=>"111001111",
  18338=>"100000000",
  18339=>"110000000",
  18340=>"011111110",
  18341=>"111111000",
  18342=>"011011111",
  18343=>"001001111",
  18344=>"111111111",
  18345=>"000111111",
  18346=>"000000111",
  18347=>"000000000",
  18348=>"000000000",
  18349=>"100001000",
  18350=>"011101111",
  18351=>"111111101",
  18352=>"000000101",
  18353=>"000000011",
  18354=>"111111110",
  18355=>"111000000",
  18356=>"111111111",
  18357=>"111111111",
  18358=>"111111111",
  18359=>"000111111",
  18360=>"000000000",
  18361=>"111110000",
  18362=>"000000111",
  18363=>"000111101",
  18364=>"111111111",
  18365=>"110100000",
  18366=>"000000000",
  18367=>"111111111",
  18368=>"010111111",
  18369=>"000000011",
  18370=>"111000000",
  18371=>"001000000",
  18372=>"000000001",
  18373=>"000000100",
  18374=>"111101000",
  18375=>"001001101",
  18376=>"000000000",
  18377=>"111111111",
  18378=>"001111110",
  18379=>"000110111",
  18380=>"000000000",
  18381=>"111101001",
  18382=>"101111111",
  18383=>"111001000",
  18384=>"010010000",
  18385=>"100111111",
  18386=>"100111111",
  18387=>"111001111",
  18388=>"111111000",
  18389=>"110000000",
  18390=>"000000000",
  18391=>"000000100",
  18392=>"111111111",
  18393=>"110000100",
  18394=>"111000000",
  18395=>"111111111",
  18396=>"100111111",
  18397=>"111111111",
  18398=>"111011111",
  18399=>"101001000",
  18400=>"000000000",
  18401=>"111000000",
  18402=>"000100111",
  18403=>"101111100",
  18404=>"000000000",
  18405=>"100111000",
  18406=>"111000000",
  18407=>"010000000",
  18408=>"000000000",
  18409=>"111101111",
  18410=>"110000111",
  18411=>"010110111",
  18412=>"000110101",
  18413=>"100100100",
  18414=>"000000110",
  18415=>"000000001",
  18416=>"100000000",
  18417=>"111111111",
  18418=>"100101101",
  18419=>"000111111",
  18420=>"110111111",
  18421=>"000000000",
  18422=>"000000111",
  18423=>"111100000",
  18424=>"111111111",
  18425=>"111000111",
  18426=>"000000000",
  18427=>"110010000",
  18428=>"000000000",
  18429=>"101111111",
  18430=>"000000100",
  18431=>"111111111",
  18432=>"010000000",
  18433=>"000010000",
  18434=>"001000101",
  18435=>"111111111",
  18436=>"000100111",
  18437=>"111000011",
  18438=>"010110010",
  18439=>"111101111",
  18440=>"111010000",
  18441=>"000000000",
  18442=>"001000111",
  18443=>"011011011",
  18444=>"110111111",
  18445=>"110000000",
  18446=>"100000000",
  18447=>"001001101",
  18448=>"000001000",
  18449=>"000011011",
  18450=>"000000000",
  18451=>"111000000",
  18452=>"000110110",
  18453=>"000000001",
  18454=>"110111111",
  18455=>"000000100",
  18456=>"000000000",
  18457=>"111111000",
  18458=>"111111000",
  18459=>"100100000",
  18460=>"111111001",
  18461=>"000000010",
  18462=>"101001000",
  18463=>"000000000",
  18464=>"011011011",
  18465=>"001001001",
  18466=>"110111110",
  18467=>"000000111",
  18468=>"011000111",
  18469=>"111111111",
  18470=>"000000000",
  18471=>"011101011",
  18472=>"110100101",
  18473=>"000000000",
  18474=>"000000101",
  18475=>"111010010",
  18476=>"111111111",
  18477=>"111111111",
  18478=>"101100010",
  18479=>"000001111",
  18480=>"001111111",
  18481=>"011001111",
  18482=>"111111110",
  18483=>"001100000",
  18484=>"111111111",
  18485=>"111111100",
  18486=>"000000000",
  18487=>"000000000",
  18488=>"000000000",
  18489=>"010000000",
  18490=>"010111111",
  18491=>"101000000",
  18492=>"000000100",
  18493=>"110111111",
  18494=>"110110110",
  18495=>"111001000",
  18496=>"111101111",
  18497=>"111001000",
  18498=>"101001101",
  18499=>"000000111",
  18500=>"100000001",
  18501=>"000000111",
  18502=>"000000111",
  18503=>"101101111",
  18504=>"111111011",
  18505=>"000001111",
  18506=>"111111100",
  18507=>"000000000",
  18508=>"001000000",
  18509=>"111111000",
  18510=>"111011111",
  18511=>"000111111",
  18512=>"011111010",
  18513=>"111001010",
  18514=>"000000111",
  18515=>"111000000",
  18516=>"001001000",
  18517=>"111110000",
  18518=>"000000000",
  18519=>"100101000",
  18520=>"000000000",
  18521=>"111100101",
  18522=>"111111110",
  18523=>"111111111",
  18524=>"111111111",
  18525=>"001001001",
  18526=>"110110011",
  18527=>"111110100",
  18528=>"000111111",
  18529=>"000010010",
  18530=>"111011010",
  18531=>"100000111",
  18532=>"111110010",
  18533=>"001001001",
  18534=>"111111011",
  18535=>"100000000",
  18536=>"000011111",
  18537=>"111101111",
  18538=>"010110000",
  18539=>"111111111",
  18540=>"111111111",
  18541=>"010010010",
  18542=>"101001001",
  18543=>"000000111",
  18544=>"000000000",
  18545=>"000000000",
  18546=>"001000000",
  18547=>"111110111",
  18548=>"110110010",
  18549=>"111111111",
  18550=>"010010111",
  18551=>"011111111",
  18552=>"000000000",
  18553=>"111111111",
  18554=>"101101100",
  18555=>"000001001",
  18556=>"111000000",
  18557=>"000001000",
  18558=>"001000000",
  18559=>"111111111",
  18560=>"111111111",
  18561=>"000000000",
  18562=>"011011000",
  18563=>"111111011",
  18564=>"111111111",
  18565=>"000000000",
  18566=>"001101011",
  18567=>"100000011",
  18568=>"000000011",
  18569=>"000001111",
  18570=>"000000010",
  18571=>"111010010",
  18572=>"100000010",
  18573=>"000000000",
  18574=>"000100000",
  18575=>"111111111",
  18576=>"101000001",
  18577=>"000000000",
  18578=>"111111000",
  18579=>"111111111",
  18580=>"111111010",
  18581=>"000100111",
  18582=>"111111111",
  18583=>"000000000",
  18584=>"100000000",
  18585=>"000000001",
  18586=>"000000000",
  18587=>"111001000",
  18588=>"110000010",
  18589=>"111111111",
  18590=>"000001101",
  18591=>"000010000",
  18592=>"111100000",
  18593=>"011000000",
  18594=>"011110110",
  18595=>"111111111",
  18596=>"001001001",
  18597=>"110110000",
  18598=>"100000000",
  18599=>"111111000",
  18600=>"101100100",
  18601=>"000000000",
  18602=>"100000000",
  18603=>"111111111",
  18604=>"100111111",
  18605=>"100100000",
  18606=>"110110110",
  18607=>"000111111",
  18608=>"111111111",
  18609=>"111011001",
  18610=>"000111010",
  18611=>"000100101",
  18612=>"001001100",
  18613=>"011011010",
  18614=>"001001001",
  18615=>"000000000",
  18616=>"000000000",
  18617=>"111111111",
  18618=>"000101101",
  18619=>"111111000",
  18620=>"000000000",
  18621=>"000000000",
  18622=>"110100111",
  18623=>"111001101",
  18624=>"000000000",
  18625=>"000000000",
  18626=>"000000000",
  18627=>"000001000",
  18628=>"000000001",
  18629=>"000000001",
  18630=>"001000100",
  18631=>"000010100",
  18632=>"000000000",
  18633=>"000000000",
  18634=>"000100100",
  18635=>"111111000",
  18636=>"001000000",
  18637=>"000000000",
  18638=>"000011111",
  18639=>"111111000",
  18640=>"110000000",
  18641=>"001000101",
  18642=>"000000111",
  18643=>"111111110",
  18644=>"010010010",
  18645=>"110111111",
  18646=>"000000000",
  18647=>"111111111",
  18648=>"111111111",
  18649=>"111111110",
  18650=>"111110110",
  18651=>"000001000",
  18652=>"001000000",
  18653=>"000000000",
  18654=>"100000000",
  18655=>"110110000",
  18656=>"001000001",
  18657=>"000000000",
  18658=>"000000000",
  18659=>"110111010",
  18660=>"000001001",
  18661=>"000000000",
  18662=>"011110000",
  18663=>"000000000",
  18664=>"111111010",
  18665=>"111100000",
  18666=>"101111001",
  18667=>"111111101",
  18668=>"100101001",
  18669=>"111000000",
  18670=>"100100111",
  18671=>"100000101",
  18672=>"111001001",
  18673=>"000000101",
  18674=>"100100111",
  18675=>"001000000",
  18676=>"111111111",
  18677=>"111101100",
  18678=>"000000000",
  18679=>"111111111",
  18680=>"111111111",
  18681=>"000010010",
  18682=>"000000000",
  18683=>"001001111",
  18684=>"110110111",
  18685=>"110110000",
  18686=>"100110000",
  18687=>"111111000",
  18688=>"110110010",
  18689=>"101111001",
  18690=>"111111011",
  18691=>"000000000",
  18692=>"000000000",
  18693=>"000000111",
  18694=>"111111111",
  18695=>"000000000",
  18696=>"000000000",
  18697=>"000000000",
  18698=>"000000000",
  18699=>"111111010",
  18700=>"101000000",
  18701=>"111111111",
  18702=>"000001101",
  18703=>"111111001",
  18704=>"000000111",
  18705=>"100100111",
  18706=>"000000000",
  18707=>"001011011",
  18708=>"000000111",
  18709=>"000111111",
  18710=>"000111110",
  18711=>"111111011",
  18712=>"111111110",
  18713=>"111111100",
  18714=>"000000000",
  18715=>"110010010",
  18716=>"111111111",
  18717=>"000000010",
  18718=>"000000000",
  18719=>"000111111",
  18720=>"100000000",
  18721=>"000000000",
  18722=>"111110000",
  18723=>"111111110",
  18724=>"000000000",
  18725=>"111111111",
  18726=>"000000001",
  18727=>"111000000",
  18728=>"110110111",
  18729=>"001000011",
  18730=>"110111010",
  18731=>"111000000",
  18732=>"110111111",
  18733=>"000000011",
  18734=>"000000111",
  18735=>"000000000",
  18736=>"011011010",
  18737=>"000110101",
  18738=>"110111111",
  18739=>"000000000",
  18740=>"010000010",
  18741=>"111101000",
  18742=>"000111100",
  18743=>"111111111",
  18744=>"111111000",
  18745=>"111101000",
  18746=>"100100101",
  18747=>"000000000",
  18748=>"111011001",
  18749=>"000000000",
  18750=>"000001001",
  18751=>"110111111",
  18752=>"011000000",
  18753=>"001001100",
  18754=>"100000110",
  18755=>"111111111",
  18756=>"000000001",
  18757=>"000000000",
  18758=>"011111110",
  18759=>"111001011",
  18760=>"111000000",
  18761=>"111111111",
  18762=>"111111111",
  18763=>"100100100",
  18764=>"001001001",
  18765=>"111110000",
  18766=>"100100001",
  18767=>"010110110",
  18768=>"110000000",
  18769=>"110111111",
  18770=>"001111101",
  18771=>"000000000",
  18772=>"000111111",
  18773=>"001001001",
  18774=>"000010000",
  18775=>"100100110",
  18776=>"110000111",
  18777=>"001011111",
  18778=>"001000100",
  18779=>"111111111",
  18780=>"110000000",
  18781=>"111111111",
  18782=>"011111101",
  18783=>"000000000",
  18784=>"000000000",
  18785=>"100000000",
  18786=>"100100100",
  18787=>"111111001",
  18788=>"100110110",
  18789=>"000000000",
  18790=>"000000000",
  18791=>"000000010",
  18792=>"000000001",
  18793=>"001111111",
  18794=>"111100101",
  18795=>"111111010",
  18796=>"010110110",
  18797=>"000101111",
  18798=>"111111110",
  18799=>"001011001",
  18800=>"000000000",
  18801=>"111111111",
  18802=>"111110110",
  18803=>"111111011",
  18804=>"000000000",
  18805=>"001111010",
  18806=>"001001000",
  18807=>"110110000",
  18808=>"111111111",
  18809=>"111110001",
  18810=>"000000000",
  18811=>"111101000",
  18812=>"001000100",
  18813=>"111111111",
  18814=>"000000001",
  18815=>"000111111",
  18816=>"000000000",
  18817=>"000000000",
  18818=>"000000111",
  18819=>"000001000",
  18820=>"111111111",
  18821=>"011111111",
  18822=>"100111111",
  18823=>"001000000",
  18824=>"000000111",
  18825=>"111111000",
  18826=>"111111111",
  18827=>"111111011",
  18828=>"000000111",
  18829=>"000000111",
  18830=>"111111000",
  18831=>"000000101",
  18832=>"000000000",
  18833=>"001001111",
  18834=>"001000001",
  18835=>"110111110",
  18836=>"111111111",
  18837=>"000011010",
  18838=>"000000000",
  18839=>"111110100",
  18840=>"000000000",
  18841=>"111111111",
  18842=>"000000000",
  18843=>"001000000",
  18844=>"000001111",
  18845=>"001010111",
  18846=>"111111111",
  18847=>"000010110",
  18848=>"111111110",
  18849=>"110110000",
  18850=>"000010000",
  18851=>"111101100",
  18852=>"111111111",
  18853=>"000000000",
  18854=>"101001101",
  18855=>"111111100",
  18856=>"111111111",
  18857=>"010011000",
  18858=>"000001111",
  18859=>"111000010",
  18860=>"111111100",
  18861=>"110000100",
  18862=>"110111101",
  18863=>"000000100",
  18864=>"100111111",
  18865=>"001011001",
  18866=>"000000011",
  18867=>"000100100",
  18868=>"111100000",
  18869=>"111000000",
  18870=>"000110000",
  18871=>"011011000",
  18872=>"000000000",
  18873=>"001011001",
  18874=>"010011111",
  18875=>"000011111",
  18876=>"001000000",
  18877=>"000000001",
  18878=>"111111000",
  18879=>"111011001",
  18880=>"110110000",
  18881=>"000000000",
  18882=>"111111111",
  18883=>"000000111",
  18884=>"000000000",
  18885=>"111101001",
  18886=>"000000000",
  18887=>"000001111",
  18888=>"100100110",
  18889=>"000000000",
  18890=>"111000000",
  18891=>"000000000",
  18892=>"000000001",
  18893=>"111111111",
  18894=>"000000010",
  18895=>"111000000",
  18896=>"001000011",
  18897=>"010111111",
  18898=>"111111011",
  18899=>"100000001",
  18900=>"000001111",
  18901=>"000000000",
  18902=>"100111111",
  18903=>"011011011",
  18904=>"000000000",
  18905=>"000000000",
  18906=>"010000110",
  18907=>"100100110",
  18908=>"111100111",
  18909=>"111111111",
  18910=>"001001111",
  18911=>"111111010",
  18912=>"001001111",
  18913=>"111111111",
  18914=>"100000000",
  18915=>"111000000",
  18916=>"111111111",
  18917=>"110111111",
  18918=>"011011111",
  18919=>"000000000",
  18920=>"111011000",
  18921=>"101001100",
  18922=>"000000000",
  18923=>"001001001",
  18924=>"110110111",
  18925=>"000001001",
  18926=>"110111111",
  18927=>"111001000",
  18928=>"111111111",
  18929=>"000111111",
  18930=>"001111111",
  18931=>"011000100",
  18932=>"000000100",
  18933=>"000000011",
  18934=>"100100100",
  18935=>"000100000",
  18936=>"000000000",
  18937=>"000000000",
  18938=>"110111110",
  18939=>"000000000",
  18940=>"011111111",
  18941=>"000001001",
  18942=>"001000000",
  18943=>"111111000",
  18944=>"011001111",
  18945=>"111111000",
  18946=>"000000100",
  18947=>"000000111",
  18948=>"111111111",
  18949=>"011001011",
  18950=>"000000000",
  18951=>"111111111",
  18952=>"101111111",
  18953=>"011000110",
  18954=>"110011001",
  18955=>"100000001",
  18956=>"001001000",
  18957=>"111111111",
  18958=>"000000110",
  18959=>"111110000",
  18960=>"111111111",
  18961=>"000000000",
  18962=>"100000000",
  18963=>"011001100",
  18964=>"110010000",
  18965=>"000000000",
  18966=>"111111111",
  18967=>"001001000",
  18968=>"111110111",
  18969=>"111111000",
  18970=>"001111101",
  18971=>"000001111",
  18972=>"111111111",
  18973=>"001000000",
  18974=>"111001111",
  18975=>"010100001",
  18976=>"111111111",
  18977=>"000000000",
  18978=>"000011111",
  18979=>"111111111",
  18980=>"001001011",
  18981=>"011011111",
  18982=>"000000000",
  18983=>"000111111",
  18984=>"000100110",
  18985=>"000000000",
  18986=>"000000100",
  18987=>"000000000",
  18988=>"000010011",
  18989=>"000000001",
  18990=>"111111111",
  18991=>"000001000",
  18992=>"111111111",
  18993=>"111111111",
  18994=>"001000000",
  18995=>"000000000",
  18996=>"111010000",
  18997=>"111001001",
  18998=>"000100110",
  18999=>"111001111",
  19000=>"111101111",
  19001=>"111111111",
  19002=>"000000111",
  19003=>"011111111",
  19004=>"000000000",
  19005=>"000000000",
  19006=>"100000110",
  19007=>"000000000",
  19008=>"110111100",
  19009=>"011101111",
  19010=>"111111111",
  19011=>"111011011",
  19012=>"001011111",
  19013=>"000000000",
  19014=>"000000000",
  19015=>"111111111",
  19016=>"011001011",
  19017=>"101000101",
  19018=>"111111111",
  19019=>"110110001",
  19020=>"110001111",
  19021=>"111000000",
  19022=>"001100111",
  19023=>"100000110",
  19024=>"000000000",
  19025=>"111111111",
  19026=>"000000110",
  19027=>"001001111",
  19028=>"000000000",
  19029=>"111001000",
  19030=>"100000001",
  19031=>"000000000",
  19032=>"001001111",
  19033=>"111111110",
  19034=>"000000000",
  19035=>"000110000",
  19036=>"111101101",
  19037=>"110011000",
  19038=>"110000000",
  19039=>"110110110",
  19040=>"111111111",
  19041=>"111111111",
  19042=>"011111010",
  19043=>"111111111",
  19044=>"110111111",
  19045=>"100111111",
  19046=>"010000111",
  19047=>"111011000",
  19048=>"000000000",
  19049=>"000000000",
  19050=>"110101111",
  19051=>"000000000",
  19052=>"011011011",
  19053=>"111111111",
  19054=>"000110000",
  19055=>"000000001",
  19056=>"111111111",
  19057=>"111001011",
  19058=>"100111111",
  19059=>"110111011",
  19060=>"111110000",
  19061=>"111111111",
  19062=>"111111111",
  19063=>"000000011",
  19064=>"011110000",
  19065=>"000000000",
  19066=>"111111111",
  19067=>"111111111",
  19068=>"011011011",
  19069=>"000000000",
  19070=>"001111000",
  19071=>"000001001",
  19072=>"000000000",
  19073=>"000111000",
  19074=>"010000000",
  19075=>"010111111",
  19076=>"111111111",
  19077=>"111000000",
  19078=>"000000010",
  19079=>"111110110",
  19080=>"111000000",
  19081=>"000000111",
  19082=>"000000100",
  19083=>"111111000",
  19084=>"011000000",
  19085=>"000000000",
  19086=>"110010111",
  19087=>"000000111",
  19088=>"111111101",
  19089=>"000111111",
  19090=>"001001111",
  19091=>"001000000",
  19092=>"111111111",
  19093=>"111111000",
  19094=>"000111111",
  19095=>"000000000",
  19096=>"000000110",
  19097=>"111111110",
  19098=>"111111110",
  19099=>"110110111",
  19100=>"000000111",
  19101=>"001000100",
  19102=>"111000001",
  19103=>"000000000",
  19104=>"110111110",
  19105=>"011001001",
  19106=>"000000111",
  19107=>"000001111",
  19108=>"111001111",
  19109=>"111110111",
  19110=>"110111000",
  19111=>"111110010",
  19112=>"000010000",
  19113=>"111111101",
  19114=>"000111111",
  19115=>"111111111",
  19116=>"100001001",
  19117=>"001111111",
  19118=>"000010000",
  19119=>"000000000",
  19120=>"000000111",
  19121=>"111111011",
  19122=>"111111111",
  19123=>"111001101",
  19124=>"000000000",
  19125=>"111011000",
  19126=>"111011000",
  19127=>"000000100",
  19128=>"000000000",
  19129=>"000000000",
  19130=>"101111111",
  19131=>"110110011",
  19132=>"000001001",
  19133=>"000000000",
  19134=>"000000000",
  19135=>"001000000",
  19136=>"111111111",
  19137=>"000000000",
  19138=>"101001001",
  19139=>"110110010",
  19140=>"111101100",
  19141=>"000000000",
  19142=>"000000000",
  19143=>"001111000",
  19144=>"101111111",
  19145=>"010001011",
  19146=>"111111111",
  19147=>"111111111",
  19148=>"001000000",
  19149=>"000111001",
  19150=>"000000101",
  19151=>"000000000",
  19152=>"000000000",
  19153=>"110111111",
  19154=>"111111111",
  19155=>"000000000",
  19156=>"001000011",
  19157=>"111111111",
  19158=>"000000000",
  19159=>"000001001",
  19160=>"000000000",
  19161=>"000000111",
  19162=>"000000000",
  19163=>"000111111",
  19164=>"000111111",
  19165=>"011000000",
  19166=>"000000000",
  19167=>"001001001",
  19168=>"000000000",
  19169=>"111000000",
  19170=>"000110000",
  19171=>"100000000",
  19172=>"000000100",
  19173=>"000000000",
  19174=>"110111101",
  19175=>"111011000",
  19176=>"100100100",
  19177=>"111111011",
  19178=>"000000000",
  19179=>"010000000",
  19180=>"000000000",
  19181=>"000000000",
  19182=>"110111000",
  19183=>"000001111",
  19184=>"111111111",
  19185=>"100101101",
  19186=>"000000000",
  19187=>"000000000",
  19188=>"000000000",
  19189=>"011011011",
  19190=>"111111101",
  19191=>"000000000",
  19192=>"000000000",
  19193=>"000000000",
  19194=>"000000001",
  19195=>"101001000",
  19196=>"000110100",
  19197=>"110000000",
  19198=>"000000000",
  19199=>"000000000",
  19200=>"111011011",
  19201=>"010000000",
  19202=>"100000000",
  19203=>"111111111",
  19204=>"000010110",
  19205=>"111011111",
  19206=>"000000000",
  19207=>"111111000",
  19208=>"000000001",
  19209=>"111111000",
  19210=>"000000100",
  19211=>"000100111",
  19212=>"111111111",
  19213=>"000000000",
  19214=>"111111111",
  19215=>"111011000",
  19216=>"111111000",
  19217=>"111111111",
  19218=>"111000010",
  19219=>"000000001",
  19220=>"111000000",
  19221=>"101000000",
  19222=>"011011111",
  19223=>"111110000",
  19224=>"011011011",
  19225=>"111000001",
  19226=>"101000100",
  19227=>"110100100",
  19228=>"000100000",
  19229=>"111011111",
  19230=>"011001111",
  19231=>"000000000",
  19232=>"001101111",
  19233=>"001001111",
  19234=>"001111111",
  19235=>"110010000",
  19236=>"000000110",
  19237=>"000000001",
  19238=>"000000100",
  19239=>"011001000",
  19240=>"100110110",
  19241=>"000000111",
  19242=>"010100101",
  19243=>"011000000",
  19244=>"000001000",
  19245=>"000000001",
  19246=>"111011000",
  19247=>"000000000",
  19248=>"111111111",
  19249=>"011011100",
  19250=>"110111111",
  19251=>"111000000",
  19252=>"111111111",
  19253=>"011011001",
  19254=>"000000000",
  19255=>"000101111",
  19256=>"000000111",
  19257=>"000000001",
  19258=>"000000000",
  19259=>"111111111",
  19260=>"110000000",
  19261=>"000000111",
  19262=>"100110111",
  19263=>"000000111",
  19264=>"111111111",
  19265=>"011001011",
  19266=>"000000000",
  19267=>"000000000",
  19268=>"000000000",
  19269=>"000000000",
  19270=>"000000000",
  19271=>"101001111",
  19272=>"000100000",
  19273=>"111000111",
  19274=>"000100000",
  19275=>"111110100",
  19276=>"011111011",
  19277=>"000000000",
  19278=>"011111110",
  19279=>"000000000",
  19280=>"100100000",
  19281=>"000000000",
  19282=>"000000000",
  19283=>"000000000",
  19284=>"001000000",
  19285=>"111110111",
  19286=>"111110001",
  19287=>"111111111",
  19288=>"111111111",
  19289=>"110111111",
  19290=>"111000111",
  19291=>"111110110",
  19292=>"000000000",
  19293=>"000000011",
  19294=>"111001000",
  19295=>"000001001",
  19296=>"011001001",
  19297=>"111111111",
  19298=>"101110111",
  19299=>"000101101",
  19300=>"000001000",
  19301=>"111111101",
  19302=>"000000000",
  19303=>"111111010",
  19304=>"111111001",
  19305=>"111111111",
  19306=>"111111111",
  19307=>"100110110",
  19308=>"000001000",
  19309=>"100111111",
  19310=>"111011011",
  19311=>"000000000",
  19312=>"111111011",
  19313=>"100111111",
  19314=>"111111110",
  19315=>"111110100",
  19316=>"100101111",
  19317=>"000000000",
  19318=>"000000110",
  19319=>"010010000",
  19320=>"110000000",
  19321=>"000101111",
  19322=>"111111110",
  19323=>"111110111",
  19324=>"111111111",
  19325=>"011000000",
  19326=>"001100100",
  19327=>"111111111",
  19328=>"111111111",
  19329=>"000000000",
  19330=>"000000000",
  19331=>"111111111",
  19332=>"000000000",
  19333=>"100000000",
  19334=>"110010001",
  19335=>"011000001",
  19336=>"111110010",
  19337=>"111111101",
  19338=>"111111010",
  19339=>"000000000",
  19340=>"111111111",
  19341=>"001111100",
  19342=>"010000000",
  19343=>"000100110",
  19344=>"111111111",
  19345=>"111111101",
  19346=>"000000000",
  19347=>"111101000",
  19348=>"100000000",
  19349=>"000110000",
  19350=>"111111111",
  19351=>"001001111",
  19352=>"111111111",
  19353=>"100100111",
  19354=>"110111111",
  19355=>"001001011",
  19356=>"001011000",
  19357=>"000000000",
  19358=>"000000000",
  19359=>"000000000",
  19360=>"111111000",
  19361=>"100000000",
  19362=>"000110111",
  19363=>"000000000",
  19364=>"000000111",
  19365=>"000001111",
  19366=>"111111111",
  19367=>"110110111",
  19368=>"000000110",
  19369=>"010000000",
  19370=>"000000111",
  19371=>"000000010",
  19372=>"000000000",
  19373=>"110110111",
  19374=>"000001011",
  19375=>"111111110",
  19376=>"001001111",
  19377=>"111010100",
  19378=>"000001111",
  19379=>"000011001",
  19380=>"110111111",
  19381=>"111111111",
  19382=>"111111111",
  19383=>"000001010",
  19384=>"001001111",
  19385=>"000000111",
  19386=>"110000000",
  19387=>"110000000",
  19388=>"000000001",
  19389=>"111111111",
  19390=>"000000111",
  19391=>"111110010",
  19392=>"000110110",
  19393=>"111111111",
  19394=>"000000000",
  19395=>"000011111",
  19396=>"000000000",
  19397=>"111011011",
  19398=>"111101101",
  19399=>"000000000",
  19400=>"100000111",
  19401=>"100100111",
  19402=>"000001001",
  19403=>"001111111",
  19404=>"000000000",
  19405=>"100111111",
  19406=>"000000001",
  19407=>"111111111",
  19408=>"111000101",
  19409=>"010000000",
  19410=>"000000000",
  19411=>"000000000",
  19412=>"110110110",
  19413=>"010000110",
  19414=>"111000000",
  19415=>"000000011",
  19416=>"000110111",
  19417=>"001111111",
  19418=>"001000000",
  19419=>"111011011",
  19420=>"111111111",
  19421=>"011111000",
  19422=>"000000001",
  19423=>"000000000",
  19424=>"000111110",
  19425=>"000001111",
  19426=>"111111111",
  19427=>"000100111",
  19428=>"001110000",
  19429=>"000000000",
  19430=>"000110111",
  19431=>"010010000",
  19432=>"000000111",
  19433=>"111111111",
  19434=>"111110000",
  19435=>"000000000",
  19436=>"011001000",
  19437=>"111111111",
  19438=>"000000000",
  19439=>"000000000",
  19440=>"101100111",
  19441=>"000000000",
  19442=>"111111111",
  19443=>"100100000",
  19444=>"001001111",
  19445=>"000110000",
  19446=>"111111111",
  19447=>"010111111",
  19448=>"011001000",
  19449=>"110110111",
  19450=>"000000111",
  19451=>"011111111",
  19452=>"110000101",
  19453=>"111111000",
  19454=>"000000100",
  19455=>"111011011",
  19456=>"000010111",
  19457=>"000001001",
  19458=>"000000110",
  19459=>"111111100",
  19460=>"111111111",
  19461=>"000000000",
  19462=>"001000000",
  19463=>"000000000",
  19464=>"111001000",
  19465=>"111111111",
  19466=>"011111111",
  19467=>"111000000",
  19468=>"111111110",
  19469=>"000011111",
  19470=>"111100110",
  19471=>"000100111",
  19472=>"011111111",
  19473=>"111111111",
  19474=>"111000000",
  19475=>"011001111",
  19476=>"011010000",
  19477=>"000000000",
  19478=>"110000000",
  19479=>"110010001",
  19480=>"110110111",
  19481=>"001000000",
  19482=>"101001001",
  19483=>"001001100",
  19484=>"000110110",
  19485=>"111111111",
  19486=>"100100000",
  19487=>"001001001",
  19488=>"000000001",
  19489=>"000000111",
  19490=>"111011010",
  19491=>"111101000",
  19492=>"000111111",
  19493=>"111110110",
  19494=>"100100111",
  19495=>"000011000",
  19496=>"110000000",
  19497=>"111000000",
  19498=>"111111111",
  19499=>"111111110",
  19500=>"000000000",
  19501=>"111100000",
  19502=>"101100000",
  19503=>"000110111",
  19504=>"100111111",
  19505=>"011000000",
  19506=>"001011011",
  19507=>"000101000",
  19508=>"001101101",
  19509=>"111011011",
  19510=>"110110001",
  19511=>"100111111",
  19512=>"100111111",
  19513=>"100100111",
  19514=>"000000000",
  19515=>"100110111",
  19516=>"000000111",
  19517=>"111101111",
  19518=>"000111111",
  19519=>"111001000",
  19520=>"100100100",
  19521=>"000111111",
  19522=>"100111000",
  19523=>"000000111",
  19524=>"000001000",
  19525=>"000000100",
  19526=>"111000000",
  19527=>"000000000",
  19528=>"001011001",
  19529=>"000000111",
  19530=>"000111111",
  19531=>"011011111",
  19532=>"000000110",
  19533=>"111111111",
  19534=>"001111111",
  19535=>"111001000",
  19536=>"011001000",
  19537=>"100100111",
  19538=>"000100110",
  19539=>"100010000",
  19540=>"000000000",
  19541=>"011011111",
  19542=>"000000111",
  19543=>"000111111",
  19544=>"000001011",
  19545=>"000000000",
  19546=>"000000000",
  19547=>"100000011",
  19548=>"000111111",
  19549=>"000000111",
  19550=>"110000000",
  19551=>"100000000",
  19552=>"000111111",
  19553=>"111000000",
  19554=>"001000000",
  19555=>"111000000",
  19556=>"001101110",
  19557=>"111000000",
  19558=>"111111001",
  19559=>"000000000",
  19560=>"111111000",
  19561=>"111111110",
  19562=>"000000000",
  19563=>"000000011",
  19564=>"010111111",
  19565=>"111000000",
  19566=>"000000000",
  19567=>"000100111",
  19568=>"100100111",
  19569=>"001001111",
  19570=>"100100000",
  19571=>"111100000",
  19572=>"000110111",
  19573=>"111111000",
  19574=>"001001111",
  19575=>"111011000",
  19576=>"101101001",
  19577=>"111101111",
  19578=>"000001001",
  19579=>"000111010",
  19580=>"111010000",
  19581=>"010011011",
  19582=>"011001111",
  19583=>"000001111",
  19584=>"111000000",
  19585=>"000000111",
  19586=>"111011111",
  19587=>"101111010",
  19588=>"000001111",
  19589=>"101000000",
  19590=>"111111111",
  19591=>"111111111",
  19592=>"111100100",
  19593=>"111000000",
  19594=>"111000000",
  19595=>"111000000",
  19596=>"000011111",
  19597=>"011000000",
  19598=>"101000111",
  19599=>"011000000",
  19600=>"111101111",
  19601=>"100100000",
  19602=>"000000000",
  19603=>"000111111",
  19604=>"111010011",
  19605=>"000000110",
  19606=>"111000101",
  19607=>"111001000",
  19608=>"000110000",
  19609=>"111111110",
  19610=>"000110000",
  19611=>"010111111",
  19612=>"000110000",
  19613=>"111000001",
  19614=>"000000001",
  19615=>"111111001",
  19616=>"000000111",
  19617=>"111111000",
  19618=>"010111111",
  19619=>"011001000",
  19620=>"111001011",
  19621=>"111011000",
  19622=>"111111011",
  19623=>"000110000",
  19624=>"000000000",
  19625=>"001000010",
  19626=>"111111001",
  19627=>"011000000",
  19628=>"111111110",
  19629=>"100011111",
  19630=>"110101110",
  19631=>"101000000",
  19632=>"111000000",
  19633=>"110111000",
  19634=>"111110010",
  19635=>"111001000",
  19636=>"000000001",
  19637=>"000000000",
  19638=>"111111111",
  19639=>"011111111",
  19640=>"000000111",
  19641=>"000111111",
  19642=>"011000000",
  19643=>"111000000",
  19644=>"000011000",
  19645=>"000000111",
  19646=>"001000000",
  19647=>"101011111",
  19648=>"000000100",
  19649=>"110100000",
  19650=>"000000000",
  19651=>"000111111",
  19652=>"000000000",
  19653=>"111000000",
  19654=>"000100000",
  19655=>"101001000",
  19656=>"100000000",
  19657=>"111001000",
  19658=>"101000100",
  19659=>"011011000",
  19660=>"111111111",
  19661=>"000000000",
  19662=>"011011001",
  19663=>"011011001",
  19664=>"000000101",
  19665=>"110000100",
  19666=>"000111111",
  19667=>"011001001",
  19668=>"011000000",
  19669=>"111001000",
  19670=>"110100000",
  19671=>"111110110",
  19672=>"001001111",
  19673=>"000000000",
  19674=>"110000000",
  19675=>"000111111",
  19676=>"110110000",
  19677=>"000001011",
  19678=>"010000000",
  19679=>"000000000",
  19680=>"000111111",
  19681=>"100000000",
  19682=>"000111111",
  19683=>"000000000",
  19684=>"000111000",
  19685=>"001000100",
  19686=>"101000000",
  19687=>"000011111",
  19688=>"011111111",
  19689=>"111111111",
  19690=>"111001000",
  19691=>"000000000",
  19692=>"111000001",
  19693=>"110000000",
  19694=>"111111101",
  19695=>"110111111",
  19696=>"111011001",
  19697=>"011011000",
  19698=>"000110111",
  19699=>"111111000",
  19700=>"001111011",
  19701=>"000000000",
  19702=>"000111111",
  19703=>"011111111",
  19704=>"111101001",
  19705=>"000000000",
  19706=>"000000000",
  19707=>"000000000",
  19708=>"000000000",
  19709=>"100100100",
  19710=>"110111111",
  19711=>"001100000",
  19712=>"000000011",
  19713=>"100110000",
  19714=>"000111111",
  19715=>"001000000",
  19716=>"000111111",
  19717=>"101111000",
  19718=>"111000000",
  19719=>"000000001",
  19720=>"110111111",
  19721=>"000011011",
  19722=>"111111111",
  19723=>"111001000",
  19724=>"111000000",
  19725=>"000000000",
  19726=>"000111110",
  19727=>"111111111",
  19728=>"000000000",
  19729=>"011010000",
  19730=>"100000000",
  19731=>"000000000",
  19732=>"111111000",
  19733=>"000010111",
  19734=>"011111111",
  19735=>"001111011",
  19736=>"111100000",
  19737=>"001111000",
  19738=>"111101111",
  19739=>"001000000",
  19740=>"000110100",
  19741=>"011111111",
  19742=>"111111111",
  19743=>"110111100",
  19744=>"000000000",
  19745=>"000000000",
  19746=>"110000000",
  19747=>"110000011",
  19748=>"111111100",
  19749=>"000001101",
  19750=>"111011000",
  19751=>"100000110",
  19752=>"110100000",
  19753=>"100000000",
  19754=>"111111000",
  19755=>"111000000",
  19756=>"000000000",
  19757=>"000110110",
  19758=>"010000000",
  19759=>"010010001",
  19760=>"000100111",
  19761=>"011011000",
  19762=>"111111110",
  19763=>"001111111",
  19764=>"000001001",
  19765=>"000000110",
  19766=>"000101000",
  19767=>"000000111",
  19768=>"101101000",
  19769=>"001111111",
  19770=>"000000000",
  19771=>"111111100",
  19772=>"111111100",
  19773=>"111110110",
  19774=>"110000000",
  19775=>"000000111",
  19776=>"111111100",
  19777=>"111000000",
  19778=>"000000010",
  19779=>"100111100",
  19780=>"000111111",
  19781=>"011011000",
  19782=>"011010000",
  19783=>"000000111",
  19784=>"000000000",
  19785=>"111111111",
  19786=>"000000000",
  19787=>"011000111",
  19788=>"000001001",
  19789=>"001000000",
  19790=>"010000000",
  19791=>"001001000",
  19792=>"000111111",
  19793=>"111111111",
  19794=>"110010000",
  19795=>"100000100",
  19796=>"000000000",
  19797=>"011011011",
  19798=>"000000000",
  19799=>"100111111",
  19800=>"111110000",
  19801=>"000011011",
  19802=>"000010011",
  19803=>"111001100",
  19804=>"111000000",
  19805=>"111111000",
  19806=>"001000000",
  19807=>"000000000",
  19808=>"000000011",
  19809=>"111111000",
  19810=>"111110011",
  19811=>"000000111",
  19812=>"100000000",
  19813=>"000000000",
  19814=>"000000000",
  19815=>"000001111",
  19816=>"100100110",
  19817=>"000111111",
  19818=>"111111110",
  19819=>"111001111",
  19820=>"100000111",
  19821=>"010011001",
  19822=>"000000000",
  19823=>"110100000",
  19824=>"000000000",
  19825=>"111111010",
  19826=>"000000111",
  19827=>"111001011",
  19828=>"000010000",
  19829=>"000000000",
  19830=>"111111111",
  19831=>"111111111",
  19832=>"000000000",
  19833=>"111111111",
  19834=>"111111001",
  19835=>"110001000",
  19836=>"111111010",
  19837=>"111001000",
  19838=>"000001001",
  19839=>"000000000",
  19840=>"000000111",
  19841=>"111001001",
  19842=>"000010011",
  19843=>"101011000",
  19844=>"111111111",
  19845=>"111111000",
  19846=>"000011011",
  19847=>"100000000",
  19848=>"110000000",
  19849=>"111110000",
  19850=>"000111111",
  19851=>"111111110",
  19852=>"000000111",
  19853=>"111001001",
  19854=>"100000000",
  19855=>"000000000",
  19856=>"000001001",
  19857=>"000000001",
  19858=>"001011011",
  19859=>"111111111",
  19860=>"001000001",
  19861=>"000000000",
  19862=>"011001111",
  19863=>"111111001",
  19864=>"101110110",
  19865=>"000111111",
  19866=>"000111111",
  19867=>"000000000",
  19868=>"010011111",
  19869=>"100000010",
  19870=>"111010000",
  19871=>"000000100",
  19872=>"000001001",
  19873=>"110110000",
  19874=>"110000000",
  19875=>"111111111",
  19876=>"111100000",
  19877=>"000111001",
  19878=>"110011000",
  19879=>"111111111",
  19880=>"001111100",
  19881=>"100110000",
  19882=>"000000000",
  19883=>"111100000",
  19884=>"100111111",
  19885=>"000000000",
  19886=>"111111111",
  19887=>"101111111",
  19888=>"111111011",
  19889=>"111000111",
  19890=>"111111111",
  19891=>"000000111",
  19892=>"111110000",
  19893=>"000000100",
  19894=>"000000100",
  19895=>"000000000",
  19896=>"000000010",
  19897=>"111000000",
  19898=>"011000010",
  19899=>"000000000",
  19900=>"001011111",
  19901=>"111111000",
  19902=>"101000000",
  19903=>"111111000",
  19904=>"111111011",
  19905=>"111110110",
  19906=>"110100000",
  19907=>"100101111",
  19908=>"111111111",
  19909=>"001011111",
  19910=>"000000000",
  19911=>"100000000",
  19912=>"000000100",
  19913=>"111000000",
  19914=>"000000001",
  19915=>"101100000",
  19916=>"000111000",
  19917=>"011011111",
  19918=>"100111111",
  19919=>"111111000",
  19920=>"111000001",
  19921=>"111010000",
  19922=>"000000100",
  19923=>"000010111",
  19924=>"110111111",
  19925=>"001011111",
  19926=>"100011111",
  19927=>"100000000",
  19928=>"111101000",
  19929=>"000000000",
  19930=>"111111010",
  19931=>"110000000",
  19932=>"000001010",
  19933=>"000110010",
  19934=>"111111111",
  19935=>"110010011",
  19936=>"111111110",
  19937=>"010111010",
  19938=>"000000000",
  19939=>"110000111",
  19940=>"111000000",
  19941=>"011110101",
  19942=>"100111000",
  19943=>"001000111",
  19944=>"000001010",
  19945=>"000111101",
  19946=>"000000001",
  19947=>"111011000",
  19948=>"111110000",
  19949=>"001000000",
  19950=>"111110100",
  19951=>"110110111",
  19952=>"011000000",
  19953=>"000011011",
  19954=>"111111111",
  19955=>"100000000",
  19956=>"011111110",
  19957=>"000000111",
  19958=>"111111111",
  19959=>"011011000",
  19960=>"000100000",
  19961=>"000000000",
  19962=>"000001110",
  19963=>"000111111",
  19964=>"000111100",
  19965=>"000110111",
  19966=>"100111111",
  19967=>"110000000",
  19968=>"111111100",
  19969=>"000000001",
  19970=>"110110110",
  19971=>"111000000",
  19972=>"111111000",
  19973=>"111100000",
  19974=>"000111111",
  19975=>"111111111",
  19976=>"111000110",
  19977=>"001001000",
  19978=>"111101111",
  19979=>"111000000",
  19980=>"010010111",
  19981=>"000000000",
  19982=>"100000000",
  19983=>"000000111",
  19984=>"000000000",
  19985=>"111111000",
  19986=>"011111111",
  19987=>"000000000",
  19988=>"000000111",
  19989=>"000000000",
  19990=>"000000000",
  19991=>"111111111",
  19992=>"001100101",
  19993=>"001000000",
  19994=>"000100100",
  19995=>"111100001",
  19996=>"001111111",
  19997=>"111111000",
  19998=>"011001001",
  19999=>"000011111",
  20000=>"101111011",
  20001=>"000000000",
  20002=>"111101101",
  20003=>"101001001",
  20004=>"100000000",
  20005=>"111010111",
  20006=>"111111000",
  20007=>"000100000",
  20008=>"111111101",
  20009=>"000000000",
  20010=>"110100111",
  20011=>"010111110",
  20012=>"000000110",
  20013=>"001011111",
  20014=>"000001000",
  20015=>"000000111",
  20016=>"111111000",
  20017=>"000000011",
  20018=>"000111111",
  20019=>"000110111",
  20020=>"001111111",
  20021=>"011011000",
  20022=>"001001000",
  20023=>"011000000",
  20024=>"010111111",
  20025=>"000000000",
  20026=>"000000000",
  20027=>"011000111",
  20028=>"111100110",
  20029=>"111111111",
  20030=>"111001000",
  20031=>"000000111",
  20032=>"001000111",
  20033=>"100000000",
  20034=>"111111111",
  20035=>"111100110",
  20036=>"011001001",
  20037=>"111001000",
  20038=>"000000100",
  20039=>"000000000",
  20040=>"101111111",
  20041=>"111111110",
  20042=>"000000111",
  20043=>"000011110",
  20044=>"101110111",
  20045=>"111000000",
  20046=>"001011001",
  20047=>"111111111",
  20048=>"111101000",
  20049=>"000000001",
  20050=>"000001111",
  20051=>"011001000",
  20052=>"001001000",
  20053=>"111111110",
  20054=>"100000000",
  20055=>"111000000",
  20056=>"001101111",
  20057=>"111111111",
  20058=>"111111001",
  20059=>"101100100",
  20060=>"111111111",
  20061=>"111011000",
  20062=>"111100000",
  20063=>"000111111",
  20064=>"001000011",
  20065=>"001000000",
  20066=>"111101000",
  20067=>"100111111",
  20068=>"011111000",
  20069=>"000000000",
  20070=>"010000110",
  20071=>"000111000",
  20072=>"110101111",
  20073=>"010000000",
  20074=>"100100111",
  20075=>"001100110",
  20076=>"111110111",
  20077=>"000000111",
  20078=>"100100111",
  20079=>"111111000",
  20080=>"000011000",
  20081=>"000000000",
  20082=>"011011000",
  20083=>"111111001",
  20084=>"000000000",
  20085=>"000000110",
  20086=>"000111111",
  20087=>"000000111",
  20088=>"001000001",
  20089=>"111100100",
  20090=>"000000000",
  20091=>"110111011",
  20092=>"111111111",
  20093=>"110100000",
  20094=>"000000000",
  20095=>"000000000",
  20096=>"100000000",
  20097=>"010010000",
  20098=>"000000111",
  20099=>"111111000",
  20100=>"011111000",
  20101=>"111000111",
  20102=>"011000000",
  20103=>"001111101",
  20104=>"111111101",
  20105=>"000000000",
  20106=>"111111101",
  20107=>"001111110",
  20108=>"001001000",
  20109=>"000000000",
  20110=>"000001111",
  20111=>"001001111",
  20112=>"000110111",
  20113=>"001000000",
  20114=>"000000010",
  20115=>"000111111",
  20116=>"111111100",
  20117=>"000000000",
  20118=>"000000001",
  20119=>"111111011",
  20120=>"011000000",
  20121=>"111111100",
  20122=>"011000000",
  20123=>"010000001",
  20124=>"111111011",
  20125=>"111111001",
  20126=>"000000111",
  20127=>"000110100",
  20128=>"001001000",
  20129=>"101000101",
  20130=>"111111001",
  20131=>"000111010",
  20132=>"011111111",
  20133=>"110111111",
  20134=>"000111111",
  20135=>"110010001",
  20136=>"100010000",
  20137=>"000000111",
  20138=>"001001000",
  20139=>"111111000",
  20140=>"000111111",
  20141=>"000100110",
  20142=>"000000000",
  20143=>"111111110",
  20144=>"000000000",
  20145=>"111001100",
  20146=>"000111000",
  20147=>"000111111",
  20148=>"110000000",
  20149=>"001111111",
  20150=>"100000101",
  20151=>"000000000",
  20152=>"011000111",
  20153=>"111111000",
  20154=>"000000000",
  20155=>"111011000",
  20156=>"000000000",
  20157=>"111001111",
  20158=>"111111111",
  20159=>"100010000",
  20160=>"011010000",
  20161=>"010001001",
  20162=>"100001000",
  20163=>"111001000",
  20164=>"000100100",
  20165=>"111010000",
  20166=>"000000111",
  20167=>"111111111",
  20168=>"001000100",
  20169=>"000000000",
  20170=>"000000000",
  20171=>"000000000",
  20172=>"101110111",
  20173=>"111111111",
  20174=>"000000001",
  20175=>"000111000",
  20176=>"000000000",
  20177=>"100000111",
  20178=>"111100100",
  20179=>"111000011",
  20180=>"101111011",
  20181=>"000100111",
  20182=>"100000010",
  20183=>"111011101",
  20184=>"111111010",
  20185=>"111100111",
  20186=>"111111101",
  20187=>"000000000",
  20188=>"111111111",
  20189=>"000100100",
  20190=>"111111000",
  20191=>"000000001",
  20192=>"000000000",
  20193=>"000011011",
  20194=>"101000000",
  20195=>"111000000",
  20196=>"111111111",
  20197=>"111111001",
  20198=>"101001001",
  20199=>"111111111",
  20200=>"111111111",
  20201=>"011011000",
  20202=>"111011000",
  20203=>"111000111",
  20204=>"111010111",
  20205=>"110110111",
  20206=>"111110111",
  20207=>"001101100",
  20208=>"000000011",
  20209=>"110111000",
  20210=>"000000001",
  20211=>"000001000",
  20212=>"110111000",
  20213=>"000000100",
  20214=>"110110000",
  20215=>"111111000",
  20216=>"001000001",
  20217=>"000001101",
  20218=>"000000000",
  20219=>"011011011",
  20220=>"111111111",
  20221=>"000111111",
  20222=>"100111111",
  20223=>"111111110",
  20224=>"111111000",
  20225=>"000000111",
  20226=>"111111011",
  20227=>"111111111",
  20228=>"001110000",
  20229=>"001011011",
  20230=>"111111000",
  20231=>"000000000",
  20232=>"000000000",
  20233=>"111111111",
  20234=>"111101101",
  20235=>"111101000",
  20236=>"000100000",
  20237=>"000000000",
  20238=>"111110110",
  20239=>"000000000",
  20240=>"000111111",
  20241=>"001000000",
  20242=>"000000000",
  20243=>"000000000",
  20244=>"000000110",
  20245=>"001000000",
  20246=>"101101111",
  20247=>"000000100",
  20248=>"111111000",
  20249=>"110101000",
  20250=>"110000000",
  20251=>"000000101",
  20252=>"110111110",
  20253=>"111000000",
  20254=>"011111111",
  20255=>"000101111",
  20256=>"011000000",
  20257=>"000000000",
  20258=>"110010000",
  20259=>"001000000",
  20260=>"000000111",
  20261=>"001100111",
  20262=>"111100110",
  20263=>"011011000",
  20264=>"000111111",
  20265=>"011110101",
  20266=>"000000000",
  20267=>"000000111",
  20268=>"111111111",
  20269=>"110000000",
  20270=>"000000011",
  20271=>"000001111",
  20272=>"011111100",
  20273=>"000000001",
  20274=>"000000000",
  20275=>"111111000",
  20276=>"000000000",
  20277=>"111111010",
  20278=>"111111000",
  20279=>"111100000",
  20280=>"111111101",
  20281=>"101111000",
  20282=>"000000000",
  20283=>"111001000",
  20284=>"111110100",
  20285=>"100100100",
  20286=>"111001110",
  20287=>"000000000",
  20288=>"000000000",
  20289=>"111111111",
  20290=>"111111111",
  20291=>"100000000",
  20292=>"100100100",
  20293=>"101001111",
  20294=>"000000000",
  20295=>"000000111",
  20296=>"101001000",
  20297=>"000100101",
  20298=>"000101111",
  20299=>"011011001",
  20300=>"000000000",
  20301=>"000000000",
  20302=>"101111111",
  20303=>"110110000",
  20304=>"011111111",
  20305=>"001000010",
  20306=>"000000000",
  20307=>"000000000",
  20308=>"000000111",
  20309=>"011011011",
  20310=>"111101001",
  20311=>"111101101",
  20312=>"111101001",
  20313=>"000000001",
  20314=>"110111000",
  20315=>"001100000",
  20316=>"111001000",
  20317=>"001000101",
  20318=>"101011000",
  20319=>"011111000",
  20320=>"111111000",
  20321=>"111111001",
  20322=>"111110000",
  20323=>"100000111",
  20324=>"000001001",
  20325=>"011111010",
  20326=>"111111000",
  20327=>"001000110",
  20328=>"000000001",
  20329=>"100111110",
  20330=>"000101111",
  20331=>"001001111",
  20332=>"111111111",
  20333=>"000000100",
  20334=>"000100110",
  20335=>"000000000",
  20336=>"000000011",
  20337=>"101111110",
  20338=>"111101101",
  20339=>"100110110",
  20340=>"000111100",
  20341=>"000000110",
  20342=>"000000110",
  20343=>"000111100",
  20344=>"000000010",
  20345=>"111111000",
  20346=>"001000000",
  20347=>"000111110",
  20348=>"000110111",
  20349=>"000000000",
  20350=>"111000000",
  20351=>"000001011",
  20352=>"000111011",
  20353=>"001000000",
  20354=>"100000000",
  20355=>"010000000",
  20356=>"000000000",
  20357=>"000000000",
  20358=>"000000000",
  20359=>"000000111",
  20360=>"000000101",
  20361=>"000000111",
  20362=>"111111111",
  20363=>"111111000",
  20364=>"000110111",
  20365=>"101111110",
  20366=>"000100111",
  20367=>"000001010",
  20368=>"000001001",
  20369=>"110111111",
  20370=>"111111000",
  20371=>"111111101",
  20372=>"111111111",
  20373=>"000000000",
  20374=>"111111111",
  20375=>"011111000",
  20376=>"011110000",
  20377=>"101111111",
  20378=>"111111000",
  20379=>"101101101",
  20380=>"000100110",
  20381=>"000000010",
  20382=>"000011111",
  20383=>"000000010",
  20384=>"111111111",
  20385=>"111111001",
  20386=>"011011111",
  20387=>"000000000",
  20388=>"001111001",
  20389=>"111111010",
  20390=>"111111101",
  20391=>"110010011",
  20392=>"000001001",
  20393=>"000000011",
  20394=>"111011000",
  20395=>"000001001",
  20396=>"000000000",
  20397=>"111100000",
  20398=>"010110000",
  20399=>"000111111",
  20400=>"111111111",
  20401=>"000111111",
  20402=>"000000111",
  20403=>"011000000",
  20404=>"100101000",
  20405=>"000000100",
  20406=>"001101111",
  20407=>"100111110",
  20408=>"000110110",
  20409=>"000000000",
  20410=>"111000000",
  20411=>"111011001",
  20412=>"011111000",
  20413=>"000001111",
  20414=>"000000111",
  20415=>"100101111",
  20416=>"100000000",
  20417=>"000000111",
  20418=>"001111111",
  20419=>"000111111",
  20420=>"000000011",
  20421=>"000000111",
  20422=>"001110110",
  20423=>"000111111",
  20424=>"111111000",
  20425=>"110111111",
  20426=>"000000111",
  20427=>"000000000",
  20428=>"111000000",
  20429=>"001000110",
  20430=>"101100110",
  20431=>"111110111",
  20432=>"000000001",
  20433=>"000001011",
  20434=>"111111010",
  20435=>"111111111",
  20436=>"000000100",
  20437=>"100110110",
  20438=>"000000000",
  20439=>"000101111",
  20440=>"101101100",
  20441=>"111001000",
  20442=>"000000000",
  20443=>"011100011",
  20444=>"000000000",
  20445=>"101111111",
  20446=>"111010011",
  20447=>"000111111",
  20448=>"110111111",
  20449=>"000000000",
  20450=>"100011000",
  20451=>"001001111",
  20452=>"111111001",
  20453=>"111111111",
  20454=>"001000000",
  20455=>"100010000",
  20456=>"111100000",
  20457=>"111001000",
  20458=>"111111000",
  20459=>"000000100",
  20460=>"000000111",
  20461=>"000000110",
  20462=>"101101000",
  20463=>"000100111",
  20464=>"111111111",
  20465=>"000010110",
  20466=>"101100100",
  20467=>"000000111",
  20468=>"001111000",
  20469=>"111111000",
  20470=>"000100001",
  20471=>"100000001",
  20472=>"111111010",
  20473=>"110011000",
  20474=>"000000000",
  20475=>"111111110",
  20476=>"111110101",
  20477=>"011000000",
  20478=>"111101001",
  20479=>"000101101",
  20480=>"000111111",
  20481=>"000000000",
  20482=>"001001001",
  20483=>"000000111",
  20484=>"010000111",
  20485=>"001000000",
  20486=>"000000000",
  20487=>"110111111",
  20488=>"011000111",
  20489=>"000000000",
  20490=>"000111000",
  20491=>"111111111",
  20492=>"001000001",
  20493=>"111111000",
  20494=>"111111100",
  20495=>"100101001",
  20496=>"011111111",
  20497=>"111111011",
  20498=>"101001111",
  20499=>"000000111",
  20500=>"000111000",
  20501=>"111111111",
  20502=>"000000000",
  20503=>"000000000",
  20504=>"000000000",
  20505=>"011101101",
  20506=>"000001111",
  20507=>"100110000",
  20508=>"000111111",
  20509=>"001000111",
  20510=>"100001001",
  20511=>"111010000",
  20512=>"111111111",
  20513=>"111111111",
  20514=>"110110101",
  20515=>"111101100",
  20516=>"110001000",
  20517=>"000000000",
  20518=>"001011111",
  20519=>"111111100",
  20520=>"000101000",
  20521=>"000000000",
  20522=>"111111111",
  20523=>"111100111",
  20524=>"111111001",
  20525=>"000000111",
  20526=>"000001000",
  20527=>"111101111",
  20528=>"000000000",
  20529=>"001000001",
  20530=>"111111111",
  20531=>"100100100",
  20532=>"111111000",
  20533=>"000000001",
  20534=>"011111101",
  20535=>"100000000",
  20536=>"110110110",
  20537=>"111111111",
  20538=>"111111111",
  20539=>"000000000",
  20540=>"000000000",
  20541=>"000000000",
  20542=>"000000000",
  20543=>"000111110",
  20544=>"000011111",
  20545=>"000111001",
  20546=>"110000000",
  20547=>"011111001",
  20548=>"000000000",
  20549=>"111101101",
  20550=>"111111111",
  20551=>"111011011",
  20552=>"111111111",
  20553=>"000000001",
  20554=>"111111111",
  20555=>"111001000",
  20556=>"111111011",
  20557=>"000001101",
  20558=>"001111111",
  20559=>"110111110",
  20560=>"000000000",
  20561=>"100100000",
  20562=>"000000000",
  20563=>"111111111",
  20564=>"000000000",
  20565=>"111011000",
  20566=>"001000111",
  20567=>"000000000",
  20568=>"000001001",
  20569=>"000000000",
  20570=>"000000001",
  20571=>"001001001",
  20572=>"111000001",
  20573=>"111111000",
  20574=>"000000111",
  20575=>"101111010",
  20576=>"000100111",
  20577=>"110110010",
  20578=>"000000000",
  20579=>"000000000",
  20580=>"111111101",
  20581=>"111010010",
  20582=>"000000001",
  20583=>"101110110",
  20584=>"000001111",
  20585=>"111111111",
  20586=>"111111101",
  20587=>"100000000",
  20588=>"011000001",
  20589=>"111101101",
  20590=>"111000000",
  20591=>"111111111",
  20592=>"100100111",
  20593=>"000100011",
  20594=>"010010000",
  20595=>"000100110",
  20596=>"110010000",
  20597=>"111111001",
  20598=>"000000000",
  20599=>"111111111",
  20600=>"000000000",
  20601=>"000000000",
  20602=>"000111111",
  20603=>"111111111",
  20604=>"000001001",
  20605=>"000000000",
  20606=>"000010000",
  20607=>"111111111",
  20608=>"001001001",
  20609=>"010000111",
  20610=>"111111111",
  20611=>"111110110",
  20612=>"111111111",
  20613=>"111111111",
  20614=>"111111111",
  20615=>"111110000",
  20616=>"001000111",
  20617=>"000000000",
  20618=>"001001111",
  20619=>"000000111",
  20620=>"110011000",
  20621=>"111111111",
  20622=>"000000000",
  20623=>"010000000",
  20624=>"001011000",
  20625=>"000000000",
  20626=>"000000000",
  20627=>"100000000",
  20628=>"010111111",
  20629=>"111111111",
  20630=>"001001001",
  20631=>"000000000",
  20632=>"001011000",
  20633=>"111111111",
  20634=>"000000100",
  20635=>"000000000",
  20636=>"000000001",
  20637=>"011111111",
  20638=>"001111111",
  20639=>"111111111",
  20640=>"001110110",
  20641=>"100000010",
  20642=>"000011011",
  20643=>"001111101",
  20644=>"100100110",
  20645=>"000100000",
  20646=>"000000000",
  20647=>"111010111",
  20648=>"111111001",
  20649=>"000011111",
  20650=>"110111111",
  20651=>"000100101",
  20652=>"111111001",
  20653=>"000100000",
  20654=>"000011101",
  20655=>"000111111",
  20656=>"000000000",
  20657=>"111111110",
  20658=>"111001111",
  20659=>"000000000",
  20660=>"100000000",
  20661=>"111001001",
  20662=>"000000000",
  20663=>"000000000",
  20664=>"101111100",
  20665=>"101000001",
  20666=>"111111111",
  20667=>"000100100",
  20668=>"110100000",
  20669=>"111111101",
  20670=>"111111111",
  20671=>"111000000",
  20672=>"000000000",
  20673=>"000100111",
  20674=>"001001001",
  20675=>"000010000",
  20676=>"100000000",
  20677=>"000000000",
  20678=>"111111111",
  20679=>"000000000",
  20680=>"000111011",
  20681=>"000011011",
  20682=>"001000000",
  20683=>"101000000",
  20684=>"111011111",
  20685=>"111101111",
  20686=>"111111111",
  20687=>"000000011",
  20688=>"111001010",
  20689=>"111111011",
  20690=>"011001000",
  20691=>"000010110",
  20692=>"000000100",
  20693=>"000000110",
  20694=>"000000000",
  20695=>"010000000",
  20696=>"000000000",
  20697=>"010110100",
  20698=>"000000000",
  20699=>"111111111",
  20700=>"011111001",
  20701=>"000011111",
  20702=>"000100110",
  20703=>"000000000",
  20704=>"110111111",
  20705=>"001010010",
  20706=>"000000000",
  20707=>"001100000",
  20708=>"010000000",
  20709=>"000100100",
  20710=>"111111111",
  20711=>"010111111",
  20712=>"000000111",
  20713=>"000000000",
  20714=>"000000100",
  20715=>"011111011",
  20716=>"111111111",
  20717=>"000011111",
  20718=>"000000111",
  20719=>"011000000",
  20720=>"010011001",
  20721=>"111111111",
  20722=>"000000000",
  20723=>"000000101",
  20724=>"111111000",
  20725=>"111111011",
  20726=>"011100111",
  20727=>"100000000",
  20728=>"000000001",
  20729=>"000000000",
  20730=>"010111110",
  20731=>"001001001",
  20732=>"001001111",
  20733=>"110110000",
  20734=>"000000000",
  20735=>"011100111",
  20736=>"110111111",
  20737=>"011011000",
  20738=>"111000000",
  20739=>"111111111",
  20740=>"110100000",
  20741=>"010000000",
  20742=>"110000000",
  20743=>"000100100",
  20744=>"001111111",
  20745=>"000000000",
  20746=>"000000000",
  20747=>"000111111",
  20748=>"111111111",
  20749=>"011111110",
  20750=>"111111111",
  20751=>"110110111",
  20752=>"110111111",
  20753=>"000000000",
  20754=>"111001000",
  20755=>"000000000",
  20756=>"011010000",
  20757=>"110111111",
  20758=>"011011011",
  20759=>"000000000",
  20760=>"001010110",
  20761=>"111111000",
  20762=>"010111111",
  20763=>"110000101",
  20764=>"111111111",
  20765=>"000111111",
  20766=>"000000000",
  20767=>"000111111",
  20768=>"110110100",
  20769=>"011111111",
  20770=>"100111111",
  20771=>"111111111",
  20772=>"111111000",
  20773=>"010110000",
  20774=>"110111111",
  20775=>"010000000",
  20776=>"000000000",
  20777=>"111111111",
  20778=>"011111000",
  20779=>"000000000",
  20780=>"111111111",
  20781=>"001001000",
  20782=>"000111000",
  20783=>"111111111",
  20784=>"110110000",
  20785=>"111111111",
  20786=>"111111010",
  20787=>"110110000",
  20788=>"000000000",
  20789=>"111101110",
  20790=>"000010110",
  20791=>"111111111",
  20792=>"000000000",
  20793=>"100000000",
  20794=>"111111111",
  20795=>"000000010",
  20796=>"001011011",
  20797=>"001111111",
  20798=>"111111111",
  20799=>"111110111",
  20800=>"111111111",
  20801=>"111111111",
  20802=>"000000000",
  20803=>"111111110",
  20804=>"111111000",
  20805=>"000111010",
  20806=>"111000001",
  20807=>"010000000",
  20808=>"000000000",
  20809=>"000111111",
  20810=>"000111000",
  20811=>"110110100",
  20812=>"111111111",
  20813=>"000001000",
  20814=>"001000001",
  20815=>"111011001",
  20816=>"011001011",
  20817=>"000001011",
  20818=>"111111111",
  20819=>"000000000",
  20820=>"000011111",
  20821=>"011011000",
  20822=>"000000000",
  20823=>"000001111",
  20824=>"111111011",
  20825=>"000000000",
  20826=>"000000001",
  20827=>"000100011",
  20828=>"001111010",
  20829=>"111111101",
  20830=>"000000110",
  20831=>"111111000",
  20832=>"000010000",
  20833=>"000000000",
  20834=>"011011111",
  20835=>"111111111",
  20836=>"110010000",
  20837=>"000000000",
  20838=>"000000000",
  20839=>"000111111",
  20840=>"011001001",
  20841=>"000010011",
  20842=>"111111111",
  20843=>"111101101",
  20844=>"000110111",
  20845=>"000100111",
  20846=>"010111011",
  20847=>"000000100",
  20848=>"000000000",
  20849=>"000000000",
  20850=>"001001011",
  20851=>"000000000",
  20852=>"000101111",
  20853=>"000110011",
  20854=>"000010111",
  20855=>"000000000",
  20856=>"101001111",
  20857=>"000000000",
  20858=>"111111111",
  20859=>"000010000",
  20860=>"111111111",
  20861=>"111111111",
  20862=>"110110110",
  20863=>"000000101",
  20864=>"111111011",
  20865=>"111111111",
  20866=>"101101101",
  20867=>"110110111",
  20868=>"000000111",
  20869=>"000101111",
  20870=>"111110000",
  20871=>"000100110",
  20872=>"000000000",
  20873=>"011000000",
  20874=>"000000111",
  20875=>"000000111",
  20876=>"000001111",
  20877=>"010110100",
  20878=>"000000100",
  20879=>"010000000",
  20880=>"000000000",
  20881=>"000000000",
  20882=>"110000110",
  20883=>"100100000",
  20884=>"111111111",
  20885=>"000000111",
  20886=>"000000001",
  20887=>"000001011",
  20888=>"111111111",
  20889=>"111111111",
  20890=>"111111111",
  20891=>"001111111",
  20892=>"011000011",
  20893=>"000100000",
  20894=>"111011001",
  20895=>"100110110",
  20896=>"111101001",
  20897=>"011011000",
  20898=>"011111111",
  20899=>"000000001",
  20900=>"001111111",
  20901=>"000000000",
  20902=>"100111110",
  20903=>"111111111",
  20904=>"000001001",
  20905=>"011111110",
  20906=>"111111011",
  20907=>"000011111",
  20908=>"000000000",
  20909=>"001111111",
  20910=>"001111111",
  20911=>"000000000",
  20912=>"110000000",
  20913=>"000000000",
  20914=>"000000000",
  20915=>"111111111",
  20916=>"000000000",
  20917=>"000000000",
  20918=>"000000001",
  20919=>"000000000",
  20920=>"000001111",
  20921=>"111111110",
  20922=>"001101111",
  20923=>"111111111",
  20924=>"111111111",
  20925=>"000000000",
  20926=>"111110111",
  20927=>"010000100",
  20928=>"000000000",
  20929=>"001000001",
  20930=>"111111000",
  20931=>"000000000",
  20932=>"000111000",
  20933=>"001111111",
  20934=>"011110100",
  20935=>"000000111",
  20936=>"000000000",
  20937=>"010000000",
  20938=>"000000001",
  20939=>"111111000",
  20940=>"000000000",
  20941=>"000000000",
  20942=>"100110000",
  20943=>"011000000",
  20944=>"111111111",
  20945=>"001001111",
  20946=>"111101000",
  20947=>"111111000",
  20948=>"111100100",
  20949=>"111001111",
  20950=>"000111111",
  20951=>"100100101",
  20952=>"000000000",
  20953=>"000000000",
  20954=>"001001001",
  20955=>"010111111",
  20956=>"000000000",
  20957=>"001011001",
  20958=>"000000000",
  20959=>"001101101",
  20960=>"100000000",
  20961=>"111111110",
  20962=>"110110110",
  20963=>"111011001",
  20964=>"100111111",
  20965=>"011001000",
  20966=>"111111111",
  20967=>"000000000",
  20968=>"001011001",
  20969=>"111111011",
  20970=>"000000011",
  20971=>"000011000",
  20972=>"000110000",
  20973=>"000000111",
  20974=>"111111000",
  20975=>"000000000",
  20976=>"000000000",
  20977=>"000000000",
  20978=>"000000010",
  20979=>"000000000",
  20980=>"000000000",
  20981=>"001001000",
  20982=>"011000000",
  20983=>"011010100",
  20984=>"000000001",
  20985=>"000000001",
  20986=>"111000000",
  20987=>"100100100",
  20988=>"011100111",
  20989=>"000000111",
  20990=>"001001000",
  20991=>"000010000",
  20992=>"111111111",
  20993=>"110100111",
  20994=>"111101111",
  20995=>"111111111",
  20996=>"111111111",
  20997=>"111100100",
  20998=>"000000000",
  20999=>"111111111",
  21000=>"100111111",
  21001=>"100100101",
  21002=>"111111111",
  21003=>"110111111",
  21004=>"100110110",
  21005=>"000000111",
  21006=>"001011010",
  21007=>"000000000",
  21008=>"000110000",
  21009=>"000101001",
  21010=>"000011001",
  21011=>"111111111",
  21012=>"000000111",
  21013=>"000111111",
  21014=>"000000000",
  21015=>"000000000",
  21016=>"000000000",
  21017=>"111001111",
  21018=>"111111111",
  21019=>"111110110",
  21020=>"111111111",
  21021=>"111110111",
  21022=>"000000000",
  21023=>"000000000",
  21024=>"111101000",
  21025=>"000000000",
  21026=>"111111111",
  21027=>"011000000",
  21028=>"000000101",
  21029=>"000110110",
  21030=>"111111010",
  21031=>"000000000",
  21032=>"001001001",
  21033=>"000000000",
  21034=>"111111111",
  21035=>"000000000",
  21036=>"001000000",
  21037=>"000000000",
  21038=>"111111000",
  21039=>"111111111",
  21040=>"111000000",
  21041=>"111100010",
  21042=>"000000000",
  21043=>"111101000",
  21044=>"000000000",
  21045=>"111111111",
  21046=>"000000000",
  21047=>"000000000",
  21048=>"000000111",
  21049=>"111000000",
  21050=>"010111111",
  21051=>"111000000",
  21052=>"000000000",
  21053=>"111111111",
  21054=>"000010010",
  21055=>"111111111",
  21056=>"111001100",
  21057=>"111111111",
  21058=>"000000001",
  21059=>"000000000",
  21060=>"000000000",
  21061=>"000000000",
  21062=>"111111111",
  21063=>"000000000",
  21064=>"000001001",
  21065=>"110000000",
  21066=>"111110000",
  21067=>"000000000",
  21068=>"101000000",
  21069=>"101101001",
  21070=>"000111111",
  21071=>"111111110",
  21072=>"110000000",
  21073=>"001000001",
  21074=>"010110110",
  21075=>"111001000",
  21076=>"001001111",
  21077=>"000000000",
  21078=>"111111110",
  21079=>"000000000",
  21080=>"000000000",
  21081=>"101000000",
  21082=>"111111111",
  21083=>"001001001",
  21084=>"111111111",
  21085=>"111111011",
  21086=>"111111011",
  21087=>"111111111",
  21088=>"100000000",
  21089=>"101101101",
  21090=>"011011011",
  21091=>"111111111",
  21092=>"000000000",
  21093=>"111101101",
  21094=>"110110111",
  21095=>"111111111",
  21096=>"000000001",
  21097=>"111111111",
  21098=>"000000000",
  21099=>"111111111",
  21100=>"000001000",
  21101=>"100000000",
  21102=>"111000100",
  21103=>"110110000",
  21104=>"000000111",
  21105=>"111111111",
  21106=>"000000000",
  21107=>"111111110",
  21108=>"111111111",
  21109=>"000000000",
  21110=>"110110111",
  21111=>"000000101",
  21112=>"100000000",
  21113=>"111100101",
  21114=>"111000000",
  21115=>"111111111",
  21116=>"000000000",
  21117=>"000000000",
  21118=>"001001111",
  21119=>"000000000",
  21120=>"000111111",
  21121=>"000000000",
  21122=>"000000000",
  21123=>"101000011",
  21124=>"111001001",
  21125=>"100111111",
  21126=>"111111110",
  21127=>"111111011",
  21128=>"000000000",
  21129=>"011111111",
  21130=>"111111111",
  21131=>"111111111",
  21132=>"000000111",
  21133=>"010010000",
  21134=>"111111111",
  21135=>"111111111",
  21136=>"011011111",
  21137=>"001101111",
  21138=>"100000000",
  21139=>"000000000",
  21140=>"111011010",
  21141=>"010111111",
  21142=>"011000000",
  21143=>"111011000",
  21144=>"011011000",
  21145=>"000000010",
  21146=>"110100101",
  21147=>"111000100",
  21148=>"000000000",
  21149=>"100000111",
  21150=>"000100111",
  21151=>"000000000",
  21152=>"000000000",
  21153=>"000011001",
  21154=>"111111111",
  21155=>"010000101",
  21156=>"001011001",
  21157=>"111111111",
  21158=>"000000000",
  21159=>"111000000",
  21160=>"000000000",
  21161=>"111111111",
  21162=>"111110111",
  21163=>"111111111",
  21164=>"111001000",
  21165=>"101001101",
  21166=>"111111111",
  21167=>"111111111",
  21168=>"000110000",
  21169=>"111111111",
  21170=>"111111111",
  21171=>"000000000",
  21172=>"000010111",
  21173=>"000010110",
  21174=>"000111010",
  21175=>"000000000",
  21176=>"000100110",
  21177=>"111111111",
  21178=>"011011000",
  21179=>"000000000",
  21180=>"111111000",
  21181=>"111001011",
  21182=>"111111000",
  21183=>"000000000",
  21184=>"011010111",
  21185=>"111000011",
  21186=>"111000111",
  21187=>"000000000",
  21188=>"011011010",
  21189=>"011000000",
  21190=>"001000000",
  21191=>"100000000",
  21192=>"000011111",
  21193=>"111101111",
  21194=>"111111111",
  21195=>"000010111",
  21196=>"010011011",
  21197=>"000111000",
  21198=>"000000000",
  21199=>"000000000",
  21200=>"111111111",
  21201=>"001011111",
  21202=>"000000000",
  21203=>"111100111",
  21204=>"111111000",
  21205=>"001111100",
  21206=>"000000000",
  21207=>"000000000",
  21208=>"000000000",
  21209=>"100110110",
  21210=>"000000000",
  21211=>"000000111",
  21212=>"000000010",
  21213=>"101111111",
  21214=>"000001111",
  21215=>"010000110",
  21216=>"111111111",
  21217=>"000010000",
  21218=>"000000000",
  21219=>"111111000",
  21220=>"111111111",
  21221=>"000111111",
  21222=>"000000000",
  21223=>"001011111",
  21224=>"111110000",
  21225=>"100101111",
  21226=>"010011011",
  21227=>"000000111",
  21228=>"111111111",
  21229=>"000000000",
  21230=>"000000111",
  21231=>"000000000",
  21232=>"111111111",
  21233=>"000000011",
  21234=>"000000000",
  21235=>"011111000",
  21236=>"000011000",
  21237=>"111111110",
  21238=>"001000000",
  21239=>"000011000",
  21240=>"000000000",
  21241=>"000000000",
  21242=>"000000000",
  21243=>"101111111",
  21244=>"000100110",
  21245=>"111111111",
  21246=>"111101101",
  21247=>"110111111",
  21248=>"000000000",
  21249=>"010000100",
  21250=>"000000000",
  21251=>"100111110",
  21252=>"111111111",
  21253=>"001111111",
  21254=>"111110111",
  21255=>"000000000",
  21256=>"110111111",
  21257=>"111111111",
  21258=>"000000000",
  21259=>"011000000",
  21260=>"001001111",
  21261=>"111011000",
  21262=>"000010000",
  21263=>"111111001",
  21264=>"111111111",
  21265=>"000011111",
  21266=>"111111111",
  21267=>"011111111",
  21268=>"010000000",
  21269=>"000000110",
  21270=>"000100110",
  21271=>"001000000",
  21272=>"111000000",
  21273=>"111111111",
  21274=>"111011111",
  21275=>"000000100",
  21276=>"111111111",
  21277=>"000000000",
  21278=>"001111111",
  21279=>"111111111",
  21280=>"000000000",
  21281=>"111001000",
  21282=>"000111111",
  21283=>"000001000",
  21284=>"000000100",
  21285=>"000000000",
  21286=>"011011001",
  21287=>"100111111",
  21288=>"111111111",
  21289=>"000000000",
  21290=>"111111111",
  21291=>"000000111",
  21292=>"001001111",
  21293=>"100001001",
  21294=>"000000000",
  21295=>"011011000",
  21296=>"001001111",
  21297=>"000000000",
  21298=>"100000000",
  21299=>"000010000",
  21300=>"000000000",
  21301=>"000000001",
  21302=>"000101000",
  21303=>"000011010",
  21304=>"000000000",
  21305=>"000000100",
  21306=>"000011111",
  21307=>"111111111",
  21308=>"000000000",
  21309=>"000000000",
  21310=>"000000100",
  21311=>"000000000",
  21312=>"111100000",
  21313=>"111111110",
  21314=>"101111101",
  21315=>"000000000",
  21316=>"000000000",
  21317=>"000000000",
  21318=>"000010110",
  21319=>"111111111",
  21320=>"110100110",
  21321=>"111110110",
  21322=>"111110100",
  21323=>"100100110",
  21324=>"111011000",
  21325=>"000000000",
  21326=>"011000000",
  21327=>"001001000",
  21328=>"000000001",
  21329=>"101001001",
  21330=>"000000000",
  21331=>"111010011",
  21332=>"111101001",
  21333=>"011011011",
  21334=>"000000000",
  21335=>"111000111",
  21336=>"110110011",
  21337=>"111111111",
  21338=>"000000000",
  21339=>"111000000",
  21340=>"000000000",
  21341=>"000000000",
  21342=>"100011011",
  21343=>"110110110",
  21344=>"000010010",
  21345=>"111111111",
  21346=>"000001001",
  21347=>"000001011",
  21348=>"000000000",
  21349=>"010010000",
  21350=>"001001000",
  21351=>"000000000",
  21352=>"001001001",
  21353=>"000000000",
  21354=>"111000000",
  21355=>"111111000",
  21356=>"000010111",
  21357=>"111110000",
  21358=>"110111110",
  21359=>"111010010",
  21360=>"000000101",
  21361=>"000100100",
  21362=>"000111111",
  21363=>"000000000",
  21364=>"000100000",
  21365=>"100111111",
  21366=>"111111111",
  21367=>"000000000",
  21368=>"111000000",
  21369=>"000000000",
  21370=>"111101111",
  21371=>"001001000",
  21372=>"110100111",
  21373=>"111111111",
  21374=>"000000000",
  21375=>"000000000",
  21376=>"000000000",
  21377=>"001001100",
  21378=>"000000000",
  21379=>"111111111",
  21380=>"100101000",
  21381=>"000010110",
  21382=>"000000000",
  21383=>"000000000",
  21384=>"111111111",
  21385=>"000001000",
  21386=>"111111111",
  21387=>"111111111",
  21388=>"111111111",
  21389=>"000000000",
  21390=>"000000111",
  21391=>"010010110",
  21392=>"000000000",
  21393=>"000000000",
  21394=>"000000000",
  21395=>"000000000",
  21396=>"001000000",
  21397=>"000000000",
  21398=>"111111011",
  21399=>"100111000",
  21400=>"000000000",
  21401=>"111111001",
  21402=>"000000000",
  21403=>"111111100",
  21404=>"000000101",
  21405=>"000000000",
  21406=>"000110000",
  21407=>"000000111",
  21408=>"100111011",
  21409=>"110100101",
  21410=>"111000000",
  21411=>"111111111",
  21412=>"011111111",
  21413=>"111111111",
  21414=>"001111111",
  21415=>"110110100",
  21416=>"000000000",
  21417=>"000000000",
  21418=>"011011001",
  21419=>"000010011",
  21420=>"111010000",
  21421=>"111111111",
  21422=>"001001111",
  21423=>"000000111",
  21424=>"111000011",
  21425=>"000001001",
  21426=>"111000000",
  21427=>"000110110",
  21428=>"000000000",
  21429=>"011000000",
  21430=>"011111111",
  21431=>"010000011",
  21432=>"111000000",
  21433=>"100100000",
  21434=>"010110110",
  21435=>"100111111",
  21436=>"000001111",
  21437=>"000011011",
  21438=>"000000000",
  21439=>"010000000",
  21440=>"110111110",
  21441=>"111111111",
  21442=>"000001000",
  21443=>"000000000",
  21444=>"111111111",
  21445=>"100111111",
  21446=>"100110000",
  21447=>"000000111",
  21448=>"011011000",
  21449=>"111100110",
  21450=>"000000000",
  21451=>"111111000",
  21452=>"000000000",
  21453=>"000000111",
  21454=>"111000000",
  21455=>"111111111",
  21456=>"000111011",
  21457=>"000001001",
  21458=>"000000100",
  21459=>"111111011",
  21460=>"000000001",
  21461=>"111011000",
  21462=>"000100101",
  21463=>"000000110",
  21464=>"111111111",
  21465=>"110000000",
  21466=>"011000011",
  21467=>"010111111",
  21468=>"000000000",
  21469=>"000000000",
  21470=>"000000000",
  21471=>"111111111",
  21472=>"111111100",
  21473=>"000000001",
  21474=>"000000010",
  21475=>"111111111",
  21476=>"011000000",
  21477=>"111111111",
  21478=>"111111111",
  21479=>"000000000",
  21480=>"001011111",
  21481=>"000000000",
  21482=>"011111111",
  21483=>"111111110",
  21484=>"000000110",
  21485=>"000000000",
  21486=>"101101011",
  21487=>"010000000",
  21488=>"000111111",
  21489=>"000000000",
  21490=>"111111111",
  21491=>"110000011",
  21492=>"010011011",
  21493=>"000000000",
  21494=>"000000000",
  21495=>"000000111",
  21496=>"000000000",
  21497=>"000001011",
  21498=>"000000010",
  21499=>"100000001",
  21500=>"000000000",
  21501=>"000000100",
  21502=>"111011111",
  21503=>"111111111",
  21504=>"111111100",
  21505=>"100111111",
  21506=>"111111000",
  21507=>"011111111",
  21508=>"110111111",
  21509=>"010011000",
  21510=>"111111000",
  21511=>"000111011",
  21512=>"000000000",
  21513=>"000000111",
  21514=>"110110010",
  21515=>"111011001",
  21516=>"111100100",
  21517=>"010111111",
  21518=>"000000000",
  21519=>"000000000",
  21520=>"000110111",
  21521=>"111000000",
  21522=>"010000000",
  21523=>"111000000",
  21524=>"100000000",
  21525=>"000000001",
  21526=>"010010111",
  21527=>"000010100",
  21528=>"010011001",
  21529=>"100111111",
  21530=>"111111111",
  21531=>"110110011",
  21532=>"111100111",
  21533=>"001111111",
  21534=>"111011011",
  21535=>"000010111",
  21536=>"010111000",
  21537=>"111111111",
  21538=>"010001001",
  21539=>"100111000",
  21540=>"011111111",
  21541=>"000001000",
  21542=>"110011111",
  21543=>"111110101",
  21544=>"001000100",
  21545=>"111000000",
  21546=>"111111111",
  21547=>"111011000",
  21548=>"111111001",
  21549=>"010111011",
  21550=>"000000101",
  21551=>"111000000",
  21552=>"001111111",
  21553=>"000001101",
  21554=>"110111111",
  21555=>"000000111",
  21556=>"000011111",
  21557=>"111100100",
  21558=>"000000000",
  21559=>"111000100",
  21560=>"111111000",
  21561=>"000000000",
  21562=>"000111100",
  21563=>"000000000",
  21564=>"101000000",
  21565=>"011010010",
  21566=>"010110000",
  21567=>"000000000",
  21568=>"100000000",
  21569=>"000100001",
  21570=>"100110011",
  21571=>"111110100",
  21572=>"110100110",
  21573=>"001011111",
  21574=>"110000000",
  21575=>"111111111",
  21576=>"001111111",
  21577=>"000110111",
  21578=>"000111111",
  21579=>"111110110",
  21580=>"100000000",
  21581=>"000000111",
  21582=>"111101000",
  21583=>"000000111",
  21584=>"000000000",
  21585=>"000001111",
  21586=>"111111100",
  21587=>"110100111",
  21588=>"100101111",
  21589=>"111101000",
  21590=>"111111111",
  21591=>"000000000",
  21592=>"000000111",
  21593=>"000000100",
  21594=>"000000000",
  21595=>"000000000",
  21596=>"111110000",
  21597=>"000111111",
  21598=>"110111111",
  21599=>"110100000",
  21600=>"010000000",
  21601=>"001001101",
  21602=>"111111010",
  21603=>"111111000",
  21604=>"000111101",
  21605=>"101001001",
  21606=>"000000000",
  21607=>"110011011",
  21608=>"111010011",
  21609=>"110000110",
  21610=>"110000111",
  21611=>"000000101",
  21612=>"110000001",
  21613=>"111000000",
  21614=>"000000111",
  21615=>"111111111",
  21616=>"111111101",
  21617=>"000100111",
  21618=>"001001001",
  21619=>"100010000",
  21620=>"111111111",
  21621=>"111111000",
  21622=>"000000000",
  21623=>"111111111",
  21624=>"000000000",
  21625=>"000111111",
  21626=>"111000000",
  21627=>"000000001",
  21628=>"100000001",
  21629=>"111111111",
  21630=>"111111110",
  21631=>"000011000",
  21632=>"111101100",
  21633=>"000000111",
  21634=>"111111111",
  21635=>"100111111",
  21636=>"110110111",
  21637=>"000000000",
  21638=>"110011001",
  21639=>"111111001",
  21640=>"000000111",
  21641=>"111110111",
  21642=>"111111111",
  21643=>"111111111",
  21644=>"001000111",
  21645=>"000000000",
  21646=>"011001000",
  21647=>"111101000",
  21648=>"000000000",
  21649=>"000000000",
  21650=>"000111111",
  21651=>"111111001",
  21652=>"001000011",
  21653=>"000111000",
  21654=>"000010010",
  21655=>"001001000",
  21656=>"111010000",
  21657=>"011111111",
  21658=>"111111011",
  21659=>"000000000",
  21660=>"010111111",
  21661=>"000010000",
  21662=>"111000000",
  21663=>"010010001",
  21664=>"011001000",
  21665=>"000001000",
  21666=>"111111000",
  21667=>"111000000",
  21668=>"111011010",
  21669=>"111111111",
  21670=>"000000000",
  21671=>"000000100",
  21672=>"100000000",
  21673=>"111000000",
  21674=>"101111111",
  21675=>"000011000",
  21676=>"000000111",
  21677=>"011011011",
  21678=>"100000100",
  21679=>"000110101",
  21680=>"111000000",
  21681=>"001100110",
  21682=>"111111010",
  21683=>"000000000",
  21684=>"001111011",
  21685=>"000000000",
  21686=>"000000000",
  21687=>"000011111",
  21688=>"111111001",
  21689=>"111111011",
  21690=>"100100110",
  21691=>"110000000",
  21692=>"000110111",
  21693=>"110100000",
  21694=>"110110001",
  21695=>"110110110",
  21696=>"000110010",
  21697=>"000000000",
  21698=>"110111111",
  21699=>"000000000",
  21700=>"101111000",
  21701=>"000000000",
  21702=>"111000001",
  21703=>"111100000",
  21704=>"111111111",
  21705=>"001001000",
  21706=>"000111010",
  21707=>"011111001",
  21708=>"000111111",
  21709=>"110100000",
  21710=>"000010011",
  21711=>"111100111",
  21712=>"100000000",
  21713=>"111111000",
  21714=>"110111000",
  21715=>"000010000",
  21716=>"111111111",
  21717=>"001001111",
  21718=>"111000000",
  21719=>"110111111",
  21720=>"000000000",
  21721=>"111111111",
  21722=>"000000100",
  21723=>"111001111",
  21724=>"010110101",
  21725=>"100111111",
  21726=>"000000001",
  21727=>"010010111",
  21728=>"000000000",
  21729=>"100111010",
  21730=>"000000000",
  21731=>"111000000",
  21732=>"111111111",
  21733=>"000000000",
  21734=>"111110010",
  21735=>"111111011",
  21736=>"000000000",
  21737=>"111111100",
  21738=>"000000101",
  21739=>"000100111",
  21740=>"110110000",
  21741=>"100000000",
  21742=>"111100000",
  21743=>"000000000",
  21744=>"111101111",
  21745=>"111000100",
  21746=>"000000000",
  21747=>"111001001",
  21748=>"000000000",
  21749=>"001011000",
  21750=>"000000110",
  21751=>"000011011",
  21752=>"111000000",
  21753=>"111111000",
  21754=>"110000111",
  21755=>"110111000",
  21756=>"000000100",
  21757=>"001000000",
  21758=>"011000111",
  21759=>"010010000",
  21760=>"111101111",
  21761=>"111111000",
  21762=>"111111000",
  21763=>"000000100",
  21764=>"100000000",
  21765=>"111011000",
  21766=>"111111111",
  21767=>"110111010",
  21768=>"111101011",
  21769=>"000100100",
  21770=>"011011011",
  21771=>"111111111",
  21772=>"000000110",
  21773=>"000000111",
  21774=>"100100111",
  21775=>"110110100",
  21776=>"000000110",
  21777=>"000000111",
  21778=>"000111111",
  21779=>"110011111",
  21780=>"000000000",
  21781=>"101111111",
  21782=>"111011111",
  21783=>"111111111",
  21784=>"111111111",
  21785=>"110111111",
  21786=>"000000000",
  21787=>"000000000",
  21788=>"000100111",
  21789=>"000000000",
  21790=>"010111111",
  21791=>"000000000",
  21792=>"111111111",
  21793=>"000001111",
  21794=>"100111111",
  21795=>"011000000",
  21796=>"001001001",
  21797=>"101100111",
  21798=>"001111111",
  21799=>"101000011",
  21800=>"011111111",
  21801=>"111111111",
  21802=>"000000111",
  21803=>"100100100",
  21804=>"100101001",
  21805=>"000000111",
  21806=>"000000000",
  21807=>"011000000",
  21808=>"001111000",
  21809=>"111000000",
  21810=>"001000000",
  21811=>"111111000",
  21812=>"010100000",
  21813=>"111111101",
  21814=>"100000000",
  21815=>"100110000",
  21816=>"111111111",
  21817=>"111100000",
  21818=>"111010110",
  21819=>"111110000",
  21820=>"111111001",
  21821=>"110010111",
  21822=>"000101111",
  21823=>"000000010",
  21824=>"101111101",
  21825=>"111100110",
  21826=>"110011000",
  21827=>"000000110",
  21828=>"001111111",
  21829=>"000110111",
  21830=>"111101000",
  21831=>"111111000",
  21832=>"111111111",
  21833=>"000000000",
  21834=>"011000101",
  21835=>"100111111",
  21836=>"000000000",
  21837=>"000000111",
  21838=>"111111110",
  21839=>"000100111",
  21840=>"100000000",
  21841=>"000000001",
  21842=>"110111111",
  21843=>"111111110",
  21844=>"000000000",
  21845=>"011111111",
  21846=>"111110111",
  21847=>"110100100",
  21848=>"110110111",
  21849=>"001001000",
  21850=>"000111110",
  21851=>"000000000",
  21852=>"000000000",
  21853=>"000000000",
  21854=>"100100000",
  21855=>"001000111",
  21856=>"111111111",
  21857=>"110111111",
  21858=>"111100100",
  21859=>"111000000",
  21860=>"000000000",
  21861=>"011111111",
  21862=>"111000000",
  21863=>"000011000",
  21864=>"001011001",
  21865=>"111001000",
  21866=>"111111111",
  21867=>"000001101",
  21868=>"000010111",
  21869=>"110100100",
  21870=>"000000111",
  21871=>"100000100",
  21872=>"111111001",
  21873=>"010111111",
  21874=>"000000000",
  21875=>"111111100",
  21876=>"001000101",
  21877=>"110100100",
  21878=>"000000000",
  21879=>"000000000",
  21880=>"111011000",
  21881=>"111001001",
  21882=>"001001001",
  21883=>"011111111",
  21884=>"111001000",
  21885=>"000000011",
  21886=>"111000000",
  21887=>"111101000",
  21888=>"110111111",
  21889=>"000000000",
  21890=>"100100111",
  21891=>"000000000",
  21892=>"000000000",
  21893=>"000000000",
  21894=>"110111001",
  21895=>"010011100",
  21896=>"111111000",
  21897=>"000010011",
  21898=>"000111001",
  21899=>"000000000",
  21900=>"000110111",
  21901=>"011011111",
  21902=>"011010111",
  21903=>"000111111",
  21904=>"000000111",
  21905=>"000100100",
  21906=>"000110100",
  21907=>"011111111",
  21908=>"110100000",
  21909=>"011011001",
  21910=>"000000000",
  21911=>"111110100",
  21912=>"111111111",
  21913=>"111111001",
  21914=>"111000000",
  21915=>"111101111",
  21916=>"001111111",
  21917=>"111111000",
  21918=>"111010110",
  21919=>"111111111",
  21920=>"111110010",
  21921=>"000010100",
  21922=>"100000111",
  21923=>"110000100",
  21924=>"111000110",
  21925=>"000111000",
  21926=>"000000000",
  21927=>"000000000",
  21928=>"011111111",
  21929=>"100100101",
  21930=>"000000000",
  21931=>"101111110",
  21932=>"001111011",
  21933=>"000000000",
  21934=>"111000001",
  21935=>"111111111",
  21936=>"110111000",
  21937=>"111111111",
  21938=>"110000001",
  21939=>"011111000",
  21940=>"011000000",
  21941=>"111111000",
  21942=>"100110111",
  21943=>"101000000",
  21944=>"000000000",
  21945=>"100111111",
  21946=>"011000000",
  21947=>"000010111",
  21948=>"011111111",
  21949=>"000011111",
  21950=>"010100100",
  21951=>"100000110",
  21952=>"000111000",
  21953=>"000000000",
  21954=>"011111000",
  21955=>"111111000",
  21956=>"100110111",
  21957=>"111100101",
  21958=>"100000011",
  21959=>"110010000",
  21960=>"111000000",
  21961=>"100000000",
  21962=>"100000000",
  21963=>"011011000",
  21964=>"000111011",
  21965=>"111110111",
  21966=>"111100100",
  21967=>"111111111",
  21968=>"111100000",
  21969=>"010010010",
  21970=>"000000000",
  21971=>"000001111",
  21972=>"011011011",
  21973=>"000000000",
  21974=>"000011000",
  21975=>"011001111",
  21976=>"000000111",
  21977=>"000000011",
  21978=>"000111111",
  21979=>"111000100",
  21980=>"011011001",
  21981=>"110111111",
  21982=>"000011000",
  21983=>"110110110",
  21984=>"111111001",
  21985=>"111011000",
  21986=>"000000110",
  21987=>"111111110",
  21988=>"100000101",
  21989=>"000100111",
  21990=>"000000000",
  21991=>"000000000",
  21992=>"011000001",
  21993=>"000111111",
  21994=>"111000111",
  21995=>"100000000",
  21996=>"001010010",
  21997=>"111110111",
  21998=>"000000000",
  21999=>"111001000",
  22000=>"111111111",
  22001=>"000000111",
  22002=>"111001111",
  22003=>"111110000",
  22004=>"111000000",
  22005=>"111000000",
  22006=>"100100000",
  22007=>"111111111",
  22008=>"111111001",
  22009=>"000000100",
  22010=>"000000000",
  22011=>"000000001",
  22012=>"000000000",
  22013=>"001001000",
  22014=>"110000000",
  22015=>"000000001",
  22016=>"100000000",
  22017=>"000000000",
  22018=>"100111111",
  22019=>"111111001",
  22020=>"001001000",
  22021=>"110100100",
  22022=>"011111111",
  22023=>"111111111",
  22024=>"111101111",
  22025=>"111101001",
  22026=>"100000111",
  22027=>"001001101",
  22028=>"111100110",
  22029=>"110110000",
  22030=>"110111101",
  22031=>"111100000",
  22032=>"110110110",
  22033=>"111111111",
  22034=>"110110111",
  22035=>"111111100",
  22036=>"010000000",
  22037=>"110111110",
  22038=>"111010010",
  22039=>"001000010",
  22040=>"100110111",
  22041=>"000000000",
  22042=>"000001000",
  22043=>"001111110",
  22044=>"111111111",
  22045=>"111100111",
  22046=>"011000000",
  22047=>"101111111",
  22048=>"111110111",
  22049=>"011001001",
  22050=>"000100111",
  22051=>"100111111",
  22052=>"001111000",
  22053=>"000000000",
  22054=>"111110110",
  22055=>"000111001",
  22056=>"111111111",
  22057=>"000000000",
  22058=>"011111111",
  22059=>"000111011",
  22060=>"001110100",
  22061=>"000000000",
  22062=>"000010011",
  22063=>"000000011",
  22064=>"111000000",
  22065=>"111111111",
  22066=>"001101111",
  22067=>"001111111",
  22068=>"000000000",
  22069=>"001001111",
  22070=>"000000000",
  22071=>"001011001",
  22072=>"000000111",
  22073=>"000000000",
  22074=>"000000001",
  22075=>"000000110",
  22076=>"000000111",
  22077=>"010111111",
  22078=>"000000001",
  22079=>"000101111",
  22080=>"110010000",
  22081=>"010111111",
  22082=>"111110111",
  22083=>"111111111",
  22084=>"001101100",
  22085=>"001001000",
  22086=>"000000100",
  22087=>"000000000",
  22088=>"001001011",
  22089=>"101101001",
  22090=>"111011000",
  22091=>"101000001",
  22092=>"111111100",
  22093=>"000111111",
  22094=>"000100111",
  22095=>"111110000",
  22096=>"110000000",
  22097=>"110110000",
  22098=>"000000101",
  22099=>"110000000",
  22100=>"000011111",
  22101=>"000000110",
  22102=>"111000000",
  22103=>"000000000",
  22104=>"000000000",
  22105=>"000000000",
  22106=>"111111011",
  22107=>"000111111",
  22108=>"001000100",
  22109=>"111111111",
  22110=>"001000111",
  22111=>"000110100",
  22112=>"111000000",
  22113=>"011111111",
  22114=>"111111111",
  22115=>"111000000",
  22116=>"100101000",
  22117=>"111111000",
  22118=>"010111110",
  22119=>"000001000",
  22120=>"001111111",
  22121=>"000000111",
  22122=>"011111111",
  22123=>"111111111",
  22124=>"000011011",
  22125=>"000110111",
  22126=>"111111111",
  22127=>"111110000",
  22128=>"000001111",
  22129=>"011011001",
  22130=>"000000111",
  22131=>"111100100",
  22132=>"000000111",
  22133=>"100000000",
  22134=>"111000000",
  22135=>"000111111",
  22136=>"110000000",
  22137=>"000111111",
  22138=>"000000001",
  22139=>"111111100",
  22140=>"001000000",
  22141=>"000111000",
  22142=>"110100111",
  22143=>"000001011",
  22144=>"101101111",
  22145=>"011011000",
  22146=>"000000111",
  22147=>"000000000",
  22148=>"000110111",
  22149=>"000000000",
  22150=>"000000110",
  22151=>"111000000",
  22152=>"000000100",
  22153=>"000000000",
  22154=>"000111111",
  22155=>"000000000",
  22156=>"111111111",
  22157=>"010000011",
  22158=>"011000000",
  22159=>"111111111",
  22160=>"111111111",
  22161=>"000111111",
  22162=>"111000000",
  22163=>"110111001",
  22164=>"011000000",
  22165=>"000000000",
  22166=>"000000000",
  22167=>"000001000",
  22168=>"110101101",
  22169=>"111001011",
  22170=>"111111111",
  22171=>"111111111",
  22172=>"000000001",
  22173=>"111111101",
  22174=>"011001001",
  22175=>"000000000",
  22176=>"000000111",
  22177=>"001011010",
  22178=>"111101000",
  22179=>"110111111",
  22180=>"000011111",
  22181=>"100111100",
  22182=>"111111111",
  22183=>"100100100",
  22184=>"000010011",
  22185=>"111100101",
  22186=>"111111111",
  22187=>"111111001",
  22188=>"111000000",
  22189=>"000111011",
  22190=>"000000011",
  22191=>"000000000",
  22192=>"111111000",
  22193=>"001000000",
  22194=>"000011011",
  22195=>"110111111",
  22196=>"110110111",
  22197=>"000000000",
  22198=>"001000000",
  22199=>"000100001",
  22200=>"000000111",
  22201=>"000000010",
  22202=>"000100110",
  22203=>"110110110",
  22204=>"110110111",
  22205=>"000100110",
  22206=>"000000101",
  22207=>"101001101",
  22208=>"000000100",
  22209=>"000001001",
  22210=>"111100100",
  22211=>"001111111",
  22212=>"111111000",
  22213=>"010000000",
  22214=>"111101000",
  22215=>"000000000",
  22216=>"010111000",
  22217=>"000000111",
  22218=>"111101111",
  22219=>"111011000",
  22220=>"111111001",
  22221=>"001000100",
  22222=>"000000111",
  22223=>"000101111",
  22224=>"000010011",
  22225=>"110000010",
  22226=>"111000000",
  22227=>"111111111",
  22228=>"111111111",
  22229=>"111000000",
  22230=>"000000000",
  22231=>"000101000",
  22232=>"111100000",
  22233=>"000000000",
  22234=>"111111000",
  22235=>"000000000",
  22236=>"111011010",
  22237=>"000001111",
  22238=>"110110110",
  22239=>"000111111",
  22240=>"111111111",
  22241=>"000010111",
  22242=>"111111010",
  22243=>"000000000",
  22244=>"000000000",
  22245=>"000110111",
  22246=>"011111110",
  22247=>"000000000",
  22248=>"100000111",
  22249=>"000100111",
  22250=>"111111011",
  22251=>"011111111",
  22252=>"111000111",
  22253=>"000000011",
  22254=>"111101000",
  22255=>"111000100",
  22256=>"111111000",
  22257=>"000000001",
  22258=>"000010011",
  22259=>"000000001",
  22260=>"000000000",
  22261=>"000111111",
  22262=>"101111111",
  22263=>"111000111",
  22264=>"111100000",
  22265=>"000000000",
  22266=>"010111111",
  22267=>"001000000",
  22268=>"000000000",
  22269=>"111000001",
  22270=>"111101000",
  22271=>"000000000",
  22272=>"000000111",
  22273=>"001000110",
  22274=>"111111111",
  22275=>"000100111",
  22276=>"111111111",
  22277=>"100001001",
  22278=>"000000000",
  22279=>"000001100",
  22280=>"000000000",
  22281=>"000000000",
  22282=>"111111111",
  22283=>"111010001",
  22284=>"000110000",
  22285=>"110000111",
  22286=>"111111111",
  22287=>"000000000",
  22288=>"000101001",
  22289=>"111110110",
  22290=>"000000101",
  22291=>"111001001",
  22292=>"011001001",
  22293=>"001000100",
  22294=>"111111111",
  22295=>"000000000",
  22296=>"101110110",
  22297=>"001000000",
  22298=>"100111111",
  22299=>"011010000",
  22300=>"000001001",
  22301=>"000000000",
  22302=>"111111100",
  22303=>"000000110",
  22304=>"000000111",
  22305=>"011111011",
  22306=>"000000110",
  22307=>"011011111",
  22308=>"000000111",
  22309=>"000100111",
  22310=>"110000111",
  22311=>"000000000",
  22312=>"111111111",
  22313=>"000010010",
  22314=>"000000000",
  22315=>"010000001",
  22316=>"010111000",
  22317=>"100100110",
  22318=>"111101111",
  22319=>"110110111",
  22320=>"011001001",
  22321=>"000000000",
  22322=>"111000110",
  22323=>"000110111",
  22324=>"111011111",
  22325=>"011010000",
  22326=>"000000111",
  22327=>"111110111",
  22328=>"001010000",
  22329=>"000000000",
  22330=>"000000000",
  22331=>"111111100",
  22332=>"000000000",
  22333=>"000111111",
  22334=>"111111100",
  22335=>"000000100",
  22336=>"111000000",
  22337=>"010011001",
  22338=>"000000000",
  22339=>"000000000",
  22340=>"000000010",
  22341=>"000000100",
  22342=>"000010000",
  22343=>"001001101",
  22344=>"000000110",
  22345=>"000000111",
  22346=>"000000111",
  22347=>"000001011",
  22348=>"000000000",
  22349=>"111111111",
  22350=>"000000011",
  22351=>"110110111",
  22352=>"001110100",
  22353=>"000100110",
  22354=>"000101000",
  22355=>"000111111",
  22356=>"000100101",
  22357=>"111111111",
  22358=>"111111111",
  22359=>"111111101",
  22360=>"000000111",
  22361=>"110110111",
  22362=>"011000111",
  22363=>"111111110",
  22364=>"100111111",
  22365=>"110000011",
  22366=>"000000101",
  22367=>"100110111",
  22368=>"111111110",
  22369=>"000000000",
  22370=>"111001001",
  22371=>"111000000",
  22372=>"111101000",
  22373=>"000000111",
  22374=>"111111000",
  22375=>"001001001",
  22376=>"000000000",
  22377=>"000111010",
  22378=>"001011000",
  22379=>"111110111",
  22380=>"000100100",
  22381=>"100111000",
  22382=>"001000000",
  22383=>"000000011",
  22384=>"101101111",
  22385=>"111101001",
  22386=>"000110111",
  22387=>"111111001",
  22388=>"111001000",
  22389=>"001000111",
  22390=>"111101111",
  22391=>"000000000",
  22392=>"011000000",
  22393=>"000000000",
  22394=>"111111000",
  22395=>"000001001",
  22396=>"000110111",
  22397=>"000010011",
  22398=>"110111000",
  22399=>"101000101",
  22400=>"001000100",
  22401=>"001111111",
  22402=>"111110000",
  22403=>"100111111",
  22404=>"101111111",
  22405=>"000000010",
  22406=>"111111111",
  22407=>"111110111",
  22408=>"001001101",
  22409=>"110111110",
  22410=>"111111100",
  22411=>"111111111",
  22412=>"101001111",
  22413=>"100111101",
  22414=>"100101111",
  22415=>"000000000",
  22416=>"000000111",
  22417=>"000010011",
  22418=>"000110111",
  22419=>"001000000",
  22420=>"000001111",
  22421=>"000000000",
  22422=>"111111111",
  22423=>"001111111",
  22424=>"111011010",
  22425=>"111111111",
  22426=>"111111111",
  22427=>"110111000",
  22428=>"001000000",
  22429=>"111001000",
  22430=>"011001001",
  22431=>"111110111",
  22432=>"100111111",
  22433=>"111011111",
  22434=>"010011111",
  22435=>"000110001",
  22436=>"010110110",
  22437=>"011111000",
  22438=>"111000000",
  22439=>"100000011",
  22440=>"111111111",
  22441=>"111010011",
  22442=>"111111111",
  22443=>"000000000",
  22444=>"000000000",
  22445=>"000000001",
  22446=>"000000101",
  22447=>"000000000",
  22448=>"111110110",
  22449=>"000000001",
  22450=>"111110000",
  22451=>"001001000",
  22452=>"111111111",
  22453=>"000000000",
  22454=>"000111100",
  22455=>"000111111",
  22456=>"100000010",
  22457=>"111111111",
  22458=>"000100000",
  22459=>"111000000",
  22460=>"110110111",
  22461=>"111111111",
  22462=>"110111111",
  22463=>"011011011",
  22464=>"000000011",
  22465=>"001111011",
  22466=>"000000011",
  22467=>"000000111",
  22468=>"000111111",
  22469=>"000000001",
  22470=>"111111000",
  22471=>"001000001",
  22472=>"000000000",
  22473=>"000001011",
  22474=>"000000100",
  22475=>"000000000",
  22476=>"000000110",
  22477=>"001010010",
  22478=>"111000111",
  22479=>"110111111",
  22480=>"101001110",
  22481=>"111110100",
  22482=>"000111111",
  22483=>"001000000",
  22484=>"000000010",
  22485=>"111001111",
  22486=>"111111100",
  22487=>"001000011",
  22488=>"000000000",
  22489=>"100100000",
  22490=>"110010010",
  22491=>"111111111",
  22492=>"100000001",
  22493=>"111111011",
  22494=>"111110000",
  22495=>"001111111",
  22496=>"000010100",
  22497=>"000001000",
  22498=>"111000001",
  22499=>"000011000",
  22500=>"010010010",
  22501=>"000000000",
  22502=>"111000000",
  22503=>"000000111",
  22504=>"010010111",
  22505=>"111111001",
  22506=>"111110010",
  22507=>"000000000",
  22508=>"110110110",
  22509=>"110110110",
  22510=>"000000111",
  22511=>"111111110",
  22512=>"000000000",
  22513=>"111110111",
  22514=>"011001111",
  22515=>"111001011",
  22516=>"000111111",
  22517=>"001000000",
  22518=>"111111111",
  22519=>"011001000",
  22520=>"000000000",
  22521=>"100110110",
  22522=>"000001000",
  22523=>"000100110",
  22524=>"111001111",
  22525=>"111111111",
  22526=>"010000000",
  22527=>"000000111",
  22528=>"001000100",
  22529=>"000000000",
  22530=>"000000100",
  22531=>"001110000",
  22532=>"111110110",
  22533=>"000000000",
  22534=>"000111111",
  22535=>"111111011",
  22536=>"111001000",
  22537=>"000001111",
  22538=>"010110000",
  22539=>"000010010",
  22540=>"000110110",
  22541=>"000000111",
  22542=>"000000001",
  22543=>"111111011",
  22544=>"110000000",
  22545=>"000010010",
  22546=>"000011111",
  22547=>"011001000",
  22548=>"100000000",
  22549=>"101101111",
  22550=>"000000110",
  22551=>"000001111",
  22552=>"100110000",
  22553=>"001001111",
  22554=>"000000111",
  22555=>"000000010",
  22556=>"000000100",
  22557=>"110111111",
  22558=>"011101001",
  22559=>"111011001",
  22560=>"011011000",
  22561=>"000000111",
  22562=>"000000000",
  22563=>"000000111",
  22564=>"000110111",
  22565=>"011011001",
  22566=>"001000000",
  22567=>"100000000",
  22568=>"011000000",
  22569=>"100100000",
  22570=>"100001111",
  22571=>"100110110",
  22572=>"000111111",
  22573=>"111111111",
  22574=>"000000000",
  22575=>"001000000",
  22576=>"111011101",
  22577=>"011111001",
  22578=>"001001111",
  22579=>"111101100",
  22580=>"000110110",
  22581=>"111110100",
  22582=>"000011111",
  22583=>"010111111",
  22584=>"111111100",
  22585=>"000000101",
  22586=>"111011011",
  22587=>"000000000",
  22588=>"111101000",
  22589=>"001000000",
  22590=>"000010110",
  22591=>"111111011",
  22592=>"000000110",
  22593=>"100110110",
  22594=>"111011000",
  22595=>"111000000",
  22596=>"110111011",
  22597=>"001000001",
  22598=>"100000001",
  22599=>"111111111",
  22600=>"001001111",
  22601=>"000000000",
  22602=>"111101111",
  22603=>"000000110",
  22604=>"111111110",
  22605=>"111011000",
  22606=>"000001011",
  22607=>"111000011",
  22608=>"000000111",
  22609=>"000000011",
  22610=>"110111011",
  22611=>"111111001",
  22612=>"011111111",
  22613=>"110110000",
  22614=>"111000000",
  22615=>"001011001",
  22616=>"110111101",
  22617=>"111101111",
  22618=>"110100000",
  22619=>"000100110",
  22620=>"100100110",
  22621=>"111010110",
  22622=>"101001111",
  22623=>"100110111",
  22624=>"001111110",
  22625=>"011001111",
  22626=>"000010000",
  22627=>"111111111",
  22628=>"111100000",
  22629=>"111001111",
  22630=>"111111111",
  22631=>"000000011",
  22632=>"000000010",
  22633=>"100000000",
  22634=>"100101001",
  22635=>"010010111",
  22636=>"001101111",
  22637=>"000000111",
  22638=>"111101111",
  22639=>"100100110",
  22640=>"001001110",
  22641=>"000001111",
  22642=>"010110101",
  22643=>"111111110",
  22644=>"000101111",
  22645=>"000000110",
  22646=>"000000001",
  22647=>"000100110",
  22648=>"000000000",
  22649=>"010010111",
  22650=>"001001111",
  22651=>"011111111",
  22652=>"011110110",
  22653=>"000010011",
  22654=>"001000111",
  22655=>"010111110",
  22656=>"000111111",
  22657=>"111111111",
  22658=>"111111100",
  22659=>"111111100",
  22660=>"000000100",
  22661=>"111101111",
  22662=>"001000000",
  22663=>"000000011",
  22664=>"001001001",
  22665=>"111111111",
  22666=>"111000000",
  22667=>"111011001",
  22668=>"001111111",
  22669=>"111111101",
  22670=>"001000000",
  22671=>"000111111",
  22672=>"111110000",
  22673=>"110111110",
  22674=>"011011011",
  22675=>"001001111",
  22676=>"001100000",
  22677=>"011011011",
  22678=>"110100100",
  22679=>"000000000",
  22680=>"101001101",
  22681=>"111111111",
  22682=>"000011011",
  22683=>"000000000",
  22684=>"111111110",
  22685=>"001000001",
  22686=>"000000001",
  22687=>"111111111",
  22688=>"111111000",
  22689=>"001000000",
  22690=>"111011100",
  22691=>"000000000",
  22692=>"000000000",
  22693=>"000001011",
  22694=>"000100000",
  22695=>"001011111",
  22696=>"101101111",
  22697=>"001001111",
  22698=>"111001101",
  22699=>"111011001",
  22700=>"101101101",
  22701=>"000000000",
  22702=>"001001011",
  22703=>"011111111",
  22704=>"010100111",
  22705=>"111000100",
  22706=>"010111010",
  22707=>"000000000",
  22708=>"000000010",
  22709=>"011011100",
  22710=>"011111111",
  22711=>"101100111",
  22712=>"000100000",
  22713=>"110111110",
  22714=>"000000000",
  22715=>"011010000",
  22716=>"000000001",
  22717=>"000000110",
  22718=>"111111000",
  22719=>"111000000",
  22720=>"000110111",
  22721=>"000000001",
  22722=>"010110110",
  22723=>"111111110",
  22724=>"011011111",
  22725=>"100000110",
  22726=>"000000000",
  22727=>"010110111",
  22728=>"000000000",
  22729=>"111111111",
  22730=>"000011000",
  22731=>"000111111",
  22732=>"111111001",
  22733=>"001001000",
  22734=>"001111011",
  22735=>"111000100",
  22736=>"000000000",
  22737=>"000000000",
  22738=>"000001011",
  22739=>"110110111",
  22740=>"111011000",
  22741=>"100100111",
  22742=>"010000100",
  22743=>"111111000",
  22744=>"111110000",
  22745=>"000000000",
  22746=>"111111111",
  22747=>"111111111",
  22748=>"110000111",
  22749=>"000000000",
  22750=>"011111110",
  22751=>"111011011",
  22752=>"000000000",
  22753=>"000011111",
  22754=>"010000110",
  22755=>"111101111",
  22756=>"001011111",
  22757=>"000000001",
  22758=>"110110110",
  22759=>"111111111",
  22760=>"011011111",
  22761=>"101001000",
  22762=>"011011011",
  22763=>"001000000",
  22764=>"100101111",
  22765=>"111111111",
  22766=>"111111000",
  22767=>"000000000",
  22768=>"110100000",
  22769=>"111110000",
  22770=>"111111101",
  22771=>"000000111",
  22772=>"100000000",
  22773=>"000000010",
  22774=>"000111111",
  22775=>"000000000",
  22776=>"111111111",
  22777=>"001011010",
  22778=>"111000001",
  22779=>"101000110",
  22780=>"100111111",
  22781=>"111111100",
  22782=>"101000001",
  22783=>"011111001",
  22784=>"000000101",
  22785=>"000010000",
  22786=>"111010110",
  22787=>"011000000",
  22788=>"111100100",
  22789=>"000000111",
  22790=>"001001000",
  22791=>"111110000",
  22792=>"000000101",
  22793=>"000000000",
  22794=>"111110110",
  22795=>"111111110",
  22796=>"100000000",
  22797=>"111110111",
  22798=>"111110111",
  22799=>"111111000",
  22800=>"000000000",
  22801=>"000100000",
  22802=>"111011011",
  22803=>"001000000",
  22804=>"000010000",
  22805=>"011001000",
  22806=>"000001011",
  22807=>"000000001",
  22808=>"001001101",
  22809=>"000100100",
  22810=>"001100000",
  22811=>"011111111",
  22812=>"000000000",
  22813=>"110111111",
  22814=>"110000010",
  22815=>"000000000",
  22816=>"000000000",
  22817=>"000001001",
  22818=>"111111110",
  22819=>"111111111",
  22820=>"111111011",
  22821=>"000000001",
  22822=>"000100110",
  22823=>"100100000",
  22824=>"011001011",
  22825=>"000111111",
  22826=>"000110000",
  22827=>"000110111",
  22828=>"111111111",
  22829=>"000001011",
  22830=>"100110000",
  22831=>"100110101",
  22832=>"111111111",
  22833=>"000000111",
  22834=>"000110011",
  22835=>"101100110",
  22836=>"000000100",
  22837=>"010000111",
  22838=>"000000111",
  22839=>"011111111",
  22840=>"000000000",
  22841=>"111001000",
  22842=>"001000001",
  22843=>"111111111",
  22844=>"111111011",
  22845=>"111101101",
  22846=>"001111110",
  22847=>"000011011",
  22848=>"111111111",
  22849=>"111111111",
  22850=>"001111111",
  22851=>"010010111",
  22852=>"000110111",
  22853=>"000000000",
  22854=>"000110111",
  22855=>"110111110",
  22856=>"111000000",
  22857=>"000000000",
  22858=>"000001101",
  22859=>"110110100",
  22860=>"111110011",
  22861=>"111111111",
  22862=>"111111111",
  22863=>"100110110",
  22864=>"111100101",
  22865=>"001000100",
  22866=>"111100000",
  22867=>"101111011",
  22868=>"111111011",
  22869=>"011011011",
  22870=>"000000000",
  22871=>"111101101",
  22872=>"000110000",
  22873=>"000000000",
  22874=>"111100000",
  22875=>"100111111",
  22876=>"000001101",
  22877=>"000000000",
  22878=>"001101000",
  22879=>"111111111",
  22880=>"111111111",
  22881=>"001001111",
  22882=>"000100101",
  22883=>"111111111",
  22884=>"100111111",
  22885=>"001000111",
  22886=>"010111110",
  22887=>"000100100",
  22888=>"000011000",
  22889=>"110000000",
  22890=>"000111111",
  22891=>"011001001",
  22892=>"110010110",
  22893=>"001001111",
  22894=>"110111111",
  22895=>"111111100",
  22896=>"010110110",
  22897=>"000000111",
  22898=>"000000000",
  22899=>"001111001",
  22900=>"110111111",
  22901=>"000000000",
  22902=>"111101111",
  22903=>"101001101",
  22904=>"111001001",
  22905=>"111111000",
  22906=>"000110010",
  22907=>"111111010",
  22908=>"111010000",
  22909=>"000000000",
  22910=>"111111111",
  22911=>"111001111",
  22912=>"010000111",
  22913=>"000000111",
  22914=>"000000000",
  22915=>"000000000",
  22916=>"110011000",
  22917=>"111111111",
  22918=>"000000000",
  22919=>"110100100",
  22920=>"000000000",
  22921=>"111000000",
  22922=>"000000111",
  22923=>"000100000",
  22924=>"111100111",
  22925=>"000010010",
  22926=>"100111110",
  22927=>"110110100",
  22928=>"000000111",
  22929=>"111111000",
  22930=>"000000111",
  22931=>"011001110",
  22932=>"111111111",
  22933=>"000110110",
  22934=>"011000010",
  22935=>"000000000",
  22936=>"001111111",
  22937=>"011011011",
  22938=>"001001000",
  22939=>"001001101",
  22940=>"111011001",
  22941=>"001111000",
  22942=>"000001000",
  22943=>"111111111",
  22944=>"111111111",
  22945=>"011010000",
  22946=>"000000011",
  22947=>"111101101",
  22948=>"111110001",
  22949=>"000100000",
  22950=>"100100110",
  22951=>"000000011",
  22952=>"110110000",
  22953=>"001010000",
  22954=>"000010011",
  22955=>"001000000",
  22956=>"100000000",
  22957=>"000000101",
  22958=>"110011001",
  22959=>"111100011",
  22960=>"111100111",
  22961=>"000111111",
  22962=>"000000000",
  22963=>"111111111",
  22964=>"000010000",
  22965=>"001001000",
  22966=>"111111000",
  22967=>"111110001",
  22968=>"001001101",
  22969=>"000110110",
  22970=>"111111111",
  22971=>"101000000",
  22972=>"001001001",
  22973=>"100110100",
  22974=>"000000000",
  22975=>"000000010",
  22976=>"111101000",
  22977=>"101000011",
  22978=>"110110010",
  22979=>"111000000",
  22980=>"111111000",
  22981=>"001000000",
  22982=>"001000010",
  22983=>"000111111",
  22984=>"111100111",
  22985=>"101000110",
  22986=>"100100101",
  22987=>"110000111",
  22988=>"000001000",
  22989=>"011000000",
  22990=>"000111000",
  22991=>"001000000",
  22992=>"111101111",
  22993=>"111100110",
  22994=>"000001111",
  22995=>"000110111",
  22996=>"011001011",
  22997=>"111111000",
  22998=>"011000000",
  22999=>"001011011",
  23000=>"000111110",
  23001=>"111111011",
  23002=>"000000000",
  23003=>"111111010",
  23004=>"001111111",
  23005=>"000000110",
  23006=>"100110110",
  23007=>"000010110",
  23008=>"111011111",
  23009=>"000000000",
  23010=>"000111000",
  23011=>"000000000",
  23012=>"111111111",
  23013=>"101100011",
  23014=>"000000000",
  23015=>"111100101",
  23016=>"001000000",
  23017=>"110110110",
  23018=>"000000111",
  23019=>"111111001",
  23020=>"101111000",
  23021=>"001001001",
  23022=>"001000000",
  23023=>"100000000",
  23024=>"001000000",
  23025=>"111000010",
  23026=>"111100000",
  23027=>"100100000",
  23028=>"111001111",
  23029=>"011001001",
  23030=>"000110110",
  23031=>"011111101",
  23032=>"010000000",
  23033=>"101000100",
  23034=>"110110110",
  23035=>"011111111",
  23036=>"011000010",
  23037=>"001000001",
  23038=>"111111111",
  23039=>"000100000",
  23040=>"000000110",
  23041=>"111000000",
  23042=>"000000110",
  23043=>"000000000",
  23044=>"100000000",
  23045=>"110000000",
  23046=>"100100100",
  23047=>"111111111",
  23048=>"111011000",
  23049=>"111011011",
  23050=>"111111111",
  23051=>"111111011",
  23052=>"111111100",
  23053=>"111011000",
  23054=>"000111111",
  23055=>"001001000",
  23056=>"100100110",
  23057=>"100111111",
  23058=>"101000011",
  23059=>"000000110",
  23060=>"111001000",
  23061=>"000000111",
  23062=>"000111111",
  23063=>"101111111",
  23064=>"110110111",
  23065=>"100111001",
  23066=>"000111011",
  23067=>"111111011",
  23068=>"111000000",
  23069=>"001000000",
  23070=>"000000000",
  23071=>"001000111",
  23072=>"111001000",
  23073=>"110111111",
  23074=>"011011111",
  23075=>"001000000",
  23076=>"111011011",
  23077=>"000100100",
  23078=>"010000010",
  23079=>"010000000",
  23080=>"000000011",
  23081=>"000000111",
  23082=>"111000000",
  23083=>"000000000",
  23084=>"111000000",
  23085=>"111001000",
  23086=>"101011001",
  23087=>"101000000",
  23088=>"111110000",
  23089=>"000000000",
  23090=>"111111101",
  23091=>"111111011",
  23092=>"011011011",
  23093=>"101100000",
  23094=>"101111010",
  23095=>"000000110",
  23096=>"101001000",
  23097=>"001000000",
  23098=>"001001101",
  23099=>"111000100",
  23100=>"111111001",
  23101=>"000011001",
  23102=>"001000000",
  23103=>"111011001",
  23104=>"101000000",
  23105=>"000000000",
  23106=>"000000000",
  23107=>"111111111",
  23108=>"111001001",
  23109=>"111111111",
  23110=>"000000000",
  23111=>"000011111",
  23112=>"000000000",
  23113=>"000000100",
  23114=>"000101111",
  23115=>"000000000",
  23116=>"111111100",
  23117=>"000000100",
  23118=>"010000000",
  23119=>"000000111",
  23120=>"000000010",
  23121=>"101000100",
  23122=>"100011001",
  23123=>"110110000",
  23124=>"000000000",
  23125=>"000001000",
  23126=>"111000000",
  23127=>"111111000",
  23128=>"000000000",
  23129=>"001000000",
  23130=>"000000000",
  23131=>"000001001",
  23132=>"000000111",
  23133=>"001001001",
  23134=>"111111111",
  23135=>"101111111",
  23136=>"011000000",
  23137=>"011001000",
  23138=>"111111111",
  23139=>"000000000",
  23140=>"110110110",
  23141=>"001000001",
  23142=>"001000111",
  23143=>"101101101",
  23144=>"111111111",
  23145=>"110111111",
  23146=>"000010000",
  23147=>"000000100",
  23148=>"100100110",
  23149=>"000000001",
  23150=>"111111111",
  23151=>"111111111",
  23152=>"000111111",
  23153=>"000100000",
  23154=>"111001000",
  23155=>"011000011",
  23156=>"111011111",
  23157=>"000000000",
  23158=>"111101101",
  23159=>"111000001",
  23160=>"011001000",
  23161=>"001000100",
  23162=>"000000010",
  23163=>"111111000",
  23164=>"100100110",
  23165=>"111111111",
  23166=>"111111011",
  23167=>"111011011",
  23168=>"111100000",
  23169=>"111111111",
  23170=>"111000000",
  23171=>"000000000",
  23172=>"111111111",
  23173=>"111111000",
  23174=>"001000000",
  23175=>"000000000",
  23176=>"111111111",
  23177=>"000000100",
  23178=>"000000000",
  23179=>"110000000",
  23180=>"111111111",
  23181=>"011000000",
  23182=>"000011000",
  23183=>"111101001",
  23184=>"111000000",
  23185=>"000010000",
  23186=>"111111111",
  23187=>"000000000",
  23188=>"000101001",
  23189=>"111111111",
  23190=>"111111000",
  23191=>"111001000",
  23192=>"010011001",
  23193=>"110111111",
  23194=>"000000000",
  23195=>"110111011",
  23196=>"000101111",
  23197=>"011011011",
  23198=>"001111000",
  23199=>"111111001",
  23200=>"000100111",
  23201=>"001111111",
  23202=>"000000000",
  23203=>"000000000",
  23204=>"000100100",
  23205=>"000011111",
  23206=>"000000000",
  23207=>"111010000",
  23208=>"000011001",
  23209=>"111000000",
  23210=>"101101000",
  23211=>"000000000",
  23212=>"111011111",
  23213=>"110111111",
  23214=>"101000111",
  23215=>"000000111",
  23216=>"000011111",
  23217=>"001001001",
  23218=>"010111111",
  23219=>"111111000",
  23220=>"101000100",
  23221=>"111001011",
  23222=>"011010011",
  23223=>"111111111",
  23224=>"000000101",
  23225=>"111111111",
  23226=>"000000000",
  23227=>"110111011",
  23228=>"000111110",
  23229=>"111000000",
  23230=>"000000000",
  23231=>"000000000",
  23232=>"001111111",
  23233=>"000000000",
  23234=>"000000000",
  23235=>"111111111",
  23236=>"100000000",
  23237=>"000000111",
  23238=>"000000000",
  23239=>"000101111",
  23240=>"000000000",
  23241=>"011011111",
  23242=>"010010000",
  23243=>"111111111",
  23244=>"111111111",
  23245=>"000000000",
  23246=>"111111101",
  23247=>"111111111",
  23248=>"111001000",
  23249=>"100000000",
  23250=>"111110111",
  23251=>"001000111",
  23252=>"110000000",
  23253=>"000000000",
  23254=>"111111111",
  23255=>"000000101",
  23256=>"000001000",
  23257=>"010111111",
  23258=>"110110000",
  23259=>"000111111",
  23260=>"001001001",
  23261=>"111000000",
  23262=>"000000000",
  23263=>"000000000",
  23264=>"111111111",
  23265=>"000000000",
  23266=>"111101111",
  23267=>"000110000",
  23268=>"000001100",
  23269=>"011010000",
  23270=>"000111111",
  23271=>"100111001",
  23272=>"100111111",
  23273=>"000000010",
  23274=>"111011001",
  23275=>"111001011",
  23276=>"011000000",
  23277=>"111111111",
  23278=>"010111111",
  23279=>"000000000",
  23280=>"001000100",
  23281=>"000000111",
  23282=>"111111111",
  23283=>"000111100",
  23284=>"111111111",
  23285=>"111111111",
  23286=>"100110000",
  23287=>"000000000",
  23288=>"111001111",
  23289=>"111101000",
  23290=>"000011111",
  23291=>"111111000",
  23292=>"011011000",
  23293=>"100000000",
  23294=>"000000000",
  23295=>"001001011",
  23296=>"000111111",
  23297=>"011010000",
  23298=>"111000011",
  23299=>"110000000",
  23300=>"000000000",
  23301=>"000000100",
  23302=>"111111101",
  23303=>"111010001",
  23304=>"111111111",
  23305=>"000111011",
  23306=>"000000000",
  23307=>"000111111",
  23308=>"000110110",
  23309=>"000000010",
  23310=>"110111111",
  23311=>"000111111",
  23312=>"111100101",
  23313=>"000000010",
  23314=>"111111000",
  23315=>"000001101",
  23316=>"000000111",
  23317=>"000000000",
  23318=>"000000111",
  23319=>"111111000",
  23320=>"110110111",
  23321=>"011111000",
  23322=>"101000000",
  23323=>"001111111",
  23324=>"000100101",
  23325=>"100000000",
  23326=>"000000101",
  23327=>"111111111",
  23328=>"000000111",
  23329=>"101001000",
  23330=>"001001111",
  23331=>"001111111",
  23332=>"000000000",
  23333=>"111111000",
  23334=>"000011011",
  23335=>"000000001",
  23336=>"110110111",
  23337=>"000111111",
  23338=>"000000000",
  23339=>"111000000",
  23340=>"010111001",
  23341=>"111011000",
  23342=>"110111000",
  23343=>"000000000",
  23344=>"011011111",
  23345=>"000010010",
  23346=>"101000100",
  23347=>"011011000",
  23348=>"101100000",
  23349=>"101000011",
  23350=>"110110000",
  23351=>"000000000",
  23352=>"111111101",
  23353=>"000000000",
  23354=>"000000111",
  23355=>"111110000",
  23356=>"110110111",
  23357=>"000000111",
  23358=>"000000000",
  23359=>"000111000",
  23360=>"000000111",
  23361=>"000000101",
  23362=>"010011111",
  23363=>"111111000",
  23364=>"111011111",
  23365=>"000000100",
  23366=>"111111111",
  23367=>"111111111",
  23368=>"010000000",
  23369=>"000000000",
  23370=>"111111111",
  23371=>"001000011",
  23372=>"111001001",
  23373=>"000111100",
  23374=>"001001111",
  23375=>"000000000",
  23376=>"000001001",
  23377=>"000000111",
  23378=>"000000111",
  23379=>"111111111",
  23380=>"000000000",
  23381=>"011011011",
  23382=>"110111000",
  23383=>"111000000",
  23384=>"000111000",
  23385=>"111111000",
  23386=>"111111000",
  23387=>"000001111",
  23388=>"111000000",
  23389=>"111000001",
  23390=>"000000000",
  23391=>"110111111",
  23392=>"000000000",
  23393=>"000000010",
  23394=>"000010000",
  23395=>"000000000",
  23396=>"111111111",
  23397=>"111111000",
  23398=>"001001000",
  23399=>"011011011",
  23400=>"000000101",
  23401=>"000000000",
  23402=>"000000000",
  23403=>"111111011",
  23404=>"111111110",
  23405=>"100000000",
  23406=>"001111111",
  23407=>"000000000",
  23408=>"000000000",
  23409=>"111111011",
  23410=>"111111111",
  23411=>"000000000",
  23412=>"000110000",
  23413=>"000000000",
  23414=>"011011000",
  23415=>"111001100",
  23416=>"111000000",
  23417=>"100111111",
  23418=>"101001000",
  23419=>"111111111",
  23420=>"000000000",
  23421=>"001000000",
  23422=>"111111000",
  23423=>"000000000",
  23424=>"100111111",
  23425=>"101001011",
  23426=>"100110111",
  23427=>"000000000",
  23428=>"110111000",
  23429=>"000010000",
  23430=>"000000000",
  23431=>"001001101",
  23432=>"111111000",
  23433=>"011000000",
  23434=>"111111010",
  23435=>"000101111",
  23436=>"111111111",
  23437=>"110110111",
  23438=>"011000000",
  23439=>"000000011",
  23440=>"000000000",
  23441=>"111100110",
  23442=>"111111111",
  23443=>"111011111",
  23444=>"001101111",
  23445=>"000000000",
  23446=>"100000100",
  23447=>"100100110",
  23448=>"111111000",
  23449=>"111000001",
  23450=>"000000111",
  23451=>"000000000",
  23452=>"000001111",
  23453=>"000000000",
  23454=>"000111010",
  23455=>"000000000",
  23456=>"111000110",
  23457=>"111011000",
  23458=>"000000010",
  23459=>"000000000",
  23460=>"100101001",
  23461=>"111111011",
  23462=>"110100000",
  23463=>"111000101",
  23464=>"111111111",
  23465=>"010010000",
  23466=>"100111111",
  23467=>"011000111",
  23468=>"000000111",
  23469=>"111001000",
  23470=>"000010000",
  23471=>"000000110",
  23472=>"111110000",
  23473=>"000000111",
  23474=>"110110000",
  23475=>"000000111",
  23476=>"111111011",
  23477=>"111111111",
  23478=>"110111010",
  23479=>"111111111",
  23480=>"000000000",
  23481=>"000111111",
  23482=>"111010010",
  23483=>"111011011",
  23484=>"111111001",
  23485=>"101110000",
  23486=>"110000010",
  23487=>"011110111",
  23488=>"000111011",
  23489=>"111111000",
  23490=>"000001001",
  23491=>"000000001",
  23492=>"000001111",
  23493=>"010110000",
  23494=>"000000000",
  23495=>"001000000",
  23496=>"000111000",
  23497=>"111000000",
  23498=>"000001000",
  23499=>"011000000",
  23500=>"001001111",
  23501=>"101000000",
  23502=>"101111111",
  23503=>"111111000",
  23504=>"000000000",
  23505=>"000111111",
  23506=>"000000110",
  23507=>"000110111",
  23508=>"000000000",
  23509=>"000000000",
  23510=>"010011111",
  23511=>"110000000",
  23512=>"111111111",
  23513=>"000010111",
  23514=>"111011010",
  23515=>"111111111",
  23516=>"000111111",
  23517=>"001110111",
  23518=>"010000000",
  23519=>"000000000",
  23520=>"110111111",
  23521=>"001001000",
  23522=>"000101111",
  23523=>"111101000",
  23524=>"110111110",
  23525=>"011100111",
  23526=>"000000111",
  23527=>"111111111",
  23528=>"000000000",
  23529=>"111111111",
  23530=>"111111000",
  23531=>"010000000",
  23532=>"100111111",
  23533=>"111111111",
  23534=>"111111000",
  23535=>"000000000",
  23536=>"000000001",
  23537=>"111111111",
  23538=>"011011111",
  23539=>"111111111",
  23540=>"000000000",
  23541=>"000000000",
  23542=>"100111111",
  23543=>"111100111",
  23544=>"000000101",
  23545=>"000001111",
  23546=>"000100110",
  23547=>"000110111",
  23548=>"111011001",
  23549=>"111111111",
  23550=>"111111111",
  23551=>"111111111",
  23552=>"000100110",
  23553=>"000000000",
  23554=>"000000000",
  23555=>"000001110",
  23556=>"111111111",
  23557=>"011000000",
  23558=>"111111111",
  23559=>"000000000",
  23560=>"000000011",
  23561=>"100111111",
  23562=>"000000000",
  23563=>"101111111",
  23564=>"111111111",
  23565=>"000101111",
  23566=>"111111100",
  23567=>"001000100",
  23568=>"000000101",
  23569=>"100100110",
  23570=>"001000110",
  23571=>"001111111",
  23572=>"000000000",
  23573=>"111111111",
  23574=>"111111111",
  23575=>"110110100",
  23576=>"000000100",
  23577=>"111111111",
  23578=>"000000111",
  23579=>"000010010",
  23580=>"000110111",
  23581=>"111111111",
  23582=>"000000000",
  23583=>"000111111",
  23584=>"111000000",
  23585=>"010110000",
  23586=>"011101001",
  23587=>"111111111",
  23588=>"000000000",
  23589=>"111101111",
  23590=>"000000000",
  23591=>"111001001",
  23592=>"001001001",
  23593=>"001011111",
  23594=>"001000000",
  23595=>"111000000",
  23596=>"000011011",
  23597=>"000000000",
  23598=>"000001000",
  23599=>"111100100",
  23600=>"000111111",
  23601=>"100111111",
  23602=>"011011111",
  23603=>"100110110",
  23604=>"100000000",
  23605=>"111001001",
  23606=>"111010000",
  23607=>"100111111",
  23608=>"110111111",
  23609=>"001001111",
  23610=>"111111111",
  23611=>"000000000",
  23612=>"111001111",
  23613=>"000000000",
  23614=>"000000000",
  23615=>"100000001",
  23616=>"111111000",
  23617=>"110110110",
  23618=>"000000000",
  23619=>"000000000",
  23620=>"101000000",
  23621=>"000011111",
  23622=>"110000000",
  23623=>"111111011",
  23624=>"000000000",
  23625=>"111111111",
  23626=>"000011000",
  23627=>"101111110",
  23628=>"011111111",
  23629=>"111111111",
  23630=>"111111000",
  23631=>"000000101",
  23632=>"111111111",
  23633=>"111111111",
  23634=>"101111000",
  23635=>"001011111",
  23636=>"000000000",
  23637=>"111111111",
  23638=>"000010111",
  23639=>"100100111",
  23640=>"000101111",
  23641=>"101000000",
  23642=>"000110111",
  23643=>"000000111",
  23644=>"011011111",
  23645=>"000001111",
  23646=>"000000000",
  23647=>"111111000",
  23648=>"000000000",
  23649=>"111011000",
  23650=>"000000000",
  23651=>"000000000",
  23652=>"100111110",
  23653=>"100100000",
  23654=>"111110111",
  23655=>"111111111",
  23656=>"000000000",
  23657=>"111111111",
  23658=>"100100100",
  23659=>"001000010",
  23660=>"110110000",
  23661=>"000000100",
  23662=>"000001001",
  23663=>"000000000",
  23664=>"000111000",
  23665=>"111000000",
  23666=>"001001000",
  23667=>"110111100",
  23668=>"000000000",
  23669=>"001000111",
  23670=>"000100100",
  23671=>"000000000",
  23672=>"000000000",
  23673=>"111111110",
  23674=>"110010100",
  23675=>"100000000",
  23676=>"100100100",
  23677=>"111111111",
  23678=>"010110110",
  23679=>"011000000",
  23680=>"111111111",
  23681=>"111111111",
  23682=>"110110110",
  23683=>"000001011",
  23684=>"001111111",
  23685=>"000000111",
  23686=>"100101101",
  23687=>"111111111",
  23688=>"111111111",
  23689=>"011011111",
  23690=>"000000000",
  23691=>"000000111",
  23692=>"000000000",
  23693=>"000000001",
  23694=>"000000000",
  23695=>"111111111",
  23696=>"000000011",
  23697=>"010000000",
  23698=>"111100100",
  23699=>"000001011",
  23700=>"111110111",
  23701=>"101111001",
  23702=>"100111111",
  23703=>"111111111",
  23704=>"000000000",
  23705=>"111100100",
  23706=>"111111111",
  23707=>"000000000",
  23708=>"000010000",
  23709=>"000000000",
  23710=>"011111111",
  23711=>"000000000",
  23712=>"111011000",
  23713=>"111110000",
  23714=>"000000000",
  23715=>"111000001",
  23716=>"011111110",
  23717=>"000001000",
  23718=>"000000111",
  23719=>"110000010",
  23720=>"010011111",
  23721=>"000000000",
  23722=>"101100000",
  23723=>"101111000",
  23724=>"001101111",
  23725=>"111011011",
  23726=>"111111101",
  23727=>"111111111",
  23728=>"011000000",
  23729=>"011001001",
  23730=>"111111111",
  23731=>"111101000",
  23732=>"111111111",
  23733=>"000000000",
  23734=>"111101001",
  23735=>"000000001",
  23736=>"001000000",
  23737=>"011001001",
  23738=>"000000000",
  23739=>"110000000",
  23740=>"000000000",
  23741=>"000001011",
  23742=>"000000000",
  23743=>"111111111",
  23744=>"110000000",
  23745=>"011111111",
  23746=>"011111111",
  23747=>"000000000",
  23748=>"000000100",
  23749=>"000000000",
  23750=>"100110111",
  23751=>"011111111",
  23752=>"000111111",
  23753=>"111011000",
  23754=>"000010111",
  23755=>"111111101",
  23756=>"000000000",
  23757=>"101111111",
  23758=>"110111011",
  23759=>"111110100",
  23760=>"100100000",
  23761=>"111101000",
  23762=>"000011000",
  23763=>"000001101",
  23764=>"100100001",
  23765=>"001100000",
  23766=>"000010010",
  23767=>"010001111",
  23768=>"100100000",
  23769=>"000000001",
  23770=>"000000101",
  23771=>"000011110",
  23772=>"000111111",
  23773=>"111111001",
  23774=>"111110100",
  23775=>"001001111",
  23776=>"000000000",
  23777=>"011000000",
  23778=>"000000000",
  23779=>"001000000",
  23780=>"111111000",
  23781=>"000000001",
  23782=>"111011011",
  23783=>"111111111",
  23784=>"111111111",
  23785=>"001001111",
  23786=>"000000000",
  23787=>"111111000",
  23788=>"000000001",
  23789=>"111000000",
  23790=>"000000000",
  23791=>"111000000",
  23792=>"000000100",
  23793=>"111111111",
  23794=>"111011111",
  23795=>"111110111",
  23796=>"111111111",
  23797=>"110000000",
  23798=>"001001000",
  23799=>"111111111",
  23800=>"101111111",
  23801=>"001011111",
  23802=>"111111111",
  23803=>"000000000",
  23804=>"001010100",
  23805=>"110111001",
  23806=>"001001111",
  23807=>"111101111",
  23808=>"111110111",
  23809=>"000010010",
  23810=>"000111111",
  23811=>"010111111",
  23812=>"000000000",
  23813=>"000001101",
  23814=>"000001001",
  23815=>"000001001",
  23816=>"000110100",
  23817=>"110110110",
  23818=>"111001001",
  23819=>"111111111",
  23820=>"000010111",
  23821=>"111111000",
  23822=>"111111111",
  23823=>"000000001",
  23824=>"111111111",
  23825=>"111111000",
  23826=>"111111111",
  23827=>"000000000",
  23828=>"000000000",
  23829=>"000000000",
  23830=>"000000000",
  23831=>"111111111",
  23832=>"000000000",
  23833=>"010011111",
  23834=>"110000000",
  23835=>"000000001",
  23836=>"100100100",
  23837=>"111111100",
  23838=>"000000000",
  23839=>"111111100",
  23840=>"001001000",
  23841=>"111111111",
  23842=>"010011000",
  23843=>"111101101",
  23844=>"000111111",
  23845=>"000000000",
  23846=>"111110111",
  23847=>"011111111",
  23848=>"100000000",
  23849=>"011000000",
  23850=>"010000100",
  23851=>"000000000",
  23852=>"110100111",
  23853=>"011011001",
  23854=>"100000000",
  23855=>"100000100",
  23856=>"000000000",
  23857=>"111111010",
  23858=>"111100110",
  23859=>"011111111",
  23860=>"000000000",
  23861=>"000000001",
  23862=>"000000000",
  23863=>"111110000",
  23864=>"000000000",
  23865=>"111111111",
  23866=>"101000111",
  23867=>"000000000",
  23868=>"000000000",
  23869=>"100000111",
  23870=>"111111101",
  23871=>"111000000",
  23872=>"000011000",
  23873=>"000000000",
  23874=>"000000000",
  23875=>"000000101",
  23876=>"001000000",
  23877=>"000000111",
  23878=>"000011111",
  23879=>"000000110",
  23880=>"000000001",
  23881=>"000000000",
  23882=>"001000000",
  23883=>"100000000",
  23884=>"011111100",
  23885=>"000100000",
  23886=>"000001011",
  23887=>"011111001",
  23888=>"001000001",
  23889=>"011010111",
  23890=>"000000000",
  23891=>"111000000",
  23892=>"111111100",
  23893=>"001001011",
  23894=>"001111111",
  23895=>"111111111",
  23896=>"000000000",
  23897=>"000000000",
  23898=>"000000000",
  23899=>"111111101",
  23900=>"100101101",
  23901=>"111111111",
  23902=>"111000000",
  23903=>"001000111",
  23904=>"111111000",
  23905=>"000000000",
  23906=>"000000010",
  23907=>"000100111",
  23908=>"011000010",
  23909=>"001000000",
  23910=>"111111111",
  23911=>"000110111",
  23912=>"001000000",
  23913=>"111111000",
  23914=>"111111110",
  23915=>"011011001",
  23916=>"111111110",
  23917=>"110110110",
  23918=>"111000000",
  23919=>"000000000",
  23920=>"000000000",
  23921=>"000000010",
  23922=>"111111111",
  23923=>"111110100",
  23924=>"000000000",
  23925=>"000000000",
  23926=>"000000010",
  23927=>"000000000",
  23928=>"000000000",
  23929=>"000010111",
  23930=>"011011000",
  23931=>"111101000",
  23932=>"110000000",
  23933=>"111111111",
  23934=>"000111111",
  23935=>"111111110",
  23936=>"111111011",
  23937=>"111111111",
  23938=>"001001011",
  23939=>"111100100",
  23940=>"101111100",
  23941=>"111111001",
  23942=>"111000000",
  23943=>"111111111",
  23944=>"100000000",
  23945=>"111110000",
  23946=>"000000000",
  23947=>"000000000",
  23948=>"101000111",
  23949=>"111100000",
  23950=>"001111111",
  23951=>"000000000",
  23952=>"000000100",
  23953=>"111111111",
  23954=>"110111111",
  23955=>"000000000",
  23956=>"001001011",
  23957=>"000000000",
  23958=>"000000000",
  23959=>"010001111",
  23960=>"110110100",
  23961=>"000000111",
  23962=>"111111110",
  23963=>"000000000",
  23964=>"111111111",
  23965=>"111111100",
  23966=>"101001001",
  23967=>"110010000",
  23968=>"001001111",
  23969=>"011011110",
  23970=>"111101111",
  23971=>"000000111",
  23972=>"000000111",
  23973=>"000000010",
  23974=>"000000000",
  23975=>"000000000",
  23976=>"000110100",
  23977=>"000011001",
  23978=>"111111111",
  23979=>"110100000",
  23980=>"000011111",
  23981=>"000000001",
  23982=>"111011011",
  23983=>"000000000",
  23984=>"100100100",
  23985=>"111111111",
  23986=>"111101111",
  23987=>"010000000",
  23988=>"111100000",
  23989=>"000000000",
  23990=>"000001101",
  23991=>"000000000",
  23992=>"000110111",
  23993=>"001111011",
  23994=>"111111111",
  23995=>"111101111",
  23996=>"100111111",
  23997=>"111111000",
  23998=>"000000000",
  23999=>"010011111",
  24000=>"000000001",
  24001=>"000000111",
  24002=>"111111010",
  24003=>"000000000",
  24004=>"000000001",
  24005=>"110100111",
  24006=>"000000000",
  24007=>"110111111",
  24008=>"000000000",
  24009=>"010111110",
  24010=>"010000000",
  24011=>"111111111",
  24012=>"111010110",
  24013=>"000010111",
  24014=>"111111101",
  24015=>"110111111",
  24016=>"000000000",
  24017=>"111001001",
  24018=>"110100000",
  24019=>"001001001",
  24020=>"111111000",
  24021=>"110100110",
  24022=>"000000000",
  24023=>"110110110",
  24024=>"111111111",
  24025=>"111110110",
  24026=>"111111101",
  24027=>"000000111",
  24028=>"111000010",
  24029=>"111001000",
  24030=>"000010000",
  24031=>"011110111",
  24032=>"000000000",
  24033=>"000000000",
  24034=>"001000000",
  24035=>"100000000",
  24036=>"111111111",
  24037=>"111011000",
  24038=>"000000000",
  24039=>"100000000",
  24040=>"000001101",
  24041=>"000000000",
  24042=>"111011001",
  24043=>"111111111",
  24044=>"111000000",
  24045=>"111111100",
  24046=>"000001001",
  24047=>"110111111",
  24048=>"111111111",
  24049=>"000100111",
  24050=>"000000000",
  24051=>"000000000",
  24052=>"111111111",
  24053=>"111111111",
  24054=>"000100110",
  24055=>"111110111",
  24056=>"111111111",
  24057=>"000000011",
  24058=>"000000000",
  24059=>"000111101",
  24060=>"011011111",
  24061=>"111110100",
  24062=>"000000000",
  24063=>"000000001",
  24064=>"111010000",
  24065=>"111101101",
  24066=>"000000111",
  24067=>"000000001",
  24068=>"001000000",
  24069=>"111000000",
  24070=>"110100100",
  24071=>"111111111",
  24072=>"101100110",
  24073=>"111111000",
  24074=>"111111101",
  24075=>"010111011",
  24076=>"100100111",
  24077=>"111111111",
  24078=>"000000000",
  24079=>"111110111",
  24080=>"000111111",
  24081=>"100000000",
  24082=>"000000111",
  24083=>"100000000",
  24084=>"110111111",
  24085=>"000000000",
  24086=>"000000000",
  24087=>"011011111",
  24088=>"000001111",
  24089=>"000100110",
  24090=>"000000000",
  24091=>"000110100",
  24092=>"111001001",
  24093=>"000000000",
  24094=>"111110111",
  24095=>"111111111",
  24096=>"111000000",
  24097=>"000000110",
  24098=>"100100000",
  24099=>"000000000",
  24100=>"111111100",
  24101=>"111111110",
  24102=>"000100111",
  24103=>"011011010",
  24104=>"010111111",
  24105=>"000000001",
  24106=>"001001101",
  24107=>"100000000",
  24108=>"000001111",
  24109=>"000000000",
  24110=>"111100110",
  24111=>"000000111",
  24112=>"000000000",
  24113=>"111111110",
  24114=>"011001000",
  24115=>"000000000",
  24116=>"000000001",
  24117=>"111011001",
  24118=>"101111111",
  24119=>"000100100",
  24120=>"000111111",
  24121=>"000000000",
  24122=>"111111111",
  24123=>"000000000",
  24124=>"000000110",
  24125=>"110111111",
  24126=>"111111111",
  24127=>"000000000",
  24128=>"100101100",
  24129=>"000000000",
  24130=>"010111111",
  24131=>"011111111",
  24132=>"011111110",
  24133=>"100111111",
  24134=>"111111000",
  24135=>"110000000",
  24136=>"000100111",
  24137=>"100000100",
  24138=>"100101111",
  24139=>"001111011",
  24140=>"000001000",
  24141=>"111111111",
  24142=>"000000110",
  24143=>"111110111",
  24144=>"000001000",
  24145=>"000000000",
  24146=>"110111111",
  24147=>"001001000",
  24148=>"111000110",
  24149=>"111011011",
  24150=>"000000000",
  24151=>"000000001",
  24152=>"111111111",
  24153=>"000000101",
  24154=>"111111111",
  24155=>"011011011",
  24156=>"111111111",
  24157=>"000000000",
  24158=>"001111111",
  24159=>"011000000",
  24160=>"111111111",
  24161=>"000110111",
  24162=>"101100000",
  24163=>"111101111",
  24164=>"111011111",
  24165=>"000000000",
  24166=>"111111110",
  24167=>"000000100",
  24168=>"111110000",
  24169=>"011010110",
  24170=>"000011000",
  24171=>"101110111",
  24172=>"111111111",
  24173=>"011010100",
  24174=>"000011001",
  24175=>"001001001",
  24176=>"000000000",
  24177=>"101101000",
  24178=>"000000000",
  24179=>"000101100",
  24180=>"111111110",
  24181=>"000100000",
  24182=>"111111111",
  24183=>"111111111",
  24184=>"110110000",
  24185=>"000000000",
  24186=>"000010011",
  24187=>"000000000",
  24188=>"001000000",
  24189=>"000000010",
  24190=>"000000111",
  24191=>"000000000",
  24192=>"111011111",
  24193=>"111111110",
  24194=>"000000111",
  24195=>"100111111",
  24196=>"111011111",
  24197=>"001000000",
  24198=>"111111111",
  24199=>"001001000",
  24200=>"100000000",
  24201=>"000100000",
  24202=>"111111111",
  24203=>"111111110",
  24204=>"111111110",
  24205=>"111111111",
  24206=>"101111111",
  24207=>"100000000",
  24208=>"111111111",
  24209=>"101101111",
  24210=>"000111111",
  24211=>"000000000",
  24212=>"111111111",
  24213=>"001001111",
  24214=>"000000000",
  24215=>"111011001",
  24216=>"111111111",
  24217=>"001101001",
  24218=>"000100000",
  24219=>"111100100",
  24220=>"000000000",
  24221=>"000000000",
  24222=>"111110111",
  24223=>"100000000",
  24224=>"000001101",
  24225=>"000000000",
  24226=>"111111111",
  24227=>"110000000",
  24228=>"110111000",
  24229=>"000111000",
  24230=>"111111110",
  24231=>"110111111",
  24232=>"000010111",
  24233=>"000000000",
  24234=>"111111111",
  24235=>"111111111",
  24236=>"000000000",
  24237=>"101111111",
  24238=>"011111111",
  24239=>"001001101",
  24240=>"100110111",
  24241=>"111001001",
  24242=>"111111111",
  24243=>"100000101",
  24244=>"011011111",
  24245=>"000010010",
  24246=>"111111111",
  24247=>"000111010",
  24248=>"101001000",
  24249=>"000100111",
  24250=>"111000001",
  24251=>"111111111",
  24252=>"000000000",
  24253=>"000000000",
  24254=>"000000001",
  24255=>"100100111",
  24256=>"000101111",
  24257=>"111111111",
  24258=>"110101111",
  24259=>"000000000",
  24260=>"000000000",
  24261=>"000000000",
  24262=>"111111010",
  24263=>"111111111",
  24264=>"111111110",
  24265=>"011001000",
  24266=>"001000000",
  24267=>"110000000",
  24268=>"000011001",
  24269=>"110000000",
  24270=>"011110111",
  24271=>"000111111",
  24272=>"010111101",
  24273=>"000110110",
  24274=>"111111001",
  24275=>"000000011",
  24276=>"111111000",
  24277=>"000100110",
  24278=>"010000000",
  24279=>"111111111",
  24280=>"111111111",
  24281=>"111111000",
  24282=>"000000000",
  24283=>"011111111",
  24284=>"111001101",
  24285=>"001100111",
  24286=>"110100100",
  24287=>"000001000",
  24288=>"111111111",
  24289=>"100000101",
  24290=>"000000000",
  24291=>"000000000",
  24292=>"000000111",
  24293=>"110100100",
  24294=>"111111000",
  24295=>"111111111",
  24296=>"100000000",
  24297=>"000000011",
  24298=>"111001011",
  24299=>"000000000",
  24300=>"000000000",
  24301=>"111000000",
  24302=>"000000011",
  24303=>"001000111",
  24304=>"000001000",
  24305=>"000000100",
  24306=>"111111111",
  24307=>"001000011",
  24308=>"111111111",
  24309=>"011011000",
  24310=>"001111111",
  24311=>"011000000",
  24312=>"000000000",
  24313=>"111111111",
  24314=>"000000011",
  24315=>"111111111",
  24316=>"101001111",
  24317=>"000001001",
  24318=>"000000000",
  24319=>"111111111",
  24320=>"000010000",
  24321=>"110111001",
  24322=>"111111111",
  24323=>"000000110",
  24324=>"111111111",
  24325=>"111111111",
  24326=>"111111000",
  24327=>"001111111",
  24328=>"111111100",
  24329=>"111100111",
  24330=>"000000000",
  24331=>"100110010",
  24332=>"111111000",
  24333=>"000000000",
  24334=>"001111111",
  24335=>"111000000",
  24336=>"000100000",
  24337=>"000111111",
  24338=>"111111011",
  24339=>"110100000",
  24340=>"111101000",
  24341=>"000000000",
  24342=>"001001001",
  24343=>"101110111",
  24344=>"111010000",
  24345=>"011010001",
  24346=>"000011111",
  24347=>"110111001",
  24348=>"000000000",
  24349=>"110110111",
  24350=>"111111111",
  24351=>"001101111",
  24352=>"000111111",
  24353=>"111000000",
  24354=>"000000000",
  24355=>"101110010",
  24356=>"100100101",
  24357=>"111111111",
  24358=>"111000001",
  24359=>"000000111",
  24360=>"111111111",
  24361=>"110000011",
  24362=>"111111111",
  24363=>"000000100",
  24364=>"111111111",
  24365=>"110100100",
  24366=>"000000000",
  24367=>"111111110",
  24368=>"101101100",
  24369=>"110100000",
  24370=>"000000000",
  24371=>"010111000",
  24372=>"000111111",
  24373=>"111001000",
  24374=>"000000000",
  24375=>"111100110",
  24376=>"000000011",
  24377=>"000010101",
  24378=>"000000000",
  24379=>"000000010",
  24380=>"000000110",
  24381=>"000000111",
  24382=>"000000000",
  24383=>"111111011",
  24384=>"000111111",
  24385=>"000111111",
  24386=>"000111011",
  24387=>"111111111",
  24388=>"111100000",
  24389=>"111001000",
  24390=>"000000011",
  24391=>"011100101",
  24392=>"111111111",
  24393=>"001001111",
  24394=>"001011111",
  24395=>"100110110",
  24396=>"110111000",
  24397=>"000010010",
  24398=>"001000000",
  24399=>"000000011",
  24400=>"110100110",
  24401=>"000000111",
  24402=>"000000000",
  24403=>"000111111",
  24404=>"011000000",
  24405=>"001001111",
  24406=>"001001001",
  24407=>"000000011",
  24408=>"001111110",
  24409=>"111101001",
  24410=>"111111111",
  24411=>"011100000",
  24412=>"000000000",
  24413=>"000000100",
  24414=>"000000000",
  24415=>"001001001",
  24416=>"000000111",
  24417=>"001000000",
  24418=>"111101011",
  24419=>"111111111",
  24420=>"100100100",
  24421=>"111101101",
  24422=>"000000000",
  24423=>"000010111",
  24424=>"001111111",
  24425=>"000001111",
  24426=>"111111111",
  24427=>"000000000",
  24428=>"000001000",
  24429=>"100100001",
  24430=>"000000000",
  24431=>"111111111",
  24432=>"100100110",
  24433=>"000111100",
  24434=>"111001011",
  24435=>"000000000",
  24436=>"111111111",
  24437=>"000000100",
  24438=>"000000000",
  24439=>"000001111",
  24440=>"000000000",
  24441=>"111111111",
  24442=>"111111100",
  24443=>"110111001",
  24444=>"011111111",
  24445=>"111111111",
  24446=>"000000011",
  24447=>"100000011",
  24448=>"011001011",
  24449=>"111101111",
  24450=>"001011011",
  24451=>"111000000",
  24452=>"010100111",
  24453=>"000000100",
  24454=>"010110111",
  24455=>"111101101",
  24456=>"111111100",
  24457=>"000000000",
  24458=>"000000001",
  24459=>"000000000",
  24460=>"111000111",
  24461=>"100100111",
  24462=>"111111111",
  24463=>"000111111",
  24464=>"000111111",
  24465=>"111111100",
  24466=>"111111111",
  24467=>"000001001",
  24468=>"000000000",
  24469=>"111101001",
  24470=>"111111111",
  24471=>"000011111",
  24472=>"000111111",
  24473=>"000000000",
  24474=>"000100110",
  24475=>"000000010",
  24476=>"110000100",
  24477=>"000000111",
  24478=>"101000000",
  24479=>"000011111",
  24480=>"000000110",
  24481=>"001011001",
  24482=>"001011011",
  24483=>"111011010",
  24484=>"000001001",
  24485=>"110110000",
  24486=>"111111111",
  24487=>"000000000",
  24488=>"111110100",
  24489=>"101111111",
  24490=>"111000000",
  24491=>"111111111",
  24492=>"000000000",
  24493=>"000000001",
  24494=>"000000011",
  24495=>"111111111",
  24496=>"000001011",
  24497=>"010000000",
  24498=>"111001001",
  24499=>"000000000",
  24500=>"111111111",
  24501=>"111111001",
  24502=>"111111111",
  24503=>"000011111",
  24504=>"011011111",
  24505=>"000010110",
  24506=>"111111111",
  24507=>"100110110",
  24508=>"000000000",
  24509=>"001011011",
  24510=>"000000000",
  24511=>"001011011",
  24512=>"000000000",
  24513=>"000000000",
  24514=>"000000000",
  24515=>"111000000",
  24516=>"001001001",
  24517=>"000100000",
  24518=>"000001111",
  24519=>"111001101",
  24520=>"011111000",
  24521=>"000001111",
  24522=>"001111111",
  24523=>"000111111",
  24524=>"011011111",
  24525=>"000000000",
  24526=>"000101111",
  24527=>"000100111",
  24528=>"000000111",
  24529=>"111111000",
  24530=>"111111101",
  24531=>"000000000",
  24532=>"111111111",
  24533=>"100111110",
  24534=>"000000000",
  24535=>"011001011",
  24536=>"000000000",
  24537=>"000000000",
  24538=>"111111111",
  24539=>"000000000",
  24540=>"110110111",
  24541=>"101111111",
  24542=>"100000000",
  24543=>"011011011",
  24544=>"000000000",
  24545=>"111111111",
  24546=>"000000111",
  24547=>"111111110",
  24548=>"001111111",
  24549=>"000100111",
  24550=>"100100110",
  24551=>"000000000",
  24552=>"000000000",
  24553=>"101000000",
  24554=>"000000000",
  24555=>"011011001",
  24556=>"111111100",
  24557=>"000100110",
  24558=>"000000000",
  24559=>"010000000",
  24560=>"000000111",
  24561=>"000001110",
  24562=>"001001001",
  24563=>"111111111",
  24564=>"000110100",
  24565=>"110110100",
  24566=>"111111111",
  24567=>"000110110",
  24568=>"100000000",
  24569=>"111011100",
  24570=>"111111111",
  24571=>"111111111",
  24572=>"000011001",
  24573=>"000000000",
  24574=>"000000000",
  24575=>"000000000",
  24576=>"101001000",
  24577=>"111111100",
  24578=>"111111111",
  24579=>"110110000",
  24580=>"110100100",
  24581=>"001001000",
  24582=>"000000000",
  24583=>"111111111",
  24584=>"111111111",
  24585=>"110111100",
  24586=>"111111010",
  24587=>"000111111",
  24588=>"000000010",
  24589=>"000000110",
  24590=>"110000000",
  24591=>"000000000",
  24592=>"000000000",
  24593=>"000000000",
  24594=>"111111111",
  24595=>"111001100",
  24596=>"111111100",
  24597=>"000100011",
  24598=>"010000000",
  24599=>"011111110",
  24600=>"101000000",
  24601=>"100101100",
  24602=>"000000000",
  24603=>"011111111",
  24604=>"111111111",
  24605=>"110010000",
  24606=>"111000000",
  24607=>"000000101",
  24608=>"000001000",
  24609=>"111111111",
  24610=>"111011000",
  24611=>"110110111",
  24612=>"000000000",
  24613=>"100000111",
  24614=>"011000011",
  24615=>"000000000",
  24616=>"111111110",
  24617=>"000000000",
  24618=>"111111100",
  24619=>"000000000",
  24620=>"000111001",
  24621=>"111000000",
  24622=>"111111111",
  24623=>"100001111",
  24624=>"001000000",
  24625=>"000101111",
  24626=>"001000000",
  24627=>"111100100",
  24628=>"111111001",
  24629=>"001001011",
  24630=>"111111111",
  24631=>"001111111",
  24632=>"000000101",
  24633=>"111111101",
  24634=>"000000000",
  24635=>"111111111",
  24636=>"111101111",
  24637=>"111010000",
  24638=>"000000000",
  24639=>"101100100",
  24640=>"111111101",
  24641=>"001011000",
  24642=>"111111111",
  24643=>"010111111",
  24644=>"011111000",
  24645=>"000100101",
  24646=>"000110111",
  24647=>"111000001",
  24648=>"100100010",
  24649=>"111111111",
  24650=>"011111111",
  24651=>"111110111",
  24652=>"100111111",
  24653=>"000111111",
  24654=>"010110111",
  24655=>"000000000",
  24656=>"011111111",
  24657=>"010010010",
  24658=>"100111111",
  24659=>"100101100",
  24660=>"111111111",
  24661=>"110010000",
  24662=>"011010011",
  24663=>"111110110",
  24664=>"100110110",
  24665=>"000000111",
  24666=>"000000011",
  24667=>"000000000",
  24668=>"011111111",
  24669=>"000000000",
  24670=>"111000000",
  24671=>"110100011",
  24672=>"000001111",
  24673=>"000000000",
  24674=>"011011000",
  24675=>"000000111",
  24676=>"011001001",
  24677=>"000000000",
  24678=>"111000111",
  24679=>"000000000",
  24680=>"110000000",
  24681=>"000010111",
  24682=>"000011011",
  24683=>"110010000",
  24684=>"111011000",
  24685=>"011111111",
  24686=>"111111111",
  24687=>"110000101",
  24688=>"100100111",
  24689=>"101001111",
  24690=>"111111101",
  24691=>"111101000",
  24692=>"001111111",
  24693=>"101000000",
  24694=>"000000000",
  24695=>"000101000",
  24696=>"000000000",
  24697=>"100000000",
  24698=>"000000000",
  24699=>"000010011",
  24700=>"111111011",
  24701=>"000000000",
  24702=>"111111111",
  24703=>"000000000",
  24704=>"101111101",
  24705=>"111111000",
  24706=>"110110111",
  24707=>"000001001",
  24708=>"011000100",
  24709=>"000000000",
  24710=>"000010000",
  24711=>"111111111",
  24712=>"000000000",
  24713=>"111111101",
  24714=>"111101000",
  24715=>"000000000",
  24716=>"111110000",
  24717=>"111111001",
  24718=>"111111111",
  24719=>"111111000",
  24720=>"111111111",
  24721=>"000000001",
  24722=>"000000000",
  24723=>"000000101",
  24724=>"001001000",
  24725=>"000000111",
  24726=>"000000001",
  24727=>"011111011",
  24728=>"111110000",
  24729=>"111111001",
  24730=>"000000000",
  24731=>"100100111",
  24732=>"000000000",
  24733=>"101101100",
  24734=>"111000000",
  24735=>"010100100",
  24736=>"000000000",
  24737=>"111111111",
  24738=>"111010001",
  24739=>"101101111",
  24740=>"111111111",
  24741=>"011010110",
  24742=>"101001011",
  24743=>"000000101",
  24744=>"111111111",
  24745=>"000000000",
  24746=>"000000000",
  24747=>"001000101",
  24748=>"001001001",
  24749=>"111111110",
  24750=>"100000000",
  24751=>"100101101",
  24752=>"000000000",
  24753=>"101111110",
  24754=>"001011001",
  24755=>"111111111",
  24756=>"111111111",
  24757=>"000010111",
  24758=>"000010111",
  24759=>"000000001",
  24760=>"110100100",
  24761=>"111111111",
  24762=>"111111111",
  24763=>"001001011",
  24764=>"000000000",
  24765=>"000000000",
  24766=>"010011111",
  24767=>"000000001",
  24768=>"000010000",
  24769=>"110000001",
  24770=>"111101110",
  24771=>"000000000",
  24772=>"110110110",
  24773=>"110100110",
  24774=>"111001011",
  24775=>"110110111",
  24776=>"001011001",
  24777=>"001000000",
  24778=>"101101111",
  24779=>"000000100",
  24780=>"010111111",
  24781=>"110010000",
  24782=>"000111111",
  24783=>"101000011",
  24784=>"011000000",
  24785=>"001000111",
  24786=>"111111111",
  24787=>"000000000",
  24788=>"110011000",
  24789=>"001111111",
  24790=>"000000010",
  24791=>"011001000",
  24792=>"100111111",
  24793=>"111111111",
  24794=>"000000000",
  24795=>"000011110",
  24796=>"111101101",
  24797=>"110110100",
  24798=>"011011111",
  24799=>"111000000",
  24800=>"000000000",
  24801=>"000010111",
  24802=>"110000010",
  24803=>"110000000",
  24804=>"110110111",
  24805=>"000000000",
  24806=>"010000000",
  24807=>"011000101",
  24808=>"000000110",
  24809=>"001111111",
  24810=>"111111011",
  24811=>"000000000",
  24812=>"111111111",
  24813=>"100000101",
  24814=>"111001011",
  24815=>"101000000",
  24816=>"111111111",
  24817=>"111100111",
  24818=>"111011011",
  24819=>"111000000",
  24820=>"000000000",
  24821=>"011010100",
  24822=>"000000000",
  24823=>"000000000",
  24824=>"111111111",
  24825=>"111111111",
  24826=>"001111111",
  24827=>"011010001",
  24828=>"001011000",
  24829=>"000000000",
  24830=>"000000000",
  24831=>"000111111",
  24832=>"000000000",
  24833=>"001000000",
  24834=>"100111111",
  24835=>"111100000",
  24836=>"000111111",
  24837=>"000101111",
  24838=>"000000000",
  24839=>"001011011",
  24840=>"000000000",
  24841=>"111111111",
  24842=>"111110110",
  24843=>"011000000",
  24844=>"101101111",
  24845=>"000000001",
  24846=>"111111111",
  24847=>"111111111",
  24848=>"000000111",
  24849=>"111101111",
  24850=>"000000000",
  24851=>"111111000",
  24852=>"000000000",
  24853=>"110011111",
  24854=>"101001000",
  24855=>"000101000",
  24856=>"111111111",
  24857=>"111111111",
  24858=>"000000000",
  24859=>"001001011",
  24860=>"111111111",
  24861=>"000000000",
  24862=>"000000000",
  24863=>"111000110",
  24864=>"001001001",
  24865=>"101101101",
  24866=>"000111010",
  24867=>"101001000",
  24868=>"001101101",
  24869=>"111111001",
  24870=>"111111110",
  24871=>"011101111",
  24872=>"000000100",
  24873=>"101111001",
  24874=>"001111111",
  24875=>"000000010",
  24876=>"000000000",
  24877=>"100100000",
  24878=>"011111111",
  24879=>"000000000",
  24880=>"000001000",
  24881=>"000001111",
  24882=>"000000000",
  24883=>"000000110",
  24884=>"010111010",
  24885=>"000000110",
  24886=>"000000011",
  24887=>"000000000",
  24888=>"000000000",
  24889=>"000010000",
  24890=>"111110110",
  24891=>"000000000",
  24892=>"111110110",
  24893=>"111111111",
  24894=>"111111111",
  24895=>"011000000",
  24896=>"100000000",
  24897=>"001100000",
  24898=>"001001100",
  24899=>"000000000",
  24900=>"011011000",
  24901=>"000011111",
  24902=>"000100100",
  24903=>"100000000",
  24904=>"111111111",
  24905=>"011000101",
  24906=>"001000100",
  24907=>"111111110",
  24908=>"111000100",
  24909=>"000000000",
  24910=>"111111111",
  24911=>"100100100",
  24912=>"100111111",
  24913=>"100111110",
  24914=>"111000000",
  24915=>"001000000",
  24916=>"100000000",
  24917=>"011111011",
  24918=>"111000000",
  24919=>"000000100",
  24920=>"110110110",
  24921=>"000000000",
  24922=>"111111111",
  24923=>"000111010",
  24924=>"110110110",
  24925=>"111111111",
  24926=>"111111111",
  24927=>"011011010",
  24928=>"000000000",
  24929=>"000000000",
  24930=>"011000000",
  24931=>"000000001",
  24932=>"100110000",
  24933=>"111111111",
  24934=>"101001001",
  24935=>"111010111",
  24936=>"111101100",
  24937=>"000100100",
  24938=>"111111111",
  24939=>"100000001",
  24940=>"100100100",
  24941=>"100000010",
  24942=>"000000001",
  24943=>"111100101",
  24944=>"111000110",
  24945=>"111011111",
  24946=>"000000111",
  24947=>"100000100",
  24948=>"000000100",
  24949=>"000000100",
  24950=>"000000001",
  24951=>"110110000",
  24952=>"000000101",
  24953=>"000100101",
  24954=>"000010000",
  24955=>"100000000",
  24956=>"101101100",
  24957=>"111100110",
  24958=>"010010000",
  24959=>"111111100",
  24960=>"000000000",
  24961=>"000000000",
  24962=>"001001000",
  24963=>"000000000",
  24964=>"000000101",
  24965=>"000000000",
  24966=>"001001111",
  24967=>"000000000",
  24968=>"000111111",
  24969=>"110100000",
  24970=>"100000001",
  24971=>"011111011",
  24972=>"111111111",
  24973=>"100111101",
  24974=>"100000000",
  24975=>"111101100",
  24976=>"000000000",
  24977=>"000000110",
  24978=>"010111111",
  24979=>"111001001",
  24980=>"000011010",
  24981=>"000000000",
  24982=>"000000000",
  24983=>"000111110",
  24984=>"110100000",
  24985=>"111111111",
  24986=>"000000111",
  24987=>"000110100",
  24988=>"000000000",
  24989=>"000000101",
  24990=>"001000000",
  24991=>"000000111",
  24992=>"000000000",
  24993=>"001001001",
  24994=>"000100111",
  24995=>"111111111",
  24996=>"110111011",
  24997=>"011111011",
  24998=>"100100000",
  24999=>"110111111",
  25000=>"111111110",
  25001=>"000000000",
  25002=>"000000000",
  25003=>"001111111",
  25004=>"000000000",
  25005=>"000000111",
  25006=>"111111111",
  25007=>"111111111",
  25008=>"111111000",
  25009=>"000111111",
  25010=>"110100111",
  25011=>"000000000",
  25012=>"111111111",
  25013=>"110110000",
  25014=>"111111111",
  25015=>"000000000",
  25016=>"000000010",
  25017=>"000000000",
  25018=>"000000100",
  25019=>"000110111",
  25020=>"111111000",
  25021=>"110010000",
  25022=>"111000000",
  25023=>"111011011",
  25024=>"100000100",
  25025=>"111111111",
  25026=>"111111111",
  25027=>"111101101",
  25028=>"001111111",
  25029=>"111100001",
  25030=>"000000100",
  25031=>"000010011",
  25032=>"111111110",
  25033=>"111111010",
  25034=>"010000111",
  25035=>"000000000",
  25036=>"111111111",
  25037=>"111111111",
  25038=>"111111000",
  25039=>"111111111",
  25040=>"100101111",
  25041=>"101100100",
  25042=>"000000000",
  25043=>"111111111",
  25044=>"100000000",
  25045=>"000000000",
  25046=>"110100000",
  25047=>"001000001",
  25048=>"000000000",
  25049=>"000000000",
  25050=>"000000111",
  25051=>"111110000",
  25052=>"001001111",
  25053=>"111000000",
  25054=>"011000000",
  25055=>"111110110",
  25056=>"000000000",
  25057=>"111100101",
  25058=>"000011111",
  25059=>"000000000",
  25060=>"111000000",
  25061=>"011111010",
  25062=>"000011011",
  25063=>"001000101",
  25064=>"111110111",
  25065=>"000110010",
  25066=>"000000000",
  25067=>"101101101",
  25068=>"001000000",
  25069=>"111111011",
  25070=>"111111111",
  25071=>"001000000",
  25072=>"101111001",
  25073=>"000001000",
  25074=>"001000000",
  25075=>"111000000",
  25076=>"100111110",
  25077=>"000000011",
  25078=>"111001000",
  25079=>"001111110",
  25080=>"111111011",
  25081=>"111111011",
  25082=>"000001001",
  25083=>"000000001",
  25084=>"000000000",
  25085=>"111111111",
  25086=>"001111111",
  25087=>"000000111",
  25088=>"001101011",
  25089=>"111111111",
  25090=>"100000000",
  25091=>"101111111",
  25092=>"001000001",
  25093=>"000000000",
  25094=>"111111111",
  25095=>"011111111",
  25096=>"111111000",
  25097=>"000101111",
  25098=>"011101000",
  25099=>"111111001",
  25100=>"011001001",
  25101=>"001100111",
  25102=>"110111111",
  25103=>"101000001",
  25104=>"001000000",
  25105=>"111111111",
  25106=>"001000010",
  25107=>"111111111",
  25108=>"110000000",
  25109=>"111101000",
  25110=>"000000010",
  25111=>"110000000",
  25112=>"000000000",
  25113=>"110111111",
  25114=>"000000000",
  25115=>"001000000",
  25116=>"000001000",
  25117=>"000000111",
  25118=>"110111001",
  25119=>"100100100",
  25120=>"001000000",
  25121=>"110100000",
  25122=>"000001111",
  25123=>"011111000",
  25124=>"101111111",
  25125=>"111111111",
  25126=>"111111111",
  25127=>"110111100",
  25128=>"111111111",
  25129=>"111111111",
  25130=>"101111000",
  25131=>"000111111",
  25132=>"111110111",
  25133=>"011111000",
  25134=>"000110111",
  25135=>"001000001",
  25136=>"000101001",
  25137=>"001000001",
  25138=>"000000100",
  25139=>"010001000",
  25140=>"001000000",
  25141=>"100000000",
  25142=>"011000000",
  25143=>"000100110",
  25144=>"110000000",
  25145=>"100100111",
  25146=>"011001111",
  25147=>"011011000",
  25148=>"111011000",
  25149=>"000000110",
  25150=>"011011111",
  25151=>"100000000",
  25152=>"111000000",
  25153=>"000011010",
  25154=>"000011111",
  25155=>"111101111",
  25156=>"001001011",
  25157=>"011000100",
  25158=>"000000000",
  25159=>"000000000",
  25160=>"010010010",
  25161=>"111000000",
  25162=>"000111101",
  25163=>"111111111",
  25164=>"100100110",
  25165=>"100000111",
  25166=>"000110110",
  25167=>"000000100",
  25168=>"000000000",
  25169=>"001001001",
  25170=>"000000000",
  25171=>"011011011",
  25172=>"111111111",
  25173=>"110000010",
  25174=>"111110111",
  25175=>"001000000",
  25176=>"111001011",
  25177=>"000000111",
  25178=>"111111110",
  25179=>"111111111",
  25180=>"111111111",
  25181=>"000100111",
  25182=>"111111111",
  25183=>"110110110",
  25184=>"000000111",
  25185=>"000000100",
  25186=>"111000011",
  25187=>"001010011",
  25188=>"111011000",
  25189=>"100111101",
  25190=>"001000111",
  25191=>"111111111",
  25192=>"100000111",
  25193=>"110111011",
  25194=>"110111111",
  25195=>"111111111",
  25196=>"111111111",
  25197=>"000000000",
  25198=>"000011111",
  25199=>"000100110",
  25200=>"100000000",
  25201=>"111111111",
  25202=>"001000000",
  25203=>"111011000",
  25204=>"001000101",
  25205=>"111000000",
  25206=>"000000000",
  25207=>"111111111",
  25208=>"000000001",
  25209=>"001000000",
  25210=>"010010000",
  25211=>"111111111",
  25212=>"000000000",
  25213=>"000000110",
  25214=>"000000110",
  25215=>"000000000",
  25216=>"000000000",
  25217=>"000000000",
  25218=>"111000001",
  25219=>"000111111",
  25220=>"111001001",
  25221=>"110111011",
  25222=>"010111111",
  25223=>"000000000",
  25224=>"000000000",
  25225=>"011011011",
  25226=>"100100000",
  25227=>"000100111",
  25228=>"000000001",
  25229=>"000101101",
  25230=>"111111111",
  25231=>"011000100",
  25232=>"000000000",
  25233=>"000000000",
  25234=>"111000001",
  25235=>"111000000",
  25236=>"001000101",
  25237=>"001000000",
  25238=>"110100111",
  25239=>"001001011",
  25240=>"001000111",
  25241=>"111000111",
  25242=>"111111111",
  25243=>"000011011",
  25244=>"100000011",
  25245=>"011001000",
  25246=>"100000000",
  25247=>"111111111",
  25248=>"110100000",
  25249=>"111000000",
  25250=>"100000011",
  25251=>"011000000",
  25252=>"111111110",
  25253=>"000000111",
  25254=>"000000000",
  25255=>"001000001",
  25256=>"010110110",
  25257=>"100111111",
  25258=>"111111000",
  25259=>"100110111",
  25260=>"111010111",
  25261=>"000011011",
  25262=>"001011111",
  25263=>"000000001",
  25264=>"000111111",
  25265=>"111101100",
  25266=>"000001000",
  25267=>"000000000",
  25268=>"111111111",
  25269=>"000110110",
  25270=>"001001111",
  25271=>"001001000",
  25272=>"000000000",
  25273=>"001000011",
  25274=>"010000000",
  25275=>"000000010",
  25276=>"001011111",
  25277=>"000000000",
  25278=>"000110000",
  25279=>"100000100",
  25280=>"111000000",
  25281=>"111001001",
  25282=>"111000000",
  25283=>"000111110",
  25284=>"001000000",
  25285=>"101001000",
  25286=>"011111111",
  25287=>"101000000",
  25288=>"011010000",
  25289=>"000111111",
  25290=>"001001011",
  25291=>"000000000",
  25292=>"111111001",
  25293=>"011001000",
  25294=>"111100111",
  25295=>"000000000",
  25296=>"111111111",
  25297=>"011011011",
  25298=>"111000111",
  25299=>"111101000",
  25300=>"101101101",
  25301=>"111111110",
  25302=>"000000010",
  25303=>"001000001",
  25304=>"000000000",
  25305=>"001001011",
  25306=>"000000111",
  25307=>"111111001",
  25308=>"011011111",
  25309=>"000000100",
  25310=>"001011111",
  25311=>"101101100",
  25312=>"011011111",
  25313=>"000000010",
  25314=>"001001011",
  25315=>"111110111",
  25316=>"001000000",
  25317=>"111111011",
  25318=>"000000000",
  25319=>"101000000",
  25320=>"110111010",
  25321=>"000000000",
  25322=>"111111111",
  25323=>"111111111",
  25324=>"000000111",
  25325=>"000000000",
  25326=>"100111111",
  25327=>"000000000",
  25328=>"000001001",
  25329=>"100000000",
  25330=>"111111111",
  25331=>"000100000",
  25332=>"111111111",
  25333=>"111011010",
  25334=>"100000011",
  25335=>"111111110",
  25336=>"001011001",
  25337=>"111111111",
  25338=>"000110111",
  25339=>"000011111",
  25340=>"111111111",
  25341=>"100100110",
  25342=>"110100111",
  25343=>"001000000",
  25344=>"000000100",
  25345=>"000000000",
  25346=>"101101111",
  25347=>"111100010",
  25348=>"111111111",
  25349=>"111000110",
  25350=>"111111111",
  25351=>"101111111",
  25352=>"010000111",
  25353=>"000000000",
  25354=>"111101000",
  25355=>"001000011",
  25356=>"000000110",
  25357=>"000000001",
  25358=>"001000000",
  25359=>"010000000",
  25360=>"000001001",
  25361=>"001011000",
  25362=>"000000000",
  25363=>"001001000",
  25364=>"001001100",
  25365=>"111111000",
  25366=>"000000000",
  25367=>"111111101",
  25368=>"000000000",
  25369=>"100000100",
  25370=>"111111011",
  25371=>"000011000",
  25372=>"101001001",
  25373=>"000001011",
  25374=>"000000000",
  25375=>"100110000",
  25376=>"111111110",
  25377=>"000001001",
  25378=>"100100111",
  25379=>"000000111",
  25380=>"000111111",
  25381=>"001001011",
  25382=>"101100111",
  25383=>"111000100",
  25384=>"011111111",
  25385=>"010011001",
  25386=>"101101001",
  25387=>"010011000",
  25388=>"111011001",
  25389=>"011000001",
  25390=>"000000000",
  25391=>"111111011",
  25392=>"000000000",
  25393=>"110000000",
  25394=>"111111110",
  25395=>"000111111",
  25396=>"000000000",
  25397=>"001001111",
  25398=>"100000011",
  25399=>"000000000",
  25400=>"111111000",
  25401=>"111110000",
  25402=>"111111010",
  25403=>"111111011",
  25404=>"000000010",
  25405=>"000000001",
  25406=>"000000000",
  25407=>"000000001",
  25408=>"010111111",
  25409=>"001100100",
  25410=>"100111001",
  25411=>"000110011",
  25412=>"001011011",
  25413=>"100111111",
  25414=>"111111111",
  25415=>"000001000",
  25416=>"000000000",
  25417=>"011011000",
  25418=>"111001011",
  25419=>"011010000",
  25420=>"011010110",
  25421=>"111111111",
  25422=>"000000000",
  25423=>"111111111",
  25424=>"001000000",
  25425=>"000110110",
  25426=>"111001001",
  25427=>"000000100",
  25428=>"000000000",
  25429=>"101100111",
  25430=>"000000000",
  25431=>"000000100",
  25432=>"111111000",
  25433=>"000000000",
  25434=>"100100100",
  25435=>"000000111",
  25436=>"001111111",
  25437=>"111111101",
  25438=>"111111011",
  25439=>"111111011",
  25440=>"111000000",
  25441=>"000000000",
  25442=>"111111011",
  25443=>"011111111",
  25444=>"011000000",
  25445=>"001000000",
  25446=>"101000000",
  25447=>"111111111",
  25448=>"011011001",
  25449=>"111111000",
  25450=>"100100101",
  25451=>"000000000",
  25452=>"111111110",
  25453=>"011000111",
  25454=>"000100111",
  25455=>"000000000",
  25456=>"111000000",
  25457=>"000010000",
  25458=>"000111111",
  25459=>"001001101",
  25460=>"100100110",
  25461=>"001111111",
  25462=>"111111010",
  25463=>"111011001",
  25464=>"000011111",
  25465=>"111000000",
  25466=>"000110000",
  25467=>"111000000",
  25468=>"000010000",
  25469=>"111111101",
  25470=>"001111111",
  25471=>"111111111",
  25472=>"111011000",
  25473=>"001001001",
  25474=>"110111111",
  25475=>"110111100",
  25476=>"000000111",
  25477=>"000000000",
  25478=>"010110110",
  25479=>"001111111",
  25480=>"000000011",
  25481=>"101100001",
  25482=>"111111011",
  25483=>"000000010",
  25484=>"000000111",
  25485=>"000000010",
  25486=>"101000000",
  25487=>"111000010",
  25488=>"111111010",
  25489=>"000000000",
  25490=>"111111111",
  25491=>"111101111",
  25492=>"111111111",
  25493=>"101111011",
  25494=>"001011111",
  25495=>"110001010",
  25496=>"111101000",
  25497=>"001011011",
  25498=>"000000000",
  25499=>"101000111",
  25500=>"000000000",
  25501=>"110111100",
  25502=>"110110110",
  25503=>"111111111",
  25504=>"110110000",
  25505=>"000100110",
  25506=>"001101111",
  25507=>"110111111",
  25508=>"100000000",
  25509=>"111111111",
  25510=>"011111011",
  25511=>"000000000",
  25512=>"001001001",
  25513=>"000111011",
  25514=>"111111111",
  25515=>"100111111",
  25516=>"110111000",
  25517=>"111101111",
  25518=>"110000000",
  25519=>"100100000",
  25520=>"100111011",
  25521=>"001011011",
  25522=>"001011000",
  25523=>"111100000",
  25524=>"111101000",
  25525=>"000000000",
  25526=>"011111111",
  25527=>"000111111",
  25528=>"100110111",
  25529=>"001011100",
  25530=>"111110110",
  25531=>"011000111",
  25532=>"111111111",
  25533=>"000000000",
  25534=>"010110000",
  25535=>"000000000",
  25536=>"000000101",
  25537=>"011111111",
  25538=>"000000000",
  25539=>"000001011",
  25540=>"011011011",
  25541=>"000000111",
  25542=>"100000000",
  25543=>"001000001",
  25544=>"000000000",
  25545=>"100000100",
  25546=>"000000000",
  25547=>"000000000",
  25548=>"011011000",
  25549=>"000000001",
  25550=>"101001001",
  25551=>"000000010",
  25552=>"001000100",
  25553=>"110111111",
  25554=>"000001111",
  25555=>"001000000",
  25556=>"011001011",
  25557=>"010000111",
  25558=>"000000000",
  25559=>"000000100",
  25560=>"100101111",
  25561=>"100110000",
  25562=>"111111000",
  25563=>"100100111",
  25564=>"000001011",
  25565=>"111001111",
  25566=>"001000000",
  25567=>"111001111",
  25568=>"001001111",
  25569=>"111111111",
  25570=>"101000000",
  25571=>"101111111",
  25572=>"111000000",
  25573=>"100000111",
  25574=>"000000000",
  25575=>"000000110",
  25576=>"001001101",
  25577=>"111000000",
  25578=>"111111001",
  25579=>"100100001",
  25580=>"001111001",
  25581=>"011000001",
  25582=>"001001001",
  25583=>"011111111",
  25584=>"111101111",
  25585=>"100000001",
  25586=>"111111111",
  25587=>"000000000",
  25588=>"111111101",
  25589=>"000101111",
  25590=>"000000011",
  25591=>"000001001",
  25592=>"000000000",
  25593=>"011001100",
  25594=>"011111111",
  25595=>"111000110",
  25596=>"111111111",
  25597=>"111000000",
  25598=>"000000001",
  25599=>"111110011",
  25600=>"110110110",
  25601=>"110100000",
  25602=>"111000100",
  25603=>"110011000",
  25604=>"111111111",
  25605=>"111011111",
  25606=>"111111110",
  25607=>"000010011",
  25608=>"111111111",
  25609=>"111111111",
  25610=>"111111011",
  25611=>"000000000",
  25612=>"111011110",
  25613=>"111111111",
  25614=>"000001111",
  25615=>"111111001",
  25616=>"001000000",
  25617=>"111111011",
  25618=>"111111111",
  25619=>"000000000",
  25620=>"000000000",
  25621=>"000000000",
  25622=>"001000110",
  25623=>"000100111",
  25624=>"001111111",
  25625=>"000000100",
  25626=>"110111100",
  25627=>"011101111",
  25628=>"000000000",
  25629=>"000000000",
  25630=>"111101000",
  25631=>"000000100",
  25632=>"000000000",
  25633=>"111011010",
  25634=>"111111110",
  25635=>"000000000",
  25636=>"000000000",
  25637=>"110011000",
  25638=>"001101111",
  25639=>"000000000",
  25640=>"000000101",
  25641=>"000010110",
  25642=>"110000111",
  25643=>"111111111",
  25644=>"000000000",
  25645=>"011011000",
  25646=>"101101101",
  25647=>"000000000",
  25648=>"011011111",
  25649=>"100110111",
  25650=>"000000100",
  25651=>"000001100",
  25652=>"001101111",
  25653=>"111111000",
  25654=>"111000111",
  25655=>"100000001",
  25656=>"111111111",
  25657=>"000110111",
  25658=>"111111111",
  25659=>"111000011",
  25660=>"000000000",
  25661=>"000000101",
  25662=>"111111011",
  25663=>"001000000",
  25664=>"000001111",
  25665=>"000000001",
  25666=>"000111111",
  25667=>"000000111",
  25668=>"000000000",
  25669=>"000000000",
  25670=>"000000100",
  25671=>"111111111",
  25672=>"111111111",
  25673=>"000110110",
  25674=>"000000000",
  25675=>"111111011",
  25676=>"000111111",
  25677=>"000000100",
  25678=>"101000000",
  25679=>"101001001",
  25680=>"110000010",
  25681=>"111111001",
  25682=>"001111111",
  25683=>"111101111",
  25684=>"101111101",
  25685=>"000000000",
  25686=>"010010110",
  25687=>"110100000",
  25688=>"000000001",
  25689=>"000000100",
  25690=>"111111110",
  25691=>"011011010",
  25692=>"000011011",
  25693=>"000000000",
  25694=>"000000011",
  25695=>"110010001",
  25696=>"111111111",
  25697=>"001001011",
  25698=>"111111001",
  25699=>"101111111",
  25700=>"111111111",
  25701=>"111111110",
  25702=>"111111111",
  25703=>"000000000",
  25704=>"110010000",
  25705=>"110111111",
  25706=>"010111111",
  25707=>"000000000",
  25708=>"111011111",
  25709=>"111111111",
  25710=>"101111111",
  25711=>"000000000",
  25712=>"000000111",
  25713=>"000000000",
  25714=>"111111000",
  25715=>"111011001",
  25716=>"011111111",
  25717=>"111001001",
  25718=>"111111000",
  25719=>"111111111",
  25720=>"000110010",
  25721=>"001000000",
  25722=>"011000001",
  25723=>"010111111",
  25724=>"011011011",
  25725=>"000000000",
  25726=>"000000000",
  25727=>"000000000",
  25728=>"111111111",
  25729=>"100111111",
  25730=>"111111111",
  25731=>"000000100",
  25732=>"010011111",
  25733=>"000100100",
  25734=>"110100101",
  25735=>"001001000",
  25736=>"001111111",
  25737=>"000000000",
  25738=>"111111111",
  25739=>"110110110",
  25740=>"011000000",
  25741=>"000000000",
  25742=>"111111000",
  25743=>"000000000",
  25744=>"111101111",
  25745=>"000000000",
  25746=>"000000000",
  25747=>"100000000",
  25748=>"111111111",
  25749=>"000101110",
  25750=>"000010110",
  25751=>"111101000",
  25752=>"001000100",
  25753=>"011011101",
  25754=>"000000111",
  25755=>"000000000",
  25756=>"110110111",
  25757=>"011001101",
  25758=>"111111111",
  25759=>"000001000",
  25760=>"111111110",
  25761=>"111110000",
  25762=>"111111111",
  25763=>"000000100",
  25764=>"000000000",
  25765=>"000111111",
  25766=>"111101111",
  25767=>"110100000",
  25768=>"000000000",
  25769=>"000101111",
  25770=>"000000000",
  25771=>"001111111",
  25772=>"011011001",
  25773=>"000000001",
  25774=>"000000100",
  25775=>"000111111",
  25776=>"000111111",
  25777=>"000100111",
  25778=>"111111111",
  25779=>"101101111",
  25780=>"101100000",
  25781=>"001001000",
  25782=>"001000000",
  25783=>"111111111",
  25784=>"000000111",
  25785=>"111111111",
  25786=>"111000000",
  25787=>"110000000",
  25788=>"000000000",
  25789=>"011111111",
  25790=>"100100000",
  25791=>"111111100",
  25792=>"111101110",
  25793=>"111111111",
  25794=>"111111111",
  25795=>"000000000",
  25796=>"010111001",
  25797=>"000000000",
  25798=>"111110001",
  25799=>"111000001",
  25800=>"000000010",
  25801=>"111111111",
  25802=>"000000000",
  25803=>"011011011",
  25804=>"111111111",
  25805=>"001001001",
  25806=>"110110110",
  25807=>"000011000",
  25808=>"111111000",
  25809=>"000101101",
  25810=>"110101101",
  25811=>"111110110",
  25812=>"111110100",
  25813=>"000001111",
  25814=>"000000001",
  25815=>"111001111",
  25816=>"000000001",
  25817=>"011111010",
  25818=>"110111111",
  25819=>"111111111",
  25820=>"100101111",
  25821=>"000000110",
  25822=>"110110111",
  25823=>"100000111",
  25824=>"101101000",
  25825=>"000000110",
  25826=>"000000000",
  25827=>"111111111",
  25828=>"110110110",
  25829=>"111110110",
  25830=>"000011111",
  25831=>"000000000",
  25832=>"000000000",
  25833=>"010000000",
  25834=>"000000000",
  25835=>"001000000",
  25836=>"000000000",
  25837=>"000000000",
  25838=>"001001001",
  25839=>"111000000",
  25840=>"000100110",
  25841=>"000000011",
  25842=>"000110111",
  25843=>"001000001",
  25844=>"111111111",
  25845=>"111000100",
  25846=>"111111100",
  25847=>"111011000",
  25848=>"001001001",
  25849=>"111111111",
  25850=>"000000000",
  25851=>"001001001",
  25852=>"000011011",
  25853=>"100110111",
  25854=>"010000000",
  25855=>"001001111",
  25856=>"111100110",
  25857=>"000001011",
  25858=>"000000111",
  25859=>"011010010",
  25860=>"000000101",
  25861=>"000000000",
  25862=>"000000000",
  25863=>"111111110",
  25864=>"111111111",
  25865=>"000000000",
  25866=>"110000000",
  25867=>"000000000",
  25868=>"111111111",
  25869=>"000000010",
  25870=>"000000110",
  25871=>"111111001",
  25872=>"000100000",
  25873=>"111000101",
  25874=>"000000000",
  25875=>"010000110",
  25876=>"000110111",
  25877=>"111111111",
  25878=>"111110000",
  25879=>"100110000",
  25880=>"111001000",
  25881=>"000000110",
  25882=>"000000101",
  25883=>"001001000",
  25884=>"110111110",
  25885=>"110111111",
  25886=>"011000000",
  25887=>"000100111",
  25888=>"100100010",
  25889=>"000000000",
  25890=>"000100111",
  25891=>"110111111",
  25892=>"110110111",
  25893=>"111000000",
  25894=>"000000000",
  25895=>"111111111",
  25896=>"110111111",
  25897=>"000000000",
  25898=>"110110010",
  25899=>"110000000",
  25900=>"100100110",
  25901=>"111001001",
  25902=>"000000000",
  25903=>"000111111",
  25904=>"000000101",
  25905=>"000010001",
  25906=>"100001110",
  25907=>"111111111",
  25908=>"010010011",
  25909=>"011111111",
  25910=>"111011000",
  25911=>"011011000",
  25912=>"111111111",
  25913=>"010000000",
  25914=>"000000000",
  25915=>"111000100",
  25916=>"000000000",
  25917=>"000010111",
  25918=>"010110111",
  25919=>"001111111",
  25920=>"000100100",
  25921=>"111011011",
  25922=>"001101111",
  25923=>"000000010",
  25924=>"010000111",
  25925=>"110110111",
  25926=>"100100111",
  25927=>"001111111",
  25928=>"000000000",
  25929=>"011001001",
  25930=>"000000001",
  25931=>"101000000",
  25932=>"111001000",
  25933=>"000000001",
  25934=>"100000110",
  25935=>"001000000",
  25936=>"100000110",
  25937=>"111101111",
  25938=>"111111001",
  25939=>"000010011",
  25940=>"000000000",
  25941=>"011011111",
  25942=>"000000000",
  25943=>"001000000",
  25944=>"101001111",
  25945=>"000000000",
  25946=>"110110110",
  25947=>"111000100",
  25948=>"000001111",
  25949=>"011011011",
  25950=>"000000000",
  25951=>"000001001",
  25952=>"000111101",
  25953=>"000000000",
  25954=>"111000000",
  25955=>"111111111",
  25956=>"111111110",
  25957=>"101101101",
  25958=>"111110111",
  25959=>"001000111",
  25960=>"000000000",
  25961=>"011000101",
  25962=>"000000001",
  25963=>"000110111",
  25964=>"000010011",
  25965=>"000000000",
  25966=>"111111111",
  25967=>"000001111",
  25968=>"000000001",
  25969=>"111110111",
  25970=>"100110010",
  25971=>"111111111",
  25972=>"110000111",
  25973=>"001001101",
  25974=>"000000101",
  25975=>"000000000",
  25976=>"000000000",
  25977=>"000111000",
  25978=>"111110100",
  25979=>"000000000",
  25980=>"111111111",
  25981=>"111111111",
  25982=>"000000000",
  25983=>"110111111",
  25984=>"001001011",
  25985=>"000000000",
  25986=>"110100000",
  25987=>"111111111",
  25988=>"000000000",
  25989=>"101111111",
  25990=>"111000010",
  25991=>"000001010",
  25992=>"000000000",
  25993=>"000011011",
  25994=>"011000000",
  25995=>"100111111",
  25996=>"100110011",
  25997=>"111111111",
  25998=>"111111110",
  25999=>"000000110",
  26000=>"001001111",
  26001=>"000000000",
  26002=>"000000100",
  26003=>"000000001",
  26004=>"111000000",
  26005=>"000000000",
  26006=>"010110010",
  26007=>"110110110",
  26008=>"111111111",
  26009=>"111111011",
  26010=>"000110011",
  26011=>"100101101",
  26012=>"111111111",
  26013=>"000110110",
  26014=>"111001000",
  26015=>"111111001",
  26016=>"001001011",
  26017=>"111010000",
  26018=>"101000100",
  26019=>"010111111",
  26020=>"111111111",
  26021=>"001000000",
  26022=>"000000111",
  26023=>"001111111",
  26024=>"001001101",
  26025=>"000000011",
  26026=>"111110110",
  26027=>"001001000",
  26028=>"000000010",
  26029=>"000111000",
  26030=>"111001001",
  26031=>"000000000",
  26032=>"000000000",
  26033=>"000111000",
  26034=>"000000000",
  26035=>"111111001",
  26036=>"001000000",
  26037=>"110110010",
  26038=>"111111110",
  26039=>"000000000",
  26040=>"000111111",
  26041=>"010111011",
  26042=>"111111011",
  26043=>"111011111",
  26044=>"011011011",
  26045=>"000000000",
  26046=>"111001000",
  26047=>"110110110",
  26048=>"011011010",
  26049=>"101101000",
  26050=>"111111110",
  26051=>"000000110",
  26052=>"011111111",
  26053=>"110110111",
  26054=>"000000000",
  26055=>"000000111",
  26056=>"000000100",
  26057=>"010000000",
  26058=>"000000111",
  26059=>"000101000",
  26060=>"000011001",
  26061=>"111111111",
  26062=>"001011001",
  26063=>"101000001",
  26064=>"101001100",
  26065=>"111111111",
  26066=>"111111110",
  26067=>"000011001",
  26068=>"000000001",
  26069=>"000000100",
  26070=>"010010010",
  26071=>"111111111",
  26072=>"111011111",
  26073=>"000000110",
  26074=>"000110110",
  26075=>"111000000",
  26076=>"011111111",
  26077=>"101101101",
  26078=>"001000011",
  26079=>"000000000",
  26080=>"000000111",
  26081=>"111010000",
  26082=>"000000011",
  26083=>"111111111",
  26084=>"111111111",
  26085=>"101100111",
  26086=>"000010011",
  26087=>"000000111",
  26088=>"100101101",
  26089=>"111100111",
  26090=>"111000000",
  26091=>"000000000",
  26092=>"111110110",
  26093=>"111111110",
  26094=>"111000000",
  26095=>"101000000",
  26096=>"111011011",
  26097=>"111111111",
  26098=>"000000100",
  26099=>"000101111",
  26100=>"001011000",
  26101=>"011000000",
  26102=>"111001111",
  26103=>"001111000",
  26104=>"000000000",
  26105=>"011011011",
  26106=>"111100110",
  26107=>"110111111",
  26108=>"000001000",
  26109=>"111010010",
  26110=>"000000100",
  26111=>"111001000",
  26112=>"110111101",
  26113=>"000000000",
  26114=>"111101001",
  26115=>"111100000",
  26116=>"000000001",
  26117=>"101001101",
  26118=>"000000000",
  26119=>"111101101",
  26120=>"011111000",
  26121=>"011111111",
  26122=>"000000000",
  26123=>"001111111",
  26124=>"100000000",
  26125=>"111111100",
  26126=>"000000100",
  26127=>"111111001",
  26128=>"000000100",
  26129=>"011000001",
  26130=>"111111111",
  26131=>"111111111",
  26132=>"000000000",
  26133=>"111101101",
  26134=>"010010000",
  26135=>"001001011",
  26136=>"100100000",
  26137=>"111101000",
  26138=>"000000100",
  26139=>"011000100",
  26140=>"110100000",
  26141=>"111111111",
  26142=>"000110100",
  26143=>"011001011",
  26144=>"000000001",
  26145=>"110111111",
  26146=>"001001111",
  26147=>"111111010",
  26148=>"000000110",
  26149=>"111101000",
  26150=>"000000000",
  26151=>"111111000",
  26152=>"111111110",
  26153=>"000001000",
  26154=>"111111101",
  26155=>"010000000",
  26156=>"000000001",
  26157=>"100001001",
  26158=>"000000001",
  26159=>"101111011",
  26160=>"000100000",
  26161=>"001001000",
  26162=>"100100100",
  26163=>"000011001",
  26164=>"100000000",
  26165=>"111100100",
  26166=>"000000111",
  26167=>"010110000",
  26168=>"000000000",
  26169=>"011111111",
  26170=>"101101111",
  26171=>"111100000",
  26172=>"000110110",
  26173=>"111111111",
  26174=>"000000001",
  26175=>"111111001",
  26176=>"011111001",
  26177=>"000000000",
  26178=>"000000000",
  26179=>"111110111",
  26180=>"111011010",
  26181=>"000000000",
  26182=>"000001011",
  26183=>"111111110",
  26184=>"111101001",
  26185=>"000000000",
  26186=>"111111111",
  26187=>"111110110",
  26188=>"000000000",
  26189=>"111111110",
  26190=>"100000111",
  26191=>"011001000",
  26192=>"111111111",
  26193=>"101101100",
  26194=>"110000110",
  26195=>"001101100",
  26196=>"111101001",
  26197=>"100000010",
  26198=>"101000100",
  26199=>"000000001",
  26200=>"001001111",
  26201=>"100100100",
  26202=>"100000111",
  26203=>"111010011",
  26204=>"000001001",
  26205=>"100000000",
  26206=>"111111111",
  26207=>"100000000",
  26208=>"110000000",
  26209=>"000000011",
  26210=>"000100100",
  26211=>"011001001",
  26212=>"111001100",
  26213=>"000110100",
  26214=>"111011110",
  26215=>"011000100",
  26216=>"110111111",
  26217=>"001101111",
  26218=>"110100110",
  26219=>"101110000",
  26220=>"000100100",
  26221=>"000000000",
  26222=>"111111111",
  26223=>"011111010",
  26224=>"011000000",
  26225=>"101101101",
  26226=>"101101111",
  26227=>"010011111",
  26228=>"000000000",
  26229=>"000010110",
  26230=>"000001001",
  26231=>"100101111",
  26232=>"010111111",
  26233=>"011111111",
  26234=>"011001000",
  26235=>"011111111",
  26236=>"110100100",
  26237=>"000100000",
  26238=>"110011100",
  26239=>"000000001",
  26240=>"000101111",
  26241=>"110111111",
  26242=>"000000011",
  26243=>"000010011",
  26244=>"000000010",
  26245=>"001000000",
  26246=>"000001000",
  26247=>"111111110",
  26248=>"100101001",
  26249=>"000000000",
  26250=>"000000000",
  26251=>"101111000",
  26252=>"000000001",
  26253=>"111111110",
  26254=>"111111001",
  26255=>"000000011",
  26256=>"000111110",
  26257=>"011111111",
  26258=>"000000010",
  26259=>"111111111",
  26260=>"000000001",
  26261=>"000000101",
  26262=>"000000001",
  26263=>"111110100",
  26264=>"001000000",
  26265=>"000100111",
  26266=>"000110111",
  26267=>"000000011",
  26268=>"001111111",
  26269=>"000110111",
  26270=>"111100011",
  26271=>"000100011",
  26272=>"001000001",
  26273=>"000000101",
  26274=>"101001100",
  26275=>"000001000",
  26276=>"111011111",
  26277=>"111101011",
  26278=>"000001000",
  26279=>"011000000",
  26280=>"000000001",
  26281=>"000000000",
  26282=>"001111111",
  26283=>"111111111",
  26284=>"010000000",
  26285=>"100110110",
  26286=>"111111111",
  26287=>"000011100",
  26288=>"000000101",
  26289=>"100110100",
  26290=>"111101111",
  26291=>"010000010",
  26292=>"000000000",
  26293=>"111000000",
  26294=>"001111001",
  26295=>"001111111",
  26296=>"110100100",
  26297=>"111100110",
  26298=>"001001001",
  26299=>"111101001",
  26300=>"111011001",
  26301=>"111111111",
  26302=>"000000001",
  26303=>"111111000",
  26304=>"000000111",
  26305=>"111010000",
  26306=>"000110111",
  26307=>"000000001",
  26308=>"111101111",
  26309=>"000000011",
  26310=>"011000000",
  26311=>"000000000",
  26312=>"110000000",
  26313=>"000000000",
  26314=>"001101100",
  26315=>"111101101",
  26316=>"111101101",
  26317=>"111111101",
  26318=>"110011111",
  26319=>"001000001",
  26320=>"111000000",
  26321=>"000000110",
  26322=>"000111111",
  26323=>"001001000",
  26324=>"100100111",
  26325=>"111111111",
  26326=>"010111111",
  26327=>"000000000",
  26328=>"000000101",
  26329=>"000110111",
  26330=>"000000000",
  26331=>"111111011",
  26332=>"110110110",
  26333=>"000000000",
  26334=>"000010111",
  26335=>"111011010",
  26336=>"000000001",
  26337=>"100110011",
  26338=>"111111000",
  26339=>"111111011",
  26340=>"111111111",
  26341=>"001001000",
  26342=>"111111111",
  26343=>"110110110",
  26344=>"000000000",
  26345=>"111111101",
  26346=>"111110111",
  26347=>"011111010",
  26348=>"010011000",
  26349=>"000000000",
  26350=>"100100100",
  26351=>"000000000",
  26352=>"111111011",
  26353=>"011000011",
  26354=>"001001111",
  26355=>"000000001",
  26356=>"000110011",
  26357=>"000011001",
  26358=>"000000011",
  26359=>"101101111",
  26360=>"111111111",
  26361=>"000000000",
  26362=>"000000000",
  26363=>"100101101",
  26364=>"000111111",
  26365=>"000000000",
  26366=>"011111111",
  26367=>"000000000",
  26368=>"011001011",
  26369=>"000000000",
  26370=>"000111111",
  26371=>"001000000",
  26372=>"011001100",
  26373=>"111100110",
  26374=>"000000100",
  26375=>"111111100",
  26376=>"111111010",
  26377=>"000000000",
  26378=>"111111111",
  26379=>"000000101",
  26380=>"001000000",
  26381=>"100101101",
  26382=>"110101111",
  26383=>"000100100",
  26384=>"001011000",
  26385=>"001000001",
  26386=>"000000101",
  26387=>"000000000",
  26388=>"000001111",
  26389=>"111011111",
  26390=>"110110110",
  26391=>"000000111",
  26392=>"111111110",
  26393=>"011010010",
  26394=>"000000111",
  26395=>"111111111",
  26396=>"001111111",
  26397=>"110000000",
  26398=>"001001001",
  26399=>"111011100",
  26400=>"100000100",
  26401=>"111011111",
  26402=>"100011111",
  26403=>"111111011",
  26404=>"011010000",
  26405=>"001111101",
  26406=>"100000100",
  26407=>"010011111",
  26408=>"111101100",
  26409=>"000001101",
  26410=>"100000000",
  26411=>"000000000",
  26412=>"111111101",
  26413=>"011111111",
  26414=>"100111110",
  26415=>"111011000",
  26416=>"111111101",
  26417=>"000000000",
  26418=>"111111111",
  26419=>"000010111",
  26420=>"010001000",
  26421=>"011111101",
  26422=>"000000000",
  26423=>"000100111",
  26424=>"000100111",
  26425=>"000000100",
  26426=>"000000000",
  26427=>"000000001",
  26428=>"000000000",
  26429=>"100110100",
  26430=>"010010000",
  26431=>"011011011",
  26432=>"000000111",
  26433=>"111111110",
  26434=>"000110000",
  26435=>"000000001",
  26436=>"111100000",
  26437=>"000000000",
  26438=>"000000000",
  26439=>"111101101",
  26440=>"000000000",
  26441=>"000000000",
  26442=>"000111111",
  26443=>"001110010",
  26444=>"000011111",
  26445=>"100110000",
  26446=>"111110111",
  26447=>"000101111",
  26448=>"001001001",
  26449=>"111011111",
  26450=>"000000000",
  26451=>"111111111",
  26452=>"110100100",
  26453=>"011011010",
  26454=>"110010010",
  26455=>"000000011",
  26456=>"000000100",
  26457=>"111111110",
  26458=>"111111100",
  26459=>"111111111",
  26460=>"001000000",
  26461=>"111111011",
  26462=>"000001101",
  26463=>"110111111",
  26464=>"110011011",
  26465=>"011011111",
  26466=>"101011011",
  26467=>"100000000",
  26468=>"100100100",
  26469=>"111111000",
  26470=>"100100000",
  26471=>"000000111",
  26472=>"000000000",
  26473=>"000000100",
  26474=>"011111111",
  26475=>"000001001",
  26476=>"000000001",
  26477=>"011001011",
  26478=>"000000000",
  26479=>"000000000",
  26480=>"000000100",
  26481=>"000000011",
  26482=>"000000001",
  26483=>"000000111",
  26484=>"011011100",
  26485=>"000000101",
  26486=>"000000000",
  26487=>"000010111",
  26488=>"000000011",
  26489=>"000000000",
  26490=>"000000111",
  26491=>"101101101",
  26492=>"011011011",
  26493=>"000001001",
  26494=>"000000000",
  26495=>"000000100",
  26496=>"110110111",
  26497=>"001000011",
  26498=>"000000111",
  26499=>"000000000",
  26500=>"000000000",
  26501=>"111111010",
  26502=>"100100110",
  26503=>"111011000",
  26504=>"000000110",
  26505=>"011011011",
  26506=>"001001111",
  26507=>"111111000",
  26508=>"111111111",
  26509=>"000101001",
  26510=>"100100111",
  26511=>"000011011",
  26512=>"001000000",
  26513=>"111110100",
  26514=>"101101111",
  26515=>"011001011",
  26516=>"111111111",
  26517=>"000010011",
  26518=>"010000110",
  26519=>"110110110",
  26520=>"111111111",
  26521=>"111010010",
  26522=>"000000000",
  26523=>"100000000",
  26524=>"111110100",
  26525=>"110111001",
  26526=>"111101101",
  26527=>"000000000",
  26528=>"001001000",
  26529=>"101111111",
  26530=>"000110001",
  26531=>"111111001",
  26532=>"000000110",
  26533=>"111111101",
  26534=>"000000000",
  26535=>"110110111",
  26536=>"110111111",
  26537=>"011101111",
  26538=>"111111011",
  26539=>"100100101",
  26540=>"111111001",
  26541=>"001001011",
  26542=>"011000000",
  26543=>"110100000",
  26544=>"110010010",
  26545=>"101101111",
  26546=>"100000100",
  26547=>"000000000",
  26548=>"111111000",
  26549=>"101001001",
  26550=>"000100110",
  26551=>"000000000",
  26552=>"000000010",
  26553=>"000000100",
  26554=>"010000000",
  26555=>"000111111",
  26556=>"001001001",
  26557=>"000000100",
  26558=>"100000001",
  26559=>"110110100",
  26560=>"000000000",
  26561=>"101001000",
  26562=>"111011111",
  26563=>"001001001",
  26564=>"111100000",
  26565=>"001000000",
  26566=>"000000000",
  26567=>"101100101",
  26568=>"000000001",
  26569=>"111111000",
  26570=>"000000001",
  26571=>"001011001",
  26572=>"110110111",
  26573=>"110111111",
  26574=>"000000011",
  26575=>"000000000",
  26576=>"111011000",
  26577=>"011011000",
  26578=>"111111001",
  26579=>"111111111",
  26580=>"100001001",
  26581=>"111110000",
  26582=>"101101101",
  26583=>"100100000",
  26584=>"100000001",
  26585=>"011001101",
  26586=>"011010000",
  26587=>"111111111",
  26588=>"111111001",
  26589=>"000000000",
  26590=>"111111111",
  26591=>"010100000",
  26592=>"000000000",
  26593=>"000000000",
  26594=>"011011000",
  26595=>"111111111",
  26596=>"000000000",
  26597=>"000000000",
  26598=>"000000000",
  26599=>"000000000",
  26600=>"000000000",
  26601=>"001111101",
  26602=>"011011110",
  26603=>"101111111",
  26604=>"111111111",
  26605=>"011011011",
  26606=>"100101001",
  26607=>"000111111",
  26608=>"101000011",
  26609=>"000000101",
  26610=>"111111111",
  26611=>"000000000",
  26612=>"111111111",
  26613=>"000000000",
  26614=>"010111111",
  26615=>"100110110",
  26616=>"001000000",
  26617=>"001001001",
  26618=>"100010110",
  26619=>"111000010",
  26620=>"001001111",
  26621=>"110111110",
  26622=>"001000000",
  26623=>"000000100",
  26624=>"001111001",
  26625=>"011101000",
  26626=>"000000000",
  26627=>"001000000",
  26628=>"111111111",
  26629=>"111111111",
  26630=>"000000000",
  26631=>"111000000",
  26632=>"000000000",
  26633=>"111010000",
  26634=>"111111111",
  26635=>"011001000",
  26636=>"111111000",
  26637=>"111111100",
  26638=>"100100100",
  26639=>"011111011",
  26640=>"000000111",
  26641=>"011011111",
  26642=>"111111111",
  26643=>"011111001",
  26644=>"000101111",
  26645=>"000001111",
  26646=>"111111111",
  26647=>"011001000",
  26648=>"111111111",
  26649=>"010010000",
  26650=>"011001101",
  26651=>"110000000",
  26652=>"000000000",
  26653=>"111111001",
  26654=>"010011000",
  26655=>"000001011",
  26656=>"100000000",
  26657=>"110110110",
  26658=>"110111000",
  26659=>"000000000",
  26660=>"111111111",
  26661=>"011111111",
  26662=>"100111101",
  26663=>"000111111",
  26664=>"110001101",
  26665=>"000000000",
  26666=>"000000000",
  26667=>"111111110",
  26668=>"111111111",
  26669=>"001010000",
  26670=>"000000001",
  26671=>"110111111",
  26672=>"111111111",
  26673=>"111011011",
  26674=>"011111111",
  26675=>"000000000",
  26676=>"011001001",
  26677=>"011000000",
  26678=>"000000000",
  26679=>"001100111",
  26680=>"000111111",
  26681=>"111111110",
  26682=>"110111110",
  26683=>"000111000",
  26684=>"001001001",
  26685=>"000000000",
  26686=>"111011000",
  26687=>"111111111",
  26688=>"000100110",
  26689=>"000000110",
  26690=>"001000001",
  26691=>"100111111",
  26692=>"000000000",
  26693=>"111111111",
  26694=>"100000000",
  26695=>"111001111",
  26696=>"111111011",
  26697=>"111111000",
  26698=>"100000110",
  26699=>"111111111",
  26700=>"000100100",
  26701=>"000000000",
  26702=>"000000000",
  26703=>"000000000",
  26704=>"000000000",
  26705=>"111111111",
  26706=>"000110111",
  26707=>"000000000",
  26708=>"000000001",
  26709=>"101111011",
  26710=>"000000000",
  26711=>"111101111",
  26712=>"111000000",
  26713=>"111111110",
  26714=>"111111111",
  26715=>"010011110",
  26716=>"110100110",
  26717=>"110110100",
  26718=>"000000100",
  26719=>"000000100",
  26720=>"000000000",
  26721=>"000000000",
  26722=>"001011111",
  26723=>"111111111",
  26724=>"100100100",
  26725=>"111111111",
  26726=>"000001011",
  26727=>"001000000",
  26728=>"000111111",
  26729=>"111111011",
  26730=>"000110111",
  26731=>"000000011",
  26732=>"000000000",
  26733=>"000000000",
  26734=>"000000001",
  26735=>"010000011",
  26736=>"111111111",
  26737=>"000000000",
  26738=>"001001001",
  26739=>"000001000",
  26740=>"000000001",
  26741=>"111110000",
  26742=>"111111111",
  26743=>"000000000",
  26744=>"111001001",
  26745=>"100000000",
  26746=>"111111001",
  26747=>"110000100",
  26748=>"111110111",
  26749=>"111101111",
  26750=>"000001000",
  26751=>"011111011",
  26752=>"000000000",
  26753=>"111111111",
  26754=>"000000000",
  26755=>"000000001",
  26756=>"000000000",
  26757=>"000000100",
  26758=>"000111111",
  26759=>"111000000",
  26760=>"111111000",
  26761=>"100111111",
  26762=>"000000000",
  26763=>"000011010",
  26764=>"000001111",
  26765=>"000000000",
  26766=>"000000100",
  26767=>"010010000",
  26768=>"000000000",
  26769=>"011011000",
  26770=>"000100100",
  26771=>"111111100",
  26772=>"101101001",
  26773=>"111000000",
  26774=>"000000000",
  26775=>"000000000",
  26776=>"001001000",
  26777=>"000000000",
  26778=>"111111111",
  26779=>"000000000",
  26780=>"001100111",
  26781=>"010111111",
  26782=>"011011111",
  26783=>"001000111",
  26784=>"011111101",
  26785=>"110100000",
  26786=>"111101111",
  26787=>"000000011",
  26788=>"000010010",
  26789=>"000001000",
  26790=>"000000000",
  26791=>"000000000",
  26792=>"111111111",
  26793=>"111111111",
  26794=>"111111111",
  26795=>"111111100",
  26796=>"000000000",
  26797=>"000011000",
  26798=>"001111111",
  26799=>"001100111",
  26800=>"111111111",
  26801=>"001000000",
  26802=>"110110110",
  26803=>"000000000",
  26804=>"111100000",
  26805=>"101000000",
  26806=>"001011000",
  26807=>"011110100",
  26808=>"111111111",
  26809=>"111000001",
  26810=>"000010111",
  26811=>"001001001",
  26812=>"111100000",
  26813=>"101111101",
  26814=>"111111001",
  26815=>"011001001",
  26816=>"000000000",
  26817=>"001000111",
  26818=>"000000100",
  26819=>"000111111",
  26820=>"111111111",
  26821=>"100110100",
  26822=>"100100111",
  26823=>"111100000",
  26824=>"000000000",
  26825=>"000000000",
  26826=>"000100111",
  26827=>"111111111",
  26828=>"000011011",
  26829=>"100111111",
  26830=>"101111111",
  26831=>"000000000",
  26832=>"000000000",
  26833=>"111111111",
  26834=>"011011000",
  26835=>"000001111",
  26836=>"000000000",
  26837=>"110110110",
  26838=>"111111111",
  26839=>"101101111",
  26840=>"000110111",
  26841=>"000110100",
  26842=>"000000000",
  26843=>"000000000",
  26844=>"000000000",
  26845=>"000000000",
  26846=>"111111111",
  26847=>"000000000",
  26848=>"111111111",
  26849=>"111111001",
  26850=>"111111111",
  26851=>"000000111",
  26852=>"110111111",
  26853=>"111111001",
  26854=>"111111111",
  26855=>"000100100",
  26856=>"000000000",
  26857=>"000000000",
  26858=>"000000110",
  26859=>"000111111",
  26860=>"010111111",
  26861=>"000111111",
  26862=>"011110111",
  26863=>"111111111",
  26864=>"000111111",
  26865=>"000101111",
  26866=>"110000000",
  26867=>"000001000",
  26868=>"000000000",
  26869=>"000001001",
  26870=>"110100011",
  26871=>"110111111",
  26872=>"000000000",
  26873=>"000000101",
  26874=>"000001001",
  26875=>"101000100",
  26876=>"000000000",
  26877=>"010110110",
  26878=>"111111001",
  26879=>"011111111",
  26880=>"001001000",
  26881=>"110100110",
  26882=>"111111111",
  26883=>"111111110",
  26884=>"111101111",
  26885=>"111100011",
  26886=>"111111111",
  26887=>"000000000",
  26888=>"000001110",
  26889=>"110000000",
  26890=>"111111111",
  26891=>"111111111",
  26892=>"000000000",
  26893=>"110111111",
  26894=>"000000000",
  26895=>"001111110",
  26896=>"111111110",
  26897=>"101101101",
  26898=>"001000000",
  26899=>"000110111",
  26900=>"111111110",
  26901=>"100000111",
  26902=>"110010111",
  26903=>"111111001",
  26904=>"011001001",
  26905=>"110110110",
  26906=>"100000000",
  26907=>"111110111",
  26908=>"100110111",
  26909=>"101111111",
  26910=>"111101001",
  26911=>"111111111",
  26912=>"000000000",
  26913=>"111111111",
  26914=>"000000000",
  26915=>"000001111",
  26916=>"111111111",
  26917=>"111101101",
  26918=>"001001001",
  26919=>"111001001",
  26920=>"111000111",
  26921=>"111111111",
  26922=>"110111111",
  26923=>"111111111",
  26924=>"000000000",
  26925=>"110111001",
  26926=>"111000111",
  26927=>"011011011",
  26928=>"111111111",
  26929=>"010000000",
  26930=>"110110000",
  26931=>"111110111",
  26932=>"000000100",
  26933=>"001000100",
  26934=>"111111111",
  26935=>"100000000",
  26936=>"000000000",
  26937=>"000000100",
  26938=>"001000111",
  26939=>"000001001",
  26940=>"111111111",
  26941=>"000111111",
  26942=>"011000011",
  26943=>"111101111",
  26944=>"100000000",
  26945=>"000000000",
  26946=>"000000000",
  26947=>"111011000",
  26948=>"001000111",
  26949=>"111111111",
  26950=>"111111001",
  26951=>"111111111",
  26952=>"010000000",
  26953=>"000000000",
  26954=>"101000001",
  26955=>"111111010",
  26956=>"111111100",
  26957=>"000000011",
  26958=>"110111111",
  26959=>"011011111",
  26960=>"111111111",
  26961=>"000001111",
  26962=>"111001111",
  26963=>"001000000",
  26964=>"111111001",
  26965=>"011011011",
  26966=>"001101111",
  26967=>"111111111",
  26968=>"111111000",
  26969=>"111111111",
  26970=>"111110000",
  26971=>"000000000",
  26972=>"100111011",
  26973=>"111100000",
  26974=>"111100000",
  26975=>"111111111",
  26976=>"000000000",
  26977=>"000000001",
  26978=>"100101100",
  26979=>"100000100",
  26980=>"111111111",
  26981=>"000000000",
  26982=>"111111111",
  26983=>"000000000",
  26984=>"110001000",
  26985=>"000000000",
  26986=>"000000000",
  26987=>"111010000",
  26988=>"010011011",
  26989=>"000111111",
  26990=>"001000000",
  26991=>"000100110",
  26992=>"111011111",
  26993=>"011011111",
  26994=>"000001000",
  26995=>"111101000",
  26996=>"111111111",
  26997=>"111011011",
  26998=>"000111110",
  26999=>"000000000",
  27000=>"101101000",
  27001=>"100111000",
  27002=>"000000000",
  27003=>"010000100",
  27004=>"001111000",
  27005=>"111001000",
  27006=>"010111111",
  27007=>"100101111",
  27008=>"001000000",
  27009=>"000100000",
  27010=>"111111111",
  27011=>"111111111",
  27012=>"111111010",
  27013=>"011011111",
  27014=>"000100110",
  27015=>"111111111",
  27016=>"101001111",
  27017=>"000110111",
  27018=>"111111101",
  27019=>"000000000",
  27020=>"111111111",
  27021=>"010011011",
  27022=>"001111111",
  27023=>"000000000",
  27024=>"000111110",
  27025=>"000000000",
  27026=>"000000000",
  27027=>"111111111",
  27028=>"001000000",
  27029=>"011000000",
  27030=>"000000000",
  27031=>"000000010",
  27032=>"000000000",
  27033=>"000000000",
  27034=>"111111111",
  27035=>"001011011",
  27036=>"000001111",
  27037=>"111010000",
  27038=>"000000110",
  27039=>"000000000",
  27040=>"000000000",
  27041=>"101101101",
  27042=>"000000001",
  27043=>"000010111",
  27044=>"000111111",
  27045=>"011111111",
  27046=>"111101111",
  27047=>"000000000",
  27048=>"110010000",
  27049=>"000000000",
  27050=>"000000000",
  27051=>"111110000",
  27052=>"111000000",
  27053=>"000000100",
  27054=>"000000000",
  27055=>"000000000",
  27056=>"111111100",
  27057=>"111111111",
  27058=>"000000000",
  27059=>"000111111",
  27060=>"111100101",
  27061=>"000000000",
  27062=>"100111111",
  27063=>"011110010",
  27064=>"000000000",
  27065=>"111111111",
  27066=>"111100000",
  27067=>"000000000",
  27068=>"011011000",
  27069=>"001001000",
  27070=>"000000111",
  27071=>"111111111",
  27072=>"000010000",
  27073=>"100000000",
  27074=>"000000000",
  27075=>"011111111",
  27076=>"000110000",
  27077=>"000111110",
  27078=>"000000001",
  27079=>"000000001",
  27080=>"000000000",
  27081=>"000001111",
  27082=>"000001111",
  27083=>"100000001",
  27084=>"000000000",
  27085=>"000000000",
  27086=>"000000000",
  27087=>"000010000",
  27088=>"000000100",
  27089=>"111111111",
  27090=>"111110111",
  27091=>"110100111",
  27092=>"000100000",
  27093=>"000000000",
  27094=>"111011000",
  27095=>"111011001",
  27096=>"001011111",
  27097=>"010110101",
  27098=>"111110111",
  27099=>"011111000",
  27100=>"000000100",
  27101=>"110101101",
  27102=>"111001111",
  27103=>"000000000",
  27104=>"010011111",
  27105=>"000000000",
  27106=>"000000000",
  27107=>"111101000",
  27108=>"000010010",
  27109=>"111100001",
  27110=>"000111111",
  27111=>"000000101",
  27112=>"110101111",
  27113=>"111011001",
  27114=>"101000110",
  27115=>"111111111",
  27116=>"100000000",
  27117=>"000001000",
  27118=>"111111111",
  27119=>"111000000",
  27120=>"111111111",
  27121=>"111111111",
  27122=>"111111111",
  27123=>"100000000",
  27124=>"000000000",
  27125=>"111110000",
  27126=>"111111111",
  27127=>"000000110",
  27128=>"101000001",
  27129=>"010111001",
  27130=>"111111011",
  27131=>"000110111",
  27132=>"000000000",
  27133=>"000000000",
  27134=>"110110100",
  27135=>"111100000",
  27136=>"100000000",
  27137=>"000000000",
  27138=>"111111111",
  27139=>"111111111",
  27140=>"111111111",
  27141=>"101000000",
  27142=>"000000000",
  27143=>"111001101",
  27144=>"111111111",
  27145=>"111111111",
  27146=>"111111111",
  27147=>"111001101",
  27148=>"000000100",
  27149=>"000000000",
  27150=>"111111001",
  27151=>"000000000",
  27152=>"000000000",
  27153=>"000000000",
  27154=>"111111111",
  27155=>"001001111",
  27156=>"000110111",
  27157=>"110111111",
  27158=>"111111111",
  27159=>"100111111",
  27160=>"000001001",
  27161=>"111011001",
  27162=>"111111000",
  27163=>"000000000",
  27164=>"001001111",
  27165=>"000000000",
  27166=>"111001001",
  27167=>"111111111",
  27168=>"111111111",
  27169=>"000000000",
  27170=>"100100100",
  27171=>"100000000",
  27172=>"001000000",
  27173=>"000101011",
  27174=>"001000000",
  27175=>"000000000",
  27176=>"101001001",
  27177=>"000000000",
  27178=>"111001001",
  27179=>"110111111",
  27180=>"001001000",
  27181=>"000111001",
  27182=>"110011001",
  27183=>"111111111",
  27184=>"000000000",
  27185=>"000000000",
  27186=>"110111011",
  27187=>"111111111",
  27188=>"100001101",
  27189=>"100000001",
  27190=>"000001100",
  27191=>"000000000",
  27192=>"010000001",
  27193=>"000000011",
  27194=>"000000000",
  27195=>"000011111",
  27196=>"000000111",
  27197=>"000000111",
  27198=>"111101101",
  27199=>"000000000",
  27200=>"001111111",
  27201=>"000000000",
  27202=>"000111111",
  27203=>"000000000",
  27204=>"000000000",
  27205=>"011011111",
  27206=>"111111000",
  27207=>"001000000",
  27208=>"000011011",
  27209=>"111111111",
  27210=>"110110110",
  27211=>"101101111",
  27212=>"111111111",
  27213=>"111101100",
  27214=>"011001000",
  27215=>"000001101",
  27216=>"000101111",
  27217=>"111011011",
  27218=>"010110110",
  27219=>"111111110",
  27220=>"000111101",
  27221=>"000000000",
  27222=>"000000000",
  27223=>"111111111",
  27224=>"111111111",
  27225=>"101000000",
  27226=>"111111111",
  27227=>"000000100",
  27228=>"110110000",
  27229=>"111111111",
  27230=>"001000000",
  27231=>"011001001",
  27232=>"111111111",
  27233=>"001000000",
  27234=>"111111111",
  27235=>"000000000",
  27236=>"111111111",
  27237=>"000000000",
  27238=>"000001111",
  27239=>"000000000",
  27240=>"011010000",
  27241=>"000000000",
  27242=>"111011010",
  27243=>"011111111",
  27244=>"111111111",
  27245=>"101000000",
  27246=>"000000000",
  27247=>"111111110",
  27248=>"000000000",
  27249=>"111001111",
  27250=>"010010000",
  27251=>"111111111",
  27252=>"000000000",
  27253=>"100110111",
  27254=>"000011111",
  27255=>"000000111",
  27256=>"000000011",
  27257=>"111111000",
  27258=>"001000000",
  27259=>"111111111",
  27260=>"100000100",
  27261=>"111010000",
  27262=>"111111111",
  27263=>"000000000",
  27264=>"111010110",
  27265=>"001111111",
  27266=>"000000000",
  27267=>"000000000",
  27268=>"011011111",
  27269=>"001000000",
  27270=>"111110000",
  27271=>"111111000",
  27272=>"111111100",
  27273=>"000001000",
  27274=>"111000001",
  27275=>"111001001",
  27276=>"000000000",
  27277=>"000000000",
  27278=>"111111111",
  27279=>"100110111",
  27280=>"111111111",
  27281=>"110111110",
  27282=>"110000000",
  27283=>"111111111",
  27284=>"111111001",
  27285=>"111111001",
  27286=>"000000000",
  27287=>"000000000",
  27288=>"111111110",
  27289=>"111111111",
  27290=>"000110111",
  27291=>"000000000",
  27292=>"111110110",
  27293=>"110010000",
  27294=>"111111111",
  27295=>"000000000",
  27296=>"000100000",
  27297=>"111111111",
  27298=>"111111111",
  27299=>"000000000",
  27300=>"000000000",
  27301=>"111000000",
  27302=>"111111101",
  27303=>"001100100",
  27304=>"000011000",
  27305=>"000000000",
  27306=>"000000000",
  27307=>"010111011",
  27308=>"111111111",
  27309=>"000000000",
  27310=>"111111111",
  27311=>"000010000",
  27312=>"000010011",
  27313=>"100111110",
  27314=>"010111010",
  27315=>"111100100",
  27316=>"111111111",
  27317=>"111000000",
  27318=>"111011001",
  27319=>"000000000",
  27320=>"111111111",
  27321=>"111111111",
  27322=>"001001111",
  27323=>"000101111",
  27324=>"111111111",
  27325=>"101111110",
  27326=>"111111111",
  27327=>"100000101",
  27328=>"000000000",
  27329=>"111111111",
  27330=>"110100100",
  27331=>"000010000",
  27332=>"111111111",
  27333=>"000000000",
  27334=>"001010000",
  27335=>"101001000",
  27336=>"111111111",
  27337=>"000100111",
  27338=>"100100101",
  27339=>"111111111",
  27340=>"000000101",
  27341=>"000000111",
  27342=>"000000101",
  27343=>"100100111",
  27344=>"000000000",
  27345=>"000000000",
  27346=>"111000000",
  27347=>"000000000",
  27348=>"001000001",
  27349=>"000000000",
  27350=>"000000111",
  27351=>"111000111",
  27352=>"100111111",
  27353=>"000000101",
  27354=>"000000000",
  27355=>"111111010",
  27356=>"111111111",
  27357=>"111111100",
  27358=>"000000000",
  27359=>"111000100",
  27360=>"011110000",
  27361=>"000011111",
  27362=>"011011000",
  27363=>"000000000",
  27364=>"000001000",
  27365=>"000000000",
  27366=>"111111111",
  27367=>"111111011",
  27368=>"000000111",
  27369=>"000000000",
  27370=>"001001001",
  27371=>"000000000",
  27372=>"111111110",
  27373=>"000000000",
  27374=>"000000000",
  27375=>"110111111",
  27376=>"011111111",
  27377=>"000000000",
  27378=>"111101110",
  27379=>"100101111",
  27380=>"011000000",
  27381=>"001001000",
  27382=>"111111000",
  27383=>"111111010",
  27384=>"111111111",
  27385=>"000000111",
  27386=>"000100111",
  27387=>"001111111",
  27388=>"111011001",
  27389=>"000000000",
  27390=>"000011000",
  27391=>"111111111",
  27392=>"000000000",
  27393=>"111001111",
  27394=>"011000000",
  27395=>"111100111",
  27396=>"111111111",
  27397=>"110001011",
  27398=>"000000001",
  27399=>"000011010",
  27400=>"111111111",
  27401=>"111111111",
  27402=>"111111111",
  27403=>"111111111",
  27404=>"000000001",
  27405=>"111111111",
  27406=>"010000000",
  27407=>"000000000",
  27408=>"000000000",
  27409=>"000100111",
  27410=>"111111111",
  27411=>"111111111",
  27412=>"010000000",
  27413=>"011000000",
  27414=>"111111101",
  27415=>"000000000",
  27416=>"000000000",
  27417=>"111111011",
  27418=>"111011111",
  27419=>"010000000",
  27420=>"110111110",
  27421=>"000000000",
  27422=>"000000000",
  27423=>"111111000",
  27424=>"100100001",
  27425=>"111111101",
  27426=>"000000000",
  27427=>"000000000",
  27428=>"111011111",
  27429=>"000000000",
  27430=>"011000011",
  27431=>"000011110",
  27432=>"000000000",
  27433=>"001000000",
  27434=>"111000000",
  27435=>"111111000",
  27436=>"000000000",
  27437=>"010110110",
  27438=>"000000000",
  27439=>"000000000",
  27440=>"001111111",
  27441=>"000000000",
  27442=>"111111111",
  27443=>"000010000",
  27444=>"000000000",
  27445=>"111111111",
  27446=>"111111111",
  27447=>"000000000",
  27448=>"111111111",
  27449=>"111000000",
  27450=>"101101111",
  27451=>"000010010",
  27452=>"100110110",
  27453=>"111111111",
  27454=>"000001001",
  27455=>"110111011",
  27456=>"100111001",
  27457=>"111111111",
  27458=>"100000100",
  27459=>"000111111",
  27460=>"100000000",
  27461=>"000001000",
  27462=>"000000100",
  27463=>"111101111",
  27464=>"111111111",
  27465=>"001000000",
  27466=>"111111111",
  27467=>"110010001",
  27468=>"000000000",
  27469=>"000000000",
  27470=>"011111111",
  27471=>"100000000",
  27472=>"001011011",
  27473=>"000000011",
  27474=>"000000011",
  27475=>"111111011",
  27476=>"111111111",
  27477=>"011011001",
  27478=>"011000000",
  27479=>"111111111",
  27480=>"000000000",
  27481=>"100100111",
  27482=>"000000000",
  27483=>"111111111",
  27484=>"000000000",
  27485=>"100000110",
  27486=>"100000000",
  27487=>"000000000",
  27488=>"111111011",
  27489=>"111111001",
  27490=>"110110000",
  27491=>"000000001",
  27492=>"000000010",
  27493=>"000000000",
  27494=>"001111000",
  27495=>"000101111",
  27496=>"001001011",
  27497=>"000000000",
  27498=>"000000100",
  27499=>"111111111",
  27500=>"000000000",
  27501=>"110111111",
  27502=>"111000000",
  27503=>"111111111",
  27504=>"111010000",
  27505=>"111000000",
  27506=>"000000000",
  27507=>"001000000",
  27508=>"100000010",
  27509=>"000000000",
  27510=>"000000000",
  27511=>"000000100",
  27512=>"000000000",
  27513=>"000000011",
  27514=>"101000000",
  27515=>"000000100",
  27516=>"000000000",
  27517=>"001000111",
  27518=>"000000100",
  27519=>"111000000",
  27520=>"100000000",
  27521=>"001000000",
  27522=>"000100100",
  27523=>"000000110",
  27524=>"000000000",
  27525=>"111111111",
  27526=>"000001000",
  27527=>"111111100",
  27528=>"111001011",
  27529=>"000000111",
  27530=>"111111111",
  27531=>"000000111",
  27532=>"101101111",
  27533=>"011111111",
  27534=>"000000000",
  27535=>"110111111",
  27536=>"000000000",
  27537=>"111000000",
  27538=>"000100100",
  27539=>"001001001",
  27540=>"000000000",
  27541=>"000010010",
  27542=>"100000000",
  27543=>"111111011",
  27544=>"111111011",
  27545=>"000000111",
  27546=>"111111111",
  27547=>"111111111",
  27548=>"000000000",
  27549=>"111111111",
  27550=>"000000011",
  27551=>"000000000",
  27552=>"111111111",
  27553=>"001001000",
  27554=>"111111111",
  27555=>"111111111",
  27556=>"111111111",
  27557=>"000000010",
  27558=>"100101111",
  27559=>"000000000",
  27560=>"000000000",
  27561=>"001000111",
  27562=>"111111111",
  27563=>"000000001",
  27564=>"000000000",
  27565=>"000100010",
  27566=>"000110111",
  27567=>"000000101",
  27568=>"110110111",
  27569=>"011111111",
  27570=>"000000000",
  27571=>"111111000",
  27572=>"100000000",
  27573=>"000000110",
  27574=>"111101111",
  27575=>"000000001",
  27576=>"100000110",
  27577=>"001011111",
  27578=>"111111111",
  27579=>"111111111",
  27580=>"000000001",
  27581=>"000000000",
  27582=>"110110000",
  27583=>"000000011",
  27584=>"111111111",
  27585=>"000000000",
  27586=>"011011111",
  27587=>"000000000",
  27588=>"111110110",
  27589=>"000100100",
  27590=>"011000000",
  27591=>"010000000",
  27592=>"000000100",
  27593=>"000000000",
  27594=>"000000000",
  27595=>"000111101",
  27596=>"111001000",
  27597=>"000000000",
  27598=>"111101111",
  27599=>"000111111",
  27600=>"000000000",
  27601=>"111100111",
  27602=>"000000000",
  27603=>"000000000",
  27604=>"000000000",
  27605=>"101000000",
  27606=>"111101111",
  27607=>"001011011",
  27608=>"011001111",
  27609=>"111111111",
  27610=>"001000000",
  27611=>"000000001",
  27612=>"111111111",
  27613=>"100100100",
  27614=>"000000000",
  27615=>"000000000",
  27616=>"011111111",
  27617=>"000001111",
  27618=>"111111111",
  27619=>"011001111",
  27620=>"111111111",
  27621=>"110111010",
  27622=>"111111000",
  27623=>"111111111",
  27624=>"001101111",
  27625=>"111111111",
  27626=>"000111111",
  27627=>"111111111",
  27628=>"111111111",
  27629=>"000100100",
  27630=>"000000000",
  27631=>"110111111",
  27632=>"111111111",
  27633=>"000001001",
  27634=>"000000000",
  27635=>"111111111",
  27636=>"000000000",
  27637=>"000000000",
  27638=>"000001001",
  27639=>"000000000",
  27640=>"111111100",
  27641=>"101111111",
  27642=>"000111111",
  27643=>"111111010",
  27644=>"111111011",
  27645=>"010000000",
  27646=>"000111000",
  27647=>"100100100",
  27648=>"011011011",
  27649=>"000100110",
  27650=>"111101101",
  27651=>"000000100",
  27652=>"001101000",
  27653=>"000000000",
  27654=>"111111111",
  27655=>"111111111",
  27656=>"111111000",
  27657=>"000110110",
  27658=>"010010000",
  27659=>"010010000",
  27660=>"110111000",
  27661=>"000000110",
  27662=>"111111000",
  27663=>"000000111",
  27664=>"001001011",
  27665=>"111111111",
  27666=>"000000000",
  27667=>"000000000",
  27668=>"110011000",
  27669=>"000000000",
  27670=>"110111000",
  27671=>"000000010",
  27672=>"000000000",
  27673=>"011011111",
  27674=>"000000010",
  27675=>"001000000",
  27676=>"001000000",
  27677=>"111111011",
  27678=>"100100100",
  27679=>"000000111",
  27680=>"000000000",
  27681=>"011001001",
  27682=>"110110000",
  27683=>"000000000",
  27684=>"111111111",
  27685=>"000000000",
  27686=>"111110111",
  27687=>"111111000",
  27688=>"000000001",
  27689=>"000000000",
  27690=>"001001000",
  27691=>"000000000",
  27692=>"111111111",
  27693=>"000111111",
  27694=>"000111111",
  27695=>"111110111",
  27696=>"111111111",
  27697=>"000000001",
  27698=>"111111110",
  27699=>"111111111",
  27700=>"000001101",
  27701=>"110010111",
  27702=>"111110000",
  27703=>"100000000",
  27704=>"111111111",
  27705=>"001001111",
  27706=>"000010111",
  27707=>"101001000",
  27708=>"100111110",
  27709=>"111111100",
  27710=>"001001001",
  27711=>"000000000",
  27712=>"110100111",
  27713=>"000101111",
  27714=>"110110111",
  27715=>"111000000",
  27716=>"000000001",
  27717=>"001011011",
  27718=>"111111000",
  27719=>"000000000",
  27720=>"011111000",
  27721=>"001000000",
  27722=>"000000110",
  27723=>"001001110",
  27724=>"000000001",
  27725=>"110000000",
  27726=>"001111000",
  27727=>"010010010",
  27728=>"000100000",
  27729=>"111111110",
  27730=>"000000001",
  27731=>"010000001",
  27732=>"101101111",
  27733=>"001000000",
  27734=>"000000000",
  27735=>"000000001",
  27736=>"001001111",
  27737=>"001000000",
  27738=>"111110000",
  27739=>"000001001",
  27740=>"000000000",
  27741=>"111011000",
  27742=>"000000000",
  27743=>"110000000",
  27744=>"111011001",
  27745=>"011111110",
  27746=>"000000000",
  27747=>"000000010",
  27748=>"110000000",
  27749=>"000011000",
  27750=>"111111000",
  27751=>"000110110",
  27752=>"100001111",
  27753=>"000000000",
  27754=>"111111110",
  27755=>"000000000",
  27756=>"010010010",
  27757=>"000000111",
  27758=>"000000000",
  27759=>"110110100",
  27760=>"011011111",
  27761=>"011001011",
  27762=>"001001001",
  27763=>"111111111",
  27764=>"000001011",
  27765=>"000000000",
  27766=>"111111000",
  27767=>"111111110",
  27768=>"000100111",
  27769=>"011111111",
  27770=>"000000000",
  27771=>"111111011",
  27772=>"000000010",
  27773=>"000000001",
  27774=>"000001000",
  27775=>"000110111",
  27776=>"001111001",
  27777=>"101100111",
  27778=>"000100111",
  27779=>"001000111",
  27780=>"001000110",
  27781=>"001111111",
  27782=>"101011110",
  27783=>"000100000",
  27784=>"111000000",
  27785=>"000000110",
  27786=>"010001000",
  27787=>"111111000",
  27788=>"000011011",
  27789=>"111111111",
  27790=>"000000000",
  27791=>"111111110",
  27792=>"000000000",
  27793=>"000111101",
  27794=>"001001001",
  27795=>"111110010",
  27796=>"111111100",
  27797=>"000010000",
  27798=>"000110110",
  27799=>"111000000",
  27800=>"111011011",
  27801=>"001000010",
  27802=>"110000001",
  27803=>"100000000",
  27804=>"100110110",
  27805=>"000110111",
  27806=>"111000000",
  27807=>"011000100",
  27808=>"000000000",
  27809=>"100111000",
  27810=>"000000000",
  27811=>"000110111",
  27812=>"111110010",
  27813=>"111000110",
  27814=>"100000000",
  27815=>"000000001",
  27816=>"000000000",
  27817=>"111111110",
  27818=>"000000000",
  27819=>"111000000",
  27820=>"111011111",
  27821=>"110100000",
  27822=>"111111111",
  27823=>"111111000",
  27824=>"111111111",
  27825=>"110111101",
  27826=>"111111010",
  27827=>"111011000",
  27828=>"000111001",
  27829=>"100000111",
  27830=>"000000010",
  27831=>"111111111",
  27832=>"010000000",
  27833=>"000110110",
  27834=>"110100000",
  27835=>"111111000",
  27836=>"011111111",
  27837=>"111111000",
  27838=>"000000001",
  27839=>"000000111",
  27840=>"000000000",
  27841=>"111111111",
  27842=>"010000000",
  27843=>"000000000",
  27844=>"000001101",
  27845=>"111111100",
  27846=>"000000111",
  27847=>"111111000",
  27848=>"000111111",
  27849=>"011001101",
  27850=>"001100100",
  27851=>"000110111",
  27852=>"000000011",
  27853=>"000111111",
  27854=>"110000110",
  27855=>"000000000",
  27856=>"111110110",
  27857=>"000110000",
  27858=>"110100100",
  27859=>"111111010",
  27860=>"111111111",
  27861=>"100000110",
  27862=>"000000000",
  27863=>"000010010",
  27864=>"000110000",
  27865=>"111111110",
  27866=>"111111110",
  27867=>"001000100",
  27868=>"011111011",
  27869=>"111001000",
  27870=>"111000000",
  27871=>"001101101",
  27872=>"001000000",
  27873=>"111111000",
  27874=>"111111000",
  27875=>"111111111",
  27876=>"111111100",
  27877=>"111010010",
  27878=>"000000111",
  27879=>"000000100",
  27880=>"001101111",
  27881=>"000010000",
  27882=>"001000111",
  27883=>"111110100",
  27884=>"111111101",
  27885=>"000000000",
  27886=>"110000000",
  27887=>"100100000",
  27888=>"000000010",
  27889=>"111111111",
  27890=>"000000110",
  27891=>"111010000",
  27892=>"111111101",
  27893=>"011000000",
  27894=>"110110111",
  27895=>"000000000",
  27896=>"011111111",
  27897=>"000000010",
  27898=>"000000000",
  27899=>"111111100",
  27900=>"110111111",
  27901=>"011011000",
  27902=>"111100000",
  27903=>"111111111",
  27904=>"111111001",
  27905=>"010110110",
  27906=>"111111011",
  27907=>"111111111",
  27908=>"000000000",
  27909=>"001000100",
  27910=>"111110110",
  27911=>"000000111",
  27912=>"110000000",
  27913=>"000000010",
  27914=>"000000001",
  27915=>"111111000",
  27916=>"000000111",
  27917=>"111110010",
  27918=>"111111111",
  27919=>"000000000",
  27920=>"001001000",
  27921=>"100000000",
  27922=>"011001001",
  27923=>"000000000",
  27924=>"000000000",
  27925=>"000000000",
  27926=>"011011000",
  27927=>"000000001",
  27928=>"011011111",
  27929=>"100000001",
  27930=>"001000000",
  27931=>"000100110",
  27932=>"000001011",
  27933=>"110100000",
  27934=>"000000000",
  27935=>"111000000",
  27936=>"000110000",
  27937=>"100000100",
  27938=>"111111111",
  27939=>"000000111",
  27940=>"111000000",
  27941=>"000000000",
  27942=>"111111011",
  27943=>"010000000",
  27944=>"111110111",
  27945=>"000001011",
  27946=>"000000000",
  27947=>"000001101",
  27948=>"000000000",
  27949=>"110110000",
  27950=>"000000000",
  27951=>"000000000",
  27952=>"000000111",
  27953=>"111000000",
  27954=>"000110110",
  27955=>"111111110",
  27956=>"000000000",
  27957=>"010000000",
  27958=>"000000000",
  27959=>"000000000",
  27960=>"000000000",
  27961=>"001000000",
  27962=>"101101111",
  27963=>"000000100",
  27964=>"000000000",
  27965=>"001000110",
  27966=>"000101101",
  27967=>"011000000",
  27968=>"000000000",
  27969=>"111111111",
  27970=>"111111111",
  27971=>"000010000",
  27972=>"001000000",
  27973=>"111111111",
  27974=>"110111111",
  27975=>"110110000",
  27976=>"000000000",
  27977=>"100000000",
  27978=>"000000000",
  27979=>"101001000",
  27980=>"000100111",
  27981=>"000111111",
  27982=>"110010111",
  27983=>"000011111",
  27984=>"000000000",
  27985=>"000000111",
  27986=>"111111110",
  27987=>"000000100",
  27988=>"000000000",
  27989=>"001011011",
  27990=>"111110110",
  27991=>"000000100",
  27992=>"001111111",
  27993=>"000000000",
  27994=>"111111000",
  27995=>"000000110",
  27996=>"101001001",
  27997=>"000110111",
  27998=>"111110100",
  27999=>"011111111",
  28000=>"001100111",
  28001=>"111011000",
  28002=>"100100000",
  28003=>"011111111",
  28004=>"000001001",
  28005=>"000000000",
  28006=>"000000000",
  28007=>"111111111",
  28008=>"000000000",
  28009=>"110110000",
  28010=>"111011001",
  28011=>"101111111",
  28012=>"111111000",
  28013=>"111111111",
  28014=>"000000000",
  28015=>"000001111",
  28016=>"110110000",
  28017=>"100000100",
  28018=>"111111111",
  28019=>"011001000",
  28020=>"100000101",
  28021=>"000101001",
  28022=>"000000000",
  28023=>"111000000",
  28024=>"111111011",
  28025=>"000000000",
  28026=>"001000000",
  28027=>"000000000",
  28028=>"110111000",
  28029=>"001010000",
  28030=>"111110010",
  28031=>"000000000",
  28032=>"001011111",
  28033=>"111111110",
  28034=>"111110110",
  28035=>"111111101",
  28036=>"011001000",
  28037=>"011000000",
  28038=>"000100100",
  28039=>"000110100",
  28040=>"111000000",
  28041=>"111111000",
  28042=>"000000000",
  28043=>"000000111",
  28044=>"000000000",
  28045=>"000100111",
  28046=>"111111001",
  28047=>"001001000",
  28048=>"000000110",
  28049=>"111111110",
  28050=>"000000111",
  28051=>"111111111",
  28052=>"100100110",
  28053=>"010111111",
  28054=>"111111111",
  28055=>"110100000",
  28056=>"111111111",
  28057=>"011111111",
  28058=>"111111111",
  28059=>"001000000",
  28060=>"000111111",
  28061=>"011111010",
  28062=>"111111111",
  28063=>"111111000",
  28064=>"000100110",
  28065=>"011000000",
  28066=>"011001011",
  28067=>"100111000",
  28068=>"001001111",
  28069=>"001001000",
  28070=>"111000000",
  28071=>"001100000",
  28072=>"111111011",
  28073=>"111000000",
  28074=>"111011000",
  28075=>"101111101",
  28076=>"000000000",
  28077=>"000000111",
  28078=>"100000011",
  28079=>"001001000",
  28080=>"000000011",
  28081=>"111110100",
  28082=>"110000000",
  28083=>"001001101",
  28084=>"111001000",
  28085=>"111111000",
  28086=>"111111111",
  28087=>"111111111",
  28088=>"111110000",
  28089=>"111111111",
  28090=>"111111011",
  28091=>"111111111",
  28092=>"001001101",
  28093=>"001001000",
  28094=>"000000000",
  28095=>"000111100",
  28096=>"111101101",
  28097=>"001001101",
  28098=>"000000000",
  28099=>"000000000",
  28100=>"001000100",
  28101=>"011000100",
  28102=>"000000110",
  28103=>"001000111",
  28104=>"000000000",
  28105=>"111111111",
  28106=>"000000000",
  28107=>"000000001",
  28108=>"000000000",
  28109=>"011110111",
  28110=>"111111110",
  28111=>"000000000",
  28112=>"000000000",
  28113=>"000010000",
  28114=>"000100000",
  28115=>"000000110",
  28116=>"101111100",
  28117=>"000000000",
  28118=>"000000000",
  28119=>"011011000",
  28120=>"000001001",
  28121=>"000000010",
  28122=>"000010000",
  28123=>"111111000",
  28124=>"000111100",
  28125=>"111111000",
  28126=>"000000000",
  28127=>"000111110",
  28128=>"001111100",
  28129=>"111011010",
  28130=>"000000000",
  28131=>"011000000",
  28132=>"111111111",
  28133=>"000101111",
  28134=>"001000100",
  28135=>"100100000",
  28136=>"111000000",
  28137=>"000000000",
  28138=>"110000100",
  28139=>"001000000",
  28140=>"000000000",
  28141=>"011010000",
  28142=>"000000100",
  28143=>"111111110",
  28144=>"000011001",
  28145=>"111111111",
  28146=>"001101110",
  28147=>"000000111",
  28148=>"000000000",
  28149=>"000110110",
  28150=>"000000000",
  28151=>"110000000",
  28152=>"000000000",
  28153=>"010110010",
  28154=>"110110110",
  28155=>"000000001",
  28156=>"111101000",
  28157=>"110111111",
  28158=>"000000100",
  28159=>"000000000",
  28160=>"101101000",
  28161=>"100000000",
  28162=>"110110111",
  28163=>"111111000",
  28164=>"001010000",
  28165=>"101001001",
  28166=>"000111111",
  28167=>"100110110",
  28168=>"111111011",
  28169=>"011000011",
  28170=>"011011000",
  28171=>"111111001",
  28172=>"000110110",
  28173=>"100100111",
  28174=>"111101111",
  28175=>"000000000",
  28176=>"110111111",
  28177=>"100001000",
  28178=>"001001011",
  28179=>"110110110",
  28180=>"000000111",
  28181=>"100000000",
  28182=>"000000000",
  28183=>"111111111",
  28184=>"100111000",
  28185=>"001100110",
  28186=>"111110111",
  28187=>"011001001",
  28188=>"000000000",
  28189=>"111000000",
  28190=>"101101100",
  28191=>"111111000",
  28192=>"111111001",
  28193=>"000000000",
  28194=>"000000000",
  28195=>"111111111",
  28196=>"000000000",
  28197=>"000110111",
  28198=>"111000000",
  28199=>"000100110",
  28200=>"001001001",
  28201=>"000000000",
  28202=>"001000000",
  28203=>"000001000",
  28204=>"111111111",
  28205=>"111111111",
  28206=>"000000000",
  28207=>"100000010",
  28208=>"110000000",
  28209=>"000000000",
  28210=>"011000000",
  28211=>"001001011",
  28212=>"001101111",
  28213=>"000100000",
  28214=>"111101111",
  28215=>"000011011",
  28216=>"111111110",
  28217=>"000000111",
  28218=>"000000000",
  28219=>"111110111",
  28220=>"011111111",
  28221=>"001001001",
  28222=>"000000000",
  28223=>"000000111",
  28224=>"101000000",
  28225=>"000000000",
  28226=>"101111111",
  28227=>"100111000",
  28228=>"111111111",
  28229=>"111111110",
  28230=>"100100000",
  28231=>"111111000",
  28232=>"110101110",
  28233=>"000011111",
  28234=>"101111000",
  28235=>"111011000",
  28236=>"111111000",
  28237=>"001011000",
  28238=>"111101001",
  28239=>"000000000",
  28240=>"000000000",
  28241=>"111001111",
  28242=>"100000000",
  28243=>"000000010",
  28244=>"000000000",
  28245=>"100000000",
  28246=>"111111011",
  28247=>"111111111",
  28248=>"111111111",
  28249=>"000000100",
  28250=>"111010000",
  28251=>"111111111",
  28252=>"000000001",
  28253=>"111111111",
  28254=>"101100100",
  28255=>"011111111",
  28256=>"000000000",
  28257=>"111111111",
  28258=>"000111111",
  28259=>"000000000",
  28260=>"111111100",
  28261=>"000000000",
  28262=>"001001011",
  28263=>"000000000",
  28264=>"000100000",
  28265=>"110111111",
  28266=>"000100100",
  28267=>"111001000",
  28268=>"100000100",
  28269=>"000000000",
  28270=>"000010001",
  28271=>"000000111",
  28272=>"110110000",
  28273=>"000000000",
  28274=>"111101111",
  28275=>"011011011",
  28276=>"000000001",
  28277=>"000000000",
  28278=>"111111111",
  28279=>"111111000",
  28280=>"111111011",
  28281=>"100100111",
  28282=>"000000000",
  28283=>"000000000",
  28284=>"100111100",
  28285=>"100110111",
  28286=>"011001000",
  28287=>"000111111",
  28288=>"000000011",
  28289=>"111001111",
  28290=>"110000000",
  28291=>"000000000",
  28292=>"100000000",
  28293=>"000000100",
  28294=>"000000000",
  28295=>"111111111",
  28296=>"111111011",
  28297=>"111100000",
  28298=>"000000000",
  28299=>"111111111",
  28300=>"000111111",
  28301=>"111111010",
  28302=>"000000101",
  28303=>"001000000",
  28304=>"100100100",
  28305=>"101000000",
  28306=>"111111101",
  28307=>"100100000",
  28308=>"110111111",
  28309=>"101000111",
  28310=>"011111111",
  28311=>"110111111",
  28312=>"001001001",
  28313=>"000000111",
  28314=>"111111111",
  28315=>"000111000",
  28316=>"000100111",
  28317=>"000000000",
  28318=>"111111111",
  28319=>"000000010",
  28320=>"000000100",
  28321=>"100000000",
  28322=>"000000000",
  28323=>"001000000",
  28324=>"000001001",
  28325=>"000000000",
  28326=>"111111111",
  28327=>"110111010",
  28328=>"100001111",
  28329=>"000000111",
  28330=>"000000110",
  28331=>"111111111",
  28332=>"001000000",
  28333=>"111111110",
  28334=>"111011001",
  28335=>"111111111",
  28336=>"000000000",
  28337=>"011011001",
  28338=>"110110110",
  28339=>"011001000",
  28340=>"111111111",
  28341=>"000000000",
  28342=>"000101100",
  28343=>"000000001",
  28344=>"000000000",
  28345=>"000000000",
  28346=>"000111001",
  28347=>"000001001",
  28348=>"111111111",
  28349=>"000000000",
  28350=>"111110110",
  28351=>"000000000",
  28352=>"100101011",
  28353=>"000001011",
  28354=>"111111111",
  28355=>"111111111",
  28356=>"000000111",
  28357=>"000000110",
  28358=>"000000000",
  28359=>"111000110",
  28360=>"111111111",
  28361=>"000000000",
  28362=>"000001001",
  28363=>"111011011",
  28364=>"111111011",
  28365=>"000110000",
  28366=>"000000001",
  28367=>"000000000",
  28368=>"100000000",
  28369=>"000000001",
  28370=>"111111111",
  28371=>"000000111",
  28372=>"101111011",
  28373=>"101111111",
  28374=>"111111111",
  28375=>"111111111",
  28376=>"101111111",
  28377=>"111111111",
  28378=>"000000000",
  28379=>"111111010",
  28380=>"101101101",
  28381=>"111100110",
  28382=>"000001111",
  28383=>"111111111",
  28384=>"111111111",
  28385=>"000011011",
  28386=>"111111000",
  28387=>"111111011",
  28388=>"000000000",
  28389=>"001001011",
  28390=>"000000000",
  28391=>"111111111",
  28392=>"000000000",
  28393=>"111111111",
  28394=>"011111111",
  28395=>"000000001",
  28396=>"101111111",
  28397=>"111111111",
  28398=>"000110000",
  28399=>"111111111",
  28400=>"000100111",
  28401=>"010111001",
  28402=>"000000111",
  28403=>"101001111",
  28404=>"111111100",
  28405=>"111111111",
  28406=>"110110010",
  28407=>"111011000",
  28408=>"000000101",
  28409=>"100110000",
  28410=>"000000000",
  28411=>"000000000",
  28412=>"011111011",
  28413=>"000000011",
  28414=>"000000000",
  28415=>"011000000",
  28416=>"111111111",
  28417=>"011010000",
  28418=>"000000000",
  28419=>"111001000",
  28420=>"000000000",
  28421=>"000000110",
  28422=>"111111111",
  28423=>"101111011",
  28424=>"111001111",
  28425=>"000000000",
  28426=>"111111111",
  28427=>"001001000",
  28428=>"110100000",
  28429=>"000000000",
  28430=>"000111111",
  28431=>"101100111",
  28432=>"111110110",
  28433=>"000000111",
  28434=>"000000000",
  28435=>"110101000",
  28436=>"000111111",
  28437=>"011111000",
  28438=>"101101100",
  28439=>"111111111",
  28440=>"000100100",
  28441=>"000110111",
  28442=>"110000000",
  28443=>"111111111",
  28444=>"000000000",
  28445=>"111100000",
  28446=>"111111110",
  28447=>"111111111",
  28448=>"000000110",
  28449=>"110111011",
  28450=>"111111111",
  28451=>"111100100",
  28452=>"110000000",
  28453=>"000000011",
  28454=>"101100000",
  28455=>"000000100",
  28456=>"101110111",
  28457=>"000000001",
  28458=>"100000000",
  28459=>"000000100",
  28460=>"111111000",
  28461=>"111011000",
  28462=>"111111000",
  28463=>"000000000",
  28464=>"001101100",
  28465=>"000000101",
  28466=>"101000000",
  28467=>"000000000",
  28468=>"111000000",
  28469=>"111111111",
  28470=>"111000000",
  28471=>"000110111",
  28472=>"111111111",
  28473=>"000000000",
  28474=>"000000001",
  28475=>"100111111",
  28476=>"011000001",
  28477=>"100000110",
  28478=>"000000011",
  28479=>"111111111",
  28480=>"000000000",
  28481=>"000000000",
  28482=>"011001001",
  28483=>"100000000",
  28484=>"000001111",
  28485=>"111010000",
  28486=>"111101111",
  28487=>"001000000",
  28488=>"000000000",
  28489=>"000100011",
  28490=>"111001000",
  28491=>"000001011",
  28492=>"101001001",
  28493=>"111111110",
  28494=>"111100100",
  28495=>"010000000",
  28496=>"111111011",
  28497=>"000000000",
  28498=>"000000111",
  28499=>"001000000",
  28500=>"001000000",
  28501=>"011010011",
  28502=>"100100000",
  28503=>"000000111",
  28504=>"000000000",
  28505=>"000000000",
  28506=>"001010000",
  28507=>"000001011",
  28508=>"111010111",
  28509=>"000000011",
  28510=>"100100101",
  28511=>"000101101",
  28512=>"001000001",
  28513=>"111111111",
  28514=>"111111011",
  28515=>"111011000",
  28516=>"101111111",
  28517=>"000000000",
  28518=>"000001001",
  28519=>"000000000",
  28520=>"000000010",
  28521=>"000000011",
  28522=>"000000000",
  28523=>"000001000",
  28524=>"111111100",
  28525=>"110101001",
  28526=>"000000000",
  28527=>"000000011",
  28528=>"001000111",
  28529=>"111111111",
  28530=>"111111111",
  28531=>"011011001",
  28532=>"001000000",
  28533=>"111111000",
  28534=>"111111111",
  28535=>"111000000",
  28536=>"000000001",
  28537=>"111100100",
  28538=>"111111111",
  28539=>"000000111",
  28540=>"000000000",
  28541=>"101000000",
  28542=>"111101111",
  28543=>"111111111",
  28544=>"111111001",
  28545=>"000001111",
  28546=>"111111111",
  28547=>"000010010",
  28548=>"000000000",
  28549=>"110110110",
  28550=>"000001001",
  28551=>"101001001",
  28552=>"111111111",
  28553=>"011111011",
  28554=>"111111111",
  28555=>"111111111",
  28556=>"000000000",
  28557=>"000000000",
  28558=>"011000000",
  28559=>"010000000",
  28560=>"111111111",
  28561=>"111111111",
  28562=>"111000000",
  28563=>"000000000",
  28564=>"111111111",
  28565=>"001011000",
  28566=>"111111111",
  28567=>"100000100",
  28568=>"111111001",
  28569=>"111011001",
  28570=>"000000000",
  28571=>"100000100",
  28572=>"011111111",
  28573=>"000000000",
  28574=>"110111000",
  28575=>"000000000",
  28576=>"000000000",
  28577=>"110111111",
  28578=>"100000111",
  28579=>"011111110",
  28580=>"000000100",
  28581=>"111000000",
  28582=>"000000000",
  28583=>"111111011",
  28584=>"000000000",
  28585=>"001000000",
  28586=>"111111111",
  28587=>"101000000",
  28588=>"011000000",
  28589=>"111111000",
  28590=>"000000100",
  28591=>"010000001",
  28592=>"111111111",
  28593=>"111111010",
  28594=>"111111111",
  28595=>"111111111",
  28596=>"100110011",
  28597=>"000000000",
  28598=>"001111111",
  28599=>"000000000",
  28600=>"000000000",
  28601=>"000011111",
  28602=>"111011111",
  28603=>"100111001",
  28604=>"111111111",
  28605=>"111111001",
  28606=>"000000100",
  28607=>"000100111",
  28608=>"000001101",
  28609=>"110111111",
  28610=>"111111111",
  28611=>"000001001",
  28612=>"000000000",
  28613=>"000000000",
  28614=>"000000000",
  28615=>"000000000",
  28616=>"001001000",
  28617=>"000000110",
  28618=>"000000000",
  28619=>"000011101",
  28620=>"000001111",
  28621=>"110100000",
  28622=>"111111111",
  28623=>"000011011",
  28624=>"000000101",
  28625=>"110111001",
  28626=>"001001000",
  28627=>"010000111",
  28628=>"111111111",
  28629=>"100110111",
  28630=>"111111011",
  28631=>"000000000",
  28632=>"000110110",
  28633=>"000000000",
  28634=>"010011011",
  28635=>"000111111",
  28636=>"000001001",
  28637=>"001001000",
  28638=>"111111000",
  28639=>"000000000",
  28640=>"000100111",
  28641=>"001001001",
  28642=>"011110100",
  28643=>"101111011",
  28644=>"110000000",
  28645=>"011111111",
  28646=>"001000111",
  28647=>"011111111",
  28648=>"011001000",
  28649=>"111111111",
  28650=>"000110111",
  28651=>"100100100",
  28652=>"000101111",
  28653=>"111000001",
  28654=>"111111111",
  28655=>"100111111",
  28656=>"000000000",
  28657=>"000000111",
  28658=>"000000000",
  28659=>"100101111",
  28660=>"111011000",
  28661=>"001111111",
  28662=>"111111000",
  28663=>"111101000",
  28664=>"000111111",
  28665=>"100000001",
  28666=>"111111111",
  28667=>"111111111",
  28668=>"111101111",
  28669=>"000000000",
  28670=>"101101111",
  28671=>"100101101",
  28672=>"111111111",
  28673=>"001000000",
  28674=>"111111101",
  28675=>"010111111",
  28676=>"011011111",
  28677=>"111000101",
  28678=>"001001101",
  28679=>"101001101",
  28680=>"111111111",
  28681=>"000000000",
  28682=>"111111111",
  28683=>"100000000",
  28684=>"111000000",
  28685=>"000100100",
  28686=>"100100101",
  28687=>"000000000",
  28688=>"000001000",
  28689=>"111111010",
  28690=>"000100100",
  28691=>"111101111",
  28692=>"111001100",
  28693=>"000000110",
  28694=>"001001111",
  28695=>"001001001",
  28696=>"000010111",
  28697=>"011011000",
  28698=>"000000000",
  28699=>"111111110",
  28700=>"111111111",
  28701=>"101101100",
  28702=>"111011000",
  28703=>"001001111",
  28704=>"100110111",
  28705=>"110110000",
  28706=>"001001000",
  28707=>"101001001",
  28708=>"111011000",
  28709=>"001000101",
  28710=>"110010111",
  28711=>"000001000",
  28712=>"111111110",
  28713=>"010010010",
  28714=>"000000111",
  28715=>"000000000",
  28716=>"001011110",
  28717=>"111111110",
  28718=>"101111111",
  28719=>"000000011",
  28720=>"000010110",
  28721=>"000011011",
  28722=>"100000011",
  28723=>"001011111",
  28724=>"000000000",
  28725=>"000001111",
  28726=>"011010000",
  28727=>"001000100",
  28728=>"000001111",
  28729=>"010010100",
  28730=>"001001111",
  28731=>"001000000",
  28732=>"111010110",
  28733=>"001000000",
  28734=>"001001111",
  28735=>"111000100",
  28736=>"001001000",
  28737=>"010011001",
  28738=>"001000000",
  28739=>"110010000",
  28740=>"010011011",
  28741=>"111011011",
  28742=>"001001001",
  28743=>"001000000",
  28744=>"000100111",
  28745=>"000000000",
  28746=>"000000100",
  28747=>"111001001",
  28748=>"000001111",
  28749=>"000000000",
  28750=>"000000000",
  28751=>"101111111",
  28752=>"001011001",
  28753=>"111111110",
  28754=>"101001111",
  28755=>"011110111",
  28756=>"000000000",
  28757=>"000000100",
  28758=>"001000001",
  28759=>"000001001",
  28760=>"100111110",
  28761=>"101000000",
  28762=>"001000000",
  28763=>"000110100",
  28764=>"000000000",
  28765=>"000000011",
  28766=>"000001111",
  28767=>"100111100",
  28768=>"000100100",
  28769=>"000000000",
  28770=>"101100100",
  28771=>"010011110",
  28772=>"000001001",
  28773=>"111101001",
  28774=>"000000001",
  28775=>"100101000",
  28776=>"000000111",
  28777=>"101101101",
  28778=>"110110001",
  28779=>"111000000",
  28780=>"111111111",
  28781=>"001111111",
  28782=>"101101111",
  28783=>"000111001",
  28784=>"001111111",
  28785=>"110111111",
  28786=>"000000101",
  28787=>"001001111",
  28788=>"000000000",
  28789=>"001101001",
  28790=>"111111110",
  28791=>"001001001",
  28792=>"000110110",
  28793=>"000000000",
  28794=>"001001001",
  28795=>"000001001",
  28796=>"100110110",
  28797=>"101111111",
  28798=>"101101001",
  28799=>"001011111",
  28800=>"001101001",
  28801=>"111111110",
  28802=>"111010000",
  28803=>"111011011",
  28804=>"000101111",
  28805=>"000000000",
  28806=>"000000001",
  28807=>"000000000",
  28808=>"101111111",
  28809=>"001101111",
  28810=>"111101111",
  28811=>"111111111",
  28812=>"101001101",
  28813=>"000000000",
  28814=>"000000101",
  28815=>"000000000",
  28816=>"111111111",
  28817=>"110111111",
  28818=>"001001111",
  28819=>"010111111",
  28820=>"110110010",
  28821=>"000000000",
  28822=>"111000000",
  28823=>"111001011",
  28824=>"000011111",
  28825=>"111100110",
  28826=>"111111111",
  28827=>"010000010",
  28828=>"111111001",
  28829=>"001011111",
  28830=>"101111111",
  28831=>"000000000",
  28832=>"110110000",
  28833=>"101101111",
  28834=>"000100110",
  28835=>"000011011",
  28836=>"001000000",
  28837=>"000111111",
  28838=>"110111111",
  28839=>"011000000",
  28840=>"001001101",
  28841=>"000010000",
  28842=>"111111111",
  28843=>"111001111",
  28844=>"001001001",
  28845=>"110110100",
  28846=>"000000100",
  28847=>"001100110",
  28848=>"110010000",
  28849=>"000000010",
  28850=>"111111110",
  28851=>"111111001",
  28852=>"010010010",
  28853=>"000000000",
  28854=>"111110010",
  28855=>"111111111",
  28856=>"000000100",
  28857=>"001000000",
  28858=>"000001001",
  28859=>"011011111",
  28860=>"000000000",
  28861=>"000000000",
  28862=>"000000100",
  28863=>"100000001",
  28864=>"101000000",
  28865=>"011000000",
  28866=>"101101001",
  28867=>"111111010",
  28868=>"100000111",
  28869=>"010000000",
  28870=>"001001111",
  28871=>"000010111",
  28872=>"000110110",
  28873=>"000000101",
  28874=>"111001111",
  28875=>"110110011",
  28876=>"000000000",
  28877=>"111111001",
  28878=>"111000000",
  28879=>"000000000",
  28880=>"000000000",
  28881=>"110110110",
  28882=>"000110110",
  28883=>"000000100",
  28884=>"000000000",
  28885=>"110011111",
  28886=>"101101000",
  28887=>"110011011",
  28888=>"000111111",
  28889=>"101101101",
  28890=>"000001000",
  28891=>"000101111",
  28892=>"111000000",
  28893=>"111110100",
  28894=>"110111110",
  28895=>"000001100",
  28896=>"001001011",
  28897=>"000100101",
  28898=>"000000000",
  28899=>"000000000",
  28900=>"111011011",
  28901=>"000001101",
  28902=>"000000101",
  28903=>"011000101",
  28904=>"110000111",
  28905=>"010011000",
  28906=>"111111111",
  28907=>"000000000",
  28908=>"011000000",
  28909=>"000110000",
  28910=>"011111100",
  28911=>"000000000",
  28912=>"111000000",
  28913=>"111011111",
  28914=>"111111111",
  28915=>"000000000",
  28916=>"000111001",
  28917=>"001001000",
  28918=>"011111111",
  28919=>"110111100",
  28920=>"011011000",
  28921=>"000000000",
  28922=>"000000000",
  28923=>"000000000",
  28924=>"110100100",
  28925=>"110110110",
  28926=>"011011000",
  28927=>"101100100",
  28928=>"010111011",
  28929=>"111011110",
  28930=>"000000000",
  28931=>"000111111",
  28932=>"000000111",
  28933=>"110010110",
  28934=>"100110111",
  28935=>"110110111",
  28936=>"001000111",
  28937=>"111001000",
  28938=>"001111111",
  28939=>"000101111",
  28940=>"000011011",
  28941=>"111111101",
  28942=>"110110110",
  28943=>"001000000",
  28944=>"001001111",
  28945=>"111111111",
  28946=>"101000000",
  28947=>"101101111",
  28948=>"100000000",
  28949=>"111001001",
  28950=>"011111100",
  28951=>"000000111",
  28952=>"111111111",
  28953=>"111110110",
  28954=>"111111110",
  28955=>"100000110",
  28956=>"010010110",
  28957=>"000000000",
  28958=>"111111111",
  28959=>"101000000",
  28960=>"001111011",
  28961=>"111111111",
  28962=>"000111111",
  28963=>"011001110",
  28964=>"111111110",
  28965=>"000000111",
  28966=>"101101111",
  28967=>"100000110",
  28968=>"101000000",
  28969=>"000000000",
  28970=>"101101110",
  28971=>"000000000",
  28972=>"000000110",
  28973=>"000000100",
  28974=>"001111100",
  28975=>"001001000",
  28976=>"110111111",
  28977=>"011001010",
  28978=>"101001011",
  28979=>"111110111",
  28980=>"001001111",
  28981=>"111111111",
  28982=>"000000000",
  28983=>"000001011",
  28984=>"000000110",
  28985=>"000000001",
  28986=>"000000111",
  28987=>"000000111",
  28988=>"111111000",
  28989=>"000000100",
  28990=>"000000000",
  28991=>"011111111",
  28992=>"010000000",
  28993=>"011001111",
  28994=>"011000011",
  28995=>"000000101",
  28996=>"101101101",
  28997=>"000010111",
  28998=>"000000000",
  28999=>"111001001",
  29000=>"111111000",
  29001=>"000000000",
  29002=>"001011111",
  29003=>"000111111",
  29004=>"101111001",
  29005=>"110110100",
  29006=>"100110110",
  29007=>"100111111",
  29008=>"110111111",
  29009=>"111111110",
  29010=>"110110111",
  29011=>"000000000",
  29012=>"000000000",
  29013=>"011011011",
  29014=>"110010000",
  29015=>"111110110",
  29016=>"011001111",
  29017=>"011111111",
  29018=>"010000000",
  29019=>"101001000",
  29020=>"010011111",
  29021=>"000000000",
  29022=>"000000011",
  29023=>"100111111",
  29024=>"000100000",
  29025=>"010000000",
  29026=>"111111110",
  29027=>"111111110",
  29028=>"100011010",
  29029=>"000000001",
  29030=>"000100000",
  29031=>"111111111",
  29032=>"110110110",
  29033=>"110111111",
  29034=>"111111111",
  29035=>"101000010",
  29036=>"111101111",
  29037=>"001101111",
  29038=>"000000010",
  29039=>"000000110",
  29040=>"111111011",
  29041=>"000000000",
  29042=>"000010010",
  29043=>"000000000",
  29044=>"111010011",
  29045=>"111111111",
  29046=>"111111010",
  29047=>"001000000",
  29048=>"000000000",
  29049=>"110111111",
  29050=>"110110010",
  29051=>"010110110",
  29052=>"101000000",
  29053=>"111101000",
  29054=>"000000000",
  29055=>"111111111",
  29056=>"110110111",
  29057=>"000001001",
  29058=>"000000110",
  29059=>"001001001",
  29060=>"111111000",
  29061=>"001111111",
  29062=>"000000000",
  29063=>"000000110",
  29064=>"111000000",
  29065=>"110100100",
  29066=>"000000001",
  29067=>"101101001",
  29068=>"001001001",
  29069=>"011111110",
  29070=>"000000111",
  29071=>"000000000",
  29072=>"010111010",
  29073=>"111111101",
  29074=>"000000010",
  29075=>"111111000",
  29076=>"111111101",
  29077=>"000000000",
  29078=>"101001100",
  29079=>"000010010",
  29080=>"000000111",
  29081=>"011001001",
  29082=>"000100111",
  29083=>"000000111",
  29084=>"000000011",
  29085=>"000011010",
  29086=>"010010010",
  29087=>"000000101",
  29088=>"000000000",
  29089=>"000010011",
  29090=>"111110110",
  29091=>"000000100",
  29092=>"011111101",
  29093=>"000111111",
  29094=>"011011011",
  29095=>"000000101",
  29096=>"000000100",
  29097=>"110110111",
  29098=>"000000000",
  29099=>"001111110",
  29100=>"001001000",
  29101=>"110110000",
  29102=>"000000100",
  29103=>"110101101",
  29104=>"111000111",
  29105=>"110100110",
  29106=>"000000001",
  29107=>"000000010",
  29108=>"000000011",
  29109=>"001001001",
  29110=>"101101101",
  29111=>"001010110",
  29112=>"011000100",
  29113=>"011000111",
  29114=>"000000000",
  29115=>"111000101",
  29116=>"000000010",
  29117=>"000000000",
  29118=>"000000110",
  29119=>"110111111",
  29120=>"110010000",
  29121=>"001001101",
  29122=>"101101101",
  29123=>"111111111",
  29124=>"001111111",
  29125=>"110110011",
  29126=>"110110010",
  29127=>"111111000",
  29128=>"111111111",
  29129=>"000000000",
  29130=>"111100011",
  29131=>"000000100",
  29132=>"000000000",
  29133=>"000000000",
  29134=>"001000010",
  29135=>"000100111",
  29136=>"111100111",
  29137=>"111110111",
  29138=>"110111010",
  29139=>"000011111",
  29140=>"000000000",
  29141=>"001101100",
  29142=>"000001001",
  29143=>"110100101",
  29144=>"110100110",
  29145=>"100111111",
  29146=>"000000000",
  29147=>"000001101",
  29148=>"110000000",
  29149=>"010010110",
  29150=>"000100111",
  29151=>"001000010",
  29152=>"100000000",
  29153=>"111111111",
  29154=>"101100111",
  29155=>"101101000",
  29156=>"110010010",
  29157=>"000001001",
  29158=>"111111000",
  29159=>"100101111",
  29160=>"000000110",
  29161=>"111110000",
  29162=>"110110000",
  29163=>"111011000",
  29164=>"000000000",
  29165=>"001011000",
  29166=>"000010000",
  29167=>"000000001",
  29168=>"000000111",
  29169=>"110010011",
  29170=>"101001101",
  29171=>"000011111",
  29172=>"111111000",
  29173=>"111100000",
  29174=>"111111000",
  29175=>"000000000",
  29176=>"111000000",
  29177=>"000011011",
  29178=>"101000110",
  29179=>"001000111",
  29180=>"000000000",
  29181=>"110111001",
  29182=>"000000000",
  29183=>"000111111",
  29184=>"110111110",
  29185=>"010010000",
  29186=>"101101111",
  29187=>"000111111",
  29188=>"010010000",
  29189=>"111000000",
  29190=>"000100111",
  29191=>"111111111",
  29192=>"101101001",
  29193=>"111111011",
  29194=>"000000000",
  29195=>"100100000",
  29196=>"000000010",
  29197=>"111000000",
  29198=>"011001000",
  29199=>"000000000",
  29200=>"000100111",
  29201=>"000000011",
  29202=>"000000111",
  29203=>"111110000",
  29204=>"000000000",
  29205=>"000000000",
  29206=>"111111111",
  29207=>"000000011",
  29208=>"000110111",
  29209=>"000000000",
  29210=>"011000000",
  29211=>"000111111",
  29212=>"111000000",
  29213=>"111101000",
  29214=>"100110110",
  29215=>"110000000",
  29216=>"111000000",
  29217=>"110100100",
  29218=>"110110110",
  29219=>"111111111",
  29220=>"111111000",
  29221=>"111111111",
  29222=>"000000000",
  29223=>"110101111",
  29224=>"111111011",
  29225=>"011010010",
  29226=>"000010000",
  29227=>"000000011",
  29228=>"101000111",
  29229=>"110000110",
  29230=>"000000000",
  29231=>"111000000",
  29232=>"110000000",
  29233=>"000000000",
  29234=>"100000000",
  29235=>"001011011",
  29236=>"111111100",
  29237=>"111110100",
  29238=>"100100111",
  29239=>"111011011",
  29240=>"000000000",
  29241=>"111111000",
  29242=>"000000000",
  29243=>"011100111",
  29244=>"111111000",
  29245=>"001011111",
  29246=>"110110011",
  29247=>"111111110",
  29248=>"001001001",
  29249=>"000100101",
  29250=>"000100110",
  29251=>"111111111",
  29252=>"000000110",
  29253=>"011001000",
  29254=>"000111111",
  29255=>"000000000",
  29256=>"001000000",
  29257=>"000000000",
  29258=>"100111101",
  29259=>"101000000",
  29260=>"111001000",
  29261=>"000000001",
  29262=>"000111111",
  29263=>"000011111",
  29264=>"000110111",
  29265=>"000000000",
  29266=>"000110000",
  29267=>"100001111",
  29268=>"100000000",
  29269=>"111111111",
  29270=>"001000000",
  29271=>"010010010",
  29272=>"000000001",
  29273=>"111100000",
  29274=>"000100000",
  29275=>"000000000",
  29276=>"010000000",
  29277=>"000111111",
  29278=>"111111101",
  29279=>"100000000",
  29280=>"000000000",
  29281=>"010110111",
  29282=>"101000000",
  29283=>"000000100",
  29284=>"000000000",
  29285=>"111111111",
  29286=>"111110110",
  29287=>"100000000",
  29288=>"111111001",
  29289=>"111010000",
  29290=>"001000000",
  29291=>"100100110",
  29292=>"000011001",
  29293=>"111101111",
  29294=>"111111111",
  29295=>"111111110",
  29296=>"000000110",
  29297=>"111000000",
  29298=>"111111111",
  29299=>"000000000",
  29300=>"011000000",
  29301=>"000110110",
  29302=>"111000000",
  29303=>"000000000",
  29304=>"000111010",
  29305=>"011001001",
  29306=>"000000010",
  29307=>"000110111",
  29308=>"001111111",
  29309=>"111111111",
  29310=>"000000000",
  29311=>"000000000",
  29312=>"101001000",
  29313=>"000000100",
  29314=>"000000000",
  29315=>"000000000",
  29316=>"001000000",
  29317=>"110000000",
  29318=>"010111111",
  29319=>"111111111",
  29320=>"000000100",
  29321=>"000000000",
  29322=>"000000000",
  29323=>"100111111",
  29324=>"000000111",
  29325=>"111111111",
  29326=>"011000000",
  29327=>"000000111",
  29328=>"110000000",
  29329=>"011000000",
  29330=>"110111111",
  29331=>"000000000",
  29332=>"111111000",
  29333=>"010110111",
  29334=>"000000000",
  29335=>"111001000",
  29336=>"010000111",
  29337=>"001000000",
  29338=>"000000010",
  29339=>"111001000",
  29340=>"000000001",
  29341=>"100000000",
  29342=>"000000000",
  29343=>"111111111",
  29344=>"011110000",
  29345=>"111100100",
  29346=>"100000000",
  29347=>"101000100",
  29348=>"100000010",
  29349=>"111000000",
  29350=>"111000000",
  29351=>"010111111",
  29352=>"001001000",
  29353=>"000000000",
  29354=>"001111111",
  29355=>"111111111",
  29356=>"000000000",
  29357=>"000110110",
  29358=>"000001001",
  29359=>"000001101",
  29360=>"000011010",
  29361=>"101000001",
  29362=>"110010010",
  29363=>"111111010",
  29364=>"000000000",
  29365=>"111111111",
  29366=>"110100110",
  29367=>"000000000",
  29368=>"000001001",
  29369=>"111111111",
  29370=>"111000000",
  29371=>"111100011",
  29372=>"111111011",
  29373=>"011011000",
  29374=>"100111111",
  29375=>"011001000",
  29376=>"111111111",
  29377=>"000000000",
  29378=>"000000000",
  29379=>"111111111",
  29380=>"000000000",
  29381=>"111000000",
  29382=>"000001111",
  29383=>"000000001",
  29384=>"000000000",
  29385=>"000010000",
  29386=>"000000000",
  29387=>"000000000",
  29388=>"111111111",
  29389=>"000110010",
  29390=>"111000000",
  29391=>"110100110",
  29392=>"100000000",
  29393=>"111000000",
  29394=>"000110111",
  29395=>"000000000",
  29396=>"000000000",
  29397=>"111110000",
  29398=>"111110100",
  29399=>"000000011",
  29400=>"000000000",
  29401=>"000000111",
  29402=>"000000000",
  29403=>"000111111",
  29404=>"111111111",
  29405=>"001001001",
  29406=>"011000000",
  29407=>"011011111",
  29408=>"111110100",
  29409=>"111111111",
  29410=>"111111111",
  29411=>"101101001",
  29412=>"000000000",
  29413=>"000000000",
  29414=>"111111111",
  29415=>"000000111",
  29416=>"111111111",
  29417=>"111000000",
  29418=>"111111111",
  29419=>"000111110",
  29420=>"000000000",
  29421=>"000100110",
  29422=>"111000100",
  29423=>"000000000",
  29424=>"000100100",
  29425=>"000000111",
  29426=>"000101111",
  29427=>"111011000",
  29428=>"111011001",
  29429=>"001000100",
  29430=>"001111111",
  29431=>"110111110",
  29432=>"101100111",
  29433=>"111010010",
  29434=>"000000000",
  29435=>"110111111",
  29436=>"100000000",
  29437=>"111000000",
  29438=>"111111111",
  29439=>"111111111",
  29440=>"000011110",
  29441=>"011111000",
  29442=>"001000000",
  29443=>"111111111",
  29444=>"000001001",
  29445=>"111100110",
  29446=>"101001101",
  29447=>"011010111",
  29448=>"000000000",
  29449=>"000000100",
  29450=>"111111111",
  29451=>"011111111",
  29452=>"001101111",
  29453=>"000000000",
  29454=>"100001111",
  29455=>"111111100",
  29456=>"111111111",
  29457=>"001011000",
  29458=>"100000111",
  29459=>"100100000",
  29460=>"000000000",
  29461=>"000000000",
  29462=>"111100100",
  29463=>"111111001",
  29464=>"000000000",
  29465=>"111000000",
  29466=>"000000000",
  29467=>"001000000",
  29468=>"101000000",
  29469=>"000000011",
  29470=>"111111111",
  29471=>"111111111",
  29472=>"000100001",
  29473=>"000000000",
  29474=>"000001111",
  29475=>"111111111",
  29476=>"000101111",
  29477=>"111111111",
  29478=>"110111111",
  29479=>"000000001",
  29480=>"111111111",
  29481=>"000000000",
  29482=>"101000000",
  29483=>"111111000",
  29484=>"000000000",
  29485=>"100100110",
  29486=>"000000000",
  29487=>"000001111",
  29488=>"111111111",
  29489=>"111111111",
  29490=>"000000000",
  29491=>"111000111",
  29492=>"000111111",
  29493=>"000001011",
  29494=>"111011011",
  29495=>"111011111",
  29496=>"000100000",
  29497=>"111000000",
  29498=>"100000000",
  29499=>"000001111",
  29500=>"110111111",
  29501=>"111111000",
  29502=>"111111011",
  29503=>"000110000",
  29504=>"111001000",
  29505=>"111111100",
  29506=>"111000001",
  29507=>"110000000",
  29508=>"000000111",
  29509=>"000000000",
  29510=>"000111111",
  29511=>"001001001",
  29512=>"010000000",
  29513=>"001000101",
  29514=>"000011111",
  29515=>"000001001",
  29516=>"101110110",
  29517=>"000000000",
  29518=>"111111111",
  29519=>"110110110",
  29520=>"100111001",
  29521=>"111111000",
  29522=>"000001000",
  29523=>"111111101",
  29524=>"000101111",
  29525=>"001000000",
  29526=>"100001001",
  29527=>"000111111",
  29528=>"011111111",
  29529=>"000000010",
  29530=>"011000000",
  29531=>"010011111",
  29532=>"111100111",
  29533=>"111111110",
  29534=>"000000000",
  29535=>"110110110",
  29536=>"001111111",
  29537=>"000000000",
  29538=>"111011001",
  29539=>"111111111",
  29540=>"111111101",
  29541=>"000000000",
  29542=>"111111111",
  29543=>"001011001",
  29544=>"000100000",
  29545=>"111111110",
  29546=>"000000000",
  29547=>"100100000",
  29548=>"000000000",
  29549=>"000000000",
  29550=>"111110111",
  29551=>"001111111",
  29552=>"111111001",
  29553=>"111111111",
  29554=>"100010111",
  29555=>"000000000",
  29556=>"111000000",
  29557=>"111111111",
  29558=>"000000000",
  29559=>"000000111",
  29560=>"000000010",
  29561=>"111101111",
  29562=>"010000000",
  29563=>"000000011",
  29564=>"111111111",
  29565=>"111111111",
  29566=>"111111110",
  29567=>"001001001",
  29568=>"000000000",
  29569=>"111111100",
  29570=>"111000000",
  29571=>"111111000",
  29572=>"011011111",
  29573=>"000100100",
  29574=>"000000110",
  29575=>"000000000",
  29576=>"000010111",
  29577=>"011111011",
  29578=>"000000000",
  29579=>"110100100",
  29580=>"111001000",
  29581=>"111110110",
  29582=>"000000001",
  29583=>"111000100",
  29584=>"110110000",
  29585=>"101110000",
  29586=>"111111111",
  29587=>"111111111",
  29588=>"000001111",
  29589=>"000000000",
  29590=>"111100101",
  29591=>"110100110",
  29592=>"000100111",
  29593=>"100100000",
  29594=>"111000000",
  29595=>"001011001",
  29596=>"111111111",
  29597=>"111111111",
  29598=>"111111111",
  29599=>"100000000",
  29600=>"000000001",
  29601=>"111111011",
  29602=>"001001000",
  29603=>"000101111",
  29604=>"111011001",
  29605=>"000000000",
  29606=>"000000000",
  29607=>"000111111",
  29608=>"000000000",
  29609=>"000000000",
  29610=>"110111111",
  29611=>"111111111",
  29612=>"000110110",
  29613=>"110110000",
  29614=>"111111111",
  29615=>"000001011",
  29616=>"000000000",
  29617=>"000000100",
  29618=>"000000111",
  29619=>"111111011",
  29620=>"000110111",
  29621=>"000101111",
  29622=>"111111101",
  29623=>"111000000",
  29624=>"011111111",
  29625=>"001011000",
  29626=>"111011010",
  29627=>"111111111",
  29628=>"111111111",
  29629=>"111111111",
  29630=>"100000000",
  29631=>"111100100",
  29632=>"111111000",
  29633=>"000000000",
  29634=>"111111110",
  29635=>"000000000",
  29636=>"111011101",
  29637=>"111100000",
  29638=>"111000111",
  29639=>"111100000",
  29640=>"000010001",
  29641=>"110010000",
  29642=>"000010011",
  29643=>"111011000",
  29644=>"100000010",
  29645=>"111000000",
  29646=>"000111111",
  29647=>"110000000",
  29648=>"111111111",
  29649=>"111111111",
  29650=>"000000110",
  29651=>"001000100",
  29652=>"100100110",
  29653=>"111011000",
  29654=>"000000000",
  29655=>"000000000",
  29656=>"000000000",
  29657=>"000111111",
  29658=>"000111111",
  29659=>"000000100",
  29660=>"011001001",
  29661=>"100101111",
  29662=>"111000000",
  29663=>"000110000",
  29664=>"111100000",
  29665=>"111111111",
  29666=>"001001111",
  29667=>"111110110",
  29668=>"111011000",
  29669=>"111001000",
  29670=>"111001000",
  29671=>"111111000",
  29672=>"000000100",
  29673=>"100100001",
  29674=>"000110010",
  29675=>"001000000",
  29676=>"000101111",
  29677=>"011011011",
  29678=>"111111111",
  29679=>"100110111",
  29680=>"111111000",
  29681=>"110110011",
  29682=>"111100100",
  29683=>"110101101",
  29684=>"000011000",
  29685=>"110001111",
  29686=>"111111111",
  29687=>"101100100",
  29688=>"000111111",
  29689=>"111011001",
  29690=>"000000100",
  29691=>"000010110",
  29692=>"000000000",
  29693=>"110110000",
  29694=>"100000100",
  29695=>"000000110",
  29696=>"100000100",
  29697=>"000100101",
  29698=>"000111111",
  29699=>"000000001",
  29700=>"000101111",
  29701=>"011011000",
  29702=>"001001111",
  29703=>"101111111",
  29704=>"111110000",
  29705=>"110111111",
  29706=>"011000111",
  29707=>"000010110",
  29708=>"001111111",
  29709=>"000000001",
  29710=>"000111111",
  29711=>"000000000",
  29712=>"110110010",
  29713=>"000000000",
  29714=>"000000010",
  29715=>"000100111",
  29716=>"000010011",
  29717=>"000000000",
  29718=>"111110110",
  29719=>"111011000",
  29720=>"111101111",
  29721=>"101000110",
  29722=>"010111101",
  29723=>"110100000",
  29724=>"111111111",
  29725=>"000000110",
  29726=>"000001111",
  29727=>"111110001",
  29728=>"000000101",
  29729=>"000111110",
  29730=>"111110111",
  29731=>"000111111",
  29732=>"110010111",
  29733=>"100110000",
  29734=>"000001010",
  29735=>"000111111",
  29736=>"111111110",
  29737=>"000000111",
  29738=>"111111111",
  29739=>"101111111",
  29740=>"000000011",
  29741=>"111111111",
  29742=>"000000111",
  29743=>"000000000",
  29744=>"000000001",
  29745=>"000000000",
  29746=>"001001000",
  29747=>"101111001",
  29748=>"000111111",
  29749=>"000001001",
  29750=>"010000001",
  29751=>"001001011",
  29752=>"000000111",
  29753=>"000000000",
  29754=>"000000000",
  29755=>"000101100",
  29756=>"000000111",
  29757=>"000010111",
  29758=>"100110110",
  29759=>"111001011",
  29760=>"111000000",
  29761=>"000000010",
  29762=>"000110111",
  29763=>"100111011",
  29764=>"110011000",
  29765=>"001111000",
  29766=>"000000000",
  29767=>"011001000",
  29768=>"000001010",
  29769=>"000000111",
  29770=>"100101100",
  29771=>"011001111",
  29772=>"001101111",
  29773=>"111111011",
  29774=>"111111101",
  29775=>"001000111",
  29776=>"000000000",
  29777=>"001000000",
  29778=>"100000000",
  29779=>"001001000",
  29780=>"011111010",
  29781=>"000000000",
  29782=>"100110111",
  29783=>"000011111",
  29784=>"000000000",
  29785=>"000000000",
  29786=>"111111000",
  29787=>"000011001",
  29788=>"010000000",
  29789=>"000000000",
  29790=>"011011111",
  29791=>"000000000",
  29792=>"000111111",
  29793=>"111000101",
  29794=>"000000000",
  29795=>"001111010",
  29796=>"111110111",
  29797=>"111000101",
  29798=>"100000000",
  29799=>"000000001",
  29800=>"000111111",
  29801=>"111100000",
  29802=>"000010111",
  29803=>"011011011",
  29804=>"001001100",
  29805=>"111111000",
  29806=>"000000000",
  29807=>"001111000",
  29808=>"000000000",
  29809=>"111000011",
  29810=>"000011111",
  29811=>"111011000",
  29812=>"101111000",
  29813=>"000000110",
  29814=>"111111000",
  29815=>"111111111",
  29816=>"000000111",
  29817=>"001000000",
  29818=>"001011011",
  29819=>"101000000",
  29820=>"000011111",
  29821=>"000010010",
  29822=>"001011000",
  29823=>"011111111",
  29824=>"000000001",
  29825=>"111000000",
  29826=>"000000011",
  29827=>"000100000",
  29828=>"100111101",
  29829=>"000000111",
  29830=>"000100100",
  29831=>"111001000",
  29832=>"111000000",
  29833=>"000011000",
  29834=>"000000111",
  29835=>"100110000",
  29836=>"011111011",
  29837=>"001000000",
  29838=>"111000111",
  29839=>"000101011",
  29840=>"000110111",
  29841=>"111111101",
  29842=>"111110110",
  29843=>"000111000",
  29844=>"001001000",
  29845=>"000001000",
  29846=>"111111011",
  29847=>"111111001",
  29848=>"011001111",
  29849=>"110110001",
  29850=>"010000110",
  29851=>"111111000",
  29852=>"111001010",
  29853=>"111110000",
  29854=>"110111110",
  29855=>"111111111",
  29856=>"001011110",
  29857=>"111100100",
  29858=>"111101000",
  29859=>"100000000",
  29860=>"011001011",
  29861=>"111101100",
  29862=>"111111000",
  29863=>"110110100",
  29864=>"000000001",
  29865=>"000111111",
  29866=>"111011000",
  29867=>"111001111",
  29868=>"111111000",
  29869=>"100111100",
  29870=>"000000111",
  29871=>"000000000",
  29872=>"111100100",
  29873=>"111111010",
  29874=>"111111000",
  29875=>"111101000",
  29876=>"000010000",
  29877=>"010000111",
  29878=>"111000000",
  29879=>"100111111",
  29880=>"001011011",
  29881=>"000010111",
  29882=>"011000001",
  29883=>"110000110",
  29884=>"011000000",
  29885=>"011111110",
  29886=>"111000000",
  29887=>"111000001",
  29888=>"000100000",
  29889=>"000000000",
  29890=>"111111000",
  29891=>"111111111",
  29892=>"000111111",
  29893=>"000101111",
  29894=>"010111111",
  29895=>"000111000",
  29896=>"111111110",
  29897=>"000011111",
  29898=>"000011001",
  29899=>"000111110",
  29900=>"100100000",
  29901=>"111111100",
  29902=>"000000000",
  29903=>"011000011",
  29904=>"111101000",
  29905=>"000000011",
  29906=>"000000000",
  29907=>"011111111",
  29908=>"110100110",
  29909=>"111111110",
  29910=>"000000011",
  29911=>"000111111",
  29912=>"000000110",
  29913=>"111111111",
  29914=>"000010111",
  29915=>"100100111",
  29916=>"011111110",
  29917=>"111111111",
  29918=>"111100000",
  29919=>"001011111",
  29920=>"101001000",
  29921=>"000000010",
  29922=>"111111100",
  29923=>"111011011",
  29924=>"010000111",
  29925=>"110110110",
  29926=>"000010011",
  29927=>"111010000",
  29928=>"000111101",
  29929=>"011000111",
  29930=>"100100111",
  29931=>"011111111",
  29932=>"110000000",
  29933=>"000000000",
  29934=>"111001101",
  29935=>"111111100",
  29936=>"111111011",
  29937=>"111110110",
  29938=>"100000110",
  29939=>"010000001",
  29940=>"000001111",
  29941=>"110000011",
  29942=>"101111001",
  29943=>"111000000",
  29944=>"000111111",
  29945=>"001111111",
  29946=>"111111111",
  29947=>"000111111",
  29948=>"000000111",
  29949=>"110001000",
  29950=>"111101101",
  29951=>"011111110",
  29952=>"000000110",
  29953=>"000000011",
  29954=>"111111001",
  29955=>"111111111",
  29956=>"000000000",
  29957=>"000001111",
  29958=>"111110000",
  29959=>"000000111",
  29960=>"011000000",
  29961=>"000000000",
  29962=>"111000000",
  29963=>"001000011",
  29964=>"001001111",
  29965=>"111101100",
  29966=>"001011000",
  29967=>"010000111",
  29968=>"111000111",
  29969=>"010001000",
  29970=>"000010001",
  29971=>"010000000",
  29972=>"000000000",
  29973=>"000111111",
  29974=>"000000011",
  29975=>"000000000",
  29976=>"001100100",
  29977=>"101001000",
  29978=>"001001011",
  29979=>"111001011",
  29980=>"100101111",
  29981=>"111111010",
  29982=>"011000000",
  29983=>"111000011",
  29984=>"110111011",
  29985=>"000000000",
  29986=>"000000000",
  29987=>"000000011",
  29988=>"000000010",
  29989=>"001000011",
  29990=>"101100111",
  29991=>"010011011",
  29992=>"000111111",
  29993=>"000000000",
  29994=>"111000011",
  29995=>"111000010",
  29996=>"000111111",
  29997=>"110100110",
  29998=>"111000000",
  29999=>"000000001",
  30000=>"111111001",
  30001=>"011111111",
  30002=>"001001111",
  30003=>"001010000",
  30004=>"111101000",
  30005=>"111000100",
  30006=>"111111001",
  30007=>"110000000",
  30008=>"000111011",
  30009=>"111000111",
  30010=>"111011111",
  30011=>"000000111",
  30012=>"100000000",
  30013=>"111111000",
  30014=>"111111111",
  30015=>"001100101",
  30016=>"111100000",
  30017=>"110100110",
  30018=>"000011111",
  30019=>"110111111",
  30020=>"100101001",
  30021=>"100010111",
  30022=>"000000010",
  30023=>"011111000",
  30024=>"000111011",
  30025=>"000111110",
  30026=>"100100001",
  30027=>"000000101",
  30028=>"011011000",
  30029=>"111000000",
  30030=>"010110110",
  30031=>"000000101",
  30032=>"111101000",
  30033=>"111011011",
  30034=>"000110111",
  30035=>"111011000",
  30036=>"000111111",
  30037=>"011110010",
  30038=>"111000111",
  30039=>"001111100",
  30040=>"000000111",
  30041=>"101111100",
  30042=>"000110110",
  30043=>"000000000",
  30044=>"110000000",
  30045=>"000100111",
  30046=>"101001111",
  30047=>"001110100",
  30048=>"000111000",
  30049=>"111111011",
  30050=>"101101111",
  30051=>"000000000",
  30052=>"000000110",
  30053=>"111111000",
  30054=>"001111111",
  30055=>"111111000",
  30056=>"100100001",
  30057=>"000111101",
  30058=>"000111101",
  30059=>"110000000",
  30060=>"001011001",
  30061=>"111011000",
  30062=>"000000000",
  30063=>"100001000",
  30064=>"111111111",
  30065=>"111111000",
  30066=>"001000111",
  30067=>"100000000",
  30068=>"111111111",
  30069=>"011111111",
  30070=>"100000110",
  30071=>"100101001",
  30072=>"111110111",
  30073=>"000111100",
  30074=>"001111111",
  30075=>"011000111",
  30076=>"111111111",
  30077=>"000000111",
  30078=>"001000001",
  30079=>"001000000",
  30080=>"011110000",
  30081=>"101101111",
  30082=>"110110000",
  30083=>"000000000",
  30084=>"000100100",
  30085=>"000000000",
  30086=>"011011101",
  30087=>"000000000",
  30088=>"111111111",
  30089=>"011110111",
  30090=>"111111011",
  30091=>"001101001",
  30092=>"111001001",
  30093=>"100100001",
  30094=>"000000000",
  30095=>"000000011",
  30096=>"111111111",
  30097=>"111000000",
  30098=>"000001000",
  30099=>"111000111",
  30100=>"000000111",
  30101=>"000000000",
  30102=>"000000000",
  30103=>"111011111",
  30104=>"101001001",
  30105=>"111111111",
  30106=>"001111111",
  30107=>"000000000",
  30108=>"000000010",
  30109=>"110111111",
  30110=>"110111111",
  30111=>"000000000",
  30112=>"011111011",
  30113=>"001010010",
  30114=>"000000111",
  30115=>"111111000",
  30116=>"000000111",
  30117=>"101111111",
  30118=>"000000000",
  30119=>"111101101",
  30120=>"000110000",
  30121=>"111111000",
  30122=>"110100101",
  30123=>"110000110",
  30124=>"000111000",
  30125=>"111110110",
  30126=>"010000100",
  30127=>"000000010",
  30128=>"111111110",
  30129=>"111011111",
  30130=>"111101111",
  30131=>"111111011",
  30132=>"111111110",
  30133=>"110111111",
  30134=>"111010111",
  30135=>"001000000",
  30136=>"111111000",
  30137=>"110010011",
  30138=>"000000000",
  30139=>"000010110",
  30140=>"000000011",
  30141=>"110000000",
  30142=>"000101000",
  30143=>"000011011",
  30144=>"000000111",
  30145=>"000000000",
  30146=>"111111000",
  30147=>"000111000",
  30148=>"100000111",
  30149=>"000010111",
  30150=>"101101000",
  30151=>"000000000",
  30152=>"011000111",
  30153=>"000100101",
  30154=>"000000101",
  30155=>"011011000",
  30156=>"111011000",
  30157=>"111011000",
  30158=>"000001111",
  30159=>"111111110",
  30160=>"000000100",
  30161=>"110000000",
  30162=>"001000011",
  30163=>"000111111",
  30164=>"011010011",
  30165=>"110110111",
  30166=>"111111111",
  30167=>"000000111",
  30168=>"101100111",
  30169=>"111000000",
  30170=>"000010000",
  30171=>"111111110",
  30172=>"000111111",
  30173=>"111000000",
  30174=>"001001000",
  30175=>"011111111",
  30176=>"011111110",
  30177=>"111000000",
  30178=>"111110110",
  30179=>"000100111",
  30180=>"111000111",
  30181=>"110111111",
  30182=>"111000111",
  30183=>"100110011",
  30184=>"000000100",
  30185=>"101000000",
  30186=>"010011111",
  30187=>"000100111",
  30188=>"100110111",
  30189=>"111100100",
  30190=>"000111111",
  30191=>"111010000",
  30192=>"111111111",
  30193=>"111111001",
  30194=>"001000001",
  30195=>"000000111",
  30196=>"000000000",
  30197=>"000111111",
  30198=>"001111111",
  30199=>"111001001",
  30200=>"110000000",
  30201=>"011000011",
  30202=>"111111100",
  30203=>"111000000",
  30204=>"100000111",
  30205=>"010000000",
  30206=>"000001001",
  30207=>"000000010",
  30208=>"110110010",
  30209=>"110111111",
  30210=>"100000001",
  30211=>"110111010",
  30212=>"111011111",
  30213=>"000000100",
  30214=>"101000001",
  30215=>"111111111",
  30216=>"001111111",
  30217=>"111111111",
  30218=>"000000000",
  30219=>"000000000",
  30220=>"001001111",
  30221=>"111111111",
  30222=>"000000001",
  30223=>"000000001",
  30224=>"110001001",
  30225=>"110111111",
  30226=>"100100100",
  30227=>"111111110",
  30228=>"111101000",
  30229=>"000000001",
  30230=>"010111111",
  30231=>"000000000",
  30232=>"110110110",
  30233=>"011011101",
  30234=>"000000000",
  30235=>"001001001",
  30236=>"001000000",
  30237=>"111111111",
  30238=>"001011011",
  30239=>"111111010",
  30240=>"110110011",
  30241=>"111111111",
  30242=>"001000101",
  30243=>"000101111",
  30244=>"111111100",
  30245=>"110110111",
  30246=>"111111111",
  30247=>"000000001",
  30248=>"000000000",
  30249=>"000000000",
  30250=>"101000100",
  30251=>"000000111",
  30252=>"101111111",
  30253=>"111111111",
  30254=>"000001101",
  30255=>"111000000",
  30256=>"111111010",
  30257=>"000000001",
  30258=>"111111000",
  30259=>"111111010",
  30260=>"000000100",
  30261=>"001011111",
  30262=>"000100001",
  30263=>"001000001",
  30264=>"011110000",
  30265=>"000000110",
  30266=>"001000001",
  30267=>"101111111",
  30268=>"000000000",
  30269=>"000000000",
  30270=>"011111111",
  30271=>"001000111",
  30272=>"011110000",
  30273=>"000111000",
  30274=>"101101111",
  30275=>"001011001",
  30276=>"010110000",
  30277=>"110000000",
  30278=>"100011111",
  30279=>"111111111",
  30280=>"000000000",
  30281=>"000000111",
  30282=>"111111001",
  30283=>"000000000",
  30284=>"010000001",
  30285=>"001011011",
  30286=>"000000000",
  30287=>"001000000",
  30288=>"111111000",
  30289=>"110111111",
  30290=>"000000000",
  30291=>"111110000",
  30292=>"010111010",
  30293=>"011011010",
  30294=>"001011001",
  30295=>"110111110",
  30296=>"000000000",
  30297=>"000000111",
  30298=>"100001111",
  30299=>"110111100",
  30300=>"000000000",
  30301=>"011011000",
  30302=>"000000110",
  30303=>"111111110",
  30304=>"000000000",
  30305=>"111110010",
  30306=>"000000111",
  30307=>"101111111",
  30308=>"000000000",
  30309=>"001111111",
  30310=>"001001111",
  30311=>"000001001",
  30312=>"111111111",
  30313=>"001101111",
  30314=>"111011000",
  30315=>"000000101",
  30316=>"010010010",
  30317=>"000000000",
  30318=>"000000111",
  30319=>"000000000",
  30320=>"000000000",
  30321=>"001000101",
  30322=>"111110101",
  30323=>"000000000",
  30324=>"000000000",
  30325=>"100100111",
  30326=>"111111101",
  30327=>"111111111",
  30328=>"000111111",
  30329=>"111011001",
  30330=>"100000111",
  30331=>"111000100",
  30332=>"100110110",
  30333=>"000000001",
  30334=>"110110111",
  30335=>"010110000",
  30336=>"111111111",
  30337=>"000000111",
  30338=>"000000111",
  30339=>"010110000",
  30340=>"010011011",
  30341=>"111101111",
  30342=>"000000000",
  30343=>"000000000",
  30344=>"000000111",
  30345=>"100101111",
  30346=>"000000000",
  30347=>"111111001",
  30348=>"001010110",
  30349=>"100111110",
  30350=>"111000100",
  30351=>"101000000",
  30352=>"101001111",
  30353=>"110110000",
  30354=>"001000100",
  30355=>"010111000",
  30356=>"111111010",
  30357=>"100101111",
  30358=>"111101100",
  30359=>"111111111",
  30360=>"000000001",
  30361=>"000000101",
  30362=>"111111111",
  30363=>"111111011",
  30364=>"000000111",
  30365=>"001000000",
  30366=>"111111101",
  30367=>"001000000",
  30368=>"111111111",
  30369=>"011111111",
  30370=>"000001000",
  30371=>"011011010",
  30372=>"111001001",
  30373=>"000001011",
  30374=>"111111111",
  30375=>"001101100",
  30376=>"000000000",
  30377=>"001000000",
  30378=>"000110111",
  30379=>"011001011",
  30380=>"000001111",
  30381=>"110110000",
  30382=>"000000001",
  30383=>"111111110",
  30384=>"010111000",
  30385=>"110111011",
  30386=>"111111110",
  30387=>"010000000",
  30388=>"000010010",
  30389=>"000111111",
  30390=>"011000000",
  30391=>"111100101",
  30392=>"000000000",
  30393=>"100100111",
  30394=>"111000000",
  30395=>"011111111",
  30396=>"110111110",
  30397=>"111001001",
  30398=>"110111111",
  30399=>"000000100",
  30400=>"110000000",
  30401=>"110110110",
  30402=>"000100100",
  30403=>"000010111",
  30404=>"001111111",
  30405=>"111101000",
  30406=>"001101000",
  30407=>"000111000",
  30408=>"000000010",
  30409=>"000000101",
  30410=>"011000000",
  30411=>"111111000",
  30412=>"011011111",
  30413=>"101001000",
  30414=>"000000000",
  30415=>"011110111",
  30416=>"111111111",
  30417=>"000010111",
  30418=>"111111110",
  30419=>"001001111",
  30420=>"001000000",
  30421=>"110110110",
  30422=>"100100111",
  30423=>"011001001",
  30424=>"111111000",
  30425=>"100110110",
  30426=>"000000111",
  30427=>"011011001",
  30428=>"111101100",
  30429=>"111111111",
  30430=>"111111110",
  30431=>"111111111",
  30432=>"000000000",
  30433=>"000010110",
  30434=>"111111010",
  30435=>"000001111",
  30436=>"111001001",
  30437=>"111111011",
  30438=>"000000000",
  30439=>"001001001",
  30440=>"101111111",
  30441=>"000011010",
  30442=>"111111111",
  30443=>"111111111",
  30444=>"101101101",
  30445=>"000000100",
  30446=>"000001111",
  30447=>"000001101",
  30448=>"111011100",
  30449=>"101100111",
  30450=>"111111001",
  30451=>"000000101",
  30452=>"111110010",
  30453=>"110110010",
  30454=>"011011001",
  30455=>"010111111",
  30456=>"001101111",
  30457=>"111111111",
  30458=>"001001000",
  30459=>"000000010",
  30460=>"000000000",
  30461=>"000000000",
  30462=>"111001000",
  30463=>"111111111",
  30464=>"111111111",
  30465=>"001000001",
  30466=>"000000000",
  30467=>"011111111",
  30468=>"111110110",
  30469=>"111111000",
  30470=>"111001111",
  30471=>"111111001",
  30472=>"100000000",
  30473=>"000001000",
  30474=>"111111111",
  30475=>"001001100",
  30476=>"000000000",
  30477=>"110000000",
  30478=>"111111011",
  30479=>"111111111",
  30480=>"010110110",
  30481=>"100100010",
  30482=>"110100000",
  30483=>"010111010",
  30484=>"101000000",
  30485=>"110110000",
  30486=>"111011011",
  30487=>"111111010",
  30488=>"110110000",
  30489=>"001101101",
  30490=>"000010111",
  30491=>"101001101",
  30492=>"100001001",
  30493=>"101101111",
  30494=>"111111111",
  30495=>"100000000",
  30496=>"111111000",
  30497=>"111111010",
  30498=>"111110010",
  30499=>"111000000",
  30500=>"111010000",
  30501=>"111111110",
  30502=>"111000100",
  30503=>"101101111",
  30504=>"111100111",
  30505=>"000000100",
  30506=>"000000100",
  30507=>"000000000",
  30508=>"111111011",
  30509=>"000000100",
  30510=>"011110110",
  30511=>"001000000",
  30512=>"110110111",
  30513=>"100000111",
  30514=>"111111111",
  30515=>"000000100",
  30516=>"110000000",
  30517=>"011011000",
  30518=>"000000110",
  30519=>"000110111",
  30520=>"000000000",
  30521=>"101000100",
  30522=>"000000001",
  30523=>"100101000",
  30524=>"000011001",
  30525=>"010010000",
  30526=>"000000001",
  30527=>"000000001",
  30528=>"000000101",
  30529=>"111111000",
  30530=>"000000000",
  30531=>"001000111",
  30532=>"111110010",
  30533=>"000101111",
  30534=>"000000000",
  30535=>"111111111",
  30536=>"000000000",
  30537=>"110111110",
  30538=>"111111110",
  30539=>"000000000",
  30540=>"111000000",
  30541=>"000000001",
  30542=>"110000000",
  30543=>"111111111",
  30544=>"011001000",
  30545=>"000101111",
  30546=>"111111110",
  30547=>"110000000",
  30548=>"000000000",
  30549=>"011011011",
  30550=>"111000000",
  30551=>"000000111",
  30552=>"111111000",
  30553=>"110111110",
  30554=>"111000000",
  30555=>"000000001",
  30556=>"000000000",
  30557=>"000000000",
  30558=>"111001000",
  30559=>"000011000",
  30560=>"111111110",
  30561=>"111001000",
  30562=>"101111110",
  30563=>"110110111",
  30564=>"100001001",
  30565=>"001000000",
  30566=>"000000001",
  30567=>"000000000",
  30568=>"010000000",
  30569=>"000110110",
  30570=>"111101101",
  30571=>"110100100",
  30572=>"110110110",
  30573=>"000001111",
  30574=>"000000101",
  30575=>"111111111",
  30576=>"010000010",
  30577=>"111111010",
  30578=>"010111111",
  30579=>"110000011",
  30580=>"000000001",
  30581=>"000000101",
  30582=>"101000000",
  30583=>"000000000",
  30584=>"101000111",
  30585=>"111111010",
  30586=>"111111111",
  30587=>"000000110",
  30588=>"111111010",
  30589=>"111111110",
  30590=>"000000001",
  30591=>"000000001",
  30592=>"000000001",
  30593=>"000000000",
  30594=>"011001011",
  30595=>"000000000",
  30596=>"111111000",
  30597=>"000100110",
  30598=>"000000000",
  30599=>"000000000",
  30600=>"001001001",
  30601=>"111111111",
  30602=>"011111111",
  30603=>"101100111",
  30604=>"111111111",
  30605=>"100000000",
  30606=>"000000000",
  30607=>"000101000",
  30608=>"001011000",
  30609=>"000111111",
  30610=>"111111111",
  30611=>"000000100",
  30612=>"111111101",
  30613=>"000000000",
  30614=>"001000000",
  30615=>"001111001",
  30616=>"000010111",
  30617=>"111111100",
  30618=>"001000010",
  30619=>"000000000",
  30620=>"000001111",
  30621=>"111011011",
  30622=>"101001000",
  30623=>"000000000",
  30624=>"010110011",
  30625=>"111111011",
  30626=>"111111011",
  30627=>"111101100",
  30628=>"000000010",
  30629=>"010110010",
  30630=>"111111111",
  30631=>"110010000",
  30632=>"000000000",
  30633=>"001010000",
  30634=>"100100000",
  30635=>"111110110",
  30636=>"000000000",
  30637=>"111000100",
  30638=>"000011111",
  30639=>"000000001",
  30640=>"111111111",
  30641=>"000000001",
  30642=>"000000000",
  30643=>"111111111",
  30644=>"000000001",
  30645=>"101101100",
  30646=>"000000000",
  30647=>"000000000",
  30648=>"111111111",
  30649=>"010000010",
  30650=>"000110000",
  30651=>"100000000",
  30652=>"100100000",
  30653=>"000000001",
  30654=>"111111111",
  30655=>"010000011",
  30656=>"010000000",
  30657=>"111111111",
  30658=>"001001000",
  30659=>"000110011",
  30660=>"000000000",
  30661=>"101000000",
  30662=>"000000000",
  30663=>"111100000",
  30664=>"000000000",
  30665=>"111100100",
  30666=>"111111111",
  30667=>"100111011",
  30668=>"111010010",
  30669=>"011111110",
  30670=>"000010000",
  30671=>"110000110",
  30672=>"111000000",
  30673=>"111111111",
  30674=>"110111110",
  30675=>"111111111",
  30676=>"001001001",
  30677=>"000000110",
  30678=>"110111011",
  30679=>"100110111",
  30680=>"000000101",
  30681=>"110111111",
  30682=>"000000000",
  30683=>"001111000",
  30684=>"111111111",
  30685=>"101000000",
  30686=>"111111000",
  30687=>"000001001",
  30688=>"101000000",
  30689=>"000111111",
  30690=>"111000000",
  30691=>"111000000",
  30692=>"000000000",
  30693=>"100000111",
  30694=>"111000000",
  30695=>"111111111",
  30696=>"010110010",
  30697=>"000000000",
  30698=>"000000111",
  30699=>"001000111",
  30700=>"111111000",
  30701=>"100111110",
  30702=>"110000100",
  30703=>"111111111",
  30704=>"001000000",
  30705=>"110111111",
  30706=>"010110111",
  30707=>"000110000",
  30708=>"000000000",
  30709=>"000100000",
  30710=>"010111110",
  30711=>"000110110",
  30712=>"110100000",
  30713=>"111111100",
  30714=>"111000000",
  30715=>"000000000",
  30716=>"111111001",
  30717=>"110110110",
  30718=>"110110000",
  30719=>"001111111",
  30720=>"001000111",
  30721=>"100100101",
  30722=>"111000000",
  30723=>"000111111",
  30724=>"011011111",
  30725=>"011000000",
  30726=>"000000000",
  30727=>"111000000",
  30728=>"110110100",
  30729=>"111111100",
  30730=>"000000111",
  30731=>"100101000",
  30732=>"000110000",
  30733=>"100111011",
  30734=>"001000011",
  30735=>"010111111",
  30736=>"110111101",
  30737=>"100100100",
  30738=>"000000111",
  30739=>"101100111",
  30740=>"000000000",
  30741=>"111111001",
  30742=>"000110100",
  30743=>"111000000",
  30744=>"111111110",
  30745=>"000000000",
  30746=>"000000111",
  30747=>"110000000",
  30748=>"000001000",
  30749=>"101000000",
  30750=>"110110110",
  30751=>"000000001",
  30752=>"000000100",
  30753=>"000000100",
  30754=>"001111111",
  30755=>"111111100",
  30756=>"000000000",
  30757=>"110111111",
  30758=>"000000101",
  30759=>"001111101",
  30760=>"000111111",
  30761=>"000111100",
  30762=>"000000000",
  30763=>"111011000",
  30764=>"110000000",
  30765=>"111111000",
  30766=>"000000100",
  30767=>"111111111",
  30768=>"000000000",
  30769=>"000000000",
  30770=>"111101000",
  30771=>"000000000",
  30772=>"011111001",
  30773=>"000000110",
  30774=>"111111111",
  30775=>"101001000",
  30776=>"111111111",
  30777=>"000000000",
  30778=>"000100000",
  30779=>"111111000",
  30780=>"111111111",
  30781=>"000000111",
  30782=>"111111000",
  30783=>"110111111",
  30784=>"011011000",
  30785=>"001001000",
  30786=>"000101111",
  30787=>"110100000",
  30788=>"110011010",
  30789=>"110110111",
  30790=>"111111000",
  30791=>"000111111",
  30792=>"000010000",
  30793=>"000101101",
  30794=>"111111110",
  30795=>"001111110",
  30796=>"000000101",
  30797=>"110000000",
  30798=>"100000000",
  30799=>"000000001",
  30800=>"100000110",
  30801=>"111111111",
  30802=>"000000000",
  30803=>"111110100",
  30804=>"111101000",
  30805=>"100100110",
  30806=>"110111111",
  30807=>"000000000",
  30808=>"011111110",
  30809=>"111111101",
  30810=>"000000000",
  30811=>"011001001",
  30812=>"111111000",
  30813=>"110000000",
  30814=>"010011110",
  30815=>"111111000",
  30816=>"011000001",
  30817=>"000000000",
  30818=>"010111111",
  30819=>"000000000",
  30820=>"111110110",
  30821=>"111111111",
  30822=>"000000000",
  30823=>"000111111",
  30824=>"111111000",
  30825=>"001000000",
  30826=>"100001111",
  30827=>"000000000",
  30828=>"001001011",
  30829=>"000110110",
  30830=>"010000000",
  30831=>"000100000",
  30832=>"110110110",
  30833=>"100001001",
  30834=>"011001001",
  30835=>"000000100",
  30836=>"101111001",
  30837=>"000111100",
  30838=>"111000000",
  30839=>"000110010",
  30840=>"111111111",
  30841=>"100100000",
  30842=>"111111100",
  30843=>"100000000",
  30844=>"000000100",
  30845=>"111100100",
  30846=>"100110100",
  30847=>"111000000",
  30848=>"010000000",
  30849=>"111111110",
  30850=>"111111110",
  30851=>"111001000",
  30852=>"111111111",
  30853=>"011000000",
  30854=>"011011000",
  30855=>"001010000",
  30856=>"000111111",
  30857=>"111111111",
  30858=>"000000000",
  30859=>"111111111",
  30860=>"110101111",
  30861=>"000000000",
  30862=>"000100000",
  30863=>"001011001",
  30864=>"101101111",
  30865=>"001000001",
  30866=>"111111000",
  30867=>"011000000",
  30868=>"001111011",
  30869=>"001000000",
  30870=>"111111000",
  30871=>"111000001",
  30872=>"101100100",
  30873=>"000111111",
  30874=>"000000000",
  30875=>"111000000",
  30876=>"111111110",
  30877=>"000000111",
  30878=>"011111111",
  30879=>"011011011",
  30880=>"110110000",
  30881=>"000011111",
  30882=>"000011111",
  30883=>"010000000",
  30884=>"000110000",
  30885=>"000111111",
  30886=>"000000001",
  30887=>"001001000",
  30888=>"000000011",
  30889=>"011000001",
  30890=>"000000000",
  30891=>"111000111",
  30892=>"110000000",
  30893=>"011010000",
  30894=>"001000000",
  30895=>"000000000",
  30896=>"000000000",
  30897=>"000001000",
  30898=>"111111111",
  30899=>"000000011",
  30900=>"000110110",
  30901=>"100000000",
  30902=>"000000000",
  30903=>"111111111",
  30904=>"000111111",
  30905=>"111101111",
  30906=>"000000010",
  30907=>"000110000",
  30908=>"110110000",
  30909=>"000000110",
  30910=>"111110000",
  30911=>"111000000",
  30912=>"111001000",
  30913=>"111000000",
  30914=>"000000000",
  30915=>"011111111",
  30916=>"000000111",
  30917=>"001000000",
  30918=>"000110110",
  30919=>"111100001",
  30920=>"010110110",
  30921=>"111000100",
  30922=>"011000100",
  30923=>"011010110",
  30924=>"000111011",
  30925=>"111111000",
  30926=>"111110000",
  30927=>"111111111",
  30928=>"101111000",
  30929=>"111000000",
  30930=>"111111000",
  30931=>"000010010",
  30932=>"000011111",
  30933=>"010000100",
  30934=>"100111111",
  30935=>"111001001",
  30936=>"000000000",
  30937=>"111110100",
  30938=>"000111111",
  30939=>"000000001",
  30940=>"001011001",
  30941=>"000000001",
  30942=>"010111111",
  30943=>"111111000",
  30944=>"000000000",
  30945=>"000000111",
  30946=>"111111110",
  30947=>"110000000",
  30948=>"010100110",
  30949=>"110110110",
  30950=>"000000010",
  30951=>"000000000",
  30952=>"111000000",
  30953=>"100111111",
  30954=>"011001011",
  30955=>"100100111",
  30956=>"001000000",
  30957=>"000000111",
  30958=>"000100000",
  30959=>"000000000",
  30960=>"111000001",
  30961=>"000001100",
  30962=>"111000111",
  30963=>"100000000",
  30964=>"111111110",
  30965=>"101011111",
  30966=>"001000001",
  30967=>"010001111",
  30968=>"000000011",
  30969=>"101000000",
  30970=>"000000111",
  30971=>"001101111",
  30972=>"011111111",
  30973=>"000000000",
  30974=>"000111111",
  30975=>"111111000",
  30976=>"001000000",
  30977=>"000000010",
  30978=>"000100000",
  30979=>"111111111",
  30980=>"000111111",
  30981=>"100100111",
  30982=>"111111111",
  30983=>"110111011",
  30984=>"111111111",
  30985=>"011001111",
  30986=>"110000000",
  30987=>"000000111",
  30988=>"111001111",
  30989=>"110110100",
  30990=>"000000000",
  30991=>"111111000",
  30992=>"000110110",
  30993=>"000000110",
  30994=>"110110000",
  30995=>"000100000",
  30996=>"000000000",
  30997=>"000100100",
  30998=>"000100000",
  30999=>"111001011",
  31000=>"000010111",
  31001=>"111111111",
  31002=>"001111110",
  31003=>"111111100",
  31004=>"010110100",
  31005=>"001000000",
  31006=>"100100000",
  31007=>"111111101",
  31008=>"100000000",
  31009=>"111111111",
  31010=>"111111000",
  31011=>"011011011",
  31012=>"111111110",
  31013=>"001000000",
  31014=>"011111111",
  31015=>"111000010",
  31016=>"000000000",
  31017=>"011111111",
  31018=>"000000111",
  31019=>"111000000",
  31020=>"111111110",
  31021=>"111110110",
  31022=>"000111000",
  31023=>"000110111",
  31024=>"001111110",
  31025=>"111110000",
  31026=>"100111001",
  31027=>"110000110",
  31028=>"000000000",
  31029=>"011111001",
  31030=>"000111001",
  31031=>"000100101",
  31032=>"011000000",
  31033=>"100111111",
  31034=>"000000110",
  31035=>"000000000",
  31036=>"110110110",
  31037=>"000000000",
  31038=>"000011111",
  31039=>"110110111",
  31040=>"110111100",
  31041=>"011111110",
  31042=>"111010000",
  31043=>"111001000",
  31044=>"000000000",
  31045=>"111111001",
  31046=>"111111110",
  31047=>"000000000",
  31048=>"000001100",
  31049=>"110000000",
  31050=>"111011111",
  31051=>"111011001",
  31052=>"000000000",
  31053=>"111111111",
  31054=>"110000100",
  31055=>"001111111",
  31056=>"111100000",
  31057=>"000111111",
  31058=>"111111111",
  31059=>"000000000",
  31060=>"000000111",
  31061=>"000000001",
  31062=>"010000000",
  31063=>"010111011",
  31064=>"101111111",
  31065=>"111111000",
  31066=>"001000001",
  31067=>"000000000",
  31068=>"111111111",
  31069=>"000000000",
  31070=>"001000000",
  31071=>"111111111",
  31072=>"000000000",
  31073=>"000111100",
  31074=>"000101000",
  31075=>"000000111",
  31076=>"000000111",
  31077=>"011011000",
  31078=>"000000110",
  31079=>"001111111",
  31080=>"011001000",
  31081=>"111000000",
  31082=>"000000000",
  31083=>"110011000",
  31084=>"111111000",
  31085=>"111110110",
  31086=>"000111110",
  31087=>"000011000",
  31088=>"111111010",
  31089=>"010000000",
  31090=>"011111000",
  31091=>"001001011",
  31092=>"111111100",
  31093=>"000111111",
  31094=>"010010000",
  31095=>"100111110",
  31096=>"000000000",
  31097=>"111111111",
  31098=>"000000111",
  31099=>"111111000",
  31100=>"111111111",
  31101=>"101111111",
  31102=>"000100100",
  31103=>"111100100",
  31104=>"000110000",
  31105=>"100100111",
  31106=>"000000111",
  31107=>"100100110",
  31108=>"110111111",
  31109=>"000000000",
  31110=>"000011011",
  31111=>"111111001",
  31112=>"011000000",
  31113=>"101111111",
  31114=>"111111111",
  31115=>"000001111",
  31116=>"111000011",
  31117=>"000011011",
  31118=>"100000000",
  31119=>"111000000",
  31120=>"111000110",
  31121=>"100000011",
  31122=>"111100000",
  31123=>"000001001",
  31124=>"111011011",
  31125=>"000010000",
  31126=>"101111111",
  31127=>"000111110",
  31128=>"011011111",
  31129=>"111000000",
  31130=>"111000000",
  31131=>"111000000",
  31132=>"111110111",
  31133=>"111111000",
  31134=>"110110111",
  31135=>"111111111",
  31136=>"110000000",
  31137=>"111111001",
  31138=>"111110000",
  31139=>"000110110",
  31140=>"111111000",
  31141=>"111100000",
  31142=>"111111001",
  31143=>"011000000",
  31144=>"111000001",
  31145=>"111101111",
  31146=>"111111010",
  31147=>"000110111",
  31148=>"111111000",
  31149=>"100001011",
  31150=>"000000100",
  31151=>"110000110",
  31152=>"111011000",
  31153=>"011010000",
  31154=>"000000000",
  31155=>"111111100",
  31156=>"000110110",
  31157=>"100111111",
  31158=>"011111111",
  31159=>"111000000",
  31160=>"000000000",
  31161=>"111111110",
  31162=>"111111110",
  31163=>"111111000",
  31164=>"001000011",
  31165=>"000000000",
  31166=>"111001011",
  31167=>"000000000",
  31168=>"000000000",
  31169=>"011100000",
  31170=>"000000000",
  31171=>"110100010",
  31172=>"000000011",
  31173=>"000100100",
  31174=>"001101111",
  31175=>"111111001",
  31176=>"000000000",
  31177=>"111011011",
  31178=>"100000000",
  31179=>"000000000",
  31180=>"001000000",
  31181=>"000000000",
  31182=>"001001000",
  31183=>"000111111",
  31184=>"000001111",
  31185=>"001111111",
  31186=>"000111110",
  31187=>"001001111",
  31188=>"001111111",
  31189=>"110111010",
  31190=>"000110111",
  31191=>"111011011",
  31192=>"000011110",
  31193=>"100100110",
  31194=>"000100111",
  31195=>"000001000",
  31196=>"110111000",
  31197=>"000000000",
  31198=>"111111011",
  31199=>"000000011",
  31200=>"000000000",
  31201=>"111000000",
  31202=>"000000000",
  31203=>"011111111",
  31204=>"001111000",
  31205=>"111111111",
  31206=>"010100110",
  31207=>"000110110",
  31208=>"001100111",
  31209=>"111111111",
  31210=>"110111111",
  31211=>"111010000",
  31212=>"100000000",
  31213=>"111111111",
  31214=>"111111111",
  31215=>"000000000",
  31216=>"111011111",
  31217=>"011000111",
  31218=>"000000001",
  31219=>"011001000",
  31220=>"000010111",
  31221=>"111000000",
  31222=>"000000000",
  31223=>"100110000",
  31224=>"111111001",
  31225=>"111001001",
  31226=>"111011000",
  31227=>"111111111",
  31228=>"000010010",
  31229=>"111111111",
  31230=>"000000110",
  31231=>"111001000",
  31232=>"000000000",
  31233=>"000111110",
  31234=>"000100111",
  31235=>"111111010",
  31236=>"111001011",
  31237=>"111100100",
  31238=>"101000101",
  31239=>"111001000",
  31240=>"000111111",
  31241=>"110000000",
  31242=>"110111111",
  31243=>"000000000",
  31244=>"001001001",
  31245=>"111111111",
  31246=>"000100110",
  31247=>"000000000",
  31248=>"001000000",
  31249=>"111111000",
  31250=>"111110011",
  31251=>"111111111",
  31252=>"000001110",
  31253=>"010111111",
  31254=>"110111111",
  31255=>"000001011",
  31256=>"000000000",
  31257=>"000000000",
  31258=>"000011011",
  31259=>"000000110",
  31260=>"000000000",
  31261=>"000000000",
  31262=>"110001100",
  31263=>"100111001",
  31264=>"111111000",
  31265=>"101101101",
  31266=>"000000000",
  31267=>"010010011",
  31268=>"111111111",
  31269=>"000000000",
  31270=>"000111000",
  31271=>"111111110",
  31272=>"110010000",
  31273=>"000000111",
  31274=>"111000101",
  31275=>"001001000",
  31276=>"000111111",
  31277=>"111000000",
  31278=>"111011010",
  31279=>"110110111",
  31280=>"000111000",
  31281=>"111110000",
  31282=>"111111111",
  31283=>"010010011",
  31284=>"000010010",
  31285=>"101101001",
  31286=>"000110111",
  31287=>"011000000",
  31288=>"111111111",
  31289=>"000001001",
  31290=>"000000001",
  31291=>"000000110",
  31292=>"000000000",
  31293=>"000000001",
  31294=>"001000000",
  31295=>"111111111",
  31296=>"111111011",
  31297=>"000011011",
  31298=>"000000000",
  31299=>"000101101",
  31300=>"111111111",
  31301=>"011111011",
  31302=>"011011111",
  31303=>"001101000",
  31304=>"010111000",
  31305=>"001001111",
  31306=>"110000000",
  31307=>"111000100",
  31308=>"000000000",
  31309=>"100000000",
  31310=>"100111110",
  31311=>"111111111",
  31312=>"111111001",
  31313=>"100100000",
  31314=>"111111111",
  31315=>"000000000",
  31316=>"111111000",
  31317=>"000000010",
  31318=>"000011111",
  31319=>"000000000",
  31320=>"000000000",
  31321=>"000000101",
  31322=>"100111111",
  31323=>"000000000",
  31324=>"000000000",
  31325=>"110111000",
  31326=>"111111100",
  31327=>"111111100",
  31328=>"010000000",
  31329=>"000111111",
  31330=>"011011011",
  31331=>"000000000",
  31332=>"000000101",
  31333=>"111111000",
  31334=>"111011011",
  31335=>"111000000",
  31336=>"001101101",
  31337=>"011111111",
  31338=>"100100000",
  31339=>"110111111",
  31340=>"000100100",
  31341=>"111111100",
  31342=>"000000000",
  31343=>"111101111",
  31344=>"000000111",
  31345=>"111111001",
  31346=>"001000011",
  31347=>"001001011",
  31348=>"000000010",
  31349=>"111111111",
  31350=>"111111111",
  31351=>"000000000",
  31352=>"000000000",
  31353=>"111000001",
  31354=>"000000000",
  31355=>"100000101",
  31356=>"000000100",
  31357=>"101000111",
  31358=>"000000000",
  31359=>"111111111",
  31360=>"001000101",
  31361=>"111111101",
  31362=>"111000000",
  31363=>"011011000",
  31364=>"111111111",
  31365=>"111010100",
  31366=>"111111110",
  31367=>"000010000",
  31368=>"011001000",
  31369=>"100010111",
  31370=>"111111111",
  31371=>"110110000",
  31372=>"111111110",
  31373=>"111111100",
  31374=>"100000000",
  31375=>"111000000",
  31376=>"000111111",
  31377=>"000000000",
  31378=>"000000010",
  31379=>"011011001",
  31380=>"000000111",
  31381=>"000111111",
  31382=>"111111111",
  31383=>"000011111",
  31384=>"000000110",
  31385=>"000000000",
  31386=>"111001000",
  31387=>"111111010",
  31388=>"111111101",
  31389=>"111100000",
  31390=>"010111011",
  31391=>"000000000",
  31392=>"000001111",
  31393=>"111111110",
  31394=>"010110010",
  31395=>"000100100",
  31396=>"110111011",
  31397=>"000010111",
  31398=>"111111111",
  31399=>"110100000",
  31400=>"000000000",
  31401=>"111110111",
  31402=>"111111001",
  31403=>"011011000",
  31404=>"000000000",
  31405=>"110110111",
  31406=>"110111000",
  31407=>"011111110",
  31408=>"000110111",
  31409=>"011001001",
  31410=>"111111111",
  31411=>"111111111",
  31412=>"111011011",
  31413=>"110000000",
  31414=>"000000110",
  31415=>"111111101",
  31416=>"001000100",
  31417=>"100000111",
  31418=>"101001001",
  31419=>"100000000",
  31420=>"001000000",
  31421=>"101101111",
  31422=>"111001101",
  31423=>"100000000",
  31424=>"000000000",
  31425=>"111111111",
  31426=>"000001111",
  31427=>"000000111",
  31428=>"000000000",
  31429=>"000001000",
  31430=>"000000000",
  31431=>"001111111",
  31432=>"100100000",
  31433=>"011111111",
  31434=>"110000000",
  31435=>"010000000",
  31436=>"000000000",
  31437=>"110010000",
  31438=>"110111110",
  31439=>"011001000",
  31440=>"111111111",
  31441=>"000000000",
  31442=>"000000000",
  31443=>"000000111",
  31444=>"111111010",
  31445=>"110111000",
  31446=>"000000000",
  31447=>"000000100",
  31448=>"111110011",
  31449=>"000000000",
  31450=>"110100100",
  31451=>"000000101",
  31452=>"000000000",
  31453=>"000110110",
  31454=>"000000000",
  31455=>"001000000",
  31456=>"000000000",
  31457=>"000000111",
  31458=>"000000000",
  31459=>"111111111",
  31460=>"101100111",
  31461=>"110110110",
  31462=>"101111111",
  31463=>"111100000",
  31464=>"000000000",
  31465=>"000000000",
  31466=>"110110110",
  31467=>"111111111",
  31468=>"000000000",
  31469=>"000000000",
  31470=>"111011001",
  31471=>"000000000",
  31472=>"011000011",
  31473=>"000000000",
  31474=>"111111001",
  31475=>"001011011",
  31476=>"101000000",
  31477=>"111011000",
  31478=>"110111111",
  31479=>"111111111",
  31480=>"111111100",
  31481=>"000000100",
  31482=>"010111111",
  31483=>"011111011",
  31484=>"111000000",
  31485=>"110000000",
  31486=>"000001000",
  31487=>"101111111",
  31488=>"111111111",
  31489=>"000001111",
  31490=>"000000000",
  31491=>"100000000",
  31492=>"111101000",
  31493=>"000110111",
  31494=>"100111111",
  31495=>"000110100",
  31496=>"000000000",
  31497=>"000000111",
  31498=>"001100100",
  31499=>"000000100",
  31500=>"110110000",
  31501=>"111100011",
  31502=>"000000001",
  31503=>"111111001",
  31504=>"010110111",
  31505=>"111111111",
  31506=>"000000000",
  31507=>"111100011",
  31508=>"111010000",
  31509=>"111100000",
  31510=>"111111111",
  31511=>"000000000",
  31512=>"000000000",
  31513=>"111111000",
  31514=>"000000000",
  31515=>"110000000",
  31516=>"110111000",
  31517=>"000000000",
  31518=>"111111110",
  31519=>"000110110",
  31520=>"111111110",
  31521=>"111111111",
  31522=>"100100111",
  31523=>"000110100",
  31524=>"000000000",
  31525=>"001111111",
  31526=>"100000000",
  31527=>"001010111",
  31528=>"100100111",
  31529=>"111111110",
  31530=>"100110110",
  31531=>"000000001",
  31532=>"110110000",
  31533=>"000010010",
  31534=>"111111100",
  31535=>"000000000",
  31536=>"000000100",
  31537=>"111111100",
  31538=>"100110110",
  31539=>"000000000",
  31540=>"010000000",
  31541=>"001000101",
  31542=>"000000000",
  31543=>"001001100",
  31544=>"010000000",
  31545=>"000000000",
  31546=>"000000111",
  31547=>"111000000",
  31548=>"110111111",
  31549=>"000000000",
  31550=>"000000000",
  31551=>"001001000",
  31552=>"110000000",
  31553=>"001001111",
  31554=>"000000000",
  31555=>"001001000",
  31556=>"000001111",
  31557=>"111101111",
  31558=>"100111111",
  31559=>"111010110",
  31560=>"110100100",
  31561=>"010011001",
  31562=>"111111110",
  31563=>"001000000",
  31564=>"110111111",
  31565=>"111110000",
  31566=>"000111111",
  31567=>"100110110",
  31568=>"000000000",
  31569=>"001111111",
  31570=>"111110110",
  31571=>"001011111",
  31572=>"000000000",
  31573=>"111011001",
  31574=>"111111110",
  31575=>"000000000",
  31576=>"100101111",
  31577=>"110110111",
  31578=>"111110000",
  31579=>"111111100",
  31580=>"110100000",
  31581=>"100000000",
  31582=>"000000111",
  31583=>"111110110",
  31584=>"000100111",
  31585=>"111100000",
  31586=>"110110111",
  31587=>"111111101",
  31588=>"111111111",
  31589=>"000000000",
  31590=>"110110110",
  31591=>"100010010",
  31592=>"111000000",
  31593=>"111100111",
  31594=>"100111110",
  31595=>"101110110",
  31596=>"001100100",
  31597=>"101111011",
  31598=>"011111111",
  31599=>"000000000",
  31600=>"000000000",
  31601=>"000000000",
  31602=>"010000101",
  31603=>"000000000",
  31604=>"011011001",
  31605=>"111101100",
  31606=>"100000100",
  31607=>"100110000",
  31608=>"111111000",
  31609=>"111111111",
  31610=>"000100101",
  31611=>"111000000",
  31612=>"000000001",
  31613=>"111111110",
  31614=>"111111111",
  31615=>"000000111",
  31616=>"001000000",
  31617=>"011011000",
  31618=>"001110111",
  31619=>"000000001",
  31620=>"111111000",
  31621=>"000000001",
  31622=>"000100111",
  31623=>"000000010",
  31624=>"001000000",
  31625=>"000000101",
  31626=>"000000000",
  31627=>"000000000",
  31628=>"111111111",
  31629=>"101111000",
  31630=>"100000000",
  31631=>"100100110",
  31632=>"111111110",
  31633=>"000000000",
  31634=>"111111111",
  31635=>"001111111",
  31636=>"111100000",
  31637=>"110000000",
  31638=>"111000000",
  31639=>"111101111",
  31640=>"001001000",
  31641=>"111001011",
  31642=>"000011111",
  31643=>"000000000",
  31644=>"000100111",
  31645=>"110110000",
  31646=>"111100000",
  31647=>"000000100",
  31648=>"111001000",
  31649=>"111110110",
  31650=>"000010100",
  31651=>"000000001",
  31652=>"011010000",
  31653=>"000000000",
  31654=>"000000100",
  31655=>"110000000",
  31656=>"000000000",
  31657=>"000000000",
  31658=>"101000000",
  31659=>"111000010",
  31660=>"010000110",
  31661=>"000000000",
  31662=>"000000000",
  31663=>"101111111",
  31664=>"100111000",
  31665=>"001111010",
  31666=>"110000000",
  31667=>"001111111",
  31668=>"000001111",
  31669=>"111000000",
  31670=>"111111111",
  31671=>"000000000",
  31672=>"111000100",
  31673=>"000100000",
  31674=>"011001001",
  31675=>"100100111",
  31676=>"111111000",
  31677=>"000001011",
  31678=>"111101111",
  31679=>"101111111",
  31680=>"111111000",
  31681=>"000000000",
  31682=>"111000111",
  31683=>"000111111",
  31684=>"000000000",
  31685=>"000000100",
  31686=>"001001100",
  31687=>"000100111",
  31688=>"000000000",
  31689=>"111101100",
  31690=>"000000000",
  31691=>"111111111",
  31692=>"111000000",
  31693=>"100110100",
  31694=>"000000000",
  31695=>"000000101",
  31696=>"000100100",
  31697=>"001110000",
  31698=>"000000111",
  31699=>"000000000",
  31700=>"000100110",
  31701=>"111111000",
  31702=>"100110100",
  31703=>"100000000",
  31704=>"110110111",
  31705=>"111111110",
  31706=>"111111111",
  31707=>"011001101",
  31708=>"000000000",
  31709=>"000000000",
  31710=>"011000000",
  31711=>"011111011",
  31712=>"110111111",
  31713=>"001001001",
  31714=>"011011011",
  31715=>"101101000",
  31716=>"100100110",
  31717=>"101101000",
  31718=>"000000000",
  31719=>"000000000",
  31720=>"000000000",
  31721=>"000000000",
  31722=>"000110110",
  31723=>"000000000",
  31724=>"000000000",
  31725=>"010001011",
  31726=>"111111111",
  31727=>"100000000",
  31728=>"101000000",
  31729=>"001000000",
  31730=>"000000000",
  31731=>"001001001",
  31732=>"000000000",
  31733=>"000000000",
  31734=>"000001001",
  31735=>"000000111",
  31736=>"000111000",
  31737=>"000100000",
  31738=>"101001111",
  31739=>"000000111",
  31740=>"111110000",
  31741=>"111111000",
  31742=>"111100110",
  31743=>"111101111",
  31744=>"111111111",
  31745=>"111111111",
  31746=>"000111000",
  31747=>"000000000",
  31748=>"111111111",
  31749=>"000010001",
  31750=>"000100000",
  31751=>"111000000",
  31752=>"111111111",
  31753=>"000000000",
  31754=>"000000111",
  31755=>"111111101",
  31756=>"001001111",
  31757=>"111111111",
  31758=>"000000100",
  31759=>"000000000",
  31760=>"101111111",
  31761=>"111100000",
  31762=>"000000000",
  31763=>"111000000",
  31764=>"000100000",
  31765=>"111111111",
  31766=>"001000111",
  31767=>"011011010",
  31768=>"100000000",
  31769=>"110000000",
  31770=>"000000000",
  31771=>"100000000",
  31772=>"000000001",
  31773=>"111111111",
  31774=>"010010011",
  31775=>"000000001",
  31776=>"011111110",
  31777=>"000001000",
  31778=>"100100010",
  31779=>"000000000",
  31780=>"111000100",
  31781=>"000000000",
  31782=>"000000000",
  31783=>"000111000",
  31784=>"111100100",
  31785=>"111000000",
  31786=>"000000000",
  31787=>"011011000",
  31788=>"000001000",
  31789=>"110110100",
  31790=>"000000000",
  31791=>"000000000",
  31792=>"001011111",
  31793=>"000000001",
  31794=>"001001000",
  31795=>"111110000",
  31796=>"011010000",
  31797=>"001000001",
  31798=>"001111100",
  31799=>"111111110",
  31800=>"111111111",
  31801=>"000001111",
  31802=>"000000000",
  31803=>"000000111",
  31804=>"000001111",
  31805=>"111111110",
  31806=>"011000000",
  31807=>"000000000",
  31808=>"100000001",
  31809=>"000111111",
  31810=>"100000000",
  31811=>"000111000",
  31812=>"111111111",
  31813=>"100011001",
  31814=>"000110111",
  31815=>"111111111",
  31816=>"001011111",
  31817=>"000000001",
  31818=>"001001000",
  31819=>"111111101",
  31820=>"100111111",
  31821=>"101101100",
  31822=>"011011011",
  31823=>"001000000",
  31824=>"110110000",
  31825=>"001111111",
  31826=>"000000100",
  31827=>"110111111",
  31828=>"000000001",
  31829=>"011011111",
  31830=>"000000111",
  31831=>"000000000",
  31832=>"000000000",
  31833=>"000000000",
  31834=>"000001000",
  31835=>"100101101",
  31836=>"111111111",
  31837=>"100000111",
  31838=>"000000000",
  31839=>"000000000",
  31840=>"100000000",
  31841=>"001000000",
  31842=>"011111111",
  31843=>"111111111",
  31844=>"100000000",
  31845=>"110111111",
  31846=>"111111111",
  31847=>"011001000",
  31848=>"000000011",
  31849=>"111010000",
  31850=>"000111111",
  31851=>"000001000",
  31852=>"111111111",
  31853=>"000000000",
  31854=>"000000000",
  31855=>"111111101",
  31856=>"001001111",
  31857=>"000111111",
  31858=>"011011001",
  31859=>"110111111",
  31860=>"000000000",
  31861=>"111111111",
  31862=>"111111111",
  31863=>"000000110",
  31864=>"000010111",
  31865=>"000111111",
  31866=>"101001001",
  31867=>"100110111",
  31868=>"001110100",
  31869=>"111111111",
  31870=>"000000000",
  31871=>"000000001",
  31872=>"000000000",
  31873=>"111111111",
  31874=>"001000000",
  31875=>"110111111",
  31876=>"000000000",
  31877=>"001001000",
  31878=>"110100111",
  31879=>"111111100",
  31880=>"111100000",
  31881=>"000111110",
  31882=>"100100110",
  31883=>"111000000",
  31884=>"111110110",
  31885=>"000000000",
  31886=>"000000001",
  31887=>"010111001",
  31888=>"111011010",
  31889=>"111111111",
  31890=>"011111111",
  31891=>"111100100",
  31892=>"001001001",
  31893=>"111111111",
  31894=>"000000000",
  31895=>"000000001",
  31896=>"000110110",
  31897=>"111111110",
  31898=>"000100000",
  31899=>"100000101",
  31900=>"000000010",
  31901=>"000010011",
  31902=>"110100000",
  31903=>"111100000",
  31904=>"000000000",
  31905=>"000000000",
  31906=>"000000001",
  31907=>"111100000",
  31908=>"001001000",
  31909=>"111111100",
  31910=>"111111111",
  31911=>"110100100",
  31912=>"000111101",
  31913=>"000000000",
  31914=>"001001001",
  31915=>"001001101",
  31916=>"101111001",
  31917=>"001001001",
  31918=>"000111000",
  31919=>"110111000",
  31920=>"100111000",
  31921=>"000000100",
  31922=>"111111111",
  31923=>"110110111",
  31924=>"000000101",
  31925=>"000011111",
  31926=>"001000000",
  31927=>"111011000",
  31928=>"000000111",
  31929=>"000000000",
  31930=>"111001000",
  31931=>"010111111",
  31932=>"001010010",
  31933=>"111111111",
  31934=>"000000000",
  31935=>"111111111",
  31936=>"110111111",
  31937=>"001001000",
  31938=>"010111111",
  31939=>"111111111",
  31940=>"000000000",
  31941=>"111111111",
  31942=>"000000000",
  31943=>"000111100",
  31944=>"001001010",
  31945=>"000000000",
  31946=>"001000111",
  31947=>"111111111",
  31948=>"000100111",
  31949=>"100000000",
  31950=>"000101111",
  31951=>"111111111",
  31952=>"000000001",
  31953=>"000101010",
  31954=>"111011000",
  31955=>"000000000",
  31956=>"111010000",
  31957=>"000000000",
  31958=>"011011001",
  31959=>"100100100",
  31960=>"111100111",
  31961=>"111101001",
  31962=>"100000000",
  31963=>"100110110",
  31964=>"000000000",
  31965=>"000011001",
  31966=>"111101001",
  31967=>"111111110",
  31968=>"000000111",
  31969=>"011000111",
  31970=>"111111110",
  31971=>"011011111",
  31972=>"100100111",
  31973=>"000000000",
  31974=>"001000110",
  31975=>"011010000",
  31976=>"000000000",
  31977=>"110110000",
  31978=>"101100100",
  31979=>"001001001",
  31980=>"010000000",
  31981=>"111111011",
  31982=>"110110000",
  31983=>"000000011",
  31984=>"000000000",
  31985=>"000110110",
  31986=>"111111111",
  31987=>"001000110",
  31988=>"111111111",
  31989=>"000000001",
  31990=>"110100111",
  31991=>"101101111",
  31992=>"111111111",
  31993=>"111111111",
  31994=>"000110000",
  31995=>"000111111",
  31996=>"001001001",
  31997=>"000100000",
  31998=>"000000000",
  31999=>"110100100",
  32000=>"011000100",
  32001=>"011011000",
  32002=>"000000000",
  32003=>"001000001",
  32004=>"000001011",
  32005=>"000000000",
  32006=>"101111110",
  32007=>"000000000",
  32008=>"101000001",
  32009=>"001100100",
  32010=>"000011011",
  32011=>"111111111",
  32012=>"100101111",
  32013=>"011111111",
  32014=>"000100101",
  32015=>"101000110",
  32016=>"000110111",
  32017=>"010011011",
  32018=>"101000000",
  32019=>"100100000",
  32020=>"111111111",
  32021=>"000101100",
  32022=>"011011000",
  32023=>"111111111",
  32024=>"110110111",
  32025=>"011010010",
  32026=>"000000001",
  32027=>"111111111",
  32028=>"100000000",
  32029=>"111111111",
  32030=>"000000000",
  32031=>"111100111",
  32032=>"011000111",
  32033=>"111111111",
  32034=>"011111111",
  32035=>"111001001",
  32036=>"111111010",
  32037=>"111111110",
  32038=>"111111101",
  32039=>"111111011",
  32040=>"101000000",
  32041=>"000000000",
  32042=>"000000101",
  32043=>"000111011",
  32044=>"000000101",
  32045=>"110111111",
  32046=>"110111100",
  32047=>"110000000",
  32048=>"101101001",
  32049=>"000000000",
  32050=>"000000000",
  32051=>"011000000",
  32052=>"000000000",
  32053=>"111011010",
  32054=>"000000101",
  32055=>"111111111",
  32056=>"000000000",
  32057=>"000111111",
  32058=>"011001111",
  32059=>"000000110",
  32060=>"111111011",
  32061=>"100101101",
  32062=>"111111111",
  32063=>"111111111",
  32064=>"000010010",
  32065=>"100110000",
  32066=>"111111111",
  32067=>"000000000",
  32068=>"111111101",
  32069=>"001001100",
  32070=>"000000000",
  32071=>"000001000",
  32072=>"111001111",
  32073=>"111111010",
  32074=>"000000000",
  32075=>"000110100",
  32076=>"000011011",
  32077=>"001100110",
  32078=>"000000111",
  32079=>"000000001",
  32080=>"000100110",
  32081=>"001001000",
  32082=>"000000110",
  32083=>"000100110",
  32084=>"110000000",
  32085=>"000000000",
  32086=>"111110100",
  32087=>"000000000",
  32088=>"111111111",
  32089=>"011010000",
  32090=>"000010011",
  32091=>"000000000",
  32092=>"000000010",
  32093=>"001000000",
  32094=>"110110001",
  32095=>"111011011",
  32096=>"111111111",
  32097=>"111001001",
  32098=>"110110100",
  32099=>"000111111",
  32100=>"111111111",
  32101=>"111111111",
  32102=>"111111111",
  32103=>"000001001",
  32104=>"011011000",
  32105=>"111001001",
  32106=>"010110111",
  32107=>"001111111",
  32108=>"001000001",
  32109=>"111101010",
  32110=>"110111101",
  32111=>"010010010",
  32112=>"111111111",
  32113=>"000000110",
  32114=>"100000100",
  32115=>"110000000",
  32116=>"111000111",
  32117=>"000100111",
  32118=>"001001001",
  32119=>"000001001",
  32120=>"000000000",
  32121=>"000001001",
  32122=>"000000000",
  32123=>"001001001",
  32124=>"100100111",
  32125=>"111111110",
  32126=>"001001111",
  32127=>"100100000",
  32128=>"000000010",
  32129=>"000110110",
  32130=>"111111100",
  32131=>"000000100",
  32132=>"111100000",
  32133=>"000000001",
  32134=>"000000111",
  32135=>"010000000",
  32136=>"011001000",
  32137=>"000011111",
  32138=>"000000100",
  32139=>"110000000",
  32140=>"000001111",
  32141=>"010010111",
  32142=>"000001111",
  32143=>"011011000",
  32144=>"100000111",
  32145=>"000000000",
  32146=>"000000001",
  32147=>"111111110",
  32148=>"001000000",
  32149=>"000000000",
  32150=>"101111111",
  32151=>"001011111",
  32152=>"000000111",
  32153=>"000000000",
  32154=>"101101100",
  32155=>"000111001",
  32156=>"111110110",
  32157=>"111111111",
  32158=>"000000000",
  32159=>"111111111",
  32160=>"101101111",
  32161=>"011011011",
  32162=>"111111001",
  32163=>"011111111",
  32164=>"000001100",
  32165=>"111111100",
  32166=>"111111000",
  32167=>"000010111",
  32168=>"000000000",
  32169=>"000000000",
  32170=>"000000000",
  32171=>"000000000",
  32172=>"000000000",
  32173=>"000101111",
  32174=>"110010110",
  32175=>"111110110",
  32176=>"000000000",
  32177=>"000000000",
  32178=>"011001000",
  32179=>"111111111",
  32180=>"000010011",
  32181=>"111111000",
  32182=>"110110110",
  32183=>"000001000",
  32184=>"001000101",
  32185=>"000010000",
  32186=>"111001000",
  32187=>"000010000",
  32188=>"100111111",
  32189=>"111000000",
  32190=>"000000000",
  32191=>"011011011",
  32192=>"111110100",
  32193=>"110111111",
  32194=>"111111111",
  32195=>"000000000",
  32196=>"000001101",
  32197=>"000000001",
  32198=>"010011111",
  32199=>"000000000",
  32200=>"100100111",
  32201=>"000000111",
  32202=>"011111111",
  32203=>"111110111",
  32204=>"000000110",
  32205=>"111111111",
  32206=>"000000000",
  32207=>"001011100",
  32208=>"000000000",
  32209=>"100100100",
  32210=>"111111111",
  32211=>"100100100",
  32212=>"111111111",
  32213=>"111110110",
  32214=>"101100100",
  32215=>"100000001",
  32216=>"000000000",
  32217=>"000000000",
  32218=>"111011001",
  32219=>"011000000",
  32220=>"111001101",
  32221=>"111111011",
  32222=>"111110111",
  32223=>"011000100",
  32224=>"000000000",
  32225=>"111111001",
  32226=>"111111111",
  32227=>"111011000",
  32228=>"000000000",
  32229=>"011011111",
  32230=>"111111101",
  32231=>"010010010",
  32232=>"000000000",
  32233=>"111111111",
  32234=>"001001001",
  32235=>"111010111",
  32236=>"111111000",
  32237=>"110100100",
  32238=>"000010110",
  32239=>"110111100",
  32240=>"100000000",
  32241=>"111100000",
  32242=>"000000000",
  32243=>"000010010",
  32244=>"111110111",
  32245=>"110111111",
  32246=>"111111101",
  32247=>"111111111",
  32248=>"111111111",
  32249=>"110110000",
  32250=>"000000000",
  32251=>"010110000",
  32252=>"111111110",
  32253=>"000000110",
  32254=>"000011001",
  32255=>"000000000",
  32256=>"010110111",
  32257=>"000000010",
  32258=>"000000000",
  32259=>"000010000",
  32260=>"110110110",
  32261=>"110010000",
  32262=>"000111111",
  32263=>"100110100",
  32264=>"010011001",
  32265=>"001000000",
  32266=>"111110111",
  32267=>"111110110",
  32268=>"000000111",
  32269=>"000111111",
  32270=>"111101000",
  32271=>"000000000",
  32272=>"001000000",
  32273=>"111111011",
  32274=>"000000111",
  32275=>"110000000",
  32276=>"000000111",
  32277=>"111100110",
  32278=>"000111101",
  32279=>"011011101",
  32280=>"000000000",
  32281=>"000000000",
  32282=>"000000010",
  32283=>"111111000",
  32284=>"100000000",
  32285=>"010000000",
  32286=>"011011111",
  32287=>"000000000",
  32288=>"111111000",
  32289=>"000000001",
  32290=>"111111111",
  32291=>"111111111",
  32292=>"000101101",
  32293=>"110111111",
  32294=>"011011000",
  32295=>"111110110",
  32296=>"000000000",
  32297=>"000001111",
  32298=>"000000000",
  32299=>"000000000",
  32300=>"001000111",
  32301=>"111111011",
  32302=>"111010000",
  32303=>"001001111",
  32304=>"011000100",
  32305=>"000000100",
  32306=>"111111111",
  32307=>"000000000",
  32308=>"000000111",
  32309=>"110111100",
  32310=>"111111111",
  32311=>"000111110",
  32312=>"111111010",
  32313=>"100011111",
  32314=>"000000000",
  32315=>"000000010",
  32316=>"000001111",
  32317=>"111111111",
  32318=>"111111111",
  32319=>"111111111",
  32320=>"000000100",
  32321=>"111101100",
  32322=>"100000000",
  32323=>"000000111",
  32324=>"011111111",
  32325=>"000111111",
  32326=>"111000000",
  32327=>"111111001",
  32328=>"000011001",
  32329=>"000000111",
  32330=>"111111000",
  32331=>"111001100",
  32332=>"111111000",
  32333=>"000111111",
  32334=>"111011000",
  32335=>"111111000",
  32336=>"111111111",
  32337=>"111111000",
  32338=>"111111000",
  32339=>"000000001",
  32340=>"000000000",
  32341=>"000000100",
  32342=>"111111111",
  32343=>"110111000",
  32344=>"000000001",
  32345=>"111000000",
  32346=>"111111111",
  32347=>"001001000",
  32348=>"000000011",
  32349=>"001000000",
  32350=>"111011000",
  32351=>"111111111",
  32352=>"000000011",
  32353=>"111011000",
  32354=>"000000000",
  32355=>"000101111",
  32356=>"100100000",
  32357=>"011000000",
  32358=>"111000000",
  32359=>"010110111",
  32360=>"101111110",
  32361=>"111000100",
  32362=>"110000000",
  32363=>"110000000",
  32364=>"110111000",
  32365=>"000000000",
  32366=>"111011000",
  32367=>"111111111",
  32368=>"000000100",
  32369=>"011010000",
  32370=>"111101001",
  32371=>"000000111",
  32372=>"000000111",
  32373=>"000000001",
  32374=>"000000011",
  32375=>"000000100",
  32376=>"000000000",
  32377=>"000000111",
  32378=>"000000111",
  32379=>"011000000",
  32380=>"001011001",
  32381=>"111111110",
  32382=>"000000100",
  32383=>"111111000",
  32384=>"000111111",
  32385=>"111011011",
  32386=>"111000001",
  32387=>"000110111",
  32388=>"000001001",
  32389=>"000000111",
  32390=>"111000001",
  32391=>"111111000",
  32392=>"110011011",
  32393=>"100000100",
  32394=>"100111111",
  32395=>"000000010",
  32396=>"000000110",
  32397=>"111101000",
  32398=>"000001111",
  32399=>"010000000",
  32400=>"111111111",
  32401=>"000001011",
  32402=>"111110111",
  32403=>"000110010",
  32404=>"000111101",
  32405=>"000001111",
  32406=>"110110000",
  32407=>"111011000",
  32408=>"000000000",
  32409=>"000000111",
  32410=>"111111110",
  32411=>"111000000",
  32412=>"011011000",
  32413=>"000000101",
  32414=>"110010000",
  32415=>"111111111",
  32416=>"110111110",
  32417=>"000000000",
  32418=>"111010111",
  32419=>"000000000",
  32420=>"000110100",
  32421=>"111111100",
  32422=>"000011111",
  32423=>"101111111",
  32424=>"010011111",
  32425=>"000101111",
  32426=>"000000000",
  32427=>"000000000",
  32428=>"111111111",
  32429=>"011011000",
  32430=>"111111011",
  32431=>"000000000",
  32432=>"000000000",
  32433=>"111111000",
  32434=>"010111000",
  32435=>"000000000",
  32436=>"011111100",
  32437=>"101101111",
  32438=>"000000111",
  32439=>"101000000",
  32440=>"011000000",
  32441=>"111111111",
  32442=>"000000101",
  32443=>"000110111",
  32444=>"000000000",
  32445=>"000100110",
  32446=>"100111111",
  32447=>"111010000",
  32448=>"001001011",
  32449=>"011111110",
  32450=>"111100100",
  32451=>"111101100",
  32452=>"001001111",
  32453=>"010010111",
  32454=>"000000000",
  32455=>"111111000",
  32456=>"000000000",
  32457=>"110110000",
  32458=>"001000100",
  32459=>"000000111",
  32460=>"010011111",
  32461=>"111111000",
  32462=>"000000000",
  32463=>"000110111",
  32464=>"001000000",
  32465=>"000000100",
  32466=>"000100110",
  32467=>"000000111",
  32468=>"000000000",
  32469=>"100000000",
  32470=>"111111111",
  32471=>"000000100",
  32472=>"000000000",
  32473=>"111111100",
  32474=>"111000000",
  32475=>"000000001",
  32476=>"111111101",
  32477=>"100111111",
  32478=>"000000000",
  32479=>"000000001",
  32480=>"111111111",
  32481=>"111100000",
  32482=>"100101101",
  32483=>"000000000",
  32484=>"011111000",
  32485=>"000100100",
  32486=>"000111111",
  32487=>"000000100",
  32488=>"110111001",
  32489=>"001000000",
  32490=>"000000111",
  32491=>"001001011",
  32492=>"000000111",
  32493=>"000100111",
  32494=>"000110111",
  32495=>"000000100",
  32496=>"111000000",
  32497=>"100111111",
  32498=>"010111111",
  32499=>"000101100",
  32500=>"000110000",
  32501=>"101110111",
  32502=>"011001011",
  32503=>"111111111",
  32504=>"000000111",
  32505=>"011000000",
  32506=>"000000110",
  32507=>"111000000",
  32508=>"100111000",
  32509=>"111111001",
  32510=>"000000011",
  32511=>"011011111",
  32512=>"000000111",
  32513=>"011011011",
  32514=>"000001011",
  32515=>"000000000",
  32516=>"111111000",
  32517=>"111101001",
  32518=>"000000111",
  32519=>"001001111",
  32520=>"000010001",
  32521=>"000000000",
  32522=>"001001111",
  32523=>"111111100",
  32524=>"000000000",
  32525=>"111111000",
  32526=>"000011011",
  32527=>"100111111",
  32528=>"000000011",
  32529=>"000001111",
  32530=>"000000011",
  32531=>"111111001",
  32532=>"111111101",
  32533=>"111111011",
  32534=>"001001001",
  32535=>"111111111",
  32536=>"000111101",
  32537=>"100001000",
  32538=>"000000000",
  32539=>"111111111",
  32540=>"001111011",
  32541=>"001001000",
  32542=>"110110111",
  32543=>"000000000",
  32544=>"111011000",
  32545=>"011011000",
  32546=>"000110000",
  32547=>"000000101",
  32548=>"100000000",
  32549=>"000000111",
  32550=>"010111110",
  32551=>"011001001",
  32552=>"111111010",
  32553=>"111110000",
  32554=>"010111111",
  32555=>"111111100",
  32556=>"100100111",
  32557=>"000100100",
  32558=>"000000000",
  32559=>"000000000",
  32560=>"111111001",
  32561=>"111111111",
  32562=>"011011011",
  32563=>"000000110",
  32564=>"110000000",
  32565=>"110110111",
  32566=>"011000010",
  32567=>"000000000",
  32568=>"011111111",
  32569=>"001000111",
  32570=>"000000000",
  32571=>"100111111",
  32572=>"000011011",
  32573=>"000110111",
  32574=>"000000000",
  32575=>"000000111",
  32576=>"000000000",
  32577=>"000010000",
  32578=>"000111111",
  32579=>"000001000",
  32580=>"111000000",
  32581=>"111111111",
  32582=>"001011111",
  32583=>"000110010",
  32584=>"111000001",
  32585=>"111111010",
  32586=>"000000000",
  32587=>"100000000",
  32588=>"000000000",
  32589=>"000111111",
  32590=>"010000000",
  32591=>"100000000",
  32592=>"011110111",
  32593=>"010010011",
  32594=>"111000000",
  32595=>"000011111",
  32596=>"000011011",
  32597=>"111111111",
  32598=>"010110111",
  32599=>"100100111",
  32600=>"111111000",
  32601=>"000000000",
  32602=>"000001010",
  32603=>"000111110",
  32604=>"100000000",
  32605=>"000001011",
  32606=>"111110000",
  32607=>"000110111",
  32608=>"011001111",
  32609=>"101001111",
  32610=>"001111111",
  32611=>"000111000",
  32612=>"111111000",
  32613=>"011011000",
  32614=>"111001111",
  32615=>"000000000",
  32616=>"001000000",
  32617=>"110111111",
  32618=>"111111110",
  32619=>"111111101",
  32620=>"110000000",
  32621=>"001000000",
  32622=>"000000000",
  32623=>"000101111",
  32624=>"000000000",
  32625=>"111110000",
  32626=>"000000001",
  32627=>"100110111",
  32628=>"111011000",
  32629=>"000000000",
  32630=>"110111111",
  32631=>"100100000",
  32632=>"010111111",
  32633=>"111000111",
  32634=>"111011001",
  32635=>"111110111",
  32636=>"111100000",
  32637=>"001001000",
  32638=>"111011011",
  32639=>"111111111",
  32640=>"010111101",
  32641=>"011011011",
  32642=>"000011111",
  32643=>"000000000",
  32644=>"000110111",
  32645=>"100101000",
  32646=>"111010011",
  32647=>"000110111",
  32648=>"000111011",
  32649=>"011001011",
  32650=>"111111010",
  32651=>"111111000",
  32652=>"111000111",
  32653=>"000111110",
  32654=>"011001000",
  32655=>"000000000",
  32656=>"100100100",
  32657=>"101011111",
  32658=>"010000001",
  32659=>"111111111",
  32660=>"111111000",
  32661=>"000010000",
  32662=>"100111110",
  32663=>"111110000",
  32664=>"000000111",
  32665=>"111111110",
  32666=>"111111111",
  32667=>"001000000",
  32668=>"000001111",
  32669=>"000000000",
  32670=>"100000000",
  32671=>"000110111",
  32672=>"011001100",
  32673=>"111110001",
  32674=>"110100100",
  32675=>"100000011",
  32676=>"000000100",
  32677=>"000110010",
  32678=>"000000000",
  32679=>"111111111",
  32680=>"000000011",
  32681=>"000000000",
  32682=>"111110011",
  32683=>"010111111",
  32684=>"000000111",
  32685=>"110000111",
  32686=>"010001001",
  32687=>"111001101",
  32688=>"110001001",
  32689=>"000000011",
  32690=>"000111111",
  32691=>"110000111",
  32692=>"111111111",
  32693=>"000000000",
  32694=>"110111101",
  32695=>"000000000",
  32696=>"000000001",
  32697=>"111111011",
  32698=>"101010000",
  32699=>"011100100",
  32700=>"110111000",
  32701=>"000000100",
  32702=>"011011010",
  32703=>"001011011",
  32704=>"111111000",
  32705=>"100000000",
  32706=>"000000000",
  32707=>"111111011",
  32708=>"010100001",
  32709=>"000000111",
  32710=>"111000011",
  32711=>"001000101",
  32712=>"100101111",
  32713=>"111111111",
  32714=>"000000000",
  32715=>"000001000",
  32716=>"000000000",
  32717=>"111000000",
  32718=>"000000000",
  32719=>"110010111",
  32720=>"111111111",
  32721=>"000000100",
  32722=>"000001111",
  32723=>"111011011",
  32724=>"000000000",
  32725=>"100000000",
  32726=>"110010011",
  32727=>"000010111",
  32728=>"000000000",
  32729=>"111111111",
  32730=>"111011000",
  32731=>"000001111",
  32732=>"100100100",
  32733=>"011111111",
  32734=>"011011011",
  32735=>"000000010",
  32736=>"111111111",
  32737=>"011011011",
  32738=>"000000011",
  32739=>"000010111",
  32740=>"111111111",
  32741=>"111111011",
  32742=>"000001111",
  32743=>"110111111",
  32744=>"111111000",
  32745=>"001111111",
  32746=>"100000000",
  32747=>"111110001",
  32748=>"111100000",
  32749=>"011111100",
  32750=>"111101000",
  32751=>"000000000",
  32752=>"000111101",
  32753=>"110111000",
  32754=>"000011000",
  32755=>"110100000",
  32756=>"010110011",
  32757=>"000110110",
  32758=>"111111111",
  32759=>"111011000",
  32760=>"000001011",
  32761=>"110000100",
  32762=>"000111111",
  32763=>"111010000",
  32764=>"110111111",
  32765=>"001001000",
  32766=>"111011011",
  32767=>"000000011",
  32768=>"111110000",
  32769=>"000000000",
  32770=>"111000111",
  32771=>"111000000",
  32772=>"000000110",
  32773=>"100111101",
  32774=>"000000000",
  32775=>"111111000",
  32776=>"000001111",
  32777=>"000111111",
  32778=>"011011011",
  32779=>"110111111",
  32780=>"000000111",
  32781=>"000000000",
  32782=>"000000000",
  32783=>"110000000",
  32784=>"000000000",
  32785=>"100111111",
  32786=>"000000000",
  32787=>"111101111",
  32788=>"000000000",
  32789=>"000000000",
  32790=>"100111101",
  32791=>"010000000",
  32792=>"000000000",
  32793=>"000011011",
  32794=>"000000111",
  32795=>"000111111",
  32796=>"001000000",
  32797=>"101111000",
  32798=>"010000000",
  32799=>"000000000",
  32800=>"111011000",
  32801=>"110101001",
  32802=>"111000101",
  32803=>"111000100",
  32804=>"001001101",
  32805=>"100000000",
  32806=>"111100111",
  32807=>"111111011",
  32808=>"000001101",
  32809=>"110010010",
  32810=>"000000000",
  32811=>"000000101",
  32812=>"000000110",
  32813=>"111111000",
  32814=>"111011011",
  32815=>"100000000",
  32816=>"011110110",
  32817=>"000000000",
  32818=>"000000011",
  32819=>"011001001",
  32820=>"111100000",
  32821=>"110010001",
  32822=>"011111001",
  32823=>"100000101",
  32824=>"000001000",
  32825=>"111111111",
  32826=>"111000011",
  32827=>"000000100",
  32828=>"011000000",
  32829=>"111111111",
  32830=>"001001111",
  32831=>"111000111",
  32832=>"100000000",
  32833=>"101000000",
  32834=>"000000000",
  32835=>"000111011",
  32836=>"110111111",
  32837=>"011111011",
  32838=>"000000000",
  32839=>"000000000",
  32840=>"111011000",
  32841=>"111000000",
  32842=>"111001101",
  32843=>"011011000",
  32844=>"101100000",
  32845=>"000000001",
  32846=>"011011111",
  32847=>"000010100",
  32848=>"000000111",
  32849=>"110111111",
  32850=>"000000000",
  32851=>"001001000",
  32852=>"000000000",
  32853=>"000100111",
  32854=>"000000100",
  32855=>"111111000",
  32856=>"100111011",
  32857=>"111101111",
  32858=>"100101111",
  32859=>"100110011",
  32860=>"011011111",
  32861=>"011111111",
  32862=>"001001000",
  32863=>"111000000",
  32864=>"111111111",
  32865=>"110010010",
  32866=>"000111111",
  32867=>"101111011",
  32868=>"000000110",
  32869=>"111100110",
  32870=>"011101100",
  32871=>"111111110",
  32872=>"111111111",
  32873=>"111101101",
  32874=>"101000000",
  32875=>"001101000",
  32876=>"110000111",
  32877=>"000000000",
  32878=>"001001000",
  32879=>"100000000",
  32880=>"011001001",
  32881=>"011101111",
  32882=>"011111111",
  32883=>"000000000",
  32884=>"000000000",
  32885=>"110100101",
  32886=>"000100111",
  32887=>"011001111",
  32888=>"110011000",
  32889=>"011111111",
  32890=>"000001100",
  32891=>"111011000",
  32892=>"110100100",
  32893=>"000000000",
  32894=>"000000000",
  32895=>"000000111",
  32896=>"000110111",
  32897=>"111001000",
  32898=>"000000111",
  32899=>"111111000",
  32900=>"111111000",
  32901=>"110000110",
  32902=>"111111111",
  32903=>"000000000",
  32904=>"000000111",
  32905=>"000000110",
  32906=>"010110000",
  32907=>"001000000",
  32908=>"111100000",
  32909=>"111111111",
  32910=>"111001001",
  32911=>"000000000",
  32912=>"111111111",
  32913=>"111111101",
  32914=>"000000001",
  32915=>"110111111",
  32916=>"000000110",
  32917=>"111111111",
  32918=>"000110010",
  32919=>"111111111",
  32920=>"000000111",
  32921=>"111110110",
  32922=>"000000000",
  32923=>"110110000",
  32924=>"111101000",
  32925=>"011011001",
  32926=>"001000000",
  32927=>"000000000",
  32928=>"101000000",
  32929=>"111111011",
  32930=>"000000000",
  32931=>"100100100",
  32932=>"000110011",
  32933=>"111111111",
  32934=>"000000111",
  32935=>"111111111",
  32936=>"001001111",
  32937=>"101001111",
  32938=>"100111111",
  32939=>"111010000",
  32940=>"111000000",
  32941=>"000000000",
  32942=>"111111101",
  32943=>"000000001",
  32944=>"111000000",
  32945=>"110110111",
  32946=>"111111000",
  32947=>"000000000",
  32948=>"000100000",
  32949=>"100111111",
  32950=>"111111111",
  32951=>"000101111",
  32952=>"110010000",
  32953=>"111101111",
  32954=>"000000001",
  32955=>"100000111",
  32956=>"000100111",
  32957=>"111000000",
  32958=>"110101001",
  32959=>"011001000",
  32960=>"001000111",
  32961=>"000000000",
  32962=>"111111111",
  32963=>"000000100",
  32964=>"111111111",
  32965=>"111111111",
  32966=>"000000000",
  32967=>"000111001",
  32968=>"000000000",
  32969=>"110011000",
  32970=>"000000000",
  32971=>"000000000",
  32972=>"111000001",
  32973=>"000000111",
  32974=>"111111111",
  32975=>"111000000",
  32976=>"110111111",
  32977=>"110110111",
  32978=>"111110000",
  32979=>"000000000",
  32980=>"011000000",
  32981=>"111001000",
  32982=>"000000111",
  32983=>"000010111",
  32984=>"100011000",
  32985=>"000000001",
  32986=>"000000000",
  32987=>"111111011",
  32988=>"000100000",
  32989=>"000101111",
  32990=>"111001111",
  32991=>"100100001",
  32992=>"000000000",
  32993=>"000100111",
  32994=>"100100111",
  32995=>"000000000",
  32996=>"001001000",
  32997=>"000100000",
  32998=>"001000011",
  32999=>"011001001",
  33000=>"000001111",
  33001=>"000001111",
  33002=>"111011111",
  33003=>"111111111",
  33004=>"000000011",
  33005=>"000100110",
  33006=>"001001111",
  33007=>"000001111",
  33008=>"111111111",
  33009=>"000000000",
  33010=>"111111000",
  33011=>"111111101",
  33012=>"100110010",
  33013=>"111000000",
  33014=>"010000000",
  33015=>"000111111",
  33016=>"000100110",
  33017=>"111110100",
  33018=>"000000111",
  33019=>"101000010",
  33020=>"100100000",
  33021=>"111010011",
  33022=>"110111111",
  33023=>"000000100",
  33024=>"000000100",
  33025=>"000000000",
  33026=>"111111100",
  33027=>"011001111",
  33028=>"110111111",
  33029=>"000000111",
  33030=>"111111111",
  33031=>"110000101",
  33032=>"111111110",
  33033=>"100111111",
  33034=>"000001111",
  33035=>"000100000",
  33036=>"000000000",
  33037=>"111111001",
  33038=>"111111111",
  33039=>"000000000",
  33040=>"111111111",
  33041=>"111111111",
  33042=>"110100111",
  33043=>"000100101",
  33044=>"000000000",
  33045=>"111111011",
  33046=>"001111001",
  33047=>"101101000",
  33048=>"111111111",
  33049=>"111110110",
  33050=>"111101000",
  33051=>"000100101",
  33052=>"110100110",
  33053=>"111111111",
  33054=>"000000000",
  33055=>"011010000",
  33056=>"000000000",
  33057=>"000011001",
  33058=>"000100000",
  33059=>"111111111",
  33060=>"010000111",
  33061=>"010111111",
  33062=>"000000000",
  33063=>"000000100",
  33064=>"000000111",
  33065=>"011011000",
  33066=>"000000000",
  33067=>"101100000",
  33068=>"000000000",
  33069=>"110110111",
  33070=>"111011000",
  33071=>"111111111",
  33072=>"011010000",
  33073=>"111001100",
  33074=>"000000000",
  33075=>"000000111",
  33076=>"000000000",
  33077=>"011111011",
  33078=>"100100100",
  33079=>"001001011",
  33080=>"100100100",
  33081=>"111001000",
  33082=>"111111101",
  33083=>"111111111",
  33084=>"000100110",
  33085=>"011010111",
  33086=>"000010101",
  33087=>"100101111",
  33088=>"000000011",
  33089=>"000000000",
  33090=>"111110111",
  33091=>"000000000",
  33092=>"000000000",
  33093=>"111101111",
  33094=>"000000000",
  33095=>"111111111",
  33096=>"110110100",
  33097=>"000000000",
  33098=>"100000001",
  33099=>"111110100",
  33100=>"100000110",
  33101=>"000000000",
  33102=>"111011110",
  33103=>"110110000",
  33104=>"000110110",
  33105=>"001001111",
  33106=>"100000000",
  33107=>"111111010",
  33108=>"000100110",
  33109=>"011011011",
  33110=>"110101001",
  33111=>"111111110",
  33112=>"000000000",
  33113=>"101111111",
  33114=>"111111111",
  33115=>"111111000",
  33116=>"000001111",
  33117=>"000000000",
  33118=>"000000111",
  33119=>"001011111",
  33120=>"100100001",
  33121=>"111101000",
  33122=>"000000011",
  33123=>"000110111",
  33124=>"000000000",
  33125=>"111111001",
  33126=>"111100000",
  33127=>"101101010",
  33128=>"111011001",
  33129=>"000000000",
  33130=>"000011010",
  33131=>"111011111",
  33132=>"110000100",
  33133=>"001111001",
  33134=>"000111111",
  33135=>"000000000",
  33136=>"000000100",
  33137=>"000000000",
  33138=>"111111111",
  33139=>"010100010",
  33140=>"000000000",
  33141=>"000100100",
  33142=>"011000111",
  33143=>"101111000",
  33144=>"000000111",
  33145=>"100110011",
  33146=>"111110110",
  33147=>"101001001",
  33148=>"111011011",
  33149=>"111111100",
  33150=>"000000000",
  33151=>"000000000",
  33152=>"111011111",
  33153=>"000010000",
  33154=>"111111111",
  33155=>"101001001",
  33156=>"100100111",
  33157=>"111111101",
  33158=>"111111011",
  33159=>"000011111",
  33160=>"000110111",
  33161=>"000100000",
  33162=>"000000000",
  33163=>"000000000",
  33164=>"110000111",
  33165=>"001000001",
  33166=>"011111111",
  33167=>"000000000",
  33168=>"000000000",
  33169=>"111011001",
  33170=>"000000001",
  33171=>"000100111",
  33172=>"111001000",
  33173=>"000111000",
  33174=>"000000100",
  33175=>"110000000",
  33176=>"000000001",
  33177=>"110010110",
  33178=>"000000000",
  33179=>"111111001",
  33180=>"101000000",
  33181=>"111111111",
  33182=>"011000000",
  33183=>"000000000",
  33184=>"000001101",
  33185=>"000100111",
  33186=>"011000100",
  33187=>"111111111",
  33188=>"111111111",
  33189=>"000001110",
  33190=>"111111111",
  33191=>"110000010",
  33192=>"000001010",
  33193=>"000000111",
  33194=>"001011111",
  33195=>"111010000",
  33196=>"000000111",
  33197=>"111001000",
  33198=>"000000100",
  33199=>"000000000",
  33200=>"100000000",
  33201=>"101111111",
  33202=>"111111001",
  33203=>"111101111",
  33204=>"111100000",
  33205=>"111111101",
  33206=>"111110101",
  33207=>"010001000",
  33208=>"000000000",
  33209=>"000000011",
  33210=>"111011111",
  33211=>"010111101",
  33212=>"000000000",
  33213=>"010000101",
  33214=>"111010011",
  33215=>"001001011",
  33216=>"001000000",
  33217=>"111111111",
  33218=>"000011010",
  33219=>"000000010",
  33220=>"111101100",
  33221=>"001011111",
  33222=>"111101011",
  33223=>"100100111",
  33224=>"000101101",
  33225=>"111111001",
  33226=>"000000111",
  33227=>"110111111",
  33228=>"000100011",
  33229=>"000000111",
  33230=>"000000000",
  33231=>"111111111",
  33232=>"001000011",
  33233=>"001111111",
  33234=>"001001000",
  33235=>"111111000",
  33236=>"110111111",
  33237=>"100000101",
  33238=>"000000000",
  33239=>"000000111",
  33240=>"111111111",
  33241=>"011111101",
  33242=>"111110000",
  33243=>"000000100",
  33244=>"000000000",
  33245=>"110000001",
  33246=>"111011011",
  33247=>"000011001",
  33248=>"000000010",
  33249=>"000000001",
  33250=>"000000000",
  33251=>"000001101",
  33252=>"111011111",
  33253=>"111000000",
  33254=>"000001000",
  33255=>"110110111",
  33256=>"011011011",
  33257=>"001111111",
  33258=>"000000000",
  33259=>"001101101",
  33260=>"011011000",
  33261=>"001000000",
  33262=>"011011001",
  33263=>"111111111",
  33264=>"000000000",
  33265=>"111111010",
  33266=>"111111111",
  33267=>"000000000",
  33268=>"111011000",
  33269=>"000000000",
  33270=>"000100100",
  33271=>"000000001",
  33272=>"111111111",
  33273=>"010000000",
  33274=>"000000111",
  33275=>"111111111",
  33276=>"000000000",
  33277=>"100100100",
  33278=>"111111011",
  33279=>"000000000",
  33280=>"110000110",
  33281=>"010111001",
  33282=>"111111111",
  33283=>"000000000",
  33284=>"111111000",
  33285=>"000000000",
  33286=>"111111011",
  33287=>"111111100",
  33288=>"000000110",
  33289=>"010000000",
  33290=>"000000000",
  33291=>"100111111",
  33292=>"111111101",
  33293=>"001111111",
  33294=>"111111000",
  33295=>"111111111",
  33296=>"111111011",
  33297=>"111111111",
  33298=>"000000000",
  33299=>"111111111",
  33300=>"111000000",
  33301=>"000010000",
  33302=>"111111001",
  33303=>"011001011",
  33304=>"111111111",
  33305=>"011111111",
  33306=>"111111111",
  33307=>"000000000",
  33308=>"011011001",
  33309=>"010000010",
  33310=>"000001111",
  33311=>"111111011",
  33312=>"110000010",
  33313=>"111001111",
  33314=>"000000000",
  33315=>"111111111",
  33316=>"000111111",
  33317=>"000111111",
  33318=>"000000000",
  33319=>"000111111",
  33320=>"111111111",
  33321=>"000000000",
  33322=>"000000000",
  33323=>"111111100",
  33324=>"111000000",
  33325=>"110110111",
  33326=>"010000000",
  33327=>"000000000",
  33328=>"000101111",
  33329=>"110111111",
  33330=>"001001001",
  33331=>"000000000",
  33332=>"010010111",
  33333=>"001001001",
  33334=>"111111111",
  33335=>"111101111",
  33336=>"111000000",
  33337=>"001111110",
  33338=>"000111111",
  33339=>"111010110",
  33340=>"000000011",
  33341=>"111111111",
  33342=>"101000000",
  33343=>"001000000",
  33344=>"000000000",
  33345=>"000010111",
  33346=>"000000010",
  33347=>"111111111",
  33348=>"100100111",
  33349=>"110100100",
  33350=>"000000000",
  33351=>"000000000",
  33352=>"000000010",
  33353=>"000000000",
  33354=>"000000000",
  33355=>"000000001",
  33356=>"111111111",
  33357=>"111000000",
  33358=>"011010110",
  33359=>"111011001",
  33360=>"000100110",
  33361=>"111111000",
  33362=>"111000110",
  33363=>"111111111",
  33364=>"000000000",
  33365=>"000010000",
  33366=>"001000111",
  33367=>"000000000",
  33368=>"000011111",
  33369=>"000000000",
  33370=>"100000000",
  33371=>"100111111",
  33372=>"000000000",
  33373=>"101111111",
  33374=>"001111111",
  33375=>"000000000",
  33376=>"000111111",
  33377=>"011001000",
  33378=>"111111000",
  33379=>"010000010",
  33380=>"000000000",
  33381=>"001000001",
  33382=>"111011000",
  33383=>"111111111",
  33384=>"110111111",
  33385=>"111000000",
  33386=>"010111111",
  33387=>"000001000",
  33388=>"101111010",
  33389=>"101111111",
  33390=>"011001111",
  33391=>"000001110",
  33392=>"110110110",
  33393=>"000000001",
  33394=>"000000000",
  33395=>"100001000",
  33396=>"000000000",
  33397=>"111111111",
  33398=>"000000000",
  33399=>"000000111",
  33400=>"111010000",
  33401=>"001001000",
  33402=>"000110111",
  33403=>"011011011",
  33404=>"000011111",
  33405=>"000000000",
  33406=>"000000000",
  33407=>"000010010",
  33408=>"111111101",
  33409=>"000000111",
  33410=>"000000000",
  33411=>"000100111",
  33412=>"011111111",
  33413=>"000000110",
  33414=>"001111111",
  33415=>"011111111",
  33416=>"010000001",
  33417=>"000000000",
  33418=>"010011111",
  33419=>"000000010",
  33420=>"111110110",
  33421=>"111000000",
  33422=>"111111111",
  33423=>"000100110",
  33424=>"111111010",
  33425=>"000000110",
  33426=>"111110000",
  33427=>"001001000",
  33428=>"010011001",
  33429=>"000000000",
  33430=>"000000000",
  33431=>"000000111",
  33432=>"001000111",
  33433=>"100100100",
  33434=>"111111011",
  33435=>"111111111",
  33436=>"001000100",
  33437=>"000000100",
  33438=>"111111111",
  33439=>"000000000",
  33440=>"110111111",
  33441=>"111111011",
  33442=>"000000000",
  33443=>"111111111",
  33444=>"000000011",
  33445=>"011000000",
  33446=>"110010110",
  33447=>"111111111",
  33448=>"111111111",
  33449=>"111111111",
  33450=>"111111111",
  33451=>"000111111",
  33452=>"001001001",
  33453=>"000111111",
  33454=>"111111111",
  33455=>"000001000",
  33456=>"000000000",
  33457=>"011001001",
  33458=>"111110110",
  33459=>"000111111",
  33460=>"111111110",
  33461=>"110000000",
  33462=>"000000111",
  33463=>"011000000",
  33464=>"000100000",
  33465=>"000000000",
  33466=>"100000111",
  33467=>"111001111",
  33468=>"001111111",
  33469=>"111110000",
  33470=>"110111111",
  33471=>"011000000",
  33472=>"000000000",
  33473=>"111111001",
  33474=>"000000110",
  33475=>"110111111",
  33476=>"111000000",
  33477=>"111000000",
  33478=>"000001101",
  33479=>"001001000",
  33480=>"000000111",
  33481=>"001000001",
  33482=>"111111111",
  33483=>"000000011",
  33484=>"011000000",
  33485=>"100111000",
  33486=>"110111111",
  33487=>"111111111",
  33488=>"111111000",
  33489=>"000000110",
  33490=>"000000000",
  33491=>"001111111",
  33492=>"111101111",
  33493=>"111111111",
  33494=>"111111000",
  33495=>"000000000",
  33496=>"111001000",
  33497=>"110110100",
  33498=>"000000000",
  33499=>"000110111",
  33500=>"111111111",
  33501=>"000000001",
  33502=>"000100000",
  33503=>"001101000",
  33504=>"111111111",
  33505=>"100010110",
  33506=>"100000000",
  33507=>"110000000",
  33508=>"000100100",
  33509=>"111111111",
  33510=>"000110010",
  33511=>"101100101",
  33512=>"111010111",
  33513=>"000000101",
  33514=>"111111000",
  33515=>"011001001",
  33516=>"111010111",
  33517=>"000000000",
  33518=>"111010000",
  33519=>"000000000",
  33520=>"000000111",
  33521=>"111100100",
  33522=>"100111111",
  33523=>"100111001",
  33524=>"001000000",
  33525=>"000000000",
  33526=>"110010000",
  33527=>"111111111",
  33528=>"111011110",
  33529=>"111111111",
  33530=>"100000000",
  33531=>"111111111",
  33532=>"001101100",
  33533=>"101000000",
  33534=>"001000000",
  33535=>"000100000",
  33536=>"111111000",
  33537=>"000000000",
  33538=>"111111111",
  33539=>"111111111",
  33540=>"111111111",
  33541=>"000000000",
  33542=>"000000001",
  33543=>"000000010",
  33544=>"111111100",
  33545=>"000000000",
  33546=>"111111111",
  33547=>"101111111",
  33548=>"100101111",
  33549=>"111111110",
  33550=>"000000011",
  33551=>"111100100",
  33552=>"011011111",
  33553=>"110110000",
  33554=>"000000000",
  33555=>"110010000",
  33556=>"000000000",
  33557=>"000011001",
  33558=>"001000000",
  33559=>"111111111",
  33560=>"111111111",
  33561=>"000000000",
  33562=>"001111111",
  33563=>"100100100",
  33564=>"000000000",
  33565=>"000000000",
  33566=>"111111111",
  33567=>"111110010",
  33568=>"000100000",
  33569=>"000111100",
  33570=>"110110000",
  33571=>"000000000",
  33572=>"111111111",
  33573=>"000000000",
  33574=>"011111110",
  33575=>"000000111",
  33576=>"100110111",
  33577=>"111111111",
  33578=>"000000100",
  33579=>"111000000",
  33580=>"100110111",
  33581=>"111111101",
  33582=>"001000000",
  33583=>"000101001",
  33584=>"000001111",
  33585=>"011000000",
  33586=>"111111110",
  33587=>"000011000",
  33588=>"101000000",
  33589=>"000000101",
  33590=>"000000000",
  33591=>"111111111",
  33592=>"111111111",
  33593=>"000000000",
  33594=>"000000000",
  33595=>"111111001",
  33596=>"000000000",
  33597=>"000000000",
  33598=>"111111101",
  33599=>"000010010",
  33600=>"101000000",
  33601=>"101111111",
  33602=>"111111111",
  33603=>"000111111",
  33604=>"000000000",
  33605=>"000111111",
  33606=>"111111111",
  33607=>"000100100",
  33608=>"000000011",
  33609=>"000000000",
  33610=>"000000111",
  33611=>"000001000",
  33612=>"101100100",
  33613=>"100100111",
  33614=>"010110110",
  33615=>"000000100",
  33616=>"101111010",
  33617=>"000000000",
  33618=>"000100111",
  33619=>"000000000",
  33620=>"000001011",
  33621=>"001011011",
  33622=>"111000100",
  33623=>"111111111",
  33624=>"111111111",
  33625=>"000110111",
  33626=>"111111111",
  33627=>"010111000",
  33628=>"110110111",
  33629=>"000000000",
  33630=>"000000000",
  33631=>"111111111",
  33632=>"110000000",
  33633=>"111111111",
  33634=>"111110111",
  33635=>"111111101",
  33636=>"000000000",
  33637=>"000011011",
  33638=>"011000000",
  33639=>"000000000",
  33640=>"101101001",
  33641=>"111000100",
  33642=>"111111111",
  33643=>"111000000",
  33644=>"000000000",
  33645=>"101111111",
  33646=>"111110100",
  33647=>"111100100",
  33648=>"111111101",
  33649=>"111111011",
  33650=>"010100100",
  33651=>"001001000",
  33652=>"111111111",
  33653=>"101101000",
  33654=>"111000000",
  33655=>"000001000",
  33656=>"111111011",
  33657=>"000000000",
  33658=>"000000101",
  33659=>"111011011",
  33660=>"100111111",
  33661=>"000000000",
  33662=>"000000000",
  33663=>"011000000",
  33664=>"011011111",
  33665=>"011111111",
  33666=>"111011001",
  33667=>"111111111",
  33668=>"000010001",
  33669=>"100100101",
  33670=>"111000100",
  33671=>"000001011",
  33672=>"000000011",
  33673=>"111000011",
  33674=>"011011011",
  33675=>"111001000",
  33676=>"101000000",
  33677=>"000000000",
  33678=>"100101111",
  33679=>"000000000",
  33680=>"111011111",
  33681=>"001000000",
  33682=>"000110110",
  33683=>"111000000",
  33684=>"000000000",
  33685=>"000010111",
  33686=>"000001001",
  33687=>"001001001",
  33688=>"100101000",
  33689=>"111111111",
  33690=>"000000101",
  33691=>"111111111",
  33692=>"111011111",
  33693=>"011000000",
  33694=>"111111001",
  33695=>"111111000",
  33696=>"000000000",
  33697=>"011001000",
  33698=>"000001111",
  33699=>"111000000",
  33700=>"111111111",
  33701=>"000110111",
  33702=>"001001111",
  33703=>"011111101",
  33704=>"000000000",
  33705=>"111011000",
  33706=>"111001001",
  33707=>"111000000",
  33708=>"000000000",
  33709=>"000001111",
  33710=>"111000110",
  33711=>"000111111",
  33712=>"011010111",
  33713=>"010000000",
  33714=>"111110111",
  33715=>"000000000",
  33716=>"111111111",
  33717=>"000010111",
  33718=>"111001111",
  33719=>"000111000",
  33720=>"000000000",
  33721=>"111111111",
  33722=>"100000000",
  33723=>"111110100",
  33724=>"000000001",
  33725=>"000000100",
  33726=>"110010000",
  33727=>"001101111",
  33728=>"000011011",
  33729=>"000011111",
  33730=>"111111111",
  33731=>"110111111",
  33732=>"111111111",
  33733=>"100000111",
  33734=>"111101000",
  33735=>"000000000",
  33736=>"111111000",
  33737=>"001001101",
  33738=>"000000010",
  33739=>"000111111",
  33740=>"000000000",
  33741=>"111011111",
  33742=>"101001001",
  33743=>"111111111",
  33744=>"111111111",
  33745=>"101101100",
  33746=>"110110111",
  33747=>"001111001",
  33748=>"000011111",
  33749=>"111111111",
  33750=>"111011000",
  33751=>"011010001",
  33752=>"001110111",
  33753=>"111010110",
  33754=>"000011011",
  33755=>"101000000",
  33756=>"000000000",
  33757=>"111110100",
  33758=>"111111111",
  33759=>"001011001",
  33760=>"110110111",
  33761=>"111101111",
  33762=>"111111011",
  33763=>"111000000",
  33764=>"100000000",
  33765=>"000000001",
  33766=>"000000111",
  33767=>"111010000",
  33768=>"000000111",
  33769=>"100000000",
  33770=>"000111111",
  33771=>"001000000",
  33772=>"000111111",
  33773=>"010010110",
  33774=>"001001001",
  33775=>"111101101",
  33776=>"000000111",
  33777=>"111111111",
  33778=>"111111101",
  33779=>"100001111",
  33780=>"000000000",
  33781=>"000110000",
  33782=>"111111011",
  33783=>"110000000",
  33784=>"111001100",
  33785=>"001001001",
  33786=>"001000000",
  33787=>"110111110",
  33788=>"000000000",
  33789=>"111111111",
  33790=>"000000110",
  33791=>"000000000",
  33792=>"111010010",
  33793=>"000000000",
  33794=>"000000000",
  33795=>"000000010",
  33796=>"111000110",
  33797=>"011110111",
  33798=>"000000001",
  33799=>"111101100",
  33800=>"000000101",
  33801=>"011111111",
  33802=>"111111001",
  33803=>"000101111",
  33804=>"000100111",
  33805=>"111111111",
  33806=>"101000000",
  33807=>"111111111",
  33808=>"000111000",
  33809=>"000000000",
  33810=>"000000000",
  33811=>"000000000",
  33812=>"000000000",
  33813=>"111111111",
  33814=>"000000000",
  33815=>"011011011",
  33816=>"110110110",
  33817=>"000001001",
  33818=>"000000010",
  33819=>"001001111",
  33820=>"111111111",
  33821=>"000101111",
  33822=>"111111000",
  33823=>"111111111",
  33824=>"000110111",
  33825=>"111111111",
  33826=>"000000000",
  33827=>"111101000",
  33828=>"000000010",
  33829=>"000000000",
  33830=>"001111111",
  33831=>"111111111",
  33832=>"110111101",
  33833=>"000000000",
  33834=>"001001001",
  33835=>"111111111",
  33836=>"111111100",
  33837=>"110111000",
  33838=>"000000010",
  33839=>"011001001",
  33840=>"111111110",
  33841=>"101000000",
  33842=>"000000000",
  33843=>"011111111",
  33844=>"111111000",
  33845=>"100100111",
  33846=>"100000000",
  33847=>"111111111",
  33848=>"011001000",
  33849=>"000000000",
  33850=>"000000000",
  33851=>"111100000",
  33852=>"101100100",
  33853=>"011000000",
  33854=>"001001111",
  33855=>"000000000",
  33856=>"111111100",
  33857=>"111111111",
  33858=>"000000000",
  33859=>"111111111",
  33860=>"000000010",
  33861=>"000000000",
  33862=>"011111110",
  33863=>"000100000",
  33864=>"001001000",
  33865=>"111111111",
  33866=>"000000110",
  33867=>"000000000",
  33868=>"111111111",
  33869=>"000001000",
  33870=>"111100101",
  33871=>"000000111",
  33872=>"000000100",
  33873=>"000000010",
  33874=>"111111111",
  33875=>"100100000",
  33876=>"111111011",
  33877=>"000000000",
  33878=>"011000000",
  33879=>"111110000",
  33880=>"111011111",
  33881=>"101100111",
  33882=>"001000000",
  33883=>"111110110",
  33884=>"111100000",
  33885=>"111101100",
  33886=>"111111111",
  33887=>"010111001",
  33888=>"101000000",
  33889=>"100000000",
  33890=>"101110111",
  33891=>"010000001",
  33892=>"000000000",
  33893=>"110110000",
  33894=>"010000111",
  33895=>"111111111",
  33896=>"000000001",
  33897=>"000000100",
  33898=>"000000000",
  33899=>"000110000",
  33900=>"111100110",
  33901=>"000000000",
  33902=>"000000000",
  33903=>"111111111",
  33904=>"000000000",
  33905=>"000011111",
  33906=>"111111111",
  33907=>"111111111",
  33908=>"011011001",
  33909=>"000100100",
  33910=>"000111111",
  33911=>"000000100",
  33912=>"000001011",
  33913=>"110111001",
  33914=>"000000000",
  33915=>"000000001",
  33916=>"111111111",
  33917=>"000001101",
  33918=>"000000000",
  33919=>"000010010",
  33920=>"111111111",
  33921=>"000000000",
  33922=>"100100100",
  33923=>"011011011",
  33924=>"000000001",
  33925=>"110101111",
  33926=>"110100000",
  33927=>"000000000",
  33928=>"110000010",
  33929=>"111111000",
  33930=>"001001000",
  33931=>"011111111",
  33932=>"100000000",
  33933=>"110110100",
  33934=>"000000000",
  33935=>"001111111",
  33936=>"000101111",
  33937=>"111111111",
  33938=>"000000000",
  33939=>"100100110",
  33940=>"000000000",
  33941=>"000000110",
  33942=>"000000000",
  33943=>"000000000",
  33944=>"100100000",
  33945=>"111000010",
  33946=>"111111111",
  33947=>"000000010",
  33948=>"010110001",
  33949=>"111110111",
  33950=>"000000000",
  33951=>"101000000",
  33952=>"011010000",
  33953=>"000000000",
  33954=>"000000000",
  33955=>"000000000",
  33956=>"000000000",
  33957=>"111111111",
  33958=>"010000000",
  33959=>"111111111",
  33960=>"001000000",
  33961=>"111111111",
  33962=>"000111111",
  33963=>"000000000",
  33964=>"000000001",
  33965=>"111111110",
  33966=>"111111111",
  33967=>"000000000",
  33968=>"000010011",
  33969=>"000000110",
  33970=>"111111110",
  33971=>"000000000",
  33972=>"001011001",
  33973=>"001111111",
  33974=>"001001111",
  33975=>"000000100",
  33976=>"110110010",
  33977=>"000111100",
  33978=>"000001000",
  33979=>"101001001",
  33980=>"000000000",
  33981=>"001001000",
  33982=>"000000000",
  33983=>"000000000",
  33984=>"001011111",
  33985=>"101111100",
  33986=>"100100110",
  33987=>"111111111",
  33988=>"000000110",
  33989=>"100000000",
  33990=>"100110111",
  33991=>"100110110",
  33992=>"000011111",
  33993=>"011011111",
  33994=>"111000000",
  33995=>"010010011",
  33996=>"000011111",
  33997=>"111111111",
  33998=>"111111111",
  33999=>"010011000",
  34000=>"111111010",
  34001=>"111111111",
  34002=>"000110010",
  34003=>"110100000",
  34004=>"000000000",
  34005=>"000111111",
  34006=>"000000000",
  34007=>"110100111",
  34008=>"000000000",
  34009=>"011011101",
  34010=>"111101000",
  34011=>"000000000",
  34012=>"011111011",
  34013=>"000000011",
  34014=>"000000000",
  34015=>"110111111",
  34016=>"000000011",
  34017=>"010011000",
  34018=>"000000011",
  34019=>"000000000",
  34020=>"000000001",
  34021=>"111100000",
  34022=>"000000000",
  34023=>"000111110",
  34024=>"000000000",
  34025=>"011001001",
  34026=>"101111111",
  34027=>"110000000",
  34028=>"111111111",
  34029=>"000000110",
  34030=>"100100001",
  34031=>"000000000",
  34032=>"010110110",
  34033=>"000100101",
  34034=>"000110111",
  34035=>"111111111",
  34036=>"111111111",
  34037=>"001000000",
  34038=>"000000011",
  34039=>"111111000",
  34040=>"100100000",
  34041=>"111001000",
  34042=>"111011111",
  34043=>"011001001",
  34044=>"111111110",
  34045=>"000010110",
  34046=>"000100111",
  34047=>"000000000",
  34048=>"111001001",
  34049=>"111100110",
  34050=>"111110111",
  34051=>"001111111",
  34052=>"111101000",
  34053=>"000000100",
  34054=>"111111111",
  34055=>"000000000",
  34056=>"000000000",
  34057=>"000000000",
  34058=>"111111111",
  34059=>"101111111",
  34060=>"011011111",
  34061=>"110111111",
  34062=>"000000010",
  34063=>"001000000",
  34064=>"000100000",
  34065=>"000000000",
  34066=>"111001111",
  34067=>"000000000",
  34068=>"000000000",
  34069=>"111111010",
  34070=>"011011110",
  34071=>"000000000",
  34072=>"000000000",
  34073=>"111111000",
  34074=>"111110000",
  34075=>"010000110",
  34076=>"000000010",
  34077=>"001000000",
  34078=>"110111111",
  34079=>"000100010",
  34080=>"001001000",
  34081=>"001001011",
  34082=>"001000000",
  34083=>"111111111",
  34084=>"111111110",
  34085=>"100100100",
  34086=>"000111111",
  34087=>"100000000",
  34088=>"000110010",
  34089=>"001001000",
  34090=>"000000011",
  34091=>"011111111",
  34092=>"111111101",
  34093=>"000000100",
  34094=>"000000000",
  34095=>"111101000",
  34096=>"000000000",
  34097=>"000100111",
  34098=>"001111001",
  34099=>"000000000",
  34100=>"011000000",
  34101=>"000000000",
  34102=>"111000000",
  34103=>"100100110",
  34104=>"000110111",
  34105=>"110111111",
  34106=>"000000000",
  34107=>"111111111",
  34108=>"111111111",
  34109=>"011011111",
  34110=>"000000000",
  34111=>"110000000",
  34112=>"000000100",
  34113=>"110011000",
  34114=>"101101111",
  34115=>"100000111",
  34116=>"011111111",
  34117=>"111011001",
  34118=>"000010000",
  34119=>"001001101",
  34120=>"111111111",
  34121=>"000000000",
  34122=>"001001101",
  34123=>"001111111",
  34124=>"110111110",
  34125=>"000110110",
  34126=>"100111110",
  34127=>"111110111",
  34128=>"000001101",
  34129=>"001001101",
  34130=>"111111111",
  34131=>"000000000",
  34132=>"000000000",
  34133=>"011011011",
  34134=>"000010100",
  34135=>"101000000",
  34136=>"101100000",
  34137=>"000000000",
  34138=>"000000000",
  34139=>"111000000",
  34140=>"111111000",
  34141=>"000000101",
  34142=>"001111111",
  34143=>"100110110",
  34144=>"001000000",
  34145=>"111000000",
  34146=>"111010011",
  34147=>"111101100",
  34148=>"000010000",
  34149=>"000000000",
  34150=>"011010011",
  34151=>"000000000",
  34152=>"000000001",
  34153=>"010111111",
  34154=>"110111011",
  34155=>"000000110",
  34156=>"000000000",
  34157=>"000001111",
  34158=>"010110111",
  34159=>"101111110",
  34160=>"111111111",
  34161=>"000000001",
  34162=>"100110111",
  34163=>"000000000",
  34164=>"011111111",
  34165=>"111111111",
  34166=>"100100111",
  34167=>"011111000",
  34168=>"111111111",
  34169=>"111111000",
  34170=>"111111111",
  34171=>"011111111",
  34172=>"101100110",
  34173=>"111111111",
  34174=>"000000000",
  34175=>"111111111",
  34176=>"111111111",
  34177=>"110110010",
  34178=>"000001000",
  34179=>"111001000",
  34180=>"111111111",
  34181=>"000000000",
  34182=>"111100111",
  34183=>"000000111",
  34184=>"111100111",
  34185=>"000000010",
  34186=>"001011111",
  34187=>"111111111",
  34188=>"111111111",
  34189=>"000000000",
  34190=>"111001000",
  34191=>"000000000",
  34192=>"111111111",
  34193=>"000111000",
  34194=>"001001011",
  34195=>"111011001",
  34196=>"111101000",
  34197=>"000000000",
  34198=>"111111111",
  34199=>"010100000",
  34200=>"000001000",
  34201=>"111111111",
  34202=>"110110000",
  34203=>"001001000",
  34204=>"000000000",
  34205=>"000000000",
  34206=>"000000000",
  34207=>"000000111",
  34208=>"101111111",
  34209=>"001000001",
  34210=>"101000000",
  34211=>"111111111",
  34212=>"111111111",
  34213=>"000010000",
  34214=>"111110110",
  34215=>"111111111",
  34216=>"000000000",
  34217=>"000000000",
  34218=>"001001101",
  34219=>"000011000",
  34220=>"000000000",
  34221=>"111111111",
  34222=>"111001111",
  34223=>"110110111",
  34224=>"100000111",
  34225=>"111111111",
  34226=>"111111111",
  34227=>"000000111",
  34228=>"001011111",
  34229=>"000000000",
  34230=>"111111111",
  34231=>"111111111",
  34232=>"001111111",
  34233=>"000000000",
  34234=>"111111111",
  34235=>"101111111",
  34236=>"111000000",
  34237=>"111110110",
  34238=>"000000000",
  34239=>"110000000",
  34240=>"000000000",
  34241=>"011000000",
  34242=>"000000000",
  34243=>"111111111",
  34244=>"000000100",
  34245=>"000100001",
  34246=>"000000000",
  34247=>"000000111",
  34248=>"001000000",
  34249=>"100000000",
  34250=>"111111111",
  34251=>"111000000",
  34252=>"000011000",
  34253=>"000000000",
  34254=>"111111011",
  34255=>"000000111",
  34256=>"111111111",
  34257=>"111111010",
  34258=>"000000000",
  34259=>"111111110",
  34260=>"100000100",
  34261=>"001000001",
  34262=>"000001011",
  34263=>"011111111",
  34264=>"000001011",
  34265=>"110110111",
  34266=>"111000000",
  34267=>"111111111",
  34268=>"000000110",
  34269=>"111111111",
  34270=>"000110111",
  34271=>"000000010",
  34272=>"010000000",
  34273=>"000000100",
  34274=>"111111111",
  34275=>"111111111",
  34276=>"000100110",
  34277=>"111000000",
  34278=>"001000000",
  34279=>"111111111",
  34280=>"111000000",
  34281=>"111111000",
  34282=>"000000000",
  34283=>"011011011",
  34284=>"001001111",
  34285=>"000000000",
  34286=>"000000100",
  34287=>"100100110",
  34288=>"000000000",
  34289=>"111100000",
  34290=>"000010111",
  34291=>"000000011",
  34292=>"000000000",
  34293=>"000000000",
  34294=>"111111111",
  34295=>"100000000",
  34296=>"111111010",
  34297=>"000000000",
  34298=>"011000000",
  34299=>"000000000",
  34300=>"011001000",
  34301=>"101001001",
  34302=>"000000000",
  34303=>"100000010",
  34304=>"111111111",
  34305=>"000000000",
  34306=>"000000110",
  34307=>"111110110",
  34308=>"111001011",
  34309=>"011010111",
  34310=>"000000000",
  34311=>"111001111",
  34312=>"000000000",
  34313=>"011111010",
  34314=>"111111111",
  34315=>"010111111",
  34316=>"000100100",
  34317=>"101000000",
  34318=>"111011111",
  34319=>"000000001",
  34320=>"100100111",
  34321=>"000111111",
  34322=>"011001000",
  34323=>"111101111",
  34324=>"000000000",
  34325=>"000000001",
  34326=>"111111011",
  34327=>"011011000",
  34328=>"000000000",
  34329=>"011111111",
  34330=>"010000000",
  34331=>"111100110",
  34332=>"000000000",
  34333=>"111111111",
  34334=>"000000100",
  34335=>"000000000",
  34336=>"110100000",
  34337=>"000101101",
  34338=>"111111111",
  34339=>"111000111",
  34340=>"000011011",
  34341=>"000000000",
  34342=>"111111111",
  34343=>"000000000",
  34344=>"111111111",
  34345=>"111111111",
  34346=>"000000001",
  34347=>"100011000",
  34348=>"111111111",
  34349=>"111100000",
  34350=>"000000001",
  34351=>"010111111",
  34352=>"101101111",
  34353=>"010110010",
  34354=>"000000000",
  34355=>"000000000",
  34356=>"111111111",
  34357=>"001111111",
  34358=>"000000111",
  34359=>"110010000",
  34360=>"010010000",
  34361=>"000000111",
  34362=>"111011010",
  34363=>"000000000",
  34364=>"111111111",
  34365=>"011101111",
  34366=>"000100100",
  34367=>"111111111",
  34368=>"001000000",
  34369=>"000100111",
  34370=>"000000000",
  34371=>"001000000",
  34372=>"111110000",
  34373=>"101111110",
  34374=>"000000000",
  34375=>"000000100",
  34376=>"111111000",
  34377=>"111111011",
  34378=>"000000000",
  34379=>"011111111",
  34380=>"011011010",
  34381=>"000000000",
  34382=>"111111111",
  34383=>"000000000",
  34384=>"000000000",
  34385=>"111111111",
  34386=>"111111000",
  34387=>"001101101",
  34388=>"000000000",
  34389=>"000000000",
  34390=>"111111111",
  34391=>"111111001",
  34392=>"000000001",
  34393=>"111111010",
  34394=>"111111110",
  34395=>"000000000",
  34396=>"000000001",
  34397=>"111111111",
  34398=>"000000000",
  34399=>"010011010",
  34400=>"000000000",
  34401=>"111111010",
  34402=>"111111111",
  34403=>"000000000",
  34404=>"110111111",
  34405=>"000111111",
  34406=>"011111111",
  34407=>"111111111",
  34408=>"000111110",
  34409=>"110111111",
  34410=>"111111110",
  34411=>"111111111",
  34412=>"111111101",
  34413=>"111111000",
  34414=>"110111111",
  34415=>"100000000",
  34416=>"011000011",
  34417=>"001011000",
  34418=>"111111111",
  34419=>"111011011",
  34420=>"000001010",
  34421=>"000011011",
  34422=>"111100000",
  34423=>"000000000",
  34424=>"011011010",
  34425=>"001000000",
  34426=>"110000000",
  34427=>"000000000",
  34428=>"110110110",
  34429=>"111111101",
  34430=>"111100111",
  34431=>"111111111",
  34432=>"110011111",
  34433=>"001111111",
  34434=>"100111111",
  34435=>"101100100",
  34436=>"000101111",
  34437=>"111101111",
  34438=>"111111110",
  34439=>"000110000",
  34440=>"111111000",
  34441=>"000111111",
  34442=>"000000000",
  34443=>"001001001",
  34444=>"111001111",
  34445=>"000000000",
  34446=>"111110000",
  34447=>"011000000",
  34448=>"111111111",
  34449=>"000011111",
  34450=>"111111111",
  34451=>"110000000",
  34452=>"000000110",
  34453=>"111111111",
  34454=>"000000000",
  34455=>"000000000",
  34456=>"110110111",
  34457=>"000000000",
  34458=>"111111111",
  34459=>"000000000",
  34460=>"011010000",
  34461=>"010000010",
  34462=>"110100110",
  34463=>"000000000",
  34464=>"111011000",
  34465=>"001011010",
  34466=>"000010111",
  34467=>"000000000",
  34468=>"000111001",
  34469=>"111011000",
  34470=>"111111111",
  34471=>"111111111",
  34472=>"000101001",
  34473=>"000000111",
  34474=>"000010000",
  34475=>"111000000",
  34476=>"111111111",
  34477=>"111111111",
  34478=>"000000000",
  34479=>"100100011",
  34480=>"110111010",
  34481=>"000000000",
  34482=>"000111010",
  34483=>"111111000",
  34484=>"001000110",
  34485=>"000000111",
  34486=>"111111111",
  34487=>"000000000",
  34488=>"000001111",
  34489=>"111111111",
  34490=>"101011000",
  34491=>"111111111",
  34492=>"110111111",
  34493=>"010011111",
  34494=>"101000100",
  34495=>"111000001",
  34496=>"110000111",
  34497=>"111111111",
  34498=>"111100000",
  34499=>"000000011",
  34500=>"111111110",
  34501=>"000000000",
  34502=>"000001000",
  34503=>"111111111",
  34504=>"111111011",
  34505=>"011011000",
  34506=>"001000100",
  34507=>"110111000",
  34508=>"001000100",
  34509=>"010011001",
  34510=>"000000000",
  34511=>"000000000",
  34512=>"111111111",
  34513=>"111111111",
  34514=>"000000000",
  34515=>"000000000",
  34516=>"000001011",
  34517=>"000000000",
  34518=>"000111111",
  34519=>"111111111",
  34520=>"110110111",
  34521=>"000100111",
  34522=>"000000111",
  34523=>"110111111",
  34524=>"000000000",
  34525=>"000000000",
  34526=>"111111111",
  34527=>"111001000",
  34528=>"000000000",
  34529=>"000000011",
  34530=>"111000000",
  34531=>"100000000",
  34532=>"001101111",
  34533=>"000000000",
  34534=>"000000111",
  34535=>"011000110",
  34536=>"100000100",
  34537=>"111011111",
  34538=>"000000000",
  34539=>"000000111",
  34540=>"000000000",
  34541=>"000000000",
  34542=>"000000001",
  34543=>"000000000",
  34544=>"000000000",
  34545=>"111111111",
  34546=>"111111001",
  34547=>"001011011",
  34548=>"000000000",
  34549=>"100100000",
  34550=>"000000000",
  34551=>"111111111",
  34552=>"111011110",
  34553=>"001111111",
  34554=>"000000000",
  34555=>"000000000",
  34556=>"000001001",
  34557=>"111101110",
  34558=>"000011101",
  34559=>"011001001",
  34560=>"000001011",
  34561=>"000001000",
  34562=>"111111000",
  34563=>"000000000",
  34564=>"000001001",
  34565=>"111111111",
  34566=>"111111111",
  34567=>"001111101",
  34568=>"011000111",
  34569=>"010111111",
  34570=>"111100100",
  34571=>"111000000",
  34572=>"000000000",
  34573=>"000000000",
  34574=>"111111111",
  34575=>"001000000",
  34576=>"110111010",
  34577=>"000000000",
  34578=>"000000000",
  34579=>"010011010",
  34580=>"000000000",
  34581=>"000000010",
  34582=>"111111111",
  34583=>"111111111",
  34584=>"000000000",
  34585=>"110111111",
  34586=>"000000101",
  34587=>"011010000",
  34588=>"111111110",
  34589=>"111011001",
  34590=>"010010000",
  34591=>"111111111",
  34592=>"111111000",
  34593=>"000000001",
  34594=>"111111010",
  34595=>"111111111",
  34596=>"111110100",
  34597=>"111110111",
  34598=>"111010011",
  34599=>"001011000",
  34600=>"100100000",
  34601=>"111111111",
  34602=>"001010110",
  34603=>"000000111",
  34604=>"000000100",
  34605=>"001001000",
  34606=>"111110110",
  34607=>"000000001",
  34608=>"011111111",
  34609=>"111101101",
  34610=>"111111111",
  34611=>"110000111",
  34612=>"111111111",
  34613=>"000000000",
  34614=>"000000000",
  34615=>"000000011",
  34616=>"000000000",
  34617=>"000000000",
  34618=>"100000000",
  34619=>"111110000",
  34620=>"000000000",
  34621=>"011001011",
  34622=>"111111111",
  34623=>"000111000",
  34624=>"000011111",
  34625=>"000001111",
  34626=>"111111111",
  34627=>"000000000",
  34628=>"000101111",
  34629=>"010010011",
  34630=>"000000000",
  34631=>"001000000",
  34632=>"100101111",
  34633=>"000000000",
  34634=>"111000000",
  34635=>"011011101",
  34636=>"111111011",
  34637=>"111011000",
  34638=>"100001001",
  34639=>"111111011",
  34640=>"111111111",
  34641=>"111001000",
  34642=>"111100100",
  34643=>"111111111",
  34644=>"111011010",
  34645=>"001001001",
  34646=>"111111001",
  34647=>"111100111",
  34648=>"100101101",
  34649=>"111111111",
  34650=>"000000000",
  34651=>"000000000",
  34652=>"000000000",
  34653=>"000000000",
  34654=>"000000111",
  34655=>"000001111",
  34656=>"010000000",
  34657=>"000000001",
  34658=>"100000001",
  34659=>"111111111",
  34660=>"111111111",
  34661=>"011001000",
  34662=>"000000111",
  34663=>"111000000",
  34664=>"111111110",
  34665=>"111110111",
  34666=>"000000000",
  34667=>"001111111",
  34668=>"111111000",
  34669=>"001000000",
  34670=>"000000000",
  34671=>"000000111",
  34672=>"100111111",
  34673=>"000000000",
  34674=>"000111111",
  34675=>"100101001",
  34676=>"111000000",
  34677=>"001011111",
  34678=>"000000000",
  34679=>"000000111",
  34680=>"000000000",
  34681=>"011010000",
  34682=>"000000100",
  34683=>"001000000",
  34684=>"111000000",
  34685=>"111111111",
  34686=>"111111000",
  34687=>"100100111",
  34688=>"100100011",
  34689=>"111011111",
  34690=>"011001001",
  34691=>"000000000",
  34692=>"000000110",
  34693=>"000000111",
  34694=>"000001011",
  34695=>"111111111",
  34696=>"111111111",
  34697=>"111111111",
  34698=>"000000000",
  34699=>"000000000",
  34700=>"111111111",
  34701=>"101111011",
  34702=>"000011111",
  34703=>"000000000",
  34704=>"000001000",
  34705=>"111111111",
  34706=>"001001001",
  34707=>"000000001",
  34708=>"111101001",
  34709=>"000000000",
  34710=>"111111111",
  34711=>"000000000",
  34712=>"011000000",
  34713=>"010010110",
  34714=>"111111011",
  34715=>"001111111",
  34716=>"011111111",
  34717=>"000110110",
  34718=>"000011001",
  34719=>"111111111",
  34720=>"111111111",
  34721=>"111111000",
  34722=>"000000000",
  34723=>"011111111",
  34724=>"011111001",
  34725=>"000000000",
  34726=>"111111111",
  34727=>"010100111",
  34728=>"111110000",
  34729=>"100000000",
  34730=>"000000001",
  34731=>"000000001",
  34732=>"000000011",
  34733=>"000000000",
  34734=>"000011111",
  34735=>"101111111",
  34736=>"000000000",
  34737=>"011011001",
  34738=>"111111111",
  34739=>"000000011",
  34740=>"000011011",
  34741=>"111000000",
  34742=>"001011101",
  34743=>"110000111",
  34744=>"111111111",
  34745=>"000000000",
  34746=>"001011111",
  34747=>"001001000",
  34748=>"111111011",
  34749=>"000000000",
  34750=>"001000000",
  34751=>"001001011",
  34752=>"111111011",
  34753=>"000000000",
  34754=>"000000000",
  34755=>"111111111",
  34756=>"000000101",
  34757=>"001001111",
  34758=>"000011001",
  34759=>"111111111",
  34760=>"010000000",
  34761=>"111111111",
  34762=>"000000000",
  34763=>"000000000",
  34764=>"000100000",
  34765=>"000000000",
  34766=>"011111110",
  34767=>"000000000",
  34768=>"100100100",
  34769=>"111111111",
  34770=>"111111001",
  34771=>"110100100",
  34772=>"111001111",
  34773=>"000000000",
  34774=>"000000000",
  34775=>"000001111",
  34776=>"000000100",
  34777=>"111111111",
  34778=>"010000011",
  34779=>"000000000",
  34780=>"011011111",
  34781=>"001000000",
  34782=>"100110111",
  34783=>"100000000",
  34784=>"000000000",
  34785=>"111111111",
  34786=>"000000000",
  34787=>"000000000",
  34788=>"111111111",
  34789=>"000000000",
  34790=>"111110011",
  34791=>"111111111",
  34792=>"011000000",
  34793=>"001111111",
  34794=>"000000111",
  34795=>"100100000",
  34796=>"110110010",
  34797=>"101000000",
  34798=>"111111000",
  34799=>"111000110",
  34800=>"000000000",
  34801=>"000000000",
  34802=>"011111011",
  34803=>"000001000",
  34804=>"011110111",
  34805=>"000000001",
  34806=>"111111111",
  34807=>"000100101",
  34808=>"111111111",
  34809=>"001000101",
  34810=>"110110110",
  34811=>"001000000",
  34812=>"110100000",
  34813=>"111001111",
  34814=>"000000000",
  34815=>"111111111",
  34816=>"111011000",
  34817=>"010010110",
  34818=>"001111111",
  34819=>"111111000",
  34820=>"110111111",
  34821=>"110000000",
  34822=>"000000000",
  34823=>"111111111",
  34824=>"111100000",
  34825=>"000100110",
  34826=>"111001111",
  34827=>"000000000",
  34828=>"001011111",
  34829=>"111000000",
  34830=>"000100111",
  34831=>"100111101",
  34832=>"000011111",
  34833=>"010111111",
  34834=>"000000000",
  34835=>"000000000",
  34836=>"000000111",
  34837=>"111101000",
  34838=>"010110110",
  34839=>"100100101",
  34840=>"110111001",
  34841=>"011110110",
  34842=>"011000000",
  34843=>"000001001",
  34844=>"000011111",
  34845=>"111111111",
  34846=>"011011010",
  34847=>"011010011",
  34848=>"000000000",
  34849=>"100000000",
  34850=>"111111000",
  34851=>"111111111",
  34852=>"000000000",
  34853=>"000100111",
  34854=>"000000000",
  34855=>"111101011",
  34856=>"111111111",
  34857=>"000000100",
  34858=>"111111111",
  34859=>"011111111",
  34860=>"111111000",
  34861=>"001011011",
  34862=>"000000000",
  34863=>"111111000",
  34864=>"111111111",
  34865=>"000000000",
  34866=>"000000100",
  34867=>"011001111",
  34868=>"000000000",
  34869=>"110100111",
  34870=>"111111000",
  34871=>"001111111",
  34872=>"111111000",
  34873=>"000001111",
  34874=>"101000001",
  34875=>"011001000",
  34876=>"111000111",
  34877=>"111000111",
  34878=>"001011010",
  34879=>"111111111",
  34880=>"000000001",
  34881=>"000000100",
  34882=>"000000000",
  34883=>"100110100",
  34884=>"111111111",
  34885=>"111100110",
  34886=>"000000111",
  34887=>"111111111",
  34888=>"100110011",
  34889=>"001001111",
  34890=>"011111000",
  34891=>"000000110",
  34892=>"000000000",
  34893=>"000001111",
  34894=>"111000000",
  34895=>"000000001",
  34896=>"000110100",
  34897=>"111111001",
  34898=>"111111111",
  34899=>"000000011",
  34900=>"000000001",
  34901=>"000000000",
  34902=>"000000000",
  34903=>"111110100",
  34904=>"001111111",
  34905=>"111000011",
  34906=>"101111111",
  34907=>"100000011",
  34908=>"010000000",
  34909=>"000100111",
  34910=>"000000111",
  34911=>"100100100",
  34912=>"000111111",
  34913=>"111011001",
  34914=>"111111111",
  34915=>"111111010",
  34916=>"000000000",
  34917=>"000000000",
  34918=>"000000001",
  34919=>"110010111",
  34920=>"111111111",
  34921=>"000000111",
  34922=>"000000000",
  34923=>"000001111",
  34924=>"000110111",
  34925=>"000000000",
  34926=>"111000111",
  34927=>"010110111",
  34928=>"000010000",
  34929=>"000011011",
  34930=>"000000011",
  34931=>"111111110",
  34932=>"000000000",
  34933=>"001000100",
  34934=>"111111000",
  34935=>"000000000",
  34936=>"000000111",
  34937=>"010000011",
  34938=>"001000000",
  34939=>"110000000",
  34940=>"110011000",
  34941=>"101101001",
  34942=>"111000000",
  34943=>"111111000",
  34944=>"000000000",
  34945=>"110111111",
  34946=>"111000000",
  34947=>"010000111",
  34948=>"111110111",
  34949=>"111011000",
  34950=>"111111111",
  34951=>"100000000",
  34952=>"001111111",
  34953=>"000000000",
  34954=>"000000000",
  34955=>"000000110",
  34956=>"111111111",
  34957=>"111111001",
  34958=>"110010000",
  34959=>"000000000",
  34960=>"111111000",
  34961=>"000100111",
  34962=>"000000000",
  34963=>"000000011",
  34964=>"110111001",
  34965=>"101111111",
  34966=>"111000000",
  34967=>"111111111",
  34968=>"000000001",
  34969=>"111010000",
  34970=>"111110110",
  34971=>"100111111",
  34972=>"100100111",
  34973=>"010000010",
  34974=>"011000111",
  34975=>"000000000",
  34976=>"111111000",
  34977=>"101000000",
  34978=>"111000100",
  34979=>"111001000",
  34980=>"110111000",
  34981=>"111111011",
  34982=>"111111111",
  34983=>"111011011",
  34984=>"000000111",
  34985=>"000000000",
  34986=>"000000111",
  34987=>"000000000",
  34988=>"111000000",
  34989=>"111111000",
  34990=>"110000000",
  34991=>"101111000",
  34992=>"000001000",
  34993=>"111110110",
  34994=>"011111111",
  34995=>"111111000",
  34996=>"100101000",
  34997=>"111101000",
  34998=>"001000111",
  34999=>"000111110",
  35000=>"111111111",
  35001=>"111000000",
  35002=>"001111111",
  35003=>"001001001",
  35004=>"111000101",
  35005=>"001001000",
  35006=>"000000000",
  35007=>"111111110",
  35008=>"000110000",
  35009=>"000000111",
  35010=>"000000000",
  35011=>"101111111",
  35012=>"001000000",
  35013=>"000011011",
  35014=>"000000111",
  35015=>"000000101",
  35016=>"111110000",
  35017=>"000000111",
  35018=>"110110110",
  35019=>"000000100",
  35020=>"010000001",
  35021=>"000111000",
  35022=>"100100000",
  35023=>"000000001",
  35024=>"000000111",
  35025=>"111111111",
  35026=>"010011010",
  35027=>"100110111",
  35028=>"100111111",
  35029=>"100111111",
  35030=>"011111111",
  35031=>"111111111",
  35032=>"111000000",
  35033=>"111001000",
  35034=>"000000011",
  35035=>"111111110",
  35036=>"000000000",
  35037=>"110000000",
  35038=>"000000000",
  35039=>"111001011",
  35040=>"000000000",
  35041=>"000101111",
  35042=>"111111111",
  35043=>"111111111",
  35044=>"000000111",
  35045=>"000000000",
  35046=>"000000011",
  35047=>"000000110",
  35048=>"111011001",
  35049=>"011011011",
  35050=>"100001111",
  35051=>"000000111",
  35052=>"000000000",
  35053=>"000000000",
  35054=>"010000000",
  35055=>"001000000",
  35056=>"000000000",
  35057=>"000110111",
  35058=>"111111111",
  35059=>"101101111",
  35060=>"001000000",
  35061=>"111001001",
  35062=>"111111100",
  35063=>"111000111",
  35064=>"000000111",
  35065=>"010000000",
  35066=>"001000111",
  35067=>"111000000",
  35068=>"111100111",
  35069=>"001001011",
  35070=>"100101111",
  35071=>"111111111",
  35072=>"111000111",
  35073=>"000011111",
  35074=>"101110000",
  35075=>"000000000",
  35076=>"000000000",
  35077=>"111100100",
  35078=>"111111111",
  35079=>"000000001",
  35080=>"111111111",
  35081=>"111111111",
  35082=>"001000101",
  35083=>"000000000",
  35084=>"001001011",
  35085=>"001000111",
  35086=>"001000100",
  35087=>"011000000",
  35088=>"110111000",
  35089=>"100100100",
  35090=>"000001111",
  35091=>"000111111",
  35092=>"000000101",
  35093=>"000000111",
  35094=>"111110001",
  35095=>"000000001",
  35096=>"000100100",
  35097=>"110110010",
  35098=>"100000111",
  35099=>"000000000",
  35100=>"000000111",
  35101=>"111111111",
  35102=>"101011111",
  35103=>"110100101",
  35104=>"100111001",
  35105=>"000000000",
  35106=>"100100000",
  35107=>"111111000",
  35108=>"001111111",
  35109=>"000000100",
  35110=>"000000101",
  35111=>"000000111",
  35112=>"000000000",
  35113=>"000000110",
  35114=>"111001001",
  35115=>"000001111",
  35116=>"000000111",
  35117=>"011111000",
  35118=>"000000111",
  35119=>"000000000",
  35120=>"010011111",
  35121=>"000111111",
  35122=>"011111111",
  35123=>"000000110",
  35124=>"111001000",
  35125=>"000000110",
  35126=>"111100000",
  35127=>"000000000",
  35128=>"001111000",
  35129=>"111100000",
  35130=>"000000111",
  35131=>"000000000",
  35132=>"111111101",
  35133=>"111111011",
  35134=>"111111000",
  35135=>"011001001",
  35136=>"000000000",
  35137=>"110011001",
  35138=>"111111011",
  35139=>"000000000",
  35140=>"000000111",
  35141=>"000100111",
  35142=>"010111111",
  35143=>"011101101",
  35144=>"111111100",
  35145=>"111111000",
  35146=>"000110011",
  35147=>"010110111",
  35148=>"011001000",
  35149=>"100101111",
  35150=>"000000111",
  35151=>"000110111",
  35152=>"100000011",
  35153=>"001101111",
  35154=>"000000010",
  35155=>"100111111",
  35156=>"000111111",
  35157=>"001000100",
  35158=>"000000000",
  35159=>"000000110",
  35160=>"111100001",
  35161=>"111000111",
  35162=>"000001000",
  35163=>"111111111",
  35164=>"001001111",
  35165=>"101111110",
  35166=>"001000000",
  35167=>"000101111",
  35168=>"001000000",
  35169=>"111111111",
  35170=>"111111001",
  35171=>"000000001",
  35172=>"001001100",
  35173=>"000111111",
  35174=>"111110100",
  35175=>"010001001",
  35176=>"011001011",
  35177=>"000010000",
  35178=>"000000000",
  35179=>"111000000",
  35180=>"001011011",
  35181=>"111101000",
  35182=>"111010011",
  35183=>"000100110",
  35184=>"111111111",
  35185=>"000000000",
  35186=>"111111010",
  35187=>"000110000",
  35188=>"111111111",
  35189=>"111111111",
  35190=>"000000000",
  35191=>"111111111",
  35192=>"000000000",
  35193=>"111111111",
  35194=>"111000000",
  35195=>"100000100",
  35196=>"111111111",
  35197=>"110011000",
  35198=>"111000010",
  35199=>"111010000",
  35200=>"001000000",
  35201=>"111110000",
  35202=>"111111001",
  35203=>"000000000",
  35204=>"000000000",
  35205=>"111010000",
  35206=>"110000000",
  35207=>"001000000",
  35208=>"111000000",
  35209=>"111111111",
  35210=>"100000000",
  35211=>"011111111",
  35212=>"111111111",
  35213=>"000000001",
  35214=>"111111111",
  35215=>"000001000",
  35216=>"111111110",
  35217=>"110000000",
  35218=>"111010000",
  35219=>"111111111",
  35220=>"111000000",
  35221=>"011110000",
  35222=>"000000100",
  35223=>"100000101",
  35224=>"111111000",
  35225=>"000000000",
  35226=>"111000000",
  35227=>"000100111",
  35228=>"110000100",
  35229=>"111000010",
  35230=>"010100111",
  35231=>"000000111",
  35232=>"111101001",
  35233=>"100111111",
  35234=>"001010111",
  35235=>"111111111",
  35236=>"000110111",
  35237=>"101111111",
  35238=>"000100000",
  35239=>"111111111",
  35240=>"011110000",
  35241=>"011101101",
  35242=>"111011001",
  35243=>"110100111",
  35244=>"010110111",
  35245=>"111111000",
  35246=>"000011111",
  35247=>"111100000",
  35248=>"111111000",
  35249=>"111100110",
  35250=>"111000101",
  35251=>"101111000",
  35252=>"000101111",
  35253=>"101011111",
  35254=>"111111111",
  35255=>"001000000",
  35256=>"111111000",
  35257=>"000000111",
  35258=>"100100101",
  35259=>"100000000",
  35260=>"111101111",
  35261=>"000110111",
  35262=>"001001000",
  35263=>"001011011",
  35264=>"100111111",
  35265=>"001000000",
  35266=>"111111111",
  35267=>"110100000",
  35268=>"100000111",
  35269=>"110111011",
  35270=>"011011011",
  35271=>"000001011",
  35272=>"011011111",
  35273=>"000101111",
  35274=>"000000000",
  35275=>"100111101",
  35276=>"111000000",
  35277=>"010111011",
  35278=>"011010000",
  35279=>"000000000",
  35280=>"000000010",
  35281=>"111111111",
  35282=>"000011011",
  35283=>"110000111",
  35284=>"011111110",
  35285=>"000001111",
  35286=>"000011111",
  35287=>"000000011",
  35288=>"000000000",
  35289=>"110010111",
  35290=>"000000111",
  35291=>"111111111",
  35292=>"100001001",
  35293=>"000000111",
  35294=>"000000000",
  35295=>"011011011",
  35296=>"000000000",
  35297=>"000010111",
  35298=>"000001101",
  35299=>"000000110",
  35300=>"100110111",
  35301=>"110000000",
  35302=>"111011000",
  35303=>"100100100",
  35304=>"000010000",
  35305=>"111111111",
  35306=>"000000100",
  35307=>"000000011",
  35308=>"000000111",
  35309=>"111111000",
  35310=>"110111111",
  35311=>"000011011",
  35312=>"000000100",
  35313=>"110000000",
  35314=>"111100000",
  35315=>"000000011",
  35316=>"111000000",
  35317=>"000000000",
  35318=>"000000100",
  35319=>"000011111",
  35320=>"000000111",
  35321=>"111000000",
  35322=>"111100100",
  35323=>"111111000",
  35324=>"000000001",
  35325=>"111111101",
  35326=>"000000001",
  35327=>"000100000",
  35328=>"001001000",
  35329=>"111111111",
  35330=>"111111111",
  35331=>"010011011",
  35332=>"000100000",
  35333=>"110011001",
  35334=>"100100111",
  35335=>"111111111",
  35336=>"111111011",
  35337=>"000001000",
  35338=>"111111111",
  35339=>"110000001",
  35340=>"011111010",
  35341=>"000000000",
  35342=>"100111110",
  35343=>"000000000",
  35344=>"110110110",
  35345=>"111111110",
  35346=>"000000000",
  35347=>"111111111",
  35348=>"000000000",
  35349=>"000000000",
  35350=>"111111111",
  35351=>"000000000",
  35352=>"001111111",
  35353=>"110011111",
  35354=>"000000011",
  35355=>"111111100",
  35356=>"110000000",
  35357=>"000100101",
  35358=>"111111110",
  35359=>"000110010",
  35360=>"111110000",
  35361=>"111111111",
  35362=>"000000110",
  35363=>"000000100",
  35364=>"000111111",
  35365=>"111100000",
  35366=>"000000000",
  35367=>"001111111",
  35368=>"000000000",
  35369=>"011101000",
  35370=>"000000000",
  35371=>"011111111",
  35372=>"101111010",
  35373=>"111111111",
  35374=>"111111111",
  35375=>"111111111",
  35376=>"110110000",
  35377=>"000000100",
  35378=>"111111100",
  35379=>"010110110",
  35380=>"001011100",
  35381=>"001001001",
  35382=>"000000000",
  35383=>"110101001",
  35384=>"110011010",
  35385=>"100000111",
  35386=>"000000101",
  35387=>"000000110",
  35388=>"111111110",
  35389=>"100000000",
  35390=>"000000110",
  35391=>"111111001",
  35392=>"110110000",
  35393=>"000001000",
  35394=>"000000000",
  35395=>"000000000",
  35396=>"000000000",
  35397=>"000000000",
  35398=>"001000101",
  35399=>"101101000",
  35400=>"111111000",
  35401=>"000000100",
  35402=>"100000000",
  35403=>"111111111",
  35404=>"011111111",
  35405=>"100111111",
  35406=>"110110111",
  35407=>"011001000",
  35408=>"001001000",
  35409=>"000000000",
  35410=>"010111011",
  35411=>"001011011",
  35412=>"111111001",
  35413=>"000000000",
  35414=>"110100000",
  35415=>"001000000",
  35416=>"000000000",
  35417=>"001000000",
  35418=>"000000000",
  35419=>"000000000",
  35420=>"110000111",
  35421=>"000110000",
  35422=>"111001001",
  35423=>"111101000",
  35424=>"111011011",
  35425=>"000100110",
  35426=>"000010110",
  35427=>"000000111",
  35428=>"111111111",
  35429=>"111111110",
  35430=>"111001001",
  35431=>"101100100",
  35432=>"011111111",
  35433=>"000111111",
  35434=>"110111111",
  35435=>"000000000",
  35436=>"001001111",
  35437=>"110110110",
  35438=>"111111111",
  35439=>"110100000",
  35440=>"111111000",
  35441=>"000001111",
  35442=>"000000000",
  35443=>"000000000",
  35444=>"100000111",
  35445=>"000001000",
  35446=>"000000000",
  35447=>"110111001",
  35448=>"000010000",
  35449=>"000000000",
  35450=>"000000110",
  35451=>"000000000",
  35452=>"110000000",
  35453=>"001000000",
  35454=>"000100111",
  35455=>"111111111",
  35456=>"111111110",
  35457=>"010000000",
  35458=>"111000000",
  35459=>"011110100",
  35460=>"000000000",
  35461=>"000000001",
  35462=>"000000001",
  35463=>"000000000",
  35464=>"111010111",
  35465=>"000000000",
  35466=>"110110111",
  35467=>"011111001",
  35468=>"110000000",
  35469=>"000000000",
  35470=>"110111111",
  35471=>"000100101",
  35472=>"100000000",
  35473=>"111111111",
  35474=>"110111111",
  35475=>"111111111",
  35476=>"000000000",
  35477=>"111111111",
  35478=>"000000000",
  35479=>"111111111",
  35480=>"100110011",
  35481=>"000000100",
  35482=>"000100000",
  35483=>"100101001",
  35484=>"000000000",
  35485=>"110110111",
  35486=>"111001001",
  35487=>"111111111",
  35488=>"000000000",
  35489=>"110111111",
  35490=>"110000000",
  35491=>"111111111",
  35492=>"000000001",
  35493=>"101111111",
  35494=>"000111011",
  35495=>"001011000",
  35496=>"100111001",
  35497=>"000000100",
  35498=>"001000000",
  35499=>"111111100",
  35500=>"001000000",
  35501=>"100000100",
  35502=>"111111111",
  35503=>"110110111",
  35504=>"000000000",
  35505=>"111111111",
  35506=>"010111110",
  35507=>"010111111",
  35508=>"110000000",
  35509=>"111111110",
  35510=>"000000000",
  35511=>"000000000",
  35512=>"000000000",
  35513=>"111111111",
  35514=>"000000000",
  35515=>"011011001",
  35516=>"110011000",
  35517=>"111001111",
  35518=>"000000000",
  35519=>"000010010",
  35520=>"110010011",
  35521=>"111111001",
  35522=>"000011001",
  35523=>"110111111",
  35524=>"101000000",
  35525=>"000101100",
  35526=>"001101101",
  35527=>"101111111",
  35528=>"111111000",
  35529=>"111111111",
  35530=>"111101101",
  35531=>"000000000",
  35532=>"111111111",
  35533=>"000111111",
  35534=>"100100010",
  35535=>"100000000",
  35536=>"111111000",
  35537=>"010000000",
  35538=>"111111101",
  35539=>"111111110",
  35540=>"111100000",
  35541=>"000001111",
  35542=>"110000000",
  35543=>"101101111",
  35544=>"111111111",
  35545=>"000000000",
  35546=>"000000011",
  35547=>"111111111",
  35548=>"111111111",
  35549=>"111011111",
  35550=>"000111111",
  35551=>"100101000",
  35552=>"111111111",
  35553=>"011011110",
  35554=>"000000000",
  35555=>"000000100",
  35556=>"000000000",
  35557=>"000000000",
  35558=>"110110111",
  35559=>"010100100",
  35560=>"000001001",
  35561=>"000000111",
  35562=>"000000011",
  35563=>"111111000",
  35564=>"111011000",
  35565=>"110111010",
  35566=>"011010010",
  35567=>"111111100",
  35568=>"010000001",
  35569=>"111100000",
  35570=>"000110110",
  35571=>"010101111",
  35572=>"101000111",
  35573=>"110111000",
  35574=>"110000000",
  35575=>"000000000",
  35576=>"000000000",
  35577=>"000000000",
  35578=>"110111111",
  35579=>"001110000",
  35580=>"000000000",
  35581=>"111111011",
  35582=>"000000000",
  35583=>"100100100",
  35584=>"000000111",
  35585=>"111111011",
  35586=>"000000000",
  35587=>"001001001",
  35588=>"110110111",
  35589=>"111011111",
  35590=>"000110110",
  35591=>"111111001",
  35592=>"110110111",
  35593=>"111000111",
  35594=>"000100000",
  35595=>"111000110",
  35596=>"100100110",
  35597=>"000000001",
  35598=>"000001000",
  35599=>"001011000",
  35600=>"100100100",
  35601=>"111101111",
  35602=>"111110000",
  35603=>"111111111",
  35604=>"101100110",
  35605=>"110010011",
  35606=>"111111111",
  35607=>"000000001",
  35608=>"001001011",
  35609=>"111111011",
  35610=>"111111111",
  35611=>"000000000",
  35612=>"111111111",
  35613=>"111110000",
  35614=>"111111111",
  35615=>"111111000",
  35616=>"110111111",
  35617=>"000000000",
  35618=>"111011000",
  35619=>"000000000",
  35620=>"111111111",
  35621=>"000011111",
  35622=>"111111111",
  35623=>"000111111",
  35624=>"111111111",
  35625=>"000000000",
  35626=>"101111111",
  35627=>"001001000",
  35628=>"111111111",
  35629=>"000000001",
  35630=>"111111000",
  35631=>"111101111",
  35632=>"001001001",
  35633=>"111011001",
  35634=>"000000000",
  35635=>"000100111",
  35636=>"000100000",
  35637=>"000000111",
  35638=>"000000000",
  35639=>"010010000",
  35640=>"001011011",
  35641=>"011011000",
  35642=>"111100111",
  35643=>"000000000",
  35644=>"000000001",
  35645=>"000000000",
  35646=>"111111111",
  35647=>"111111100",
  35648=>"111111111",
  35649=>"111111111",
  35650=>"111111111",
  35651=>"000000000",
  35652=>"100110111",
  35653=>"111010010",
  35654=>"111110110",
  35655=>"111111111",
  35656=>"000000000",
  35657=>"001000000",
  35658=>"100000000",
  35659=>"000000000",
  35660=>"011000000",
  35661=>"000000010",
  35662=>"111110000",
  35663=>"011111111",
  35664=>"000000000",
  35665=>"111111111",
  35666=>"000000000",
  35667=>"000000000",
  35668=>"000000000",
  35669=>"111110110",
  35670=>"000000000",
  35671=>"100000000",
  35672=>"100100100",
  35673=>"000100000",
  35674=>"100100011",
  35675=>"000111111",
  35676=>"111111111",
  35677=>"111111111",
  35678=>"000000001",
  35679=>"000000000",
  35680=>"111111111",
  35681=>"000000000",
  35682=>"110111111",
  35683=>"000100000",
  35684=>"111111111",
  35685=>"000000000",
  35686=>"111111111",
  35687=>"000000001",
  35688=>"000000000",
  35689=>"111000000",
  35690=>"111111001",
  35691=>"000010010",
  35692=>"000001001",
  35693=>"000000000",
  35694=>"000000000",
  35695=>"111000000",
  35696=>"111111111",
  35697=>"111111111",
  35698=>"000000010",
  35699=>"011000100",
  35700=>"100110100",
  35701=>"000000101",
  35702=>"110010000",
  35703=>"000000110",
  35704=>"111111110",
  35705=>"000010110",
  35706=>"111111111",
  35707=>"001111101",
  35708=>"011001000",
  35709=>"111111000",
  35710=>"000100000",
  35711=>"000000000",
  35712=>"000000000",
  35713=>"000000000",
  35714=>"000000000",
  35715=>"000100101",
  35716=>"100111111",
  35717=>"111110111",
  35718=>"111111111",
  35719=>"000111110",
  35720=>"000000000",
  35721=>"111101100",
  35722=>"001001001",
  35723=>"000000000",
  35724=>"101000000",
  35725=>"111110110",
  35726=>"000000000",
  35727=>"110010000",
  35728=>"000000000",
  35729=>"100000000",
  35730=>"000000000",
  35731=>"110110100",
  35732=>"000111111",
  35733=>"000111111",
  35734=>"000000000",
  35735=>"101001100",
  35736=>"111111111",
  35737=>"000000000",
  35738=>"000000000",
  35739=>"000000110",
  35740=>"000000000",
  35741=>"011100000",
  35742=>"000000000",
  35743=>"000000001",
  35744=>"111100111",
  35745=>"110110000",
  35746=>"111101111",
  35747=>"111111111",
  35748=>"111111001",
  35749=>"001011000",
  35750=>"000000000",
  35751=>"111111111",
  35752=>"000111011",
  35753=>"011001110",
  35754=>"000000000",
  35755=>"000000011",
  35756=>"000000000",
  35757=>"110110000",
  35758=>"111111100",
  35759=>"000000000",
  35760=>"000000000",
  35761=>"000111101",
  35762=>"000000000",
  35763=>"000000000",
  35764=>"010110110",
  35765=>"000001000",
  35766=>"000000000",
  35767=>"111011000",
  35768=>"000001000",
  35769=>"111111001",
  35770=>"111000000",
  35771=>"111111111",
  35772=>"111111011",
  35773=>"111111111",
  35774=>"010111111",
  35775=>"111111111",
  35776=>"110111111",
  35777=>"111111111",
  35778=>"111100000",
  35779=>"111111001",
  35780=>"111111111",
  35781=>"111111111",
  35782=>"000000111",
  35783=>"111111111",
  35784=>"000000000",
  35785=>"100110100",
  35786=>"000000000",
  35787=>"111111000",
  35788=>"011010000",
  35789=>"111111111",
  35790=>"000101001",
  35791=>"100100000",
  35792=>"111001111",
  35793=>"111110000",
  35794=>"111111111",
  35795=>"110110111",
  35796=>"000000000",
  35797=>"001101111",
  35798=>"111111000",
  35799=>"100000001",
  35800=>"111111111",
  35801=>"111111111",
  35802=>"000000000",
  35803=>"101001000",
  35804=>"000001001",
  35805=>"000000000",
  35806=>"000000100",
  35807=>"000000001",
  35808=>"111111111",
  35809=>"111111111",
  35810=>"000000000",
  35811=>"110101100",
  35812=>"111110111",
  35813=>"111111110",
  35814=>"000001000",
  35815=>"000000000",
  35816=>"100000000",
  35817=>"010011010",
  35818=>"111110100",
  35819=>"000001111",
  35820=>"000100111",
  35821=>"011011111",
  35822=>"111111000",
  35823=>"000000000",
  35824=>"111000111",
  35825=>"000110001",
  35826=>"011111000",
  35827=>"111001000",
  35828=>"000100111",
  35829=>"101111111",
  35830=>"111101111",
  35831=>"000000100",
  35832=>"110001001",
  35833=>"111111111",
  35834=>"111101111",
  35835=>"011111011",
  35836=>"011000001",
  35837=>"100110000",
  35838=>"000000000",
  35839=>"000000000",
  35840=>"000000000",
  35841=>"000000000",
  35842=>"000100111",
  35843=>"011011011",
  35844=>"000000111",
  35845=>"111011101",
  35846=>"000000000",
  35847=>"000000111",
  35848=>"000000111",
  35849=>"011111111",
  35850=>"111111111",
  35851=>"111100000",
  35852=>"000110111",
  35853=>"101001001",
  35854=>"110111100",
  35855=>"000001111",
  35856=>"111100111",
  35857=>"000111111",
  35858=>"000000100",
  35859=>"111111111",
  35860=>"000000000",
  35861=>"000101111",
  35862=>"011111110",
  35863=>"010010001",
  35864=>"100100111",
  35865=>"111101001",
  35866=>"000000000",
  35867=>"111001100",
  35868=>"000000000",
  35869=>"100100101",
  35870=>"000101111",
  35871=>"000110111",
  35872=>"000000000",
  35873=>"111100000",
  35874=>"111111111",
  35875=>"000000000",
  35876=>"000000000",
  35877=>"111111111",
  35878=>"000000111",
  35879=>"000001111",
  35880=>"000000000",
  35881=>"000000000",
  35882=>"000000000",
  35883=>"111110100",
  35884=>"000000101",
  35885=>"100111111",
  35886=>"111111111",
  35887=>"111100100",
  35888=>"111111111",
  35889=>"000000000",
  35890=>"110110100",
  35891=>"010011000",
  35892=>"011111111",
  35893=>"110110110",
  35894=>"011000000",
  35895=>"111111111",
  35896=>"111111000",
  35897=>"111111111",
  35898=>"111111001",
  35899=>"111101000",
  35900=>"111100000",
  35901=>"000000000",
  35902=>"000000011",
  35903=>"100110110",
  35904=>"011000000",
  35905=>"011010000",
  35906=>"111001110",
  35907=>"100100100",
  35908=>"111101111",
  35909=>"011111000",
  35910=>"101000001",
  35911=>"111111111",
  35912=>"111110101",
  35913=>"011111111",
  35914=>"001000000",
  35915=>"000000111",
  35916=>"010111111",
  35917=>"000111111",
  35918=>"111001111",
  35919=>"111101000",
  35920=>"111111111",
  35921=>"000001000",
  35922=>"111111000",
  35923=>"000000000",
  35924=>"111111000",
  35925=>"010111110",
  35926=>"111100000",
  35927=>"111100000",
  35928=>"001011111",
  35929=>"111000000",
  35930=>"111111111",
  35931=>"100000100",
  35932=>"000000000",
  35933=>"000000000",
  35934=>"000000100",
  35935=>"010000000",
  35936=>"000000000",
  35937=>"000000001",
  35938=>"011111100",
  35939=>"000000000",
  35940=>"000000000",
  35941=>"111010010",
  35942=>"111111001",
  35943=>"111111111",
  35944=>"000000000",
  35945=>"000000111",
  35946=>"111100111",
  35947=>"000001101",
  35948=>"000000111",
  35949=>"011111111",
  35950=>"111000000",
  35951=>"001001011",
  35952=>"111011001",
  35953=>"000000000",
  35954=>"011001001",
  35955=>"000010000",
  35956=>"011000010",
  35957=>"111111111",
  35958=>"000000000",
  35959=>"100000000",
  35960=>"111111011",
  35961=>"110110111",
  35962=>"111111100",
  35963=>"000000000",
  35964=>"100100100",
  35965=>"001000000",
  35966=>"001000000",
  35967=>"111011111",
  35968=>"000000011",
  35969=>"111111111",
  35970=>"111011011",
  35971=>"000100100",
  35972=>"111111111",
  35973=>"111111111",
  35974=>"000110111",
  35975=>"000111111",
  35976=>"101111111",
  35977=>"111100000",
  35978=>"000000100",
  35979=>"000100111",
  35980=>"001111111",
  35981=>"111111111",
  35982=>"100100100",
  35983=>"001001001",
  35984=>"111111110",
  35985=>"111011011",
  35986=>"110111110",
  35987=>"110000100",
  35988=>"111111101",
  35989=>"101101111",
  35990=>"111111000",
  35991=>"111110111",
  35992=>"011111010",
  35993=>"111011011",
  35994=>"111100100",
  35995=>"111000101",
  35996=>"000000000",
  35997=>"100000000",
  35998=>"111111111",
  35999=>"111000000",
  36000=>"111000000",
  36001=>"111111000",
  36002=>"111111111",
  36003=>"001111111",
  36004=>"000000000",
  36005=>"111110111",
  36006=>"110110001",
  36007=>"001001001",
  36008=>"000000001",
  36009=>"000000000",
  36010=>"111100000",
  36011=>"000000101",
  36012=>"111111011",
  36013=>"111100001",
  36014=>"110111111",
  36015=>"001000000",
  36016=>"000000000",
  36017=>"100111111",
  36018=>"010111111",
  36019=>"000000000",
  36020=>"000000000",
  36021=>"000000000",
  36022=>"000000000",
  36023=>"111111110",
  36024=>"111111111",
  36025=>"011000000",
  36026=>"000111111",
  36027=>"000000001",
  36028=>"101000000",
  36029=>"000001111",
  36030=>"001000001",
  36031=>"000000010",
  36032=>"000000011",
  36033=>"111111000",
  36034=>"001001011",
  36035=>"111111000",
  36036=>"111110111",
  36037=>"001111111",
  36038=>"000100111",
  36039=>"000000011",
  36040=>"001001001",
  36041=>"100101011",
  36042=>"110110100",
  36043=>"000000000",
  36044=>"100000001",
  36045=>"111111111",
  36046=>"111111100",
  36047=>"101111001",
  36048=>"001111111",
  36049=>"000000000",
  36050=>"100000000",
  36051=>"111110000",
  36052=>"111111001",
  36053=>"111111111",
  36054=>"000000000",
  36055=>"111111011",
  36056=>"111111110",
  36057=>"100110111",
  36058=>"000000000",
  36059=>"000000000",
  36060=>"000000101",
  36061=>"100011101",
  36062=>"111111111",
  36063=>"100000000",
  36064=>"000000000",
  36065=>"000111111",
  36066=>"000000000",
  36067=>"000101101",
  36068=>"000011000",
  36069=>"000000100",
  36070=>"111101111",
  36071=>"111111101",
  36072=>"110111111",
  36073=>"110110110",
  36074=>"000111111",
  36075=>"111110000",
  36076=>"001000000",
  36077=>"111000101",
  36078=>"000010110",
  36079=>"100000101",
  36080=>"001000100",
  36081=>"111111111",
  36082=>"111111111",
  36083=>"000000000",
  36084=>"101000101",
  36085=>"110000001",
  36086=>"010011100",
  36087=>"000000111",
  36088=>"111111111",
  36089=>"100110110",
  36090=>"000100001",
  36091=>"000000000",
  36092=>"011001000",
  36093=>"000011111",
  36094=>"000111111",
  36095=>"000000001",
  36096=>"000000111",
  36097=>"101101101",
  36098=>"110100000",
  36099=>"111111101",
  36100=>"001011001",
  36101=>"000011000",
  36102=>"111111111",
  36103=>"101100100",
  36104=>"011100111",
  36105=>"001011011",
  36106=>"011000100",
  36107=>"011111111",
  36108=>"100100000",
  36109=>"111111111",
  36110=>"000100000",
  36111=>"011111000",
  36112=>"100100111",
  36113=>"001111100",
  36114=>"111111000",
  36115=>"000110111",
  36116=>"000000001",
  36117=>"000011111",
  36118=>"111111111",
  36119=>"001001111",
  36120=>"010010000",
  36121=>"000000100",
  36122=>"111000000",
  36123=>"000000111",
  36124=>"011111111",
  36125=>"000110111",
  36126=>"000000000",
  36127=>"000000111",
  36128=>"110100111",
  36129=>"111010110",
  36130=>"011000000",
  36131=>"001000000",
  36132=>"110000000",
  36133=>"111100101",
  36134=>"000010110",
  36135=>"000000110",
  36136=>"000000000",
  36137=>"111111111",
  36138=>"101110000",
  36139=>"000000000",
  36140=>"111000000",
  36141=>"001001110",
  36142=>"000111111",
  36143=>"111000000",
  36144=>"000001101",
  36145=>"100000000",
  36146=>"111111000",
  36147=>"000111111",
  36148=>"111101001",
  36149=>"111111101",
  36150=>"010000000",
  36151=>"111111111",
  36152=>"011011001",
  36153=>"111000000",
  36154=>"101001000",
  36155=>"000000000",
  36156=>"100000001",
  36157=>"000000000",
  36158=>"000000000",
  36159=>"100000000",
  36160=>"000000001",
  36161=>"111111111",
  36162=>"111011010",
  36163=>"001000011",
  36164=>"011100111",
  36165=>"001111111",
  36166=>"000101111",
  36167=>"000000000",
  36168=>"001111111",
  36169=>"000111111",
  36170=>"010000000",
  36171=>"000000110",
  36172=>"001000000",
  36173=>"110000000",
  36174=>"111110111",
  36175=>"110110000",
  36176=>"111110000",
  36177=>"011111110",
  36178=>"001000111",
  36179=>"000000000",
  36180=>"000111111",
  36181=>"000001001",
  36182=>"111000010",
  36183=>"000000000",
  36184=>"000000100",
  36185=>"000000111",
  36186=>"111111100",
  36187=>"001111111",
  36188=>"101111111",
  36189=>"011011111",
  36190=>"001101000",
  36191=>"111111001",
  36192=>"000010011",
  36193=>"000111111",
  36194=>"011011111",
  36195=>"101000001",
  36196=>"111111110",
  36197=>"100111001",
  36198=>"000011111",
  36199=>"111101111",
  36200=>"001000110",
  36201=>"110000000",
  36202=>"001001011",
  36203=>"000000010",
  36204=>"010110111",
  36205=>"011111111",
  36206=>"000000000",
  36207=>"110110000",
  36208=>"011001000",
  36209=>"000111111",
  36210=>"000000111",
  36211=>"000111001",
  36212=>"111011000",
  36213=>"011111111",
  36214=>"000000000",
  36215=>"000001111",
  36216=>"000000000",
  36217=>"000100000",
  36218=>"110110111",
  36219=>"111000000",
  36220=>"111011111",
  36221=>"100101111",
  36222=>"000111011",
  36223=>"100010000",
  36224=>"111100110",
  36225=>"000010011",
  36226=>"110010000",
  36227=>"000011111",
  36228=>"000000000",
  36229=>"111111011",
  36230=>"000000000",
  36231=>"000000000",
  36232=>"000010000",
  36233=>"111111111",
  36234=>"000000111",
  36235=>"011011011",
  36236=>"111111111",
  36237=>"100101111",
  36238=>"000001111",
  36239=>"000000001",
  36240=>"111111111",
  36241=>"111001101",
  36242=>"111111000",
  36243=>"000000100",
  36244=>"111111111",
  36245=>"000001001",
  36246=>"000000000",
  36247=>"000000100",
  36248=>"001011100",
  36249=>"000110011",
  36250=>"111000000",
  36251=>"100100111",
  36252=>"111001001",
  36253=>"000000010",
  36254=>"011000001",
  36255=>"101000000",
  36256=>"000001011",
  36257=>"000100110",
  36258=>"001000000",
  36259=>"000111001",
  36260=>"000000101",
  36261=>"101111111",
  36262=>"000000000",
  36263=>"111110010",
  36264=>"011011111",
  36265=>"111111111",
  36266=>"111100111",
  36267=>"000000100",
  36268=>"000000000",
  36269=>"111111011",
  36270=>"000000111",
  36271=>"000000111",
  36272=>"100000000",
  36273=>"110110111",
  36274=>"101101111",
  36275=>"111111111",
  36276=>"011011111",
  36277=>"000000000",
  36278=>"000000111",
  36279=>"111111111",
  36280=>"111111000",
  36281=>"100000100",
  36282=>"000000001",
  36283=>"111111111",
  36284=>"111111000",
  36285=>"100100000",
  36286=>"111111111",
  36287=>"111111001",
  36288=>"000000000",
  36289=>"010000111",
  36290=>"111010111",
  36291=>"001001000",
  36292=>"001101110",
  36293=>"000010100",
  36294=>"110100000",
  36295=>"000111011",
  36296=>"101000000",
  36297=>"001000000",
  36298=>"000000000",
  36299=>"111111000",
  36300=>"110000000",
  36301=>"000000001",
  36302=>"111110000",
  36303=>"001000000",
  36304=>"011001000",
  36305=>"011001011",
  36306=>"101111111",
  36307=>"000000000",
  36308=>"111000101",
  36309=>"000001111",
  36310=>"000000111",
  36311=>"101111111",
  36312=>"000000111",
  36313=>"111101000",
  36314=>"000111111",
  36315=>"000000001",
  36316=>"111111110",
  36317=>"001001000",
  36318=>"111111000",
  36319=>"101001011",
  36320=>"000010011",
  36321=>"111011000",
  36322=>"000000000",
  36323=>"001001001",
  36324=>"000000000",
  36325=>"001110110",
  36326=>"011001010",
  36327=>"000000000",
  36328=>"110000011",
  36329=>"000001000",
  36330=>"001000101",
  36331=>"010111111",
  36332=>"111100111",
  36333=>"011011000",
  36334=>"111111000",
  36335=>"111100100",
  36336=>"000000000",
  36337=>"111000000",
  36338=>"111100000",
  36339=>"000000000",
  36340=>"101110111",
  36341=>"111111000",
  36342=>"000000111",
  36343=>"100100000",
  36344=>"001111011",
  36345=>"101100100",
  36346=>"100000000",
  36347=>"111110110",
  36348=>"111111100",
  36349=>"111100001",
  36350=>"111000000",
  36351=>"110100100",
  36352=>"001001000",
  36353=>"111110101",
  36354=>"001111111",
  36355=>"111111001",
  36356=>"110000100",
  36357=>"100000000",
  36358=>"111001000",
  36359=>"111111111",
  36360=>"001001111",
  36361=>"000000000",
  36362=>"101001111",
  36363=>"000000000",
  36364=>"110110000",
  36365=>"010100100",
  36366=>"000001001",
  36367=>"110000100",
  36368=>"000111000",
  36369=>"111011000",
  36370=>"111111111",
  36371=>"000000111",
  36372=>"000000100",
  36373=>"000110110",
  36374=>"111111000",
  36375=>"001001000",
  36376=>"110111001",
  36377=>"111111111",
  36378=>"000111111",
  36379=>"000011000",
  36380=>"111101000",
  36381=>"111100100",
  36382=>"110100101",
  36383=>"000000111",
  36384=>"100011000",
  36385=>"111111111",
  36386=>"000110110",
  36387=>"000011000",
  36388=>"000001111",
  36389=>"000000000",
  36390=>"100000000",
  36391=>"001101111",
  36392=>"111111011",
  36393=>"000000000",
  36394=>"111001111",
  36395=>"110110111",
  36396=>"111111010",
  36397=>"111000000",
  36398=>"011000000",
  36399=>"000000000",
  36400=>"011011000",
  36401=>"110111011",
  36402=>"110000000",
  36403=>"000000001",
  36404=>"111111110",
  36405=>"110111111",
  36406=>"001000000",
  36407=>"110111110",
  36408=>"000111100",
  36409=>"000000000",
  36410=>"000000100",
  36411=>"000001011",
  36412=>"000000000",
  36413=>"010000111",
  36414=>"111011010",
  36415=>"000111000",
  36416=>"000001011",
  36417=>"101111001",
  36418=>"101100111",
  36419=>"000000000",
  36420=>"000000110",
  36421=>"110000000",
  36422=>"000000001",
  36423=>"111001001",
  36424=>"000000000",
  36425=>"000001111",
  36426=>"011000111",
  36427=>"110111101",
  36428=>"111111011",
  36429=>"000000000",
  36430=>"001111111",
  36431=>"111111010",
  36432=>"000000111",
  36433=>"001000000",
  36434=>"111111011",
  36435=>"111011001",
  36436=>"111111111",
  36437=>"000100000",
  36438=>"111111101",
  36439=>"110100000",
  36440=>"100101111",
  36441=>"111101100",
  36442=>"000000111",
  36443=>"011000000",
  36444=>"100000011",
  36445=>"111011000",
  36446=>"000000000",
  36447=>"011111111",
  36448=>"000000011",
  36449=>"010010111",
  36450=>"111010011",
  36451=>"111000011",
  36452=>"000110110",
  36453=>"000000000",
  36454=>"000000000",
  36455=>"111101100",
  36456=>"011111111",
  36457=>"000000011",
  36458=>"111111111",
  36459=>"000100101",
  36460=>"110100000",
  36461=>"000000000",
  36462=>"000000000",
  36463=>"111111111",
  36464=>"100000000",
  36465=>"000000000",
  36466=>"101101111",
  36467=>"111100000",
  36468=>"000000011",
  36469=>"110000000",
  36470=>"000110111",
  36471=>"111111001",
  36472=>"011111000",
  36473=>"111000000",
  36474=>"111111111",
  36475=>"000000000",
  36476=>"001001011",
  36477=>"011111100",
  36478=>"000000001",
  36479=>"100000000",
  36480=>"000000000",
  36481=>"000110000",
  36482=>"111001101",
  36483=>"011011011",
  36484=>"000000000",
  36485=>"110111111",
  36486=>"000000000",
  36487=>"000010111",
  36488=>"111011111",
  36489=>"011001111",
  36490=>"001001111",
  36491=>"111111111",
  36492=>"000001111",
  36493=>"110110110",
  36494=>"101000000",
  36495=>"111000001",
  36496=>"111000011",
  36497=>"111001001",
  36498=>"000000000",
  36499=>"111111100",
  36500=>"000000000",
  36501=>"000000110",
  36502=>"000000000",
  36503=>"001111111",
  36504=>"100000000",
  36505=>"000000001",
  36506=>"010110111",
  36507=>"111001111",
  36508=>"110000110",
  36509=>"001000000",
  36510=>"001000110",
  36511=>"010011000",
  36512=>"001011000",
  36513=>"001111111",
  36514=>"000000010",
  36515=>"000000101",
  36516=>"110110010",
  36517=>"000010110",
  36518=>"110000000",
  36519=>"100110110",
  36520=>"000111111",
  36521=>"111101001",
  36522=>"101001000",
  36523=>"000111111",
  36524=>"000000000",
  36525=>"000000000",
  36526=>"000000100",
  36527=>"111000000",
  36528=>"000111110",
  36529=>"001100000",
  36530=>"111111111",
  36531=>"111100011",
  36532=>"110000000",
  36533=>"000111111",
  36534=>"111100111",
  36535=>"111111111",
  36536=>"111111110",
  36537=>"111111000",
  36538=>"111111111",
  36539=>"100000100",
  36540=>"000000000",
  36541=>"001011100",
  36542=>"111111111",
  36543=>"011011000",
  36544=>"111111111",
  36545=>"111110111",
  36546=>"111001100",
  36547=>"111111000",
  36548=>"111010010",
  36549=>"000000000",
  36550=>"100000111",
  36551=>"000010000",
  36552=>"110000000",
  36553=>"001000000",
  36554=>"010110100",
  36555=>"000000000",
  36556=>"111110000",
  36557=>"001000000",
  36558=>"100111111",
  36559=>"100000100",
  36560=>"100000000",
  36561=>"000000000",
  36562=>"000000000",
  36563=>"111000000",
  36564=>"111110100",
  36565=>"100100110",
  36566=>"011000000",
  36567=>"001001001",
  36568=>"000010000",
  36569=>"000001001",
  36570=>"000000000",
  36571=>"001111110",
  36572=>"011000000",
  36573=>"000000000",
  36574=>"000111111",
  36575=>"111111111",
  36576=>"011001001",
  36577=>"001111111",
  36578=>"011001011",
  36579=>"000000110",
  36580=>"110111111",
  36581=>"000000000",
  36582=>"000010000",
  36583=>"000000111",
  36584=>"000000000",
  36585=>"001111111",
  36586=>"000000111",
  36587=>"100000000",
  36588=>"111111011",
  36589=>"111001000",
  36590=>"001001111",
  36591=>"111111111",
  36592=>"110000111",
  36593=>"010000000",
  36594=>"111101000",
  36595=>"000000010",
  36596=>"000101110",
  36597=>"111011011",
  36598=>"000000001",
  36599=>"111111000",
  36600=>"111111111",
  36601=>"110110111",
  36602=>"000000111",
  36603=>"111000000",
  36604=>"111011000",
  36605=>"001011011",
  36606=>"001111000",
  36607=>"000001000",
  36608=>"011011110",
  36609=>"011000000",
  36610=>"111111111",
  36611=>"100111111",
  36612=>"000011111",
  36613=>"101111111",
  36614=>"000111111",
  36615=>"111111101",
  36616=>"001011011",
  36617=>"000000100",
  36618=>"110110000",
  36619=>"110111000",
  36620=>"110110110",
  36621=>"001001000",
  36622=>"000001001",
  36623=>"110100000",
  36624=>"011110110",
  36625=>"011001000",
  36626=>"000100111",
  36627=>"111111111",
  36628=>"111110111",
  36629=>"110000000",
  36630=>"111110100",
  36631=>"110000000",
  36632=>"111011111",
  36633=>"111111111",
  36634=>"000000000",
  36635=>"110010111",
  36636=>"111111010",
  36637=>"000010000",
  36638=>"001001100",
  36639=>"000000001",
  36640=>"000000000",
  36641=>"011001000",
  36642=>"010000000",
  36643=>"100001000",
  36644=>"001101100",
  36645=>"000000101",
  36646=>"111011011",
  36647=>"000000000",
  36648=>"000100111",
  36649=>"011010110",
  36650=>"000110110",
  36651=>"000001001",
  36652=>"000110000",
  36653=>"011011011",
  36654=>"000000111",
  36655=>"000011011",
  36656=>"110100000",
  36657=>"000100111",
  36658=>"111111111",
  36659=>"000000110",
  36660=>"111000000",
  36661=>"001000100",
  36662=>"000000111",
  36663=>"001000000",
  36664=>"000111110",
  36665=>"000110101",
  36666=>"000010110",
  36667=>"111000100",
  36668=>"110000000",
  36669=>"000100111",
  36670=>"111111111",
  36671=>"111001101",
  36672=>"000000000",
  36673=>"001111001",
  36674=>"000000100",
  36675=>"001001001",
  36676=>"111111111",
  36677=>"011000000",
  36678=>"111111100",
  36679=>"001000000",
  36680=>"110111001",
  36681=>"000000000",
  36682=>"000000100",
  36683=>"110000000",
  36684=>"100100100",
  36685=>"000000000",
  36686=>"000000000",
  36687=>"000001111",
  36688=>"000010110",
  36689=>"000110100",
  36690=>"000000000",
  36691=>"000000000",
  36692=>"000111000",
  36693=>"111111111",
  36694=>"001111111",
  36695=>"101100000",
  36696=>"111111111",
  36697=>"111000000",
  36698=>"111110000",
  36699=>"111111110",
  36700=>"000000000",
  36701=>"000110111",
  36702=>"010111111",
  36703=>"001001001",
  36704=>"100000000",
  36705=>"111001000",
  36706=>"011011011",
  36707=>"111111100",
  36708=>"111110000",
  36709=>"110000000",
  36710=>"100000000",
  36711=>"011111000",
  36712=>"001001001",
  36713=>"001000000",
  36714=>"111000000",
  36715=>"000000000",
  36716=>"110110100",
  36717=>"001001001",
  36718=>"100111101",
  36719=>"111111101",
  36720=>"000011111",
  36721=>"111001011",
  36722=>"111111111",
  36723=>"000111111",
  36724=>"111111100",
  36725=>"111011111",
  36726=>"110001000",
  36727=>"111111000",
  36728=>"111111110",
  36729=>"000111011",
  36730=>"111000000",
  36731=>"001001000",
  36732=>"100000000",
  36733=>"111111111",
  36734=>"001010000",
  36735=>"111111111",
  36736=>"111111000",
  36737=>"111111110",
  36738=>"110110111",
  36739=>"000000001",
  36740=>"001000000",
  36741=>"111111100",
  36742=>"111100111",
  36743=>"000111101",
  36744=>"111110111",
  36745=>"011111000",
  36746=>"000000000",
  36747=>"111111111",
  36748=>"100000101",
  36749=>"011000010",
  36750=>"111111111",
  36751=>"000000000",
  36752=>"001001001",
  36753=>"000000000",
  36754=>"000000000",
  36755=>"011000100",
  36756=>"010111010",
  36757=>"111110000",
  36758=>"111000001",
  36759=>"100110111",
  36760=>"110001000",
  36761=>"000100110",
  36762=>"110111111",
  36763=>"111001001",
  36764=>"010010000",
  36765=>"110110111",
  36766=>"000001111",
  36767=>"000000000",
  36768=>"100100110",
  36769=>"001101111",
  36770=>"110111111",
  36771=>"000000011",
  36772=>"000110000",
  36773=>"111111111",
  36774=>"111000111",
  36775=>"000000110",
  36776=>"111111101",
  36777=>"011011001",
  36778=>"011011111",
  36779=>"000111111",
  36780=>"000000000",
  36781=>"000000011",
  36782=>"011001000",
  36783=>"001111111",
  36784=>"001000000",
  36785=>"001111111",
  36786=>"110111111",
  36787=>"000000000",
  36788=>"001000101",
  36789=>"000001011",
  36790=>"011111111",
  36791=>"111011001",
  36792=>"000100111",
  36793=>"001011000",
  36794=>"111111100",
  36795=>"000000001",
  36796=>"111000000",
  36797=>"111111011",
  36798=>"000000010",
  36799=>"011010011",
  36800=>"000000000",
  36801=>"111000000",
  36802=>"111010000",
  36803=>"011010000",
  36804=>"011111000",
  36805=>"000001011",
  36806=>"000000101",
  36807=>"111000001",
  36808=>"000001000",
  36809=>"111111011",
  36810=>"110111011",
  36811=>"101000000",
  36812=>"111111001",
  36813=>"110111011",
  36814=>"001000100",
  36815=>"110000111",
  36816=>"111111111",
  36817=>"111110111",
  36818=>"001000000",
  36819=>"011011011",
  36820=>"000001000",
  36821=>"111111100",
  36822=>"000000000",
  36823=>"011001001",
  36824=>"111111000",
  36825=>"000000000",
  36826=>"000100111",
  36827=>"000000111",
  36828=>"100000000",
  36829=>"000000000",
  36830=>"011000111",
  36831=>"011111011",
  36832=>"111111100",
  36833=>"000110111",
  36834=>"000000000",
  36835=>"011000000",
  36836=>"110110011",
  36837=>"111000000",
  36838=>"000001111",
  36839=>"000000000",
  36840=>"000000000",
  36841=>"111100000",
  36842=>"000000000",
  36843=>"111011001",
  36844=>"000000000",
  36845=>"000110010",
  36846=>"001111111",
  36847=>"010000000",
  36848=>"000000111",
  36849=>"111111111",
  36850=>"010111111",
  36851=>"110100000",
  36852=>"110111111",
  36853=>"111010111",
  36854=>"111111111",
  36855=>"000000000",
  36856=>"111111000",
  36857=>"110110110",
  36858=>"110000000",
  36859=>"000000000",
  36860=>"000000000",
  36861=>"000000100",
  36862=>"111111000",
  36863=>"000000101",
  36864=>"000000000",
  36865=>"001011010",
  36866=>"100000101",
  36867=>"111111100",
  36868=>"111111111",
  36869=>"110110100",
  36870=>"011111011",
  36871=>"111111111",
  36872=>"000000000",
  36873=>"111111111",
  36874=>"111111111",
  36875=>"110110110",
  36876=>"110110111",
  36877=>"110100100",
  36878=>"000000011",
  36879=>"000000001",
  36880=>"111111111",
  36881=>"000111101",
  36882=>"000000000",
  36883=>"000000000",
  36884=>"000000011",
  36885=>"000000111",
  36886=>"000100000",
  36887=>"011011001",
  36888=>"100100100",
  36889=>"111111100",
  36890=>"101111110",
  36891=>"000001000",
  36892=>"001000000",
  36893=>"110010000",
  36894=>"101001001",
  36895=>"100100100",
  36896=>"110111001",
  36897=>"111111110",
  36898=>"000000000",
  36899=>"000000000",
  36900=>"000000001",
  36901=>"111011011",
  36902=>"000000110",
  36903=>"111000100",
  36904=>"111111110",
  36905=>"100000000",
  36906=>"111111111",
  36907=>"000000000",
  36908=>"111111111",
  36909=>"000111010",
  36910=>"000000000",
  36911=>"000010011",
  36912=>"101100101",
  36913=>"011011011",
  36914=>"001011011",
  36915=>"100000101",
  36916=>"101000000",
  36917=>"110010000",
  36918=>"101000000",
  36919=>"100110100",
  36920=>"000000111",
  36921=>"010011011",
  36922=>"011111111",
  36923=>"001111111",
  36924=>"111100100",
  36925=>"111000000",
  36926=>"000100001",
  36927=>"111111111",
  36928=>"011000011",
  36929=>"101101001",
  36930=>"110000111",
  36931=>"100100101",
  36932=>"111001001",
  36933=>"000000110",
  36934=>"000110010",
  36935=>"000000000",
  36936=>"001011001",
  36937=>"111111111",
  36938=>"110110000",
  36939=>"001000001",
  36940=>"111111111",
  36941=>"111111000",
  36942=>"000010110",
  36943=>"000000100",
  36944=>"110110000",
  36945=>"101100000",
  36946=>"000000000",
  36947=>"011001110",
  36948=>"011000000",
  36949=>"111111001",
  36950=>"111111111",
  36951=>"111111111",
  36952=>"011000110",
  36953=>"101000101",
  36954=>"000000000",
  36955=>"001110111",
  36956=>"000000000",
  36957=>"000000101",
  36958=>"111110110",
  36959=>"110010000",
  36960=>"000011111",
  36961=>"000000000",
  36962=>"011011000",
  36963=>"101111111",
  36964=>"111111110",
  36965=>"001001111",
  36966=>"111111111",
  36967=>"000000000",
  36968=>"101111110",
  36969=>"001000000",
  36970=>"010000111",
  36971=>"100011001",
  36972=>"111111110",
  36973=>"000001011",
  36974=>"100000100",
  36975=>"000111010",
  36976=>"011011111",
  36977=>"111101111",
  36978=>"110111111",
  36979=>"111111111",
  36980=>"111111110",
  36981=>"110111111",
  36982=>"001001111",
  36983=>"011111111",
  36984=>"000000000",
  36985=>"000000000",
  36986=>"000000000",
  36987=>"001101100",
  36988=>"111111101",
  36989=>"111111101",
  36990=>"000100000",
  36991=>"010000001",
  36992=>"000000000",
  36993=>"111111111",
  36994=>"011111001",
  36995=>"111111011",
  36996=>"010110110",
  36997=>"010000011",
  36998=>"001001111",
  36999=>"111010111",
  37000=>"000110111",
  37001=>"111000000",
  37002=>"111111111",
  37003=>"011000010",
  37004=>"110011001",
  37005=>"000000000",
  37006=>"000000000",
  37007=>"010011011",
  37008=>"101000101",
  37009=>"111011010",
  37010=>"011011110",
  37011=>"111111010",
  37012=>"111111111",
  37013=>"000000000",
  37014=>"010111111",
  37015=>"111100100",
  37016=>"100000000",
  37017=>"000000000",
  37018=>"100101111",
  37019=>"100100101",
  37020=>"110110000",
  37021=>"010000011",
  37022=>"111110000",
  37023=>"111111111",
  37024=>"100010000",
  37025=>"101000000",
  37026=>"111111111",
  37027=>"111111111",
  37028=>"000000000",
  37029=>"100110111",
  37030=>"000000111",
  37031=>"110110110",
  37032=>"111000101",
  37033=>"001001000",
  37034=>"010010010",
  37035=>"000000000",
  37036=>"111111000",
  37037=>"110100001",
  37038=>"111000000",
  37039=>"001001111",
  37040=>"111010000",
  37041=>"111000000",
  37042=>"011011010",
  37043=>"111001000",
  37044=>"000000000",
  37045=>"000000000",
  37046=>"001111111",
  37047=>"000000010",
  37048=>"110110101",
  37049=>"111111111",
  37050=>"000000000",
  37051=>"110110010",
  37052=>"111111000",
  37053=>"111111010",
  37054=>"100100100",
  37055=>"000001000",
  37056=>"000000100",
  37057=>"111110111",
  37058=>"111111111",
  37059=>"101001000",
  37060=>"000000000",
  37061=>"000000011",
  37062=>"100000110",
  37063=>"000000100",
  37064=>"010110111",
  37065=>"011000100",
  37066=>"010000000",
  37067=>"010111111",
  37068=>"100000000",
  37069=>"001001001",
  37070=>"001000001",
  37071=>"011000000",
  37072=>"000000000",
  37073=>"000000000",
  37074=>"001001000",
  37075=>"000000000",
  37076=>"000100100",
  37077=>"100100110",
  37078=>"000000000",
  37079=>"011000110",
  37080=>"110110111",
  37081=>"111001111",
  37082=>"111111111",
  37083=>"100111111",
  37084=>"100000100",
  37085=>"000000000",
  37086=>"001100101",
  37087=>"010010000",
  37088=>"000001011",
  37089=>"000000011",
  37090=>"100100110",
  37091=>"000000000",
  37092=>"110101100",
  37093=>"011011100",
  37094=>"000100100",
  37095=>"111111111",
  37096=>"111111011",
  37097=>"111111110",
  37098=>"000000000",
  37099=>"110111100",
  37100=>"100000000",
  37101=>"100000000",
  37102=>"000000110",
  37103=>"110111111",
  37104=>"111110100",
  37105=>"010000000",
  37106=>"111111010",
  37107=>"111000000",
  37108=>"111111111",
  37109=>"111111001",
  37110=>"011111011",
  37111=>"111100000",
  37112=>"010000000",
  37113=>"000000000",
  37114=>"111000001",
  37115=>"101101001",
  37116=>"010011111",
  37117=>"110011011",
  37118=>"000001001",
  37119=>"010110110",
  37120=>"111000000",
  37121=>"111001101",
  37122=>"111111111",
  37123=>"010010000",
  37124=>"001000000",
  37125=>"010010110",
  37126=>"111111100",
  37127=>"111001001",
  37128=>"000000000",
  37129=>"111000000",
  37130=>"000000000",
  37131=>"111111111",
  37132=>"101000001",
  37133=>"001000010",
  37134=>"111111011",
  37135=>"111100000",
  37136=>"000000000",
  37137=>"111100000",
  37138=>"001001001",
  37139=>"011111111",
  37140=>"000000010",
  37141=>"011111111",
  37142=>"010011111",
  37143=>"011001001",
  37144=>"000001111",
  37145=>"111100100",
  37146=>"000000000",
  37147=>"010000110",
  37148=>"110000000",
  37149=>"110110000",
  37150=>"000000000",
  37151=>"111011110",
  37152=>"100100001",
  37153=>"101111111",
  37154=>"000000000",
  37155=>"111110000",
  37156=>"110110100",
  37157=>"000000101",
  37158=>"000000001",
  37159=>"000000110",
  37160=>"000011111",
  37161=>"000000000",
  37162=>"100110111",
  37163=>"000000000",
  37164=>"111000010",
  37165=>"110100000",
  37166=>"000001000",
  37167=>"000000000",
  37168=>"000100000",
  37169=>"010010000",
  37170=>"111111101",
  37171=>"100111111",
  37172=>"000000000",
  37173=>"001010000",
  37174=>"111111100",
  37175=>"000111110",
  37176=>"110010010",
  37177=>"101001001",
  37178=>"000000000",
  37179=>"111111100",
  37180=>"111010111",
  37181=>"111111111",
  37182=>"111111000",
  37183=>"110110000",
  37184=>"101100000",
  37185=>"100101111",
  37186=>"110111111",
  37187=>"000000101",
  37188=>"010110111",
  37189=>"000000000",
  37190=>"010111111",
  37191=>"110110010",
  37192=>"101101101",
  37193=>"000000000",
  37194=>"111111110",
  37195=>"001000000",
  37196=>"000000000",
  37197=>"110100011",
  37198=>"110101000",
  37199=>"110110110",
  37200=>"011001111",
  37201=>"100000101",
  37202=>"011011011",
  37203=>"000000000",
  37204=>"000110110",
  37205=>"001001011",
  37206=>"110110111",
  37207=>"101111111",
  37208=>"110100110",
  37209=>"001000101",
  37210=>"000000010",
  37211=>"000000000",
  37212=>"000011011",
  37213=>"000000000",
  37214=>"000010110",
  37215=>"111111000",
  37216=>"000001101",
  37217=>"000000100",
  37218=>"110110110",
  37219=>"111101111",
  37220=>"100100010",
  37221=>"011000000",
  37222=>"001000110",
  37223=>"110111110",
  37224=>"100000100",
  37225=>"100000000",
  37226=>"010010000",
  37227=>"000110010",
  37228=>"110100100",
  37229=>"000000100",
  37230=>"010111111",
  37231=>"111110111",
  37232=>"000000000",
  37233=>"111101001",
  37234=>"111000010",
  37235=>"000000000",
  37236=>"000000000",
  37237=>"011111111",
  37238=>"001111111",
  37239=>"111111010",
  37240=>"001000000",
  37241=>"101000000",
  37242=>"100000000",
  37243=>"000000000",
  37244=>"100100000",
  37245=>"000000010",
  37246=>"000100110",
  37247=>"000111011",
  37248=>"110110110",
  37249=>"111111111",
  37250=>"000011010",
  37251=>"000000001",
  37252=>"000000000",
  37253=>"000000111",
  37254=>"000000111",
  37255=>"000000000",
  37256=>"100000100",
  37257=>"000011111",
  37258=>"000110111",
  37259=>"000000000",
  37260=>"111000111",
  37261=>"110100100",
  37262=>"111111010",
  37263=>"111001001",
  37264=>"000000101",
  37265=>"000100100",
  37266=>"111101000",
  37267=>"001000100",
  37268=>"111000000",
  37269=>"000000000",
  37270=>"001001101",
  37271=>"111000000",
  37272=>"000000111",
  37273=>"111010000",
  37274=>"101100101",
  37275=>"110100111",
  37276=>"111111111",
  37277=>"011111111",
  37278=>"000000000",
  37279=>"111111011",
  37280=>"000000000",
  37281=>"010011000",
  37282=>"111000000",
  37283=>"110000111",
  37284=>"101100011",
  37285=>"001001011",
  37286=>"101001000",
  37287=>"011011000",
  37288=>"110110110",
  37289=>"011010010",
  37290=>"010011111",
  37291=>"111001000",
  37292=>"111111111",
  37293=>"001100001",
  37294=>"000000000",
  37295=>"000000100",
  37296=>"000000000",
  37297=>"111101000",
  37298=>"110110010",
  37299=>"000011010",
  37300=>"011000000",
  37301=>"110111110",
  37302=>"111110100",
  37303=>"111111111",
  37304=>"110110110",
  37305=>"011111111",
  37306=>"110110110",
  37307=>"000000001",
  37308=>"010000000",
  37309=>"010001111",
  37310=>"101001001",
  37311=>"111111111",
  37312=>"000000000",
  37313=>"001000000",
  37314=>"000001000",
  37315=>"000000111",
  37316=>"111000111",
  37317=>"000111111",
  37318=>"000000011",
  37319=>"000000000",
  37320=>"000000001",
  37321=>"000000000",
  37322=>"111100110",
  37323=>"111000111",
  37324=>"111111111",
  37325=>"000000010",
  37326=>"100111000",
  37327=>"111111111",
  37328=>"111111101",
  37329=>"111111111",
  37330=>"000000100",
  37331=>"100000100",
  37332=>"111110110",
  37333=>"111000000",
  37334=>"000010000",
  37335=>"011011000",
  37336=>"001000100",
  37337=>"100100000",
  37338=>"000000101",
  37339=>"011000010",
  37340=>"011111010",
  37341=>"010000000",
  37342=>"001000100",
  37343=>"011001111",
  37344=>"001001000",
  37345=>"000000011",
  37346=>"010010010",
  37347=>"111111010",
  37348=>"111110110",
  37349=>"101001001",
  37350=>"111100110",
  37351=>"001000000",
  37352=>"110010011",
  37353=>"000000000",
  37354=>"011111111",
  37355=>"111110100",
  37356=>"111111111",
  37357=>"001001100",
  37358=>"100100110",
  37359=>"111111111",
  37360=>"000000000",
  37361=>"000000000",
  37362=>"000000000",
  37363=>"001000101",
  37364=>"001001101",
  37365=>"100100000",
  37366=>"110111111",
  37367=>"000111000",
  37368=>"110000111",
  37369=>"011011001",
  37370=>"101000000",
  37371=>"000010110",
  37372=>"000000111",
  37373=>"110110111",
  37374=>"100000000",
  37375=>"000000000",
  37376=>"001001001",
  37377=>"101111110",
  37378=>"111111111",
  37379=>"001001001",
  37380=>"100001111",
  37381=>"001111000",
  37382=>"110110111",
  37383=>"111111111",
  37384=>"000001001",
  37385=>"111111111",
  37386=>"111100101",
  37387=>"011000000",
  37388=>"000000000",
  37389=>"110001011",
  37390=>"001000111",
  37391=>"111111111",
  37392=>"100000100",
  37393=>"111111011",
  37394=>"111111111",
  37395=>"111111111",
  37396=>"111000100",
  37397=>"000000000",
  37398=>"111111111",
  37399=>"111110111",
  37400=>"110111111",
  37401=>"000000000",
  37402=>"000000010",
  37403=>"001111111",
  37404=>"111111011",
  37405=>"000000111",
  37406=>"100001011",
  37407=>"000000000",
  37408=>"111111111",
  37409=>"000000000",
  37410=>"111111111",
  37411=>"001001000",
  37412=>"011000000",
  37413=>"010010010",
  37414=>"000000000",
  37415=>"111000000",
  37416=>"111111111",
  37417=>"111111100",
  37418=>"111111111",
  37419=>"110000100",
  37420=>"000000000",
  37421=>"111111000",
  37422=>"000000011",
  37423=>"000000000",
  37424=>"011001111",
  37425=>"100110111",
  37426=>"111111111",
  37427=>"111111111",
  37428=>"111111111",
  37429=>"010000000",
  37430=>"011000001",
  37431=>"100000000",
  37432=>"111111111",
  37433=>"111000110",
  37434=>"101111111",
  37435=>"111111001",
  37436=>"011000011",
  37437=>"111000111",
  37438=>"111000001",
  37439=>"111111000",
  37440=>"000000000",
  37441=>"000111111",
  37442=>"010010011",
  37443=>"111111111",
  37444=>"000000000",
  37445=>"000000000",
  37446=>"111111111",
  37447=>"000000000",
  37448=>"000000001",
  37449=>"111011001",
  37450=>"111001000",
  37451=>"111111111",
  37452=>"001000101",
  37453=>"000000011",
  37454=>"010000000",
  37455=>"000000111",
  37456=>"111111111",
  37457=>"110110000",
  37458=>"000000000",
  37459=>"111111111",
  37460=>"000100111",
  37461=>"110000000",
  37462=>"111011111",
  37463=>"111111111",
  37464=>"111111111",
  37465=>"111101101",
  37466=>"010010011",
  37467=>"000000000",
  37468=>"111111000",
  37469=>"000011010",
  37470=>"110000100",
  37471=>"011011111",
  37472=>"111000000",
  37473=>"000000000",
  37474=>"000100111",
  37475=>"111111111",
  37476=>"001000000",
  37477=>"001000000",
  37478=>"011111111",
  37479=>"000000000",
  37480=>"100000011",
  37481=>"000111111",
  37482=>"110000000",
  37483=>"111111111",
  37484=>"011111101",
  37485=>"000000010",
  37486=>"000000111",
  37487=>"100000000",
  37488=>"011111010",
  37489=>"000001001",
  37490=>"000000001",
  37491=>"100000110",
  37492=>"000000110",
  37493=>"000000100",
  37494=>"000000000",
  37495=>"100000000",
  37496=>"111111111",
  37497=>"100000101",
  37498=>"000000000",
  37499=>"000000000",
  37500=>"000000000",
  37501=>"111011011",
  37502=>"100100110",
  37503=>"100000000",
  37504=>"111001000",
  37505=>"111000001",
  37506=>"000000000",
  37507=>"111111111",
  37508=>"100111100",
  37509=>"101000111",
  37510=>"111010000",
  37511=>"111111100",
  37512=>"111111111",
  37513=>"000001001",
  37514=>"111111111",
  37515=>"111111111",
  37516=>"000000000",
  37517=>"000000000",
  37518=>"111100010",
  37519=>"000000000",
  37520=>"001001000",
  37521=>"111110000",
  37522=>"111100100",
  37523=>"111111111",
  37524=>"111111111",
  37525=>"001001000",
  37526=>"000000000",
  37527=>"000000000",
  37528=>"000000000",
  37529=>"111111000",
  37530=>"001101101",
  37531=>"000000000",
  37532=>"111111111",
  37533=>"111000000",
  37534=>"010000011",
  37535=>"000001001",
  37536=>"000000111",
  37537=>"000000111",
  37538=>"000000000",
  37539=>"000111011",
  37540=>"100100000",
  37541=>"111101101",
  37542=>"000000000",
  37543=>"110111100",
  37544=>"111101110",
  37545=>"111101000",
  37546=>"111111111",
  37547=>"101100000",
  37548=>"010000111",
  37549=>"100011111",
  37550=>"000000001",
  37551=>"000000010",
  37552=>"000000000",
  37553=>"111100111",
  37554=>"000010110",
  37555=>"111111000",
  37556=>"000010111",
  37557=>"111110110",
  37558=>"011000000",
  37559=>"111111111",
  37560=>"110110110",
  37561=>"000000111",
  37562=>"100100000",
  37563=>"111101000",
  37564=>"000000000",
  37565=>"001111111",
  37566=>"111111111",
  37567=>"111111111",
  37568=>"111111111",
  37569=>"000000001",
  37570=>"110110000",
  37571=>"111111111",
  37572=>"111111001",
  37573=>"100100000",
  37574=>"000000000",
  37575=>"000000011",
  37576=>"000000000",
  37577=>"000000001",
  37578=>"111001111",
  37579=>"000000000",
  37580=>"000001001",
  37581=>"001000000",
  37582=>"111111011",
  37583=>"111111111",
  37584=>"000011011",
  37585=>"000000010",
  37586=>"000000111",
  37587=>"000000000",
  37588=>"001000001",
  37589=>"000000001",
  37590=>"000000000",
  37591=>"111111111",
  37592=>"111001111",
  37593=>"101001001",
  37594=>"001000001",
  37595=>"111000000",
  37596=>"000100100",
  37597=>"000000000",
  37598=>"000000000",
  37599=>"000000000",
  37600=>"100111011",
  37601=>"000000000",
  37602=>"000000000",
  37603=>"101111111",
  37604=>"000000000",
  37605=>"001000000",
  37606=>"000000000",
  37607=>"011001111",
  37608=>"111111111",
  37609=>"100100000",
  37610=>"000000000",
  37611=>"111111110",
  37612=>"111111011",
  37613=>"000010000",
  37614=>"000111111",
  37615=>"111111010",
  37616=>"111000000",
  37617=>"110110111",
  37618=>"000010110",
  37619=>"010000000",
  37620=>"000000000",
  37621=>"000000101",
  37622=>"011111111",
  37623=>"111110111",
  37624=>"111100000",
  37625=>"000000000",
  37626=>"110111011",
  37627=>"000000000",
  37628=>"001000001",
  37629=>"001000000",
  37630=>"111011011",
  37631=>"100000000",
  37632=>"100100111",
  37633=>"110111111",
  37634=>"111101111",
  37635=>"000000000",
  37636=>"100101111",
  37637=>"111111111",
  37638=>"000000110",
  37639=>"111100110",
  37640=>"111111111",
  37641=>"100000000",
  37642=>"000000000",
  37643=>"111111111",
  37644=>"010011010",
  37645=>"000000001",
  37646=>"000101111",
  37647=>"000000000",
  37648=>"000001001",
  37649=>"000001001",
  37650=>"110111111",
  37651=>"111111111",
  37652=>"011111111",
  37653=>"000000000",
  37654=>"001001000",
  37655=>"110100100",
  37656=>"110100000",
  37657=>"010111101",
  37658=>"000001000",
  37659=>"100000010",
  37660=>"000000000",
  37661=>"111111111",
  37662=>"111111111",
  37663=>"001000000",
  37664=>"001000000",
  37665=>"000100000",
  37666=>"111111100",
  37667=>"111001011",
  37668=>"001001110",
  37669=>"000000000",
  37670=>"001000000",
  37671=>"000100000",
  37672=>"011011110",
  37673=>"001001000",
  37674=>"100000000",
  37675=>"111111111",
  37676=>"110111001",
  37677=>"000110111",
  37678=>"111110111",
  37679=>"111111110",
  37680=>"111111111",
  37681=>"010000001",
  37682=>"100101001",
  37683=>"111111110",
  37684=>"111111111",
  37685=>"111111111",
  37686=>"000000000",
  37687=>"000000000",
  37688=>"000000000",
  37689=>"110110000",
  37690=>"111111110",
  37691=>"000000001",
  37692=>"111111111",
  37693=>"111110111",
  37694=>"100000000",
  37695=>"001000000",
  37696=>"000100000",
  37697=>"111111111",
  37698=>"100100111",
  37699=>"000000000",
  37700=>"001000000",
  37701=>"001001111",
  37702=>"011010111",
  37703=>"100111111",
  37704=>"111111000",
  37705=>"111111001",
  37706=>"111001001",
  37707=>"001001010",
  37708=>"010010000",
  37709=>"111111100",
  37710=>"101100101",
  37711=>"101100110",
  37712=>"011000000",
  37713=>"111111111",
  37714=>"000000000",
  37715=>"000011111",
  37716=>"000000111",
  37717=>"000000000",
  37718=>"000000000",
  37719=>"111111011",
  37720=>"111111111",
  37721=>"000000000",
  37722=>"111111100",
  37723=>"000000000",
  37724=>"001000000",
  37725=>"001000000",
  37726=>"100100100",
  37727=>"000000000",
  37728=>"000000000",
  37729=>"011001000",
  37730=>"111100100",
  37731=>"000000110",
  37732=>"111111111",
  37733=>"000000100",
  37734=>"111111110",
  37735=>"000000000",
  37736=>"000001000",
  37737=>"011001011",
  37738=>"101000000",
  37739=>"000101101",
  37740=>"110110110",
  37741=>"100110000",
  37742=>"000000000",
  37743=>"000001000",
  37744=>"000000000",
  37745=>"100110111",
  37746=>"000000000",
  37747=>"111111111",
  37748=>"110111111",
  37749=>"000000000",
  37750=>"011001000",
  37751=>"111111001",
  37752=>"111111111",
  37753=>"011010111",
  37754=>"001000011",
  37755=>"110110100",
  37756=>"011001000",
  37757=>"110111110",
  37758=>"000000000",
  37759=>"111001000",
  37760=>"111011111",
  37761=>"000000000",
  37762=>"000000000",
  37763=>"000000000",
  37764=>"000000000",
  37765=>"000000000",
  37766=>"000001000",
  37767=>"000010010",
  37768=>"111001001",
  37769=>"111110100",
  37770=>"001111111",
  37771=>"101111111",
  37772=>"000100000",
  37773=>"000000000",
  37774=>"101000111",
  37775=>"011011000",
  37776=>"000000000",
  37777=>"111111111",
  37778=>"000000001",
  37779=>"111111111",
  37780=>"111000000",
  37781=>"000110111",
  37782=>"111111111",
  37783=>"000000110",
  37784=>"110101111",
  37785=>"011001000",
  37786=>"111111111",
  37787=>"111111111",
  37788=>"000000001",
  37789=>"111111110",
  37790=>"111010000",
  37791=>"000000000",
  37792=>"010011011",
  37793=>"000000000",
  37794=>"111000111",
  37795=>"000000001",
  37796=>"101000011",
  37797=>"100111111",
  37798=>"111111100",
  37799=>"000000001",
  37800=>"100000011",
  37801=>"010011011",
  37802=>"101001011",
  37803=>"100000000",
  37804=>"101101001",
  37805=>"111111111",
  37806=>"111111111",
  37807=>"000000000",
  37808=>"111111111",
  37809=>"000110001",
  37810=>"111111111",
  37811=>"111111111",
  37812=>"000000000",
  37813=>"000000000",
  37814=>"111100110",
  37815=>"001000000",
  37816=>"100000100",
  37817=>"000010111",
  37818=>"001011000",
  37819=>"111111111",
  37820=>"000000111",
  37821=>"111111111",
  37822=>"000000000",
  37823=>"110110011",
  37824=>"001001001",
  37825=>"001011011",
  37826=>"111111111",
  37827=>"111111111",
  37828=>"111101111",
  37829=>"110110000",
  37830=>"110110000",
  37831=>"000111011",
  37832=>"111111111",
  37833=>"111000011",
  37834=>"000000001",
  37835=>"111101011",
  37836=>"000000000",
  37837=>"000000000",
  37838=>"001000000",
  37839=>"000111111",
  37840=>"000000000",
  37841=>"001111100",
  37842=>"111111000",
  37843=>"011000111",
  37844=>"000000111",
  37845=>"111011101",
  37846=>"000000000",
  37847=>"011011011",
  37848=>"000000000",
  37849=>"110110001",
  37850=>"000000110",
  37851=>"111101111",
  37852=>"000011000",
  37853=>"000000000",
  37854=>"111011011",
  37855=>"000010000",
  37856=>"111100001",
  37857=>"000000100",
  37858=>"001000000",
  37859=>"000000111",
  37860=>"111111110",
  37861=>"110000000",
  37862=>"111111111",
  37863=>"110000000",
  37864=>"100000111",
  37865=>"111110100",
  37866=>"011010010",
  37867=>"111101111",
  37868=>"111111111",
  37869=>"100110100",
  37870=>"000111111",
  37871=>"111000000",
  37872=>"000000000",
  37873=>"001001011",
  37874=>"011001101",
  37875=>"000000000",
  37876=>"000000111",
  37877=>"000000000",
  37878=>"111111001",
  37879=>"110011001",
  37880=>"001000011",
  37881=>"001010010",
  37882=>"110110111",
  37883=>"100110111",
  37884=>"000000000",
  37885=>"010110111",
  37886=>"110000100",
  37887=>"100000110",
  37888=>"000000010",
  37889=>"000000000",
  37890=>"000000000",
  37891=>"111000000",
  37892=>"000000000",
  37893=>"000000000",
  37894=>"000000000",
  37895=>"111111111",
  37896=>"000000110",
  37897=>"000100100",
  37898=>"010010000",
  37899=>"000000000",
  37900=>"000000000",
  37901=>"101111111",
  37902=>"010000000",
  37903=>"111111111",
  37904=>"111111001",
  37905=>"000000000",
  37906=>"000000000",
  37907=>"011111110",
  37908=>"111000000",
  37909=>"111110100",
  37910=>"111111111",
  37911=>"110011001",
  37912=>"111111001",
  37913=>"111110000",
  37914=>"111011111",
  37915=>"000000000",
  37916=>"111101111",
  37917=>"000000111",
  37918=>"111111111",
  37919=>"000000000",
  37920=>"000010010",
  37921=>"110110011",
  37922=>"111110000",
  37923=>"111000000",
  37924=>"100111110",
  37925=>"000001000",
  37926=>"000010000",
  37927=>"011111111",
  37928=>"111111111",
  37929=>"110000000",
  37930=>"111111110",
  37931=>"100000000",
  37932=>"111111000",
  37933=>"111001000",
  37934=>"000000000",
  37935=>"100000011",
  37936=>"111110111",
  37937=>"111000000",
  37938=>"100110110",
  37939=>"000000000",
  37940=>"000000000",
  37941=>"000011001",
  37942=>"111111010",
  37943=>"101111111",
  37944=>"000000000",
  37945=>"111111000",
  37946=>"000000000",
  37947=>"111111111",
  37948=>"101100111",
  37949=>"000011011",
  37950=>"000000000",
  37951=>"111110000",
  37952=>"000000000",
  37953=>"011011111",
  37954=>"000110111",
  37955=>"111010000",
  37956=>"000000000",
  37957=>"110110110",
  37958=>"111000000",
  37959=>"000000000",
  37960=>"000000100",
  37961=>"000100111",
  37962=>"110000111",
  37963=>"000000000",
  37964=>"101000100",
  37965=>"001000000",
  37966=>"000000111",
  37967=>"111111111",
  37968=>"111111111",
  37969=>"100000000",
  37970=>"000000000",
  37971=>"100100000",
  37972=>"000000111",
  37973=>"111111010",
  37974=>"100110110",
  37975=>"000000000",
  37976=>"000000100",
  37977=>"111101111",
  37978=>"111111110",
  37979=>"001000000",
  37980=>"111111110",
  37981=>"111111111",
  37982=>"100100000",
  37983=>"000000000",
  37984=>"111111111",
  37985=>"000100100",
  37986=>"110000000",
  37987=>"000000110",
  37988=>"000000100",
  37989=>"000000000",
  37990=>"000011000",
  37991=>"111111110",
  37992=>"000000000",
  37993=>"110110111",
  37994=>"010010011",
  37995=>"111001111",
  37996=>"001000000",
  37997=>"110111011",
  37998=>"111011001",
  37999=>"111111100",
  38000=>"000000000",
  38001=>"111111111",
  38002=>"000000111",
  38003=>"110000000",
  38004=>"011001001",
  38005=>"111110000",
  38006=>"100111111",
  38007=>"001000111",
  38008=>"000000000",
  38009=>"001111111",
  38010=>"011111010",
  38011=>"000000010",
  38012=>"011011011",
  38013=>"010111110",
  38014=>"010000000",
  38015=>"000000011",
  38016=>"111011001",
  38017=>"000000000",
  38018=>"111111001",
  38019=>"000011111",
  38020=>"111110000",
  38021=>"000000111",
  38022=>"111111111",
  38023=>"000111110",
  38024=>"111111010",
  38025=>"111111111",
  38026=>"000000000",
  38027=>"000000000",
  38028=>"111111111",
  38029=>"110010010",
  38030=>"111101111",
  38031=>"000000000",
  38032=>"110110000",
  38033=>"000000111",
  38034=>"111101000",
  38035=>"111100101",
  38036=>"110000000",
  38037=>"000000000",
  38038=>"100000100",
  38039=>"000101111",
  38040=>"111111011",
  38041=>"000110111",
  38042=>"000000000",
  38043=>"000100111",
  38044=>"000000000",
  38045=>"000001111",
  38046=>"110111111",
  38047=>"011000000",
  38048=>"111000000",
  38049=>"111111111",
  38050=>"001111100",
  38051=>"000000000",
  38052=>"000100100",
  38053=>"101101111",
  38054=>"010111111",
  38055=>"000001011",
  38056=>"111000000",
  38057=>"110001111",
  38058=>"000000000",
  38059=>"100000111",
  38060=>"010000000",
  38061=>"111001001",
  38062=>"111010000",
  38063=>"001000000",
  38064=>"000000111",
  38065=>"011000000",
  38066=>"111110111",
  38067=>"110000010",
  38068=>"000001000",
  38069=>"000000000",
  38070=>"110111110",
  38071=>"111111111",
  38072=>"001111100",
  38073=>"000000000",
  38074=>"001111111",
  38075=>"101111111",
  38076=>"000000000",
  38077=>"011011001",
  38078=>"111111111",
  38079=>"000000000",
  38080=>"111111111",
  38081=>"111111100",
  38082=>"000111111",
  38083=>"111111111",
  38084=>"110110000",
  38085=>"010000000",
  38086=>"000000000",
  38087=>"111111110",
  38088=>"000000000",
  38089=>"000000000",
  38090=>"100001111",
  38091=>"000000000",
  38092=>"011100000",
  38093=>"111111111",
  38094=>"111011111",
  38095=>"000000000",
  38096=>"000000000",
  38097=>"000000000",
  38098=>"000000000",
  38099=>"011011000",
  38100=>"101000111",
  38101=>"110100100",
  38102=>"000100000",
  38103=>"001000001",
  38104=>"111111110",
  38105=>"000000000",
  38106=>"000000000",
  38107=>"111111111",
  38108=>"011011111",
  38109=>"111111111",
  38110=>"000000000",
  38111=>"000001001",
  38112=>"111111111",
  38113=>"110111111",
  38114=>"111111110",
  38115=>"000000000",
  38116=>"011111011",
  38117=>"100000000",
  38118=>"010111111",
  38119=>"000010100",
  38120=>"000000000",
  38121=>"111111111",
  38122=>"000000100",
  38123=>"000000000",
  38124=>"010111111",
  38125=>"000111111",
  38126=>"000000111",
  38127=>"000000000",
  38128=>"111111111",
  38129=>"100111101",
  38130=>"111011001",
  38131=>"111111001",
  38132=>"000000000",
  38133=>"000000001",
  38134=>"100100111",
  38135=>"010010000",
  38136=>"000011111",
  38137=>"111110111",
  38138=>"000000000",
  38139=>"000000000",
  38140=>"110100011",
  38141=>"111001111",
  38142=>"111100100",
  38143=>"111111100",
  38144=>"110010000",
  38145=>"111111110",
  38146=>"111111111",
  38147=>"000111011",
  38148=>"000000000",
  38149=>"011111010",
  38150=>"000000000",
  38151=>"011111001",
  38152=>"111011111",
  38153=>"000000010",
  38154=>"000000000",
  38155=>"010011001",
  38156=>"001001111",
  38157=>"000111001",
  38158=>"000000100",
  38159=>"111000000",
  38160=>"000000111",
  38161=>"000000000",
  38162=>"000100111",
  38163=>"000000001",
  38164=>"111100000",
  38165=>"000000010",
  38166=>"110110100",
  38167=>"000001001",
  38168=>"111111111",
  38169=>"111111100",
  38170=>"000000000",
  38171=>"110010000",
  38172=>"111111111",
  38173=>"111111000",
  38174=>"000111111",
  38175=>"010111111",
  38176=>"101101001",
  38177=>"000001111",
  38178=>"000110111",
  38179=>"110111100",
  38180=>"111111111",
  38181=>"000000000",
  38182=>"111111111",
  38183=>"100111100",
  38184=>"111011111",
  38185=>"111010111",
  38186=>"111111000",
  38187=>"000111111",
  38188=>"111000000",
  38189=>"111111000",
  38190=>"000111001",
  38191=>"000000000",
  38192=>"111101100",
  38193=>"011111111",
  38194=>"111111011",
  38195=>"111000000",
  38196=>"001100000",
  38197=>"111111110",
  38198=>"111111110",
  38199=>"111111110",
  38200=>"000110000",
  38201=>"000111111",
  38202=>"000000000",
  38203=>"000000111",
  38204=>"100100110",
  38205=>"000001001",
  38206=>"100000000",
  38207=>"000000000",
  38208=>"000000000",
  38209=>"111111111",
  38210=>"111101001",
  38211=>"000000000",
  38212=>"100111111",
  38213=>"111111110",
  38214=>"111000000",
  38215=>"000000001",
  38216=>"111000000",
  38217=>"000000000",
  38218=>"111010000",
  38219=>"111111100",
  38220=>"000110000",
  38221=>"000000111",
  38222=>"110000000",
  38223=>"101111111",
  38224=>"000000000",
  38225=>"000000000",
  38226=>"111110111",
  38227=>"111000000",
  38228=>"000000000",
  38229=>"001000001",
  38230=>"111111011",
  38231=>"110000000",
  38232=>"000000111",
  38233=>"000000000",
  38234=>"000000000",
  38235=>"110111100",
  38236=>"011111111",
  38237=>"000100110",
  38238=>"000000010",
  38239=>"111111111",
  38240=>"011111111",
  38241=>"000000010",
  38242=>"100110011",
  38243=>"000000000",
  38244=>"000000000",
  38245=>"001000000",
  38246=>"000000000",
  38247=>"000000001",
  38248=>"110111111",
  38249=>"000000000",
  38250=>"010110111",
  38251=>"000000000",
  38252=>"011011111",
  38253=>"011111111",
  38254=>"000000000",
  38255=>"100100100",
  38256=>"110100000",
  38257=>"111111011",
  38258=>"111111110",
  38259=>"101000000",
  38260=>"001000000",
  38261=>"000011111",
  38262=>"111001000",
  38263=>"100000000",
  38264=>"111000000",
  38265=>"000100100",
  38266=>"111111111",
  38267=>"111110100",
  38268=>"111000000",
  38269=>"100000000",
  38270=>"000011111",
  38271=>"111011000",
  38272=>"000111111",
  38273=>"111001000",
  38274=>"111111011",
  38275=>"010011111",
  38276=>"000000010",
  38277=>"000010111",
  38278=>"111101111",
  38279=>"000000110",
  38280=>"000001111",
  38281=>"011010110",
  38282=>"111011111",
  38283=>"111111000",
  38284=>"111111111",
  38285=>"000111101",
  38286=>"111111111",
  38287=>"010000110",
  38288=>"001000000",
  38289=>"100000000",
  38290=>"011111000",
  38291=>"111001001",
  38292=>"011001111",
  38293=>"000000011",
  38294=>"000111111",
  38295=>"000000110",
  38296=>"000000000",
  38297=>"101001111",
  38298=>"111111001",
  38299=>"100000000",
  38300=>"111011000",
  38301=>"000000110",
  38302=>"000000000",
  38303=>"111111100",
  38304=>"111000000",
  38305=>"100111111",
  38306=>"011111101",
  38307=>"111011111",
  38308=>"111111011",
  38309=>"111001010",
  38310=>"000000001",
  38311=>"111111111",
  38312=>"000000000",
  38313=>"110111101",
  38314=>"111111111",
  38315=>"000000001",
  38316=>"000000000",
  38317=>"111010010",
  38318=>"111001111",
  38319=>"011011000",
  38320=>"000000000",
  38321=>"111111111",
  38322=>"101101000",
  38323=>"000110111",
  38324=>"111111100",
  38325=>"111111100",
  38326=>"010111111",
  38327=>"111001000",
  38328=>"000000000",
  38329=>"011011111",
  38330=>"000000000",
  38331=>"100010010",
  38332=>"111111111",
  38333=>"111111001",
  38334=>"000000000",
  38335=>"100101001",
  38336=>"111011001",
  38337=>"000000000",
  38338=>"111111111",
  38339=>"111000111",
  38340=>"000000000",
  38341=>"111001011",
  38342=>"111111111",
  38343=>"000000000",
  38344=>"110000000",
  38345=>"100110010",
  38346=>"000000001",
  38347=>"001001001",
  38348=>"000001001",
  38349=>"100000000",
  38350=>"111111111",
  38351=>"111111111",
  38352=>"111111111",
  38353=>"111111001",
  38354=>"000000000",
  38355=>"001000000",
  38356=>"000000000",
  38357=>"100100111",
  38358=>"001000000",
  38359=>"000001011",
  38360=>"001000000",
  38361=>"000000000",
  38362=>"100111111",
  38363=>"100010111",
  38364=>"000001011",
  38365=>"000111011",
  38366=>"000100111",
  38367=>"000000000",
  38368=>"000111011",
  38369=>"000000000",
  38370=>"011111111",
  38371=>"000000011",
  38372=>"000000001",
  38373=>"011011001",
  38374=>"010111110",
  38375=>"111100000",
  38376=>"011001001",
  38377=>"000000000",
  38378=>"100000011",
  38379=>"111111111",
  38380=>"000000000",
  38381=>"000000000",
  38382=>"000000000",
  38383=>"000100100",
  38384=>"001000001",
  38385=>"111111100",
  38386=>"111111000",
  38387=>"000000000",
  38388=>"110000000",
  38389=>"000111010",
  38390=>"111000000",
  38391=>"011000000",
  38392=>"000000000",
  38393=>"001000000",
  38394=>"000000000",
  38395=>"111111000",
  38396=>"000000111",
  38397=>"111101000",
  38398=>"000100000",
  38399=>"110010010",
  38400=>"111111010",
  38401=>"001000000",
  38402=>"000000000",
  38403=>"111010011",
  38404=>"000000011",
  38405=>"000000000",
  38406=>"000000000",
  38407=>"000000000",
  38408=>"010010011",
  38409=>"000000000",
  38410=>"100110111",
  38411=>"111111111",
  38412=>"001011111",
  38413=>"011000000",
  38414=>"000100111",
  38415=>"111111001",
  38416=>"000000001",
  38417=>"000000010",
  38418=>"100100000",
  38419=>"000000000",
  38420=>"011111011",
  38421=>"111111111",
  38422=>"000000011",
  38423=>"111111111",
  38424=>"111111111",
  38425=>"001011010",
  38426=>"001000000",
  38427=>"111111011",
  38428=>"111111111",
  38429=>"000001001",
  38430=>"011111111",
  38431=>"100010011",
  38432=>"000000111",
  38433=>"111101000",
  38434=>"000011011",
  38435=>"110110000",
  38436=>"111111111",
  38437=>"110110111",
  38438=>"111111111",
  38439=>"111111110",
  38440=>"111110000",
  38441=>"000000000",
  38442=>"000000000",
  38443=>"000000000",
  38444=>"000000000",
  38445=>"000000110",
  38446=>"111111111",
  38447=>"011001000",
  38448=>"000000000",
  38449=>"000000000",
  38450=>"111110100",
  38451=>"110110000",
  38452=>"001111000",
  38453=>"111010010",
  38454=>"000000000",
  38455=>"010010000",
  38456=>"001000010",
  38457=>"000000111",
  38458=>"111111111",
  38459=>"011111111",
  38460=>"000000000",
  38461=>"111111001",
  38462=>"000111011",
  38463=>"100100000",
  38464=>"100111010",
  38465=>"110111100",
  38466=>"000110100",
  38467=>"000100111",
  38468=>"111111111",
  38469=>"000000000",
  38470=>"111111111",
  38471=>"111111111",
  38472=>"001001000",
  38473=>"011000000",
  38474=>"111111111",
  38475=>"000000000",
  38476=>"000010010",
  38477=>"001011011",
  38478=>"000000000",
  38479=>"000000111",
  38480=>"000001011",
  38481=>"000000000",
  38482=>"000011111",
  38483=>"111111111",
  38484=>"000000000",
  38485=>"111110111",
  38486=>"001011000",
  38487=>"000000000",
  38488=>"000000000",
  38489=>"100101111",
  38490=>"000000000",
  38491=>"001001111",
  38492=>"100111111",
  38493=>"111111001",
  38494=>"111111111",
  38495=>"111111111",
  38496=>"101000000",
  38497=>"100110110",
  38498=>"111001001",
  38499=>"100000111",
  38500=>"000000100",
  38501=>"000010010",
  38502=>"000010000",
  38503=>"111101101",
  38504=>"111101111",
  38505=>"111011111",
  38506=>"000000000",
  38507=>"111111110",
  38508=>"000100100",
  38509=>"000000001",
  38510=>"111111111",
  38511=>"111110000",
  38512=>"111111000",
  38513=>"000000000",
  38514=>"111111111",
  38515=>"110111111",
  38516=>"110110000",
  38517=>"000000000",
  38518=>"001000001",
  38519=>"111111111",
  38520=>"000000000",
  38521=>"000000110",
  38522=>"111110111",
  38523=>"000100111",
  38524=>"110110110",
  38525=>"000000000",
  38526=>"100000011",
  38527=>"111000001",
  38528=>"000100000",
  38529=>"011111111",
  38530=>"001001001",
  38531=>"000000000",
  38532=>"000111110",
  38533=>"000000111",
  38534=>"110000111",
  38535=>"100100111",
  38536=>"111111111",
  38537=>"110110100",
  38538=>"100101111",
  38539=>"011000111",
  38540=>"111111111",
  38541=>"111111111",
  38542=>"010010000",
  38543=>"101111111",
  38544=>"000100110",
  38545=>"000000000",
  38546=>"100111111",
  38547=>"000110111",
  38548=>"000100110",
  38549=>"111111101",
  38550=>"000000000",
  38551=>"000000000",
  38552=>"000001011",
  38553=>"000000000",
  38554=>"111111111",
  38555=>"011101100",
  38556=>"111111111",
  38557=>"000000000",
  38558=>"011011111",
  38559=>"111111011",
  38560=>"000000000",
  38561=>"000000000",
  38562=>"111001111",
  38563=>"100111010",
  38564=>"000000000",
  38565=>"000111111",
  38566=>"111111111",
  38567=>"000000000",
  38568=>"111111000",
  38569=>"000000000",
  38570=>"000000000",
  38571=>"000000011",
  38572=>"000000000",
  38573=>"110110111",
  38574=>"000000100",
  38575=>"000000000",
  38576=>"111111111",
  38577=>"111111011",
  38578=>"111111111",
  38579=>"000000000",
  38580=>"111011000",
  38581=>"111111111",
  38582=>"001000000",
  38583=>"100110000",
  38584=>"101111111",
  38585=>"001000000",
  38586=>"000011011",
  38587=>"000000000",
  38588=>"111111111",
  38589=>"011011000",
  38590=>"000000000",
  38591=>"111111111",
  38592=>"000111111",
  38593=>"000001001",
  38594=>"111011111",
  38595=>"000000000",
  38596=>"000000000",
  38597=>"111100100",
  38598=>"111111111",
  38599=>"111111110",
  38600=>"000000000",
  38601=>"111111111",
  38602=>"000000110",
  38603=>"110111111",
  38604=>"000001011",
  38605=>"101101000",
  38606=>"100100100",
  38607=>"000100111",
  38608=>"111110011",
  38609=>"011000000",
  38610=>"000011011",
  38611=>"000000111",
  38612=>"000110110",
  38613=>"111111111",
  38614=>"000000000",
  38615=>"010110111",
  38616=>"111111111",
  38617=>"011011010",
  38618=>"000000000",
  38619=>"111111111",
  38620=>"111011001",
  38621=>"001011011",
  38622=>"111111000",
  38623=>"001101001",
  38624=>"011000001",
  38625=>"111101111",
  38626=>"100110111",
  38627=>"111111000",
  38628=>"110110010",
  38629=>"111111000",
  38630=>"000000000",
  38631=>"000001011",
  38632=>"111111111",
  38633=>"000000001",
  38634=>"111111111",
  38635=>"000000100",
  38636=>"110110111",
  38637=>"000000000",
  38638=>"110111111",
  38639=>"111001111",
  38640=>"000000000",
  38641=>"100100000",
  38642=>"001000101",
  38643=>"000000000",
  38644=>"111111110",
  38645=>"111111111",
  38646=>"001001011",
  38647=>"111111111",
  38648=>"110110110",
  38649=>"100000000",
  38650=>"000000000",
  38651=>"110110110",
  38652=>"111011011",
  38653=>"100000000",
  38654=>"000100000",
  38655=>"000011111",
  38656=>"011010000",
  38657=>"000100110",
  38658=>"111110110",
  38659=>"010000000",
  38660=>"111111100",
  38661=>"111011001",
  38662=>"000000110",
  38663=>"000001000",
  38664=>"000000000",
  38665=>"111101001",
  38666=>"110111111",
  38667=>"101100000",
  38668=>"000000110",
  38669=>"010000000",
  38670=>"111111111",
  38671=>"110000000",
  38672=>"000111111",
  38673=>"001001001",
  38674=>"000010011",
  38675=>"111111111",
  38676=>"111111111",
  38677=>"000000000",
  38678=>"000000001",
  38679=>"100111111",
  38680=>"110100000",
  38681=>"111000000",
  38682=>"000111111",
  38683=>"111000111",
  38684=>"111111111",
  38685=>"001001111",
  38686=>"000000000",
  38687=>"001001011",
  38688=>"000100000",
  38689=>"000000000",
  38690=>"000000000",
  38691=>"111110000",
  38692=>"001011001",
  38693=>"001111111",
  38694=>"000000011",
  38695=>"011111111",
  38696=>"111111111",
  38697=>"110000000",
  38698=>"000111111",
  38699=>"000000000",
  38700=>"111111100",
  38701=>"001011111",
  38702=>"111000111",
  38703=>"000000101",
  38704=>"000000000",
  38705=>"000101111",
  38706=>"000000110",
  38707=>"101000000",
  38708=>"000000000",
  38709=>"111111111",
  38710=>"000100111",
  38711=>"111011111",
  38712=>"000000000",
  38713=>"110111111",
  38714=>"000000000",
  38715=>"000000111",
  38716=>"000000000",
  38717=>"010011111",
  38718=>"000111111",
  38719=>"111111011",
  38720=>"000000000",
  38721=>"000000000",
  38722=>"000111011",
  38723=>"101101101",
  38724=>"000000000",
  38725=>"111000000",
  38726=>"111011111",
  38727=>"111111111",
  38728=>"000011000",
  38729=>"000000110",
  38730=>"111100000",
  38731=>"111100100",
  38732=>"000000000",
  38733=>"000011011",
  38734=>"001111110",
  38735=>"000000000",
  38736=>"111111101",
  38737=>"000000111",
  38738=>"000100111",
  38739=>"000000001",
  38740=>"111000011",
  38741=>"011011011",
  38742=>"000000111",
  38743=>"110000000",
  38744=>"111111011",
  38745=>"111100000",
  38746=>"010110111",
  38747=>"111111111",
  38748=>"011000000",
  38749=>"000000000",
  38750=>"000000111",
  38751=>"111111111",
  38752=>"001000100",
  38753=>"000000011",
  38754=>"011111101",
  38755=>"001111111",
  38756=>"000000000",
  38757=>"000000000",
  38758=>"000000100",
  38759=>"001111111",
  38760=>"001000110",
  38761=>"000000110",
  38762=>"000000011",
  38763=>"111111010",
  38764=>"001101111",
  38765=>"000100111",
  38766=>"111110010",
  38767=>"011111111",
  38768=>"111111111",
  38769=>"000000111",
  38770=>"111111111",
  38771=>"111111111",
  38772=>"000000000",
  38773=>"100111000",
  38774=>"000000000",
  38775=>"100111110",
  38776=>"000000000",
  38777=>"000000000",
  38778=>"000000000",
  38779=>"100110011",
  38780=>"010110111",
  38781=>"111110100",
  38782=>"000000110",
  38783=>"000000000",
  38784=>"000000100",
  38785=>"101000111",
  38786=>"001001000",
  38787=>"000000000",
  38788=>"011000011",
  38789=>"000000000",
  38790=>"111111110",
  38791=>"111110111",
  38792=>"000000010",
  38793=>"111111111",
  38794=>"111111111",
  38795=>"111111111",
  38796=>"111001111",
  38797=>"111111111",
  38798=>"000111011",
  38799=>"111111111",
  38800=>"000000000",
  38801=>"111111111",
  38802=>"011111111",
  38803=>"000000000",
  38804=>"110110111",
  38805=>"000000000",
  38806=>"000000000",
  38807=>"001000010",
  38808=>"000000001",
  38809=>"111110111",
  38810=>"000000000",
  38811=>"000000000",
  38812=>"100000000",
  38813=>"111111111",
  38814=>"111011000",
  38815=>"000010000",
  38816=>"111111000",
  38817=>"011000000",
  38818=>"000000000",
  38819=>"010110111",
  38820=>"000100110",
  38821=>"000000100",
  38822=>"111000000",
  38823=>"001111111",
  38824=>"011111100",
  38825=>"000000000",
  38826=>"101001001",
  38827=>"000000000",
  38828=>"000000000",
  38829=>"111111111",
  38830=>"001101100",
  38831=>"110111000",
  38832=>"111111110",
  38833=>"111001111",
  38834=>"110100000",
  38835=>"111111111",
  38836=>"000011001",
  38837=>"000000111",
  38838=>"000111110",
  38839=>"111000000",
  38840=>"010011011",
  38841=>"111111111",
  38842=>"111111111",
  38843=>"111111011",
  38844=>"100000000",
  38845=>"111111001",
  38846=>"000000010",
  38847=>"000000100",
  38848=>"110110111",
  38849=>"101111111",
  38850=>"000000110",
  38851=>"000000000",
  38852=>"000000000",
  38853=>"000000000",
  38854=>"111000000",
  38855=>"000000000",
  38856=>"000000000",
  38857=>"100111000",
  38858=>"001000111",
  38859=>"000010000",
  38860=>"000000011",
  38861=>"000000000",
  38862=>"000000000",
  38863=>"100100010",
  38864=>"111110100",
  38865=>"000000001",
  38866=>"000000000",
  38867=>"001001101",
  38868=>"000101111",
  38869=>"000111000",
  38870=>"000000111",
  38871=>"100100000",
  38872=>"000010000",
  38873=>"000000000",
  38874=>"001011001",
  38875=>"111110000",
  38876=>"000000010",
  38877=>"011010000",
  38878=>"111111111",
  38879=>"001001111",
  38880=>"100100100",
  38881=>"111111100",
  38882=>"111111100",
  38883=>"011011000",
  38884=>"110111000",
  38885=>"111101111",
  38886=>"010110110",
  38887=>"000010000",
  38888=>"111111011",
  38889=>"000000010",
  38890=>"111111000",
  38891=>"111111111",
  38892=>"000001111",
  38893=>"010000000",
  38894=>"000000000",
  38895=>"100111111",
  38896=>"000000111",
  38897=>"111111111",
  38898=>"111110111",
  38899=>"111111110",
  38900=>"111111111",
  38901=>"001000000",
  38902=>"111111001",
  38903=>"100000000",
  38904=>"000111111",
  38905=>"000110100",
  38906=>"000000001",
  38907=>"000000111",
  38908=>"111111000",
  38909=>"100100100",
  38910=>"000000000",
  38911=>"101101100",
  38912=>"000000000",
  38913=>"111111110",
  38914=>"000000111",
  38915=>"000000100",
  38916=>"000000000",
  38917=>"001000111",
  38918=>"000000000",
  38919=>"111111111",
  38920=>"010000000",
  38921=>"000000111",
  38922=>"000000000",
  38923=>"000000100",
  38924=>"000110010",
  38925=>"100000000",
  38926=>"011001001",
  38927=>"110111000",
  38928=>"111111110",
  38929=>"001001111",
  38930=>"000000000",
  38931=>"000000000",
  38932=>"111111000",
  38933=>"100101111",
  38934=>"111000000",
  38935=>"010111001",
  38936=>"111111111",
  38937=>"001001111",
  38938=>"000000000",
  38939=>"000000000",
  38940=>"000111111",
  38941=>"111111000",
  38942=>"000000011",
  38943=>"111111111",
  38944=>"011011000",
  38945=>"111111100",
  38946=>"100000001",
  38947=>"000000000",
  38948=>"011011000",
  38949=>"110111111",
  38950=>"111100000",
  38951=>"000000000",
  38952=>"000000111",
  38953=>"100000110",
  38954=>"000111111",
  38955=>"111110100",
  38956=>"000111111",
  38957=>"000110111",
  38958=>"001001000",
  38959=>"000000010",
  38960=>"000000000",
  38961=>"011111111",
  38962=>"000000000",
  38963=>"111111111",
  38964=>"000111111",
  38965=>"111111111",
  38966=>"010111111",
  38967=>"000001111",
  38968=>"000000001",
  38969=>"110000000",
  38970=>"000110111",
  38971=>"000000000",
  38972=>"000100111",
  38973=>"001000000",
  38974=>"111111011",
  38975=>"001000000",
  38976=>"000000000",
  38977=>"000000000",
  38978=>"000110110",
  38979=>"111111011",
  38980=>"000011000",
  38981=>"111111111",
  38982=>"000000101",
  38983=>"101111111",
  38984=>"000000011",
  38985=>"000000110",
  38986=>"111000000",
  38987=>"011011111",
  38988=>"111110100",
  38989=>"000000111",
  38990=>"110000000",
  38991=>"111111111",
  38992=>"111111010",
  38993=>"000000011",
  38994=>"100111111",
  38995=>"110100111",
  38996=>"000000000",
  38997=>"000001001",
  38998=>"101000000",
  38999=>"111111111",
  39000=>"110111000",
  39001=>"111000000",
  39002=>"101000100",
  39003=>"111110000",
  39004=>"111111111",
  39005=>"000111001",
  39006=>"000000110",
  39007=>"000001110",
  39008=>"000000000",
  39009=>"110111110",
  39010=>"111111111",
  39011=>"101000111",
  39012=>"000001001",
  39013=>"001011111",
  39014=>"111001000",
  39015=>"000000000",
  39016=>"000000111",
  39017=>"111111111",
  39018=>"111111001",
  39019=>"001011111",
  39020=>"111111111",
  39021=>"111000000",
  39022=>"111011111",
  39023=>"000000100",
  39024=>"111001111",
  39025=>"000000111",
  39026=>"001111000",
  39027=>"110100101",
  39028=>"000000000",
  39029=>"111111110",
  39030=>"000000011",
  39031=>"000000000",
  39032=>"000000000",
  39033=>"000000000",
  39034=>"000000000",
  39035=>"000000000",
  39036=>"110111011",
  39037=>"000101100",
  39038=>"111111000",
  39039=>"110100100",
  39040=>"111011000",
  39041=>"111111101",
  39042=>"111011001",
  39043=>"001001001",
  39044=>"000000110",
  39045=>"001000001",
  39046=>"111111110",
  39047=>"111000000",
  39048=>"000000000",
  39049=>"000000000",
  39050=>"110110000",
  39051=>"000000001",
  39052=>"000000000",
  39053=>"111111111",
  39054=>"000000111",
  39055=>"000111111",
  39056=>"000111111",
  39057=>"010110110",
  39058=>"111001000",
  39059=>"111111111",
  39060=>"111111000",
  39061=>"000111111",
  39062=>"011000000",
  39063=>"111000011",
  39064=>"000000000",
  39065=>"000001101",
  39066=>"000000000",
  39067=>"000000000",
  39068=>"101000000",
  39069=>"111001000",
  39070=>"111111000",
  39071=>"110110000",
  39072=>"111111110",
  39073=>"111000000",
  39074=>"000001111",
  39075=>"000000000",
  39076=>"111001001",
  39077=>"111001000",
  39078=>"111111111",
  39079=>"111111111",
  39080=>"111111111",
  39081=>"100100111",
  39082=>"000000000",
  39083=>"001000000",
  39084=>"111111110",
  39085=>"000000100",
  39086=>"010110010",
  39087=>"000100111",
  39088=>"111010110",
  39089=>"100100000",
  39090=>"111111110",
  39091=>"010000000",
  39092=>"000000000",
  39093=>"111111000",
  39094=>"110111000",
  39095=>"100000100",
  39096=>"101000000",
  39097=>"000000111",
  39098=>"100100100",
  39099=>"000000000",
  39100=>"011000100",
  39101=>"110110000",
  39102=>"111011000",
  39103=>"000000000",
  39104=>"000000111",
  39105=>"000000000",
  39106=>"000001000",
  39107=>"110000001",
  39108=>"000100111",
  39109=>"000000111",
  39110=>"111111111",
  39111=>"000000111",
  39112=>"000000000",
  39113=>"101111111",
  39114=>"000000000",
  39115=>"000001001",
  39116=>"100000101",
  39117=>"100000111",
  39118=>"111111111",
  39119=>"001001111",
  39120=>"000000000",
  39121=>"110111000",
  39122=>"000000000",
  39123=>"000000000",
  39124=>"101001001",
  39125=>"111001000",
  39126=>"000000000",
  39127=>"000111011",
  39128=>"000001111",
  39129=>"010000000",
  39130=>"000000111",
  39131=>"000000111",
  39132=>"111001000",
  39133=>"001000000",
  39134=>"010010111",
  39135=>"000000011",
  39136=>"111111000",
  39137=>"000100111",
  39138=>"111000101",
  39139=>"000000000",
  39140=>"001011000",
  39141=>"000000001",
  39142=>"111010111",
  39143=>"000000000",
  39144=>"000111110",
  39145=>"111010001",
  39146=>"111110100",
  39147=>"100000100",
  39148=>"000000000",
  39149=>"111000000",
  39150=>"111111111",
  39151=>"000000000",
  39152=>"000000000",
  39153=>"111111111",
  39154=>"111000000",
  39155=>"001000000",
  39156=>"000101111",
  39157=>"000000001",
  39158=>"001111111",
  39159=>"111000111",
  39160=>"111111100",
  39161=>"111111001",
  39162=>"111000000",
  39163=>"010010000",
  39164=>"110111101",
  39165=>"111000111",
  39166=>"111111100",
  39167=>"000111111",
  39168=>"101000110",
  39169=>"100100100",
  39170=>"100100111",
  39171=>"000000100",
  39172=>"111111111",
  39173=>"000011000",
  39174=>"000000000",
  39175=>"111011001",
  39176=>"111100100",
  39177=>"000100111",
  39178=>"001000000",
  39179=>"000000000",
  39180=>"101101111",
  39181=>"011101001",
  39182=>"111100110",
  39183=>"111111010",
  39184=>"011111000",
  39185=>"000000111",
  39186=>"010111111",
  39187=>"111010000",
  39188=>"000100000",
  39189=>"111001110",
  39190=>"000000111",
  39191=>"000001111",
  39192=>"000000011",
  39193=>"000011111",
  39194=>"111111111",
  39195=>"000000000",
  39196=>"000111111",
  39197=>"001000000",
  39198=>"000111111",
  39199=>"000000111",
  39200=>"000001011",
  39201=>"111111000",
  39202=>"100000000",
  39203=>"001001111",
  39204=>"101100100",
  39205=>"111001001",
  39206=>"000001001",
  39207=>"111100111",
  39208=>"001000000",
  39209=>"000111000",
  39210=>"111111111",
  39211=>"111111011",
  39212=>"000000100",
  39213=>"001001001",
  39214=>"000000000",
  39215=>"000000111",
  39216=>"000000110",
  39217=>"000000111",
  39218=>"000000000",
  39219=>"000111000",
  39220=>"111000000",
  39221=>"111110000",
  39222=>"111111110",
  39223=>"111111111",
  39224=>"000000111",
  39225=>"111000001",
  39226=>"111001000",
  39227=>"111111011",
  39228=>"101100101",
  39229=>"101101100",
  39230=>"100111111",
  39231=>"111111110",
  39232=>"111000000",
  39233=>"111110000",
  39234=>"011110110",
  39235=>"111111111",
  39236=>"000010100",
  39237=>"000001111",
  39238=>"110111000",
  39239=>"000000000",
  39240=>"111111110",
  39241=>"111111000",
  39242=>"011111000",
  39243=>"111111101",
  39244=>"011111100",
  39245=>"100111111",
  39246=>"111100000",
  39247=>"000111111",
  39248=>"111111111",
  39249=>"000000111",
  39250=>"110010111",
  39251=>"000111111",
  39252=>"100111000",
  39253=>"001011011",
  39254=>"111011000",
  39255=>"111111111",
  39256=>"111111111",
  39257=>"000000000",
  39258=>"100110110",
  39259=>"001000000",
  39260=>"001001001",
  39261=>"000110111",
  39262=>"000000111",
  39263=>"000111111",
  39264=>"000000011",
  39265=>"001111111",
  39266=>"110100111",
  39267=>"111111111",
  39268=>"100101001",
  39269=>"111111111",
  39270=>"111000000",
  39271=>"011011111",
  39272=>"111111111",
  39273=>"111000000",
  39274=>"111111000",
  39275=>"101000000",
  39276=>"000000110",
  39277=>"111111000",
  39278=>"000000000",
  39279=>"111111111",
  39280=>"100111111",
  39281=>"111110000",
  39282=>"101001100",
  39283=>"110000000",
  39284=>"000000000",
  39285=>"000110110",
  39286=>"001001101",
  39287=>"000000111",
  39288=>"000000110",
  39289=>"000101111",
  39290=>"111111111",
  39291=>"111011001",
  39292=>"111111000",
  39293=>"111001000",
  39294=>"010011111",
  39295=>"111111111",
  39296=>"000000000",
  39297=>"000111111",
  39298=>"110111111",
  39299=>"001111111",
  39300=>"100000000",
  39301=>"000111100",
  39302=>"110111111",
  39303=>"011011111",
  39304=>"000110111",
  39305=>"100000111",
  39306=>"000000000",
  39307=>"011000000",
  39308=>"001000111",
  39309=>"001001111",
  39310=>"000001000",
  39311=>"111111111",
  39312=>"110110111",
  39313=>"000000001",
  39314=>"000000011",
  39315=>"110111011",
  39316=>"111000000",
  39317=>"000000000",
  39318=>"000000111",
  39319=>"000000001",
  39320=>"000111111",
  39321=>"101011000",
  39322=>"111000000",
  39323=>"000111111",
  39324=>"111111001",
  39325=>"000111111",
  39326=>"111000001",
  39327=>"000000101",
  39328=>"000000111",
  39329=>"100111111",
  39330=>"101001001",
  39331=>"111001001",
  39332=>"111000000",
  39333=>"000111110",
  39334=>"000000001",
  39335=>"000000000",
  39336=>"000100000",
  39337=>"000000111",
  39338=>"011001101",
  39339=>"111111111",
  39340=>"111111111",
  39341=>"000000000",
  39342=>"000000111",
  39343=>"111111111",
  39344=>"111111000",
  39345=>"111111111",
  39346=>"111111111",
  39347=>"101000000",
  39348=>"000000000",
  39349=>"111000000",
  39350=>"111111111",
  39351=>"001011010",
  39352=>"111001000",
  39353=>"111000000",
  39354=>"000000111",
  39355=>"010111110",
  39356=>"101001001",
  39357=>"001000000",
  39358=>"000000000",
  39359=>"100000001",
  39360=>"111000000",
  39361=>"111000000",
  39362=>"000101101",
  39363=>"111111100",
  39364=>"001101100",
  39365=>"111001001",
  39366=>"111000000",
  39367=>"000110111",
  39368=>"000000000",
  39369=>"000000001",
  39370=>"101111101",
  39371=>"111111111",
  39372=>"111000000",
  39373=>"001000011",
  39374=>"100000100",
  39375=>"111110000",
  39376=>"000000111",
  39377=>"101100000",
  39378=>"000011111",
  39379=>"111111111",
  39380=>"000011111",
  39381=>"000000000",
  39382=>"111111000",
  39383=>"000000000",
  39384=>"101101000",
  39385=>"011000000",
  39386=>"000110100",
  39387=>"000000000",
  39388=>"000111111",
  39389=>"111111001",
  39390=>"111011111",
  39391=>"100100000",
  39392=>"111000001",
  39393=>"011100110",
  39394=>"000000110",
  39395=>"011000001",
  39396=>"001100111",
  39397=>"000000100",
  39398=>"000111111",
  39399=>"111011111",
  39400=>"000000000",
  39401=>"111000000",
  39402=>"000000000",
  39403=>"111111111",
  39404=>"111111111",
  39405=>"001000000",
  39406=>"000111111",
  39407=>"111000111",
  39408=>"111111111",
  39409=>"111111111",
  39410=>"000000000",
  39411=>"000000000",
  39412=>"001000000",
  39413=>"110000110",
  39414=>"110100000",
  39415=>"111001111",
  39416=>"111001000",
  39417=>"001001101",
  39418=>"110111011",
  39419=>"001000000",
  39420=>"001000000",
  39421=>"100100111",
  39422=>"001000111",
  39423=>"000000011",
  39424=>"000000001",
  39425=>"111111111",
  39426=>"111000000",
  39427=>"111001000",
  39428=>"011001101",
  39429=>"000000001",
  39430=>"000000000",
  39431=>"111111111",
  39432=>"000111110",
  39433=>"111000000",
  39434=>"011001000",
  39435=>"111111111",
  39436=>"111111111",
  39437=>"000000000",
  39438=>"011011011",
  39439=>"010110111",
  39440=>"110111111",
  39441=>"000100111",
  39442=>"001101111",
  39443=>"000011111",
  39444=>"010000000",
  39445=>"001101000",
  39446=>"111111111",
  39447=>"110111111",
  39448=>"111001011",
  39449=>"100100000",
  39450=>"011011001",
  39451=>"111011000",
  39452=>"111101001",
  39453=>"011000000",
  39454=>"000001011",
  39455=>"000000111",
  39456=>"000000111",
  39457=>"000000000",
  39458=>"000000000",
  39459=>"101000000",
  39460=>"011011000",
  39461=>"011001001",
  39462=>"000000110",
  39463=>"011111110",
  39464=>"111101111",
  39465=>"011010000",
  39466=>"111111111",
  39467=>"110111011",
  39468=>"000000000",
  39469=>"100000001",
  39470=>"100110110",
  39471=>"001000011",
  39472=>"000000000",
  39473=>"111101111",
  39474=>"111111111",
  39475=>"001001001",
  39476=>"000110111",
  39477=>"000000000",
  39478=>"111111111",
  39479=>"000000000",
  39480=>"000000000",
  39481=>"111011000",
  39482=>"111111011",
  39483=>"111111111",
  39484=>"111110110",
  39485=>"001001001",
  39486=>"000000100",
  39487=>"000000001",
  39488=>"110111011",
  39489=>"000110110",
  39490=>"001000000",
  39491=>"010011111",
  39492=>"110110110",
  39493=>"000001111",
  39494=>"111011000",
  39495=>"111111110",
  39496=>"011001011",
  39497=>"111111110",
  39498=>"000000000",
  39499=>"111111111",
  39500=>"000000100",
  39501=>"100110000",
  39502=>"111111100",
  39503=>"111111000",
  39504=>"100110000",
  39505=>"000000000",
  39506=>"111111111",
  39507=>"001111111",
  39508=>"000000001",
  39509=>"010111001",
  39510=>"000000000",
  39511=>"100000000",
  39512=>"000000001",
  39513=>"111111111",
  39514=>"011111110",
  39515=>"110010000",
  39516=>"100000000",
  39517=>"000000011",
  39518=>"110110000",
  39519=>"110100001",
  39520=>"101111110",
  39521=>"000010100",
  39522=>"111111011",
  39523=>"111111110",
  39524=>"111010000",
  39525=>"111101101",
  39526=>"010000000",
  39527=>"111111111",
  39528=>"111100000",
  39529=>"000000001",
  39530=>"011011010",
  39531=>"000000110",
  39532=>"100000000",
  39533=>"000000000",
  39534=>"000000000",
  39535=>"111111111",
  39536=>"000000001",
  39537=>"100100101",
  39538=>"100100110",
  39539=>"100001111",
  39540=>"000001001",
  39541=>"100100110",
  39542=>"110111010",
  39543=>"000000000",
  39544=>"100100101",
  39545=>"011001011",
  39546=>"000000001",
  39547=>"111111111",
  39548=>"110110110",
  39549=>"100000000",
  39550=>"110111111",
  39551=>"000000100",
  39552=>"000000000",
  39553=>"110000000",
  39554=>"111111111",
  39555=>"110111100",
  39556=>"000000000",
  39557=>"011011111",
  39558=>"001000000",
  39559=>"110000000",
  39560=>"111001111",
  39561=>"000000001",
  39562=>"110111110",
  39563=>"000100011",
  39564=>"011011011",
  39565=>"000000000",
  39566=>"110111111",
  39567=>"111110110",
  39568=>"111111111",
  39569=>"111111110",
  39570=>"111010011",
  39571=>"000000000",
  39572=>"000000000",
  39573=>"010111111",
  39574=>"111111010",
  39575=>"000000000",
  39576=>"100000000",
  39577=>"111111111",
  39578=>"101100100",
  39579=>"011010010",
  39580=>"110000000",
  39581=>"100001000",
  39582=>"111111111",
  39583=>"000110110",
  39584=>"000000000",
  39585=>"010000000",
  39586=>"111111001",
  39587=>"110111111",
  39588=>"100110111",
  39589=>"010000000",
  39590=>"110111111",
  39591=>"000000010",
  39592=>"000011001",
  39593=>"100110111",
  39594=>"111111111",
  39595=>"000000000",
  39596=>"000110110",
  39597=>"101111000",
  39598=>"111111111",
  39599=>"011011011",
  39600=>"000000111",
  39601=>"001101101",
  39602=>"111111111",
  39603=>"000000000",
  39604=>"000001111",
  39605=>"000000000",
  39606=>"111000000",
  39607=>"111111000",
  39608=>"000001111",
  39609=>"111101111",
  39610=>"000111101",
  39611=>"110110000",
  39612=>"000010011",
  39613=>"000000000",
  39614=>"111111011",
  39615=>"011001001",
  39616=>"111110000",
  39617=>"111000000",
  39618=>"000000000",
  39619=>"000000000",
  39620=>"000000000",
  39621=>"000000000",
  39622=>"111000000",
  39623=>"111111000",
  39624=>"000000000",
  39625=>"111111111",
  39626=>"101001011",
  39627=>"111111001",
  39628=>"000100100",
  39629=>"000111111",
  39630=>"110110110",
  39631=>"000000111",
  39632=>"000000000",
  39633=>"000001000",
  39634=>"111111011",
  39635=>"111111111",
  39636=>"111000001",
  39637=>"000000000",
  39638=>"001000001",
  39639=>"010111001",
  39640=>"000000000",
  39641=>"000000000",
  39642=>"011000111",
  39643=>"000111011",
  39644=>"111001011",
  39645=>"101100000",
  39646=>"000000000",
  39647=>"110101111",
  39648=>"000000000",
  39649=>"111111111",
  39650=>"000000111",
  39651=>"010111111",
  39652=>"110100000",
  39653=>"010111000",
  39654=>"011011000",
  39655=>"000000001",
  39656=>"111111111",
  39657=>"000000101",
  39658=>"000000001",
  39659=>"111111111",
  39660=>"111111111",
  39661=>"011111011",
  39662=>"111111111",
  39663=>"000000000",
  39664=>"001000001",
  39665=>"100110111",
  39666=>"011111111",
  39667=>"111101111",
  39668=>"110111111",
  39669=>"000000001",
  39670=>"111001111",
  39671=>"000100100",
  39672=>"001001111",
  39673=>"111111111",
  39674=>"000000000",
  39675=>"000000110",
  39676=>"001001111",
  39677=>"001000000",
  39678=>"000010000",
  39679=>"011100111",
  39680=>"000000000",
  39681=>"110111111",
  39682=>"111111111",
  39683=>"111111111",
  39684=>"000000000",
  39685=>"000000000",
  39686=>"011111010",
  39687=>"000011111",
  39688=>"000010000",
  39689=>"000111111",
  39690=>"111011000",
  39691=>"111111111",
  39692=>"111111111",
  39693=>"000000000",
  39694=>"111001000",
  39695=>"000110111",
  39696=>"111111111",
  39697=>"000000000",
  39698=>"001111111",
  39699=>"001000000",
  39700=>"011011001",
  39701=>"001001000",
  39702=>"000000000",
  39703=>"000001001",
  39704=>"110110000",
  39705=>"000000001",
  39706=>"111000110",
  39707=>"000010011",
  39708=>"100100100",
  39709=>"111111001",
  39710=>"110111111",
  39711=>"110110000",
  39712=>"000000000",
  39713=>"000000000",
  39714=>"001001000",
  39715=>"111111111",
  39716=>"000110000",
  39717=>"100000001",
  39718=>"000000101",
  39719=>"001000110",
  39720=>"111001011",
  39721=>"111111111",
  39722=>"111000010",
  39723=>"111111111",
  39724=>"001011000",
  39725=>"100100000",
  39726=>"111111000",
  39727=>"111111111",
  39728=>"110111111",
  39729=>"000000000",
  39730=>"000000000",
  39731=>"011011011",
  39732=>"000011000",
  39733=>"100110111",
  39734=>"000000001",
  39735=>"000111111",
  39736=>"001100100",
  39737=>"111111111",
  39738=>"010010000",
  39739=>"011000001",
  39740=>"000000001",
  39741=>"110110000",
  39742=>"000000001",
  39743=>"000000001",
  39744=>"000011111",
  39745=>"110000010",
  39746=>"111111001",
  39747=>"000000000",
  39748=>"111111110",
  39749=>"000000000",
  39750=>"000000000",
  39751=>"101101001",
  39752=>"000000000",
  39753=>"010010000",
  39754=>"001000010",
  39755=>"000100100",
  39756=>"010010010",
  39757=>"000000000",
  39758=>"111111101",
  39759=>"011111101",
  39760=>"000110111",
  39761=>"000000100",
  39762=>"000010000",
  39763=>"000000000",
  39764=>"111111111",
  39765=>"011011011",
  39766=>"010010011",
  39767=>"000111111",
  39768=>"000000000",
  39769=>"001001000",
  39770=>"111011000",
  39771=>"110111001",
  39772=>"000000000",
  39773=>"111011111",
  39774=>"111111111",
  39775=>"000000000",
  39776=>"111111111",
  39777=>"111111101",
  39778=>"000100100",
  39779=>"000100100",
  39780=>"001001111",
  39781=>"000000000",
  39782=>"011000000",
  39783=>"101001001",
  39784=>"000011001",
  39785=>"100000000",
  39786=>"111111000",
  39787=>"011011111",
  39788=>"110000001",
  39789=>"000011111",
  39790=>"111111111",
  39791=>"110010010",
  39792=>"110110100",
  39793=>"010111111",
  39794=>"000000000",
  39795=>"111011000",
  39796=>"110111101",
  39797=>"100000000",
  39798=>"100001111",
  39799=>"000001001",
  39800=>"111000000",
  39801=>"000010000",
  39802=>"111011000",
  39803=>"001001011",
  39804=>"000000010",
  39805=>"111111111",
  39806=>"000111111",
  39807=>"100000101",
  39808=>"011011011",
  39809=>"110111111",
  39810=>"101111111",
  39811=>"010111111",
  39812=>"000110111",
  39813=>"000000100",
  39814=>"111111111",
  39815=>"000111111",
  39816=>"000000000",
  39817=>"000000000",
  39818=>"111100111",
  39819=>"111111111",
  39820=>"000000111",
  39821=>"001001110",
  39822=>"011111111",
  39823=>"000010011",
  39824=>"010010000",
  39825=>"110111110",
  39826=>"111111010",
  39827=>"100100100",
  39828=>"000100111",
  39829=>"111100111",
  39830=>"111111111",
  39831=>"010010000",
  39832=>"111111001",
  39833=>"100100001",
  39834=>"000001011",
  39835=>"000000111",
  39836=>"110101111",
  39837=>"111111111",
  39838=>"111101001",
  39839=>"000011001",
  39840=>"010000000",
  39841=>"111111111",
  39842=>"011001000",
  39843=>"000000000",
  39844=>"000000000",
  39845=>"101111111",
  39846=>"111010000",
  39847=>"010011111",
  39848=>"000000000",
  39849=>"000000000",
  39850=>"000000000",
  39851=>"000000000",
  39852=>"111111111",
  39853=>"000111111",
  39854=>"000110110",
  39855=>"000000000",
  39856=>"111111111",
  39857=>"000000000",
  39858=>"100100000",
  39859=>"001000100",
  39860=>"010011000",
  39861=>"000110110",
  39862=>"000000100",
  39863=>"000010000",
  39864=>"000000000",
  39865=>"000011000",
  39866=>"100000001",
  39867=>"000000000",
  39868=>"000000000",
  39869=>"111101001",
  39870=>"111111000",
  39871=>"110110010",
  39872=>"000000000",
  39873=>"000000000",
  39874=>"000000000",
  39875=>"111111111",
  39876=>"001000000",
  39877=>"000011111",
  39878=>"111111111",
  39879=>"110111111",
  39880=>"000111111",
  39881=>"110000000",
  39882=>"111111111",
  39883=>"111000101",
  39884=>"010000000",
  39885=>"000000000",
  39886=>"100111001",
  39887=>"110110111",
  39888=>"111110110",
  39889=>"111111011",
  39890=>"000010110",
  39891=>"000000101",
  39892=>"011111011",
  39893=>"110111110",
  39894=>"000000111",
  39895=>"001001111",
  39896=>"100100111",
  39897=>"110000100",
  39898=>"000001001",
  39899=>"110110000",
  39900=>"001011111",
  39901=>"111111011",
  39902=>"111001000",
  39903=>"000110111",
  39904=>"111111111",
  39905=>"001000000",
  39906=>"011111110",
  39907=>"010011001",
  39908=>"011111111",
  39909=>"011001011",
  39910=>"100110010",
  39911=>"000111111",
  39912=>"001000111",
  39913=>"000000001",
  39914=>"011011011",
  39915=>"101101100",
  39916=>"001000000",
  39917=>"000110000",
  39918=>"111110110",
  39919=>"110111011",
  39920=>"001000000",
  39921=>"011111111",
  39922=>"111111011",
  39923=>"000111110",
  39924=>"001001001",
  39925=>"000000001",
  39926=>"001111111",
  39927=>"111101111",
  39928=>"000101111",
  39929=>"010010110",
  39930=>"001001111",
  39931=>"000010000",
  39932=>"111100000",
  39933=>"000100111",
  39934=>"111111000",
  39935=>"000101111",
  39936=>"110111101",
  39937=>"111111111",
  39938=>"111111111",
  39939=>"111111111",
  39940=>"110011111",
  39941=>"110010110",
  39942=>"000111000",
  39943=>"110000111",
  39944=>"111111001",
  39945=>"111111111",
  39946=>"001111111",
  39947=>"001000000",
  39948=>"000111011",
  39949=>"111110100",
  39950=>"011000000",
  39951=>"000000000",
  39952=>"111111000",
  39953=>"000001101",
  39954=>"111111000",
  39955=>"000000000",
  39956=>"010111111",
  39957=>"110111111",
  39958=>"110000000",
  39959=>"011111000",
  39960=>"011011111",
  39961=>"001011111",
  39962=>"000011111",
  39963=>"001111111",
  39964=>"110000000",
  39965=>"001001000",
  39966=>"011110100",
  39967=>"111111110",
  39968=>"001000000",
  39969=>"000000001",
  39970=>"000100100",
  39971=>"111110010",
  39972=>"111000000",
  39973=>"111110000",
  39974=>"101000000",
  39975=>"100000000",
  39976=>"000000000",
  39977=>"001111111",
  39978=>"000000111",
  39979=>"000111111",
  39980=>"111111101",
  39981=>"101101001",
  39982=>"001000000",
  39983=>"000000000",
  39984=>"000000000",
  39985=>"000000000",
  39986=>"001111111",
  39987=>"010000000",
  39988=>"111001000",
  39989=>"000000001",
  39990=>"011001000",
  39991=>"001110000",
  39992=>"110111111",
  39993=>"110110111",
  39994=>"011101111",
  39995=>"000000000",
  39996=>"000000101",
  39997=>"000000001",
  39998=>"000000010",
  39999=>"111111111",
  40000=>"011001110",
  40001=>"101101101",
  40002=>"000101111",
  40003=>"010000000",
  40004=>"000011111",
  40005=>"111100110",
  40006=>"111111101",
  40007=>"000000111",
  40008=>"000000000",
  40009=>"111000000",
  40010=>"000000000",
  40011=>"000000000",
  40012=>"111011111",
  40013=>"000000111",
  40014=>"000000000",
  40015=>"111111111",
  40016=>"010111111",
  40017=>"111011000",
  40018=>"111001000",
  40019=>"110000011",
  40020=>"101000000",
  40021=>"111111000",
  40022=>"111111111",
  40023=>"100000000",
  40024=>"011000000",
  40025=>"111100000",
  40026=>"111111001",
  40027=>"100110110",
  40028=>"011110111",
  40029=>"101000000",
  40030=>"010000111",
  40031=>"000000001",
  40032=>"001001000",
  40033=>"000011101",
  40034=>"111111111",
  40035=>"000000000",
  40036=>"000111111",
  40037=>"000000110",
  40038=>"000000000",
  40039=>"111110000",
  40040=>"011111111",
  40041=>"000000000",
  40042=>"111111111",
  40043=>"000000000",
  40044=>"111100000",
  40045=>"100100000",
  40046=>"111000101",
  40047=>"011101000",
  40048=>"001000000",
  40049=>"000000000",
  40050=>"100100101",
  40051=>"000000001",
  40052=>"111111000",
  40053=>"000000000",
  40054=>"000000111",
  40055=>"111001000",
  40056=>"011111111",
  40057=>"000000011",
  40058=>"111100000",
  40059=>"000000000",
  40060=>"001001000",
  40061=>"000000000",
  40062=>"111111110",
  40063=>"000000000",
  40064=>"111111101",
  40065=>"111000000",
  40066=>"111011001",
  40067=>"111100000",
  40068=>"000111111",
  40069=>"111101000",
  40070=>"010010010",
  40071=>"001000000",
  40072=>"001001001",
  40073=>"001000010",
  40074=>"001000000",
  40075=>"111001000",
  40076=>"000111111",
  40077=>"111111111",
  40078=>"110100110",
  40079=>"000111000",
  40080=>"001101101",
  40081=>"000000000",
  40082=>"001000000",
  40083=>"111111000",
  40084=>"111111000",
  40085=>"000000000",
  40086=>"110110110",
  40087=>"111100111",
  40088=>"000101111",
  40089=>"000000000",
  40090=>"001001111",
  40091=>"111101111",
  40092=>"010111111",
  40093=>"111100101",
  40094=>"000000001",
  40095=>"111010000",
  40096=>"000000000",
  40097=>"000011001",
  40098=>"000000000",
  40099=>"111111100",
  40100=>"000111111",
  40101=>"000001000",
  40102=>"001111111",
  40103=>"100100100",
  40104=>"001000111",
  40105=>"111111000",
  40106=>"110000000",
  40107=>"101001000",
  40108=>"111111111",
  40109=>"011011111",
  40110=>"110100111",
  40111=>"011000000",
  40112=>"001111101",
  40113=>"100110111",
  40114=>"101101001",
  40115=>"001000000",
  40116=>"000000100",
  40117=>"100000100",
  40118=>"000000000",
  40119=>"111111111",
  40120=>"111111111",
  40121=>"111111000",
  40122=>"111000000",
  40123=>"111111111",
  40124=>"100000000",
  40125=>"111111111",
  40126=>"111000100",
  40127=>"001001000",
  40128=>"111111000",
  40129=>"111111111",
  40130=>"000000000",
  40131=>"111111011",
  40132=>"111111111",
  40133=>"111111011",
  40134=>"011001000",
  40135=>"000000000",
  40136=>"100000111",
  40137=>"000000000",
  40138=>"000000000",
  40139=>"100100111",
  40140=>"011110010",
  40141=>"000100111",
  40142=>"001011011",
  40143=>"011000001",
  40144=>"111111000",
  40145=>"001000000",
  40146=>"111111000",
  40147=>"000001000",
  40148=>"000000000",
  40149=>"110110110",
  40150=>"111111111",
  40151=>"000000000",
  40152=>"000000000",
  40153=>"000000101",
  40154=>"111111111",
  40155=>"111111111",
  40156=>"000000101",
  40157=>"000110111",
  40158=>"000000111",
  40159=>"111111111",
  40160=>"000001111",
  40161=>"001001001",
  40162=>"000000000",
  40163=>"001011000",
  40164=>"000000000",
  40165=>"100111111",
  40166=>"110000110",
  40167=>"000111110",
  40168=>"111111111",
  40169=>"000000001",
  40170=>"000000101",
  40171=>"000111111",
  40172=>"011111111",
  40173=>"111000000",
  40174=>"000000001",
  40175=>"111111111",
  40176=>"100111011",
  40177=>"000111111",
  40178=>"111000000",
  40179=>"001111111",
  40180=>"010111111",
  40181=>"000000110",
  40182=>"111111000",
  40183=>"111010000",
  40184=>"000111000",
  40185=>"110111111",
  40186=>"000000000",
  40187=>"000000111",
  40188=>"001001111",
  40189=>"010000001",
  40190=>"111101000",
  40191=>"111111011",
  40192=>"111010001",
  40193=>"100111101",
  40194=>"111110000",
  40195=>"000000101",
  40196=>"111000000",
  40197=>"000101101",
  40198=>"111111111",
  40199=>"000000000",
  40200=>"001110111",
  40201=>"111000000",
  40202=>"111111111",
  40203=>"000000111",
  40204=>"101001101",
  40205=>"001000111",
  40206=>"000000111",
  40207=>"000100000",
  40208=>"010000000",
  40209=>"000111111",
  40210=>"111111111",
  40211=>"101101111",
  40212=>"011111111",
  40213=>"000111111",
  40214=>"011011001",
  40215=>"000000000",
  40216=>"000000001",
  40217=>"010000000",
  40218=>"001001111",
  40219=>"000111001",
  40220=>"000000100",
  40221=>"110111111",
  40222=>"000110000",
  40223=>"001111101",
  40224=>"011001001",
  40225=>"111001100",
  40226=>"111100000",
  40227=>"111111100",
  40228=>"000000110",
  40229=>"010111111",
  40230=>"001011111",
  40231=>"111100111",
  40232=>"000000000",
  40233=>"000111000",
  40234=>"000111111",
  40235=>"000000000",
  40236=>"000000000",
  40237=>"000000000",
  40238=>"111001111",
  40239=>"111111000",
  40240=>"001000000",
  40241=>"000000000",
  40242=>"000000000",
  40243=>"111111100",
  40244=>"110111100",
  40245=>"101101000",
  40246=>"000000000",
  40247=>"111101000",
  40248=>"111111000",
  40249=>"000000111",
  40250=>"000000001",
  40251=>"111111111",
  40252=>"111111011",
  40253=>"000011011",
  40254=>"000110111",
  40255=>"111111111",
  40256=>"011000000",
  40257=>"000000001",
  40258=>"000000000",
  40259=>"111111000",
  40260=>"101100111",
  40261=>"111010111",
  40262=>"111000000",
  40263=>"001011000",
  40264=>"101000000",
  40265=>"110001111",
  40266=>"110110111",
  40267=>"011000000",
  40268=>"001000000",
  40269=>"000111111",
  40270=>"000110111",
  40271=>"001001000",
  40272=>"011011001",
  40273=>"100010011",
  40274=>"111111111",
  40275=>"011000111",
  40276=>"111000111",
  40277=>"000011011",
  40278=>"111000000",
  40279=>"001001001",
  40280=>"100101111",
  40281=>"001001111",
  40282=>"111100000",
  40283=>"110000000",
  40284=>"000001111",
  40285=>"011000000",
  40286=>"000000001",
  40287=>"011111000",
  40288=>"111000000",
  40289=>"001101111",
  40290=>"000001000",
  40291=>"101101111",
  40292=>"011011000",
  40293=>"111100000",
  40294=>"111111000",
  40295=>"111111111",
  40296=>"110110110",
  40297=>"000010110",
  40298=>"011000000",
  40299=>"010000100",
  40300=>"001001001",
  40301=>"111011111",
  40302=>"111111100",
  40303=>"111111000",
  40304=>"000000000",
  40305=>"101000000",
  40306=>"000000000",
  40307=>"000000000",
  40308=>"111111000",
  40309=>"111111111",
  40310=>"111000000",
  40311=>"111110000",
  40312=>"111111001",
  40313=>"111111111",
  40314=>"000000000",
  40315=>"100111111",
  40316=>"101000000",
  40317=>"111111111",
  40318=>"111111000",
  40319=>"111000000",
  40320=>"011111111",
  40321=>"111111111",
  40322=>"000100000",
  40323=>"000001001",
  40324=>"111000000",
  40325=>"110100110",
  40326=>"000000111",
  40327=>"001111111",
  40328=>"111111101",
  40329=>"111011010",
  40330=>"000000111",
  40331=>"000101111",
  40332=>"000000111",
  40333=>"110110000",
  40334=>"111111111",
  40335=>"111111111",
  40336=>"111111111",
  40337=>"111000000",
  40338=>"111101111",
  40339=>"111111000",
  40340=>"000001101",
  40341=>"110110000",
  40342=>"110111110",
  40343=>"001000000",
  40344=>"100111111",
  40345=>"111111111",
  40346=>"000000000",
  40347=>"000101111",
  40348=>"000011011",
  40349=>"111101101",
  40350=>"001001000",
  40351=>"000111111",
  40352=>"000000001",
  40353=>"101100101",
  40354=>"100000000",
  40355=>"000000111",
  40356=>"110010000",
  40357=>"100101100",
  40358=>"001001000",
  40359=>"001000000",
  40360=>"000100000",
  40361=>"011000000",
  40362=>"111111111",
  40363=>"000000000",
  40364=>"000000000",
  40365=>"101111111",
  40366=>"110111111",
  40367=>"111111111",
  40368=>"111111001",
  40369=>"011100100",
  40370=>"100111111",
  40371=>"000000000",
  40372=>"001100111",
  40373=>"000000101",
  40374=>"111011001",
  40375=>"000100101",
  40376=>"000000111",
  40377=>"000000000",
  40378=>"111010110",
  40379=>"000000000",
  40380=>"001101111",
  40381=>"000010111",
  40382=>"001001001",
  40383=>"101111110",
  40384=>"001111111",
  40385=>"011001000",
  40386=>"111101101",
  40387=>"000111100",
  40388=>"111111111",
  40389=>"011011011",
  40390=>"001000000",
  40391=>"001001111",
  40392=>"000000000",
  40393=>"110000000",
  40394=>"111111011",
  40395=>"111001011",
  40396=>"001111000",
  40397=>"011000011",
  40398=>"111101110",
  40399=>"000000101",
  40400=>"110111111",
  40401=>"000011011",
  40402=>"000110110",
  40403=>"000000111",
  40404=>"000100000",
  40405=>"111111000",
  40406=>"000000011",
  40407=>"000110110",
  40408=>"000000110",
  40409=>"000000001",
  40410=>"101100111",
  40411=>"000000000",
  40412=>"000001000",
  40413=>"000000101",
  40414=>"000000101",
  40415=>"110110000",
  40416=>"000000111",
  40417=>"000000110",
  40418=>"000000001",
  40419=>"111101000",
  40420=>"000000101",
  40421=>"110110010",
  40422=>"101101001",
  40423=>"000000000",
  40424=>"001001001",
  40425=>"111000000",
  40426=>"000111111",
  40427=>"001000000",
  40428=>"111111111",
  40429=>"100000000",
  40430=>"000000000",
  40431=>"000000000",
  40432=>"000000000",
  40433=>"000111011",
  40434=>"111111111",
  40435=>"111111111",
  40436=>"111011000",
  40437=>"001000000",
  40438=>"111000000",
  40439=>"110000000",
  40440=>"001111101",
  40441=>"000110000",
  40442=>"001000000",
  40443=>"111000000",
  40444=>"100111111",
  40445=>"000110111",
  40446=>"001001000",
  40447=>"000000000",
  40448=>"000100000",
  40449=>"111111111",
  40450=>"111111111",
  40451=>"010000010",
  40452=>"001000100",
  40453=>"010010010",
  40454=>"111111110",
  40455=>"011001000",
  40456=>"010100111",
  40457=>"111111011",
  40458=>"001111111",
  40459=>"000110110",
  40460=>"000000000",
  40461=>"000101011",
  40462=>"110100000",
  40463=>"110110110",
  40464=>"001001000",
  40465=>"000000000",
  40466=>"111111100",
  40467=>"111100000",
  40468=>"110100111",
  40469=>"000000000",
  40470=>"000000010",
  40471=>"111111111",
  40472=>"000001000",
  40473=>"111111111",
  40474=>"000000000",
  40475=>"100100111",
  40476=>"001000001",
  40477=>"111111111",
  40478=>"100101000",
  40479=>"000000101",
  40480=>"000000000",
  40481=>"111111110",
  40482=>"100000000",
  40483=>"111101000",
  40484=>"000000100",
  40485=>"111110110",
  40486=>"111111111",
  40487=>"000011011",
  40488=>"000011001",
  40489=>"000000000",
  40490=>"111111111",
  40491=>"001101111",
  40492=>"011001111",
  40493=>"111111010",
  40494=>"111111000",
  40495=>"000000001",
  40496=>"111111111",
  40497=>"111111111",
  40498=>"001000100",
  40499=>"000111111",
  40500=>"100000000",
  40501=>"011011111",
  40502=>"000000000",
  40503=>"110110110",
  40504=>"000000000",
  40505=>"000000000",
  40506=>"000011011",
  40507=>"111111111",
  40508=>"111111111",
  40509=>"111111111",
  40510=>"111110110",
  40511=>"000000000",
  40512=>"000001000",
  40513=>"111111001",
  40514=>"000010110",
  40515=>"010000000",
  40516=>"100000100",
  40517=>"111011001",
  40518=>"111000000",
  40519=>"000000000",
  40520=>"011001000",
  40521=>"111111111",
  40522=>"000011111",
  40523=>"000000000",
  40524=>"000000000",
  40525=>"100000111",
  40526=>"111111111",
  40527=>"000000000",
  40528=>"000000000",
  40529=>"011111101",
  40530=>"010010000",
  40531=>"111111111",
  40532=>"100100100",
  40533=>"000000000",
  40534=>"001000000",
  40535=>"100111111",
  40536=>"000000000",
  40537=>"111111111",
  40538=>"111111010",
  40539=>"100110000",
  40540=>"111111111",
  40541=>"110110111",
  40542=>"000000000",
  40543=>"011011011",
  40544=>"111111111",
  40545=>"111111111",
  40546=>"111001111",
  40547=>"111011000",
  40548=>"111101000",
  40549=>"000111111",
  40550=>"111111000",
  40551=>"000100100",
  40552=>"101001001",
  40553=>"000000000",
  40554=>"000000000",
  40555=>"110110100",
  40556=>"111111111",
  40557=>"111111111",
  40558=>"101101000",
  40559=>"001000010",
  40560=>"110111111",
  40561=>"000010011",
  40562=>"111101001",
  40563=>"000000000",
  40564=>"101000100",
  40565=>"101000111",
  40566=>"111111010",
  40567=>"000111111",
  40568=>"110111111",
  40569=>"000000000",
  40570=>"111111111",
  40571=>"111111111",
  40572=>"000000000",
  40573=>"111111111",
  40574=>"101000000",
  40575=>"000000000",
  40576=>"001000000",
  40577=>"000101111",
  40578=>"000111111",
  40579=>"111111100",
  40580=>"111111111",
  40581=>"000000111",
  40582=>"111111111",
  40583=>"000000000",
  40584=>"110111111",
  40585=>"001011010",
  40586=>"000000000",
  40587=>"000000111",
  40588=>"000001000",
  40589=>"000000000",
  40590=>"111111011",
  40591=>"100110000",
  40592=>"000000000",
  40593=>"111111111",
  40594=>"000000111",
  40595=>"000000000",
  40596=>"111111111",
  40597=>"000000000",
  40598=>"000111111",
  40599=>"000000000",
  40600=>"000000000",
  40601=>"111111111",
  40602=>"000100000",
  40603=>"000000000",
  40604=>"000000001",
  40605=>"111101101",
  40606=>"100100001",
  40607=>"000000011",
  40608=>"010011000",
  40609=>"010001000",
  40610=>"000100100",
  40611=>"000000000",
  40612=>"111110000",
  40613=>"100111111",
  40614=>"000011011",
  40615=>"111111000",
  40616=>"000000000",
  40617=>"110111111",
  40618=>"000010110",
  40619=>"000000000",
  40620=>"000000000",
  40621=>"111111111",
  40622=>"101101111",
  40623=>"011001001",
  40624=>"000000000",
  40625=>"111110000",
  40626=>"011111011",
  40627=>"111111111",
  40628=>"111111111",
  40629=>"000001000",
  40630=>"111000111",
  40631=>"111111111",
  40632=>"000011111",
  40633=>"011000011",
  40634=>"110100100",
  40635=>"000010110",
  40636=>"000000001",
  40637=>"110110110",
  40638=>"111001011",
  40639=>"000010111",
  40640=>"011111111",
  40641=>"000000100",
  40642=>"011011011",
  40643=>"110111111",
  40644=>"111111111",
  40645=>"111111111",
  40646=>"111111111",
  40647=>"000000000",
  40648=>"111101000",
  40649=>"001000110",
  40650=>"000000000",
  40651=>"110000000",
  40652=>"001001001",
  40653=>"111111111",
  40654=>"010111111",
  40655=>"111100100",
  40656=>"111111111",
  40657=>"011111111",
  40658=>"111111110",
  40659=>"000101111",
  40660=>"110111111",
  40661=>"111111111",
  40662=>"000000000",
  40663=>"000000111",
  40664=>"111111111",
  40665=>"111111001",
  40666=>"011111111",
  40667=>"000000000",
  40668=>"000000001",
  40669=>"000000000",
  40670=>"000000000",
  40671=>"100100001",
  40672=>"010111011",
  40673=>"000000000",
  40674=>"111110010",
  40675=>"000000000",
  40676=>"000000000",
  40677=>"000000010",
  40678=>"111111111",
  40679=>"110111000",
  40680=>"011000000",
  40681=>"100000000",
  40682=>"111000000",
  40683=>"111111111",
  40684=>"111111000",
  40685=>"111111111",
  40686=>"100000001",
  40687=>"111111111",
  40688=>"100111101",
  40689=>"111110110",
  40690=>"000000000",
  40691=>"000000000",
  40692=>"000011001",
  40693=>"110110100",
  40694=>"001111111",
  40695=>"000000001",
  40696=>"000000000",
  40697=>"111111111",
  40698=>"110111111",
  40699=>"111111110",
  40700=>"100000000",
  40701=>"111111101",
  40702=>"110111111",
  40703=>"000000000",
  40704=>"000000000",
  40705=>"111111111",
  40706=>"000000000",
  40707=>"000000000",
  40708=>"000000000",
  40709=>"011000000",
  40710=>"000000111",
  40711=>"111011111",
  40712=>"000000000",
  40713=>"000000000",
  40714=>"010111010",
  40715=>"000000000",
  40716=>"001001001",
  40717=>"011011111",
  40718=>"111111000",
  40719=>"111111000",
  40720=>"000000101",
  40721=>"000000000",
  40722=>"111111111",
  40723=>"000000000",
  40724=>"001010111",
  40725=>"000110100",
  40726=>"000000000",
  40727=>"001111111",
  40728=>"111011101",
  40729=>"000000110",
  40730=>"100000000",
  40731=>"000010111",
  40732=>"000000000",
  40733=>"000000000",
  40734=>"011111111",
  40735=>"000000111",
  40736=>"000000000",
  40737=>"000010000",
  40738=>"000000011",
  40739=>"000011111",
  40740=>"110100110",
  40741=>"000000000",
  40742=>"000000000",
  40743=>"000000000",
  40744=>"111101100",
  40745=>"000000000",
  40746=>"000010000",
  40747=>"011011000",
  40748=>"111111111",
  40749=>"100000000",
  40750=>"111000010",
  40751=>"111111111",
  40752=>"000011010",
  40753=>"010000000",
  40754=>"000001000",
  40755=>"111111110",
  40756=>"000000011",
  40757=>"000000000",
  40758=>"000100100",
  40759=>"011111011",
  40760=>"000000000",
  40761=>"111111101",
  40762=>"000000100",
  40763=>"111110111",
  40764=>"110111010",
  40765=>"100000000",
  40766=>"001101100",
  40767=>"111111111",
  40768=>"000000000",
  40769=>"000111000",
  40770=>"110111110",
  40771=>"101101101",
  40772=>"000000000",
  40773=>"000000000",
  40774=>"111100000",
  40775=>"111111111",
  40776=>"000000000",
  40777=>"000000111",
  40778=>"010111111",
  40779=>"111111111",
  40780=>"110110110",
  40781=>"111111111",
  40782=>"000000000",
  40783=>"111111111",
  40784=>"011011010",
  40785=>"000111110",
  40786=>"010010111",
  40787=>"111111111",
  40788=>"111001001",
  40789=>"011010010",
  40790=>"110010011",
  40791=>"000000000",
  40792=>"000000000",
  40793=>"010111111",
  40794=>"111011011",
  40795=>"000011001",
  40796=>"111111111",
  40797=>"111110000",
  40798=>"111111111",
  40799=>"100100100",
  40800=>"010010111",
  40801=>"000010000",
  40802=>"111111000",
  40803=>"111110000",
  40804=>"111101011",
  40805=>"000000000",
  40806=>"000101111",
  40807=>"111100000",
  40808=>"111100000",
  40809=>"000000000",
  40810=>"011000000",
  40811=>"111111111",
  40812=>"000000000",
  40813=>"000000000",
  40814=>"000101111",
  40815=>"010111010",
  40816=>"111111111",
  40817=>"000111110",
  40818=>"110111111",
  40819=>"110111111",
  40820=>"010010110",
  40821=>"111101111",
  40822=>"000010011",
  40823=>"000011111",
  40824=>"111101111",
  40825=>"000010000",
  40826=>"100000000",
  40827=>"111111111",
  40828=>"111111111",
  40829=>"111111111",
  40830=>"000000000",
  40831=>"000000001",
  40832=>"000100101",
  40833=>"111111100",
  40834=>"110000111",
  40835=>"000000000",
  40836=>"111111111",
  40837=>"111000000",
  40838=>"111110101",
  40839=>"011111101",
  40840=>"111010000",
  40841=>"000000010",
  40842=>"000000000",
  40843=>"000000000",
  40844=>"111101111",
  40845=>"111111001",
  40846=>"101111111",
  40847=>"111111111",
  40848=>"000100100",
  40849=>"011011011",
  40850=>"010000000",
  40851=>"010010000",
  40852=>"100110011",
  40853=>"010110000",
  40854=>"111111111",
  40855=>"000000000",
  40856=>"011000100",
  40857=>"111101000",
  40858=>"000000000",
  40859=>"100001001",
  40860=>"000110000",
  40861=>"100000000",
  40862=>"000000000",
  40863=>"000000000",
  40864=>"100110110",
  40865=>"100000001",
  40866=>"000001001",
  40867=>"000000000",
  40868=>"000000111",
  40869=>"111111111",
  40870=>"011001011",
  40871=>"000000000",
  40872=>"111111011",
  40873=>"111111111",
  40874=>"000000000",
  40875=>"000000000",
  40876=>"111111100",
  40877=>"000110000",
  40878=>"000111101",
  40879=>"000010000",
  40880=>"000111111",
  40881=>"111111000",
  40882=>"000000000",
  40883=>"000000000",
  40884=>"000001001",
  40885=>"111111111",
  40886=>"000001011",
  40887=>"101000000",
  40888=>"111000000",
  40889=>"000011110",
  40890=>"100110111",
  40891=>"001001000",
  40892=>"001000000",
  40893=>"111111111",
  40894=>"000000001",
  40895=>"111000000",
  40896=>"000000000",
  40897=>"000000001",
  40898=>"111111111",
  40899=>"011011011",
  40900=>"111111101",
  40901=>"111111011",
  40902=>"000000000",
  40903=>"001001001",
  40904=>"000000000",
  40905=>"101111111",
  40906=>"000000000",
  40907=>"000000111",
  40908=>"111111010",
  40909=>"000111111",
  40910=>"000000100",
  40911=>"000000000",
  40912=>"011000000",
  40913=>"111111111",
  40914=>"001001000",
  40915=>"000000000",
  40916=>"111111111",
  40917=>"110110000",
  40918=>"101111111",
  40919=>"011000001",
  40920=>"111111111",
  40921=>"000000000",
  40922=>"001111100",
  40923=>"110111000",
  40924=>"111110110",
  40925=>"000000000",
  40926=>"011000100",
  40927=>"100100000",
  40928=>"000000000",
  40929=>"111001111",
  40930=>"111111111",
  40931=>"000111110",
  40932=>"010000111",
  40933=>"100110000",
  40934=>"000101101",
  40935=>"001000111",
  40936=>"000000110",
  40937=>"000000000",
  40938=>"111111110",
  40939=>"111100000",
  40940=>"000001001",
  40941=>"111111111",
  40942=>"001000000",
  40943=>"111110001",
  40944=>"111111110",
  40945=>"111111111",
  40946=>"111111111",
  40947=>"011000000",
  40948=>"000001000",
  40949=>"110000000",
  40950=>"111111111",
  40951=>"100100000",
  40952=>"011001001",
  40953=>"110111111",
  40954=>"111111101",
  40955=>"111111000",
  40956=>"111100000",
  40957=>"000000000",
  40958=>"000100000",
  40959=>"111111111",
  40960=>"111111011",
  40961=>"000000000",
  40962=>"000000000",
  40963=>"111110000",
  40964=>"000011000",
  40965=>"111101100",
  40966=>"000000000",
  40967=>"101000000",
  40968=>"011001001",
  40969=>"111111000",
  40970=>"000000000",
  40971=>"011011111",
  40972=>"001111111",
  40973=>"011000011",
  40974=>"111111011",
  40975=>"000110110",
  40976=>"000000101",
  40977=>"111011000",
  40978=>"111111111",
  40979=>"110111110",
  40980=>"111001000",
  40981=>"111000000",
  40982=>"100010000",
  40983=>"111111011",
  40984=>"110110110",
  40985=>"001001011",
  40986=>"111111111",
  40987=>"000110110",
  40988=>"100100000",
  40989=>"000101111",
  40990=>"000000111",
  40991=>"000100111",
  40992=>"111110110",
  40993=>"101000000",
  40994=>"000000010",
  40995=>"111111111",
  40996=>"111111111",
  40997=>"001000000",
  40998=>"101000000",
  40999=>"101011011",
  41000=>"000100111",
  41001=>"000010010",
  41002=>"000110111",
  41003=>"000000000",
  41004=>"111111111",
  41005=>"000000000",
  41006=>"111000000",
  41007=>"011000000",
  41008=>"000010111",
  41009=>"000000000",
  41010=>"000000011",
  41011=>"111011011",
  41012=>"111111111",
  41013=>"011111110",
  41014=>"100000000",
  41015=>"000000011",
  41016=>"000011111",
  41017=>"000100100",
  41018=>"111111111",
  41019=>"111111000",
  41020=>"000000000",
  41021=>"000000000",
  41022=>"111111111",
  41023=>"000000000",
  41024=>"000100111",
  41025=>"111101101",
  41026=>"111011001",
  41027=>"111011000",
  41028=>"011000000",
  41029=>"111111011",
  41030=>"111101101",
  41031=>"000000111",
  41032=>"000000110",
  41033=>"111101111",
  41034=>"111000000",
  41035=>"010010010",
  41036=>"010110000",
  41037=>"110110100",
  41038=>"111101000",
  41039=>"011111111",
  41040=>"000000000",
  41041=>"001001000",
  41042=>"000000000",
  41043=>"000000000",
  41044=>"100110111",
  41045=>"010011111",
  41046=>"000000111",
  41047=>"011010000",
  41048=>"000011111",
  41049=>"111000000",
  41050=>"000000000",
  41051=>"000000000",
  41052=>"000000000",
  41053=>"111111110",
  41054=>"000100000",
  41055=>"000000000",
  41056=>"000000000",
  41057=>"000111111",
  41058=>"111111111",
  41059=>"111111111",
  41060=>"000000000",
  41061=>"001100110",
  41062=>"110111111",
  41063=>"000000000",
  41064=>"000000000",
  41065=>"000000000",
  41066=>"111111111",
  41067=>"111111111",
  41068=>"001011111",
  41069=>"000001001",
  41070=>"000000010",
  41071=>"111111110",
  41072=>"000101001",
  41073=>"110111111",
  41074=>"111111111",
  41075=>"001000000",
  41076=>"000000010",
  41077=>"111111110",
  41078=>"000000000",
  41079=>"000000000",
  41080=>"100100111",
  41081=>"000100101",
  41082=>"101111111",
  41083=>"111111100",
  41084=>"001000000",
  41085=>"111110000",
  41086=>"101101111",
  41087=>"111011011",
  41088=>"000000000",
  41089=>"000111111",
  41090=>"111111111",
  41091=>"000011011",
  41092=>"001111111",
  41093=>"000011111",
  41094=>"111111111",
  41095=>"000000000",
  41096=>"111111111",
  41097=>"111001000",
  41098=>"111111111",
  41099=>"100000000",
  41100=>"011111111",
  41101=>"111111111",
  41102=>"000101001",
  41103=>"110111111",
  41104=>"111111111",
  41105=>"000000000",
  41106=>"010100100",
  41107=>"111011010",
  41108=>"110000000",
  41109=>"000000110",
  41110=>"111111111",
  41111=>"011011111",
  41112=>"000010010",
  41113=>"001000000",
  41114=>"101111110",
  41115=>"000000000",
  41116=>"000111111",
  41117=>"111111111",
  41118=>"000100000",
  41119=>"000000000",
  41120=>"111111111",
  41121=>"001101001",
  41122=>"111111111",
  41123=>"000000000",
  41124=>"001001111",
  41125=>"000111111",
  41126=>"000000000",
  41127=>"011111011",
  41128=>"011000000",
  41129=>"000000000",
  41130=>"000000000",
  41131=>"011011111",
  41132=>"000111010",
  41133=>"111111110",
  41134=>"111111111",
  41135=>"000000001",
  41136=>"000001111",
  41137=>"111011101",
  41138=>"111111011",
  41139=>"000000000",
  41140=>"010000000",
  41141=>"000000000",
  41142=>"001111001",
  41143=>"111111111",
  41144=>"000000010",
  41145=>"111111011",
  41146=>"100111011",
  41147=>"100100010",
  41148=>"111111111",
  41149=>"000000000",
  41150=>"111111110",
  41151=>"110100000",
  41152=>"111101000",
  41153=>"000111000",
  41154=>"000000000",
  41155=>"110110010",
  41156=>"111111111",
  41157=>"000011000",
  41158=>"000000000",
  41159=>"010010000",
  41160=>"000000000",
  41161=>"000001000",
  41162=>"000111111",
  41163=>"000000000",
  41164=>"000001001",
  41165=>"000011111",
  41166=>"000000000",
  41167=>"110110110",
  41168=>"011100110",
  41169=>"001000000",
  41170=>"111000000",
  41171=>"000000000",
  41172=>"111111011",
  41173=>"100110100",
  41174=>"011000000",
  41175=>"000001011",
  41176=>"111001011",
  41177=>"000011011",
  41178=>"111111111",
  41179=>"111111111",
  41180=>"001001111",
  41181=>"010010111",
  41182=>"111111111",
  41183=>"000100100",
  41184=>"000110111",
  41185=>"000001000",
  41186=>"000000000",
  41187=>"000000000",
  41188=>"000000100",
  41189=>"001001001",
  41190=>"011000000",
  41191=>"101001101",
  41192=>"111111111",
  41193=>"010000000",
  41194=>"000111111",
  41195=>"000001100",
  41196=>"001000111",
  41197=>"000000110",
  41198=>"000111111",
  41199=>"111000000",
  41200=>"000010011",
  41201=>"010000000",
  41202=>"011101111",
  41203=>"111111111",
  41204=>"111111011",
  41205=>"001000000",
  41206=>"111000000",
  41207=>"000000000",
  41208=>"000000000",
  41209=>"110110111",
  41210=>"000000111",
  41211=>"111111111",
  41212=>"010001111",
  41213=>"000000000",
  41214=>"000000000",
  41215=>"111111111",
  41216=>"000000000",
  41217=>"001100100",
  41218=>"111101001",
  41219=>"000000000",
  41220=>"111111100",
  41221=>"000000000",
  41222=>"111111110",
  41223=>"011111111",
  41224=>"000000111",
  41225=>"111101111",
  41226=>"000000001",
  41227=>"000000001",
  41228=>"111111111",
  41229=>"011101001",
  41230=>"000000011",
  41231=>"001001000",
  41232=>"000100100",
  41233=>"111111000",
  41234=>"111111111",
  41235=>"000111000",
  41236=>"111000000",
  41237=>"111111111",
  41238=>"011111110",
  41239=>"110000010",
  41240=>"000000110",
  41241=>"000000100",
  41242=>"000000111",
  41243=>"000111111",
  41244=>"000000000",
  41245=>"110010111",
  41246=>"000000000",
  41247=>"111000111",
  41248=>"011111111",
  41249=>"011111000",
  41250=>"000000000",
  41251=>"000111111",
  41252=>"101000000",
  41253=>"111011011",
  41254=>"111111111",
  41255=>"000100000",
  41256=>"000000000",
  41257=>"111110000",
  41258=>"100100111",
  41259=>"000110111",
  41260=>"000000000",
  41261=>"010011111",
  41262=>"111100000",
  41263=>"000000000",
  41264=>"100110111",
  41265=>"000110110",
  41266=>"000000000",
  41267=>"001111010",
  41268=>"000000000",
  41269=>"111111111",
  41270=>"110000110",
  41271=>"000000000",
  41272=>"100000000",
  41273=>"011111111",
  41274=>"010010000",
  41275=>"001000000",
  41276=>"000000110",
  41277=>"100110111",
  41278=>"000000000",
  41279=>"000100010",
  41280=>"000000000",
  41281=>"100101111",
  41282=>"000000110",
  41283=>"000000110",
  41284=>"111111111",
  41285=>"010111111",
  41286=>"000000001",
  41287=>"111110110",
  41288=>"000000000",
  41289=>"111001000",
  41290=>"000100110",
  41291=>"110110010",
  41292=>"001010111",
  41293=>"011000000",
  41294=>"000100110",
  41295=>"110111111",
  41296=>"000110110",
  41297=>"100110100",
  41298=>"000111111",
  41299=>"111000100",
  41300=>"000000000",
  41301=>"111111011",
  41302=>"000000000",
  41303=>"100100111",
  41304=>"000011001",
  41305=>"000000110",
  41306=>"110011001",
  41307=>"111111111",
  41308=>"010000000",
  41309=>"111111000",
  41310=>"010110110",
  41311=>"111111111",
  41312=>"011110011",
  41313=>"111111011",
  41314=>"110110111",
  41315=>"001000110",
  41316=>"000000000",
  41317=>"000000000",
  41318=>"000110111",
  41319=>"000000000",
  41320=>"001001000",
  41321=>"001000000",
  41322=>"100100000",
  41323=>"001111111",
  41324=>"010011110",
  41325=>"000000000",
  41326=>"000000000",
  41327=>"000000100",
  41328=>"000000000",
  41329=>"000101000",
  41330=>"111111011",
  41331=>"100000000",
  41332=>"000001111",
  41333=>"000000000",
  41334=>"100100100",
  41335=>"100000110",
  41336=>"000010111",
  41337=>"001011011",
  41338=>"110000110",
  41339=>"100110110",
  41340=>"100100100",
  41341=>"000100111",
  41342=>"000000011",
  41343=>"111111111",
  41344=>"001000000",
  41345=>"011111011",
  41346=>"100110110",
  41347=>"110000000",
  41348=>"000111111",
  41349=>"101101111",
  41350=>"100111111",
  41351=>"000101000",
  41352=>"010000110",
  41353=>"000010000",
  41354=>"011111111",
  41355=>"000000000",
  41356=>"110111111",
  41357=>"111110110",
  41358=>"111111111",
  41359=>"011111011",
  41360=>"000000000",
  41361=>"110110000",
  41362=>"000000000",
  41363=>"000010010",
  41364=>"000000001",
  41365=>"011011000",
  41366=>"001001000",
  41367=>"100100100",
  41368=>"000000000",
  41369=>"000000000",
  41370=>"000000000",
  41371=>"000010110",
  41372=>"000000010",
  41373=>"000000000",
  41374=>"111111111",
  41375=>"000000000",
  41376=>"001100111",
  41377=>"100100111",
  41378=>"111010000",
  41379=>"110011000",
  41380=>"000001111",
  41381=>"000110000",
  41382=>"000000011",
  41383=>"001000000",
  41384=>"000000000",
  41385=>"000000000",
  41386=>"110111100",
  41387=>"111111111",
  41388=>"111111111",
  41389=>"010111111",
  41390=>"000100000",
  41391=>"000110111",
  41392=>"001001001",
  41393=>"011111111",
  41394=>"000000000",
  41395=>"000000000",
  41396=>"000100101",
  41397=>"000000000",
  41398=>"000000000",
  41399=>"000000010",
  41400=>"110010110",
  41401=>"111111110",
  41402=>"100100110",
  41403=>"000000000",
  41404=>"000000110",
  41405=>"111111111",
  41406=>"111000000",
  41407=>"001111100",
  41408=>"000000000",
  41409=>"000001011",
  41410=>"000000110",
  41411=>"000110000",
  41412=>"000000011",
  41413=>"000100111",
  41414=>"010011000",
  41415=>"000000000",
  41416=>"000000111",
  41417=>"000001000",
  41418=>"000011011",
  41419=>"011011011",
  41420=>"011010000",
  41421=>"000000000",
  41422=>"111101001",
  41423=>"110111100",
  41424=>"111000100",
  41425=>"000001111",
  41426=>"000000101",
  41427=>"011111101",
  41428=>"100100111",
  41429=>"111111110",
  41430=>"000011011",
  41431=>"101101000",
  41432=>"111111111",
  41433=>"111111110",
  41434=>"001000000",
  41435=>"000000000",
  41436=>"000001000",
  41437=>"111111011",
  41438=>"110111001",
  41439=>"000110100",
  41440=>"000000000",
  41441=>"111010000",
  41442=>"111111100",
  41443=>"100111011",
  41444=>"001000111",
  41445=>"111111111",
  41446=>"001001001",
  41447=>"000000111",
  41448=>"111111100",
  41449=>"001000000",
  41450=>"010111111",
  41451=>"111111111",
  41452=>"101111111",
  41453=>"100111011",
  41454=>"111111101",
  41455=>"111001000",
  41456=>"100000100",
  41457=>"011111111",
  41458=>"000000000",
  41459=>"100000000",
  41460=>"000111111",
  41461=>"000000000",
  41462=>"000000110",
  41463=>"001111111",
  41464=>"011001001",
  41465=>"110010011",
  41466=>"011011001",
  41467=>"000000000",
  41468=>"111111111",
  41469=>"000000100",
  41470=>"100000000",
  41471=>"000000000",
  41472=>"001111011",
  41473=>"111111010",
  41474=>"000000000",
  41475=>"110100000",
  41476=>"010000100",
  41477=>"000000000",
  41478=>"000000100",
  41479=>"000000000",
  41480=>"111100000",
  41481=>"001001001",
  41482=>"111011011",
  41483=>"111000011",
  41484=>"000000000",
  41485=>"000111110",
  41486=>"010111111",
  41487=>"000100100",
  41488=>"001001000",
  41489=>"111111101",
  41490=>"111001000",
  41491=>"100111111",
  41492=>"001000000",
  41493=>"100100000",
  41494=>"000000000",
  41495=>"111111001",
  41496=>"111111110",
  41497=>"110110110",
  41498=>"000000000",
  41499=>"000010000",
  41500=>"000000000",
  41501=>"000000111",
  41502=>"110110000",
  41503=>"001000111",
  41504=>"000011010",
  41505=>"111111110",
  41506=>"100110110",
  41507=>"010111000",
  41508=>"111001111",
  41509=>"111111111",
  41510=>"111111111",
  41511=>"000111100",
  41512=>"110110000",
  41513=>"000000000",
  41514=>"011000000",
  41515=>"000010010",
  41516=>"011111111",
  41517=>"011011011",
  41518=>"111111110",
  41519=>"000111111",
  41520=>"110111111",
  41521=>"000000100",
  41522=>"111110000",
  41523=>"111111111",
  41524=>"111111011",
  41525=>"101101001",
  41526=>"010111000",
  41527=>"000011000",
  41528=>"011111011",
  41529=>"000000000",
  41530=>"000000000",
  41531=>"000000000",
  41532=>"000000000",
  41533=>"000011011",
  41534=>"000011011",
  41535=>"100111000",
  41536=>"010000000",
  41537=>"001111110",
  41538=>"000010010",
  41539=>"010010010",
  41540=>"100101110",
  41541=>"001100111",
  41542=>"010010010",
  41543=>"000000000",
  41544=>"011111011",
  41545=>"101100101",
  41546=>"010111111",
  41547=>"110110110",
  41548=>"100100110",
  41549=>"100000101",
  41550=>"111111000",
  41551=>"000000100",
  41552=>"000000000",
  41553=>"000111111",
  41554=>"000110011",
  41555=>"111111111",
  41556=>"000000000",
  41557=>"011111111",
  41558=>"101011111",
  41559=>"111111010",
  41560=>"001011111",
  41561=>"000000000",
  41562=>"000000000",
  41563=>"111100000",
  41564=>"011111111",
  41565=>"000000000",
  41566=>"010111110",
  41567=>"110110010",
  41568=>"000000100",
  41569=>"101111000",
  41570=>"111110111",
  41571=>"111111100",
  41572=>"110111011",
  41573=>"000000000",
  41574=>"010011111",
  41575=>"110111111",
  41576=>"000001111",
  41577=>"000000000",
  41578=>"111100111",
  41579=>"111111111",
  41580=>"000000010",
  41581=>"000000000",
  41582=>"000000000",
  41583=>"111111111",
  41584=>"000000000",
  41585=>"000000111",
  41586=>"011011011",
  41587=>"100111111",
  41588=>"000110111",
  41589=>"111111011",
  41590=>"001111111",
  41591=>"011011011",
  41592=>"000111110",
  41593=>"000000000",
  41594=>"000001000",
  41595=>"000000000",
  41596=>"101000000",
  41597=>"000110110",
  41598=>"000011001",
  41599=>"000000000",
  41600=>"000100100",
  41601=>"000010111",
  41602=>"000100111",
  41603=>"000000101",
  41604=>"111101100",
  41605=>"000000000",
  41606=>"110011011",
  41607=>"000011111",
  41608=>"101001000",
  41609=>"000000000",
  41610=>"111101100",
  41611=>"000000000",
  41612=>"100111001",
  41613=>"111010010",
  41614=>"000011010",
  41615=>"011111111",
  41616=>"000000001",
  41617=>"011111001",
  41618=>"100000001",
  41619=>"111111111",
  41620=>"000001000",
  41621=>"111111111",
  41622=>"001001011",
  41623=>"000000000",
  41624=>"000001100",
  41625=>"111111111",
  41626=>"000010111",
  41627=>"010000000",
  41628=>"000010000",
  41629=>"111111111",
  41630=>"111011111",
  41631=>"000000000",
  41632=>"000000010",
  41633=>"000110010",
  41634=>"100110111",
  41635=>"111000000",
  41636=>"010110011",
  41637=>"110110111",
  41638=>"000000000",
  41639=>"110010111",
  41640=>"111111011",
  41641=>"111111111",
  41642=>"111101111",
  41643=>"001000001",
  41644=>"000000010",
  41645=>"001011001",
  41646=>"000111111",
  41647=>"000100000",
  41648=>"000000000",
  41649=>"000101101",
  41650=>"000000000",
  41651=>"000000000",
  41652=>"111111110",
  41653=>"000011111",
  41654=>"111111111",
  41655=>"111111111",
  41656=>"000110010",
  41657=>"000000000",
  41658=>"011000000",
  41659=>"000110010",
  41660=>"001001101",
  41661=>"011111111",
  41662=>"000000000",
  41663=>"111100000",
  41664=>"000000111",
  41665=>"000000000",
  41666=>"111000000",
  41667=>"000010010",
  41668=>"101101111",
  41669=>"000011001",
  41670=>"000010111",
  41671=>"000000010",
  41672=>"010010010",
  41673=>"011011010",
  41674=>"010000111",
  41675=>"001111111",
  41676=>"000000000",
  41677=>"000001111",
  41678=>"000111000",
  41679=>"111110110",
  41680=>"000000000",
  41681=>"011011000",
  41682=>"111111000",
  41683=>"111001111",
  41684=>"101101111",
  41685=>"100010000",
  41686=>"000000000",
  41687=>"111111111",
  41688=>"111111111",
  41689=>"111011000",
  41690=>"111111111",
  41691=>"111010010",
  41692=>"000001000",
  41693=>"000010010",
  41694=>"000000000",
  41695=>"000001001",
  41696=>"101000000",
  41697=>"011011111",
  41698=>"101001111",
  41699=>"110111011",
  41700=>"111100100",
  41701=>"010011010",
  41702=>"111011111",
  41703=>"110010000",
  41704=>"000111111",
  41705=>"101110011",
  41706=>"111111000",
  41707=>"011111000",
  41708=>"100000000",
  41709=>"101000111",
  41710=>"111101101",
  41711=>"000011010",
  41712=>"000001000",
  41713=>"011111100",
  41714=>"000000000",
  41715=>"010011000",
  41716=>"011110100",
  41717=>"000011011",
  41718=>"110000000",
  41719=>"111000000",
  41720=>"000000000",
  41721=>"110000000",
  41722=>"000000000",
  41723=>"010111101",
  41724=>"111001110",
  41725=>"110000011",
  41726=>"111000100",
  41727=>"111011000",
  41728=>"000000000",
  41729=>"011011000",
  41730=>"000000000",
  41731=>"000011110",
  41732=>"011010000",
  41733=>"101111111",
  41734=>"000000000",
  41735=>"000000001",
  41736=>"111011111",
  41737=>"000110110",
  41738=>"110110110",
  41739=>"000000000",
  41740=>"000000000",
  41741=>"000001111",
  41742=>"010011110",
  41743=>"000000000",
  41744=>"000000100",
  41745=>"000011001",
  41746=>"000000000",
  41747=>"010010111",
  41748=>"011111000",
  41749=>"100100001",
  41750=>"001001001",
  41751=>"010010000",
  41752=>"111111111",
  41753=>"111000111",
  41754=>"000000000",
  41755=>"100000000",
  41756=>"110000000",
  41757=>"001001111",
  41758=>"111111111",
  41759=>"111111111",
  41760=>"010111001",
  41761=>"010110111",
  41762=>"111111011",
  41763=>"100100000",
  41764=>"000000000",
  41765=>"111111111",
  41766=>"101111111",
  41767=>"111000101",
  41768=>"000110100",
  41769=>"000000000",
  41770=>"010010011",
  41771=>"000000011",
  41772=>"011111111",
  41773=>"110010111",
  41774=>"000000000",
  41775=>"011011011",
  41776=>"111111111",
  41777=>"000000110",
  41778=>"001000000",
  41779=>"001101111",
  41780=>"000000000",
  41781=>"111111011",
  41782=>"100000000",
  41783=>"100111001",
  41784=>"000000000",
  41785=>"011011000",
  41786=>"001011111",
  41787=>"111111111",
  41788=>"111011000",
  41789=>"000000000",
  41790=>"101100000",
  41791=>"000000010",
  41792=>"000000000",
  41793=>"000010000",
  41794=>"000100111",
  41795=>"000000000",
  41796=>"001010000",
  41797=>"000001011",
  41798=>"011011000",
  41799=>"000001011",
  41800=>"101111111",
  41801=>"001011000",
  41802=>"011011111",
  41803=>"000010000",
  41804=>"011011111",
  41805=>"010111111",
  41806=>"011000000",
  41807=>"110111111",
  41808=>"010000000",
  41809=>"000100000",
  41810=>"111100000",
  41811=>"111111111",
  41812=>"111111111",
  41813=>"111111111",
  41814=>"101011111",
  41815=>"001011111",
  41816=>"000000000",
  41817=>"000000000",
  41818=>"110111100",
  41819=>"010010011",
  41820=>"000000000",
  41821=>"001111111",
  41822=>"111111001",
  41823=>"001011001",
  41824=>"111111111",
  41825=>"111111111",
  41826=>"011010010",
  41827=>"100001011",
  41828=>"111111001",
  41829=>"111111111",
  41830=>"111011011",
  41831=>"000010000",
  41832=>"011011001",
  41833=>"000000000",
  41834=>"000110011",
  41835=>"000111101",
  41836=>"111111001",
  41837=>"010010111",
  41838=>"011111111",
  41839=>"000000000",
  41840=>"001001001",
  41841=>"001011111",
  41842=>"000001111",
  41843=>"111111101",
  41844=>"100000100",
  41845=>"011011011",
  41846=>"111000000",
  41847=>"111111111",
  41848=>"111111111",
  41849=>"111111111",
  41850=>"111111111",
  41851=>"000000000",
  41852=>"000000000",
  41853=>"000110110",
  41854=>"101100100",
  41855=>"100110110",
  41856=>"111001001",
  41857=>"011111010",
  41858=>"100101101",
  41859=>"001111111",
  41860=>"111111111",
  41861=>"000000000",
  41862=>"111011001",
  41863=>"000011111",
  41864=>"000000000",
  41865=>"000000000",
  41866=>"111111011",
  41867=>"000000100",
  41868=>"001000111",
  41869=>"100000110",
  41870=>"000000000",
  41871=>"111111111",
  41872=>"111111111",
  41873=>"111111111",
  41874=>"111101100",
  41875=>"111011001",
  41876=>"000000000",
  41877=>"111101111",
  41878=>"100100110",
  41879=>"110000000",
  41880=>"000011111",
  41881=>"111111011",
  41882=>"000000000",
  41883=>"000111000",
  41884=>"111011111",
  41885=>"000000000",
  41886=>"111111111",
  41887=>"000000010",
  41888=>"111111111",
  41889=>"111000001",
  41890=>"010110010",
  41891=>"000000011",
  41892=>"010110010",
  41893=>"001111111",
  41894=>"000000000",
  41895=>"111000000",
  41896=>"000000000",
  41897=>"000100101",
  41898=>"111101111",
  41899=>"100111110",
  41900=>"101000000",
  41901=>"000111011",
  41902=>"000000111",
  41903=>"000010000",
  41904=>"000010010",
  41905=>"101101011",
  41906=>"001111110",
  41907=>"001000001",
  41908=>"010000000",
  41909=>"000110110",
  41910=>"010010000",
  41911=>"111111100",
  41912=>"000000000",
  41913=>"000000000",
  41914=>"100100111",
  41915=>"000010000",
  41916=>"101001000",
  41917=>"110111111",
  41918=>"001001000",
  41919=>"011011001",
  41920=>"000000000",
  41921=>"000000010",
  41922=>"000000000",
  41923=>"000000000",
  41924=>"010011010",
  41925=>"000110010",
  41926=>"010111111",
  41927=>"011000110",
  41928=>"000000000",
  41929=>"111111111",
  41930=>"111111111",
  41931=>"000000111",
  41932=>"100111011",
  41933=>"000010000",
  41934=>"000010000",
  41935=>"001000100",
  41936=>"100101101",
  41937=>"010111000",
  41938=>"111111011",
  41939=>"111111111",
  41940=>"011011111",
  41941=>"111110110",
  41942=>"000110101",
  41943=>"000000000",
  41944=>"000010010",
  41945=>"000110110",
  41946=>"111111000",
  41947=>"000000111",
  41948=>"100101101",
  41949=>"111111000",
  41950=>"111111010",
  41951=>"111001001",
  41952=>"000110000",
  41953=>"111111011",
  41954=>"000000010",
  41955=>"111000000",
  41956=>"111111111",
  41957=>"111111101",
  41958=>"000110110",
  41959=>"111111111",
  41960=>"010111110",
  41961=>"111111111",
  41962=>"000000000",
  41963=>"111001000",
  41964=>"011011000",
  41965=>"000010010",
  41966=>"000000000",
  41967=>"110111010",
  41968=>"000000000",
  41969=>"111111000",
  41970=>"010111111",
  41971=>"011011010",
  41972=>"000000000",
  41973=>"111111111",
  41974=>"111010000",
  41975=>"000000000",
  41976=>"011010010",
  41977=>"000110100",
  41978=>"011011011",
  41979=>"001000000",
  41980=>"000000000",
  41981=>"111111111",
  41982=>"011011011",
  41983=>"111001111",
  41984=>"001001001",
  41985=>"010000100",
  41986=>"100000001",
  41987=>"111111011",
  41988=>"000001011",
  41989=>"011000100",
  41990=>"000000110",
  41991=>"101000111",
  41992=>"011111110",
  41993=>"000100000",
  41994=>"111011001",
  41995=>"111000000",
  41996=>"000100000",
  41997=>"111110110",
  41998=>"001000000",
  41999=>"100100000",
  42000=>"000000000",
  42001=>"000000000",
  42002=>"111111001",
  42003=>"111111111",
  42004=>"111011001",
  42005=>"111111111",
  42006=>"111011111",
  42007=>"100110110",
  42008=>"100001000",
  42009=>"000110111",
  42010=>"111111110",
  42011=>"110110111",
  42012=>"000000000",
  42013=>"000000111",
  42014=>"011011011",
  42015=>"000000111",
  42016=>"000000001",
  42017=>"001000111",
  42018=>"111000000",
  42019=>"000000000",
  42020=>"111000100",
  42021=>"000000100",
  42022=>"111001000",
  42023=>"011000111",
  42024=>"111111111",
  42025=>"001011111",
  42026=>"111111111",
  42027=>"111111111",
  42028=>"110111111",
  42029=>"000001001",
  42030=>"011011011",
  42031=>"111000000",
  42032=>"000000111",
  42033=>"000000000",
  42034=>"000010000",
  42035=>"000000100",
  42036=>"000011011",
  42037=>"100100100",
  42038=>"011111111",
  42039=>"100100000",
  42040=>"011001001",
  42041=>"110110111",
  42042=>"111111111",
  42043=>"111001000",
  42044=>"111111111",
  42045=>"000111111",
  42046=>"000000000",
  42047=>"101001000",
  42048=>"100111111",
  42049=>"010011011",
  42050=>"000011011",
  42051=>"000000111",
  42052=>"111001111",
  42053=>"000100110",
  42054=>"011000000",
  42055=>"111111111",
  42056=>"011011011",
  42057=>"000010111",
  42058=>"111111011",
  42059=>"010010000",
  42060=>"111111111",
  42061=>"110010111",
  42062=>"110000100",
  42063=>"001101111",
  42064=>"111100111",
  42065=>"000000111",
  42066=>"111110100",
  42067=>"100110000",
  42068=>"000000101",
  42069=>"000010111",
  42070=>"111111000",
  42071=>"000000000",
  42072=>"111111111",
  42073=>"000000100",
  42074=>"111011011",
  42075=>"111100001",
  42076=>"000000000",
  42077=>"111100100",
  42078=>"100111111",
  42079=>"000010011",
  42080=>"111111111",
  42081=>"000000000",
  42082=>"111111111",
  42083=>"000000000",
  42084=>"111111111",
  42085=>"000000001",
  42086=>"111011111",
  42087=>"011000000",
  42088=>"111000000",
  42089=>"011000000",
  42090=>"000000000",
  42091=>"110110100",
  42092=>"000001111",
  42093=>"111111111",
  42094=>"000000000",
  42095=>"111001000",
  42096=>"000000011",
  42097=>"111111111",
  42098=>"111111000",
  42099=>"111111111",
  42100=>"111111111",
  42101=>"000000100",
  42102=>"111111111",
  42103=>"000000011",
  42104=>"000000111",
  42105=>"111100000",
  42106=>"001000000",
  42107=>"000000100",
  42108=>"111111111",
  42109=>"000000001",
  42110=>"111001001",
  42111=>"000000000",
  42112=>"001000000",
  42113=>"000000000",
  42114=>"000000001",
  42115=>"011111000",
  42116=>"110000000",
  42117=>"111001011",
  42118=>"000010000",
  42119=>"000000000",
  42120=>"111110010",
  42121=>"001000111",
  42122=>"000000000",
  42123=>"000000000",
  42124=>"000000011",
  42125=>"111111000",
  42126=>"000000000",
  42127=>"001111111",
  42128=>"000011001",
  42129=>"000011111",
  42130=>"100000000",
  42131=>"001111111",
  42132=>"100000000",
  42133=>"000100000",
  42134=>"011001111",
  42135=>"000001001",
  42136=>"111011111",
  42137=>"000100110",
  42138=>"000000000",
  42139=>"000000000",
  42140=>"111011000",
  42141=>"011011000",
  42142=>"000110110",
  42143=>"000000000",
  42144=>"100000000",
  42145=>"111000000",
  42146=>"011011111",
  42147=>"000000111",
  42148=>"000011000",
  42149=>"111011111",
  42150=>"111001001",
  42151=>"110000000",
  42152=>"111111100",
  42153=>"000000000",
  42154=>"000000000",
  42155=>"100111111",
  42156=>"010000000",
  42157=>"100001011",
  42158=>"111111000",
  42159=>"011011011",
  42160=>"000111011",
  42161=>"100100100",
  42162=>"001101000",
  42163=>"011000111",
  42164=>"110100100",
  42165=>"011110110",
  42166=>"000001001",
  42167=>"111011111",
  42168=>"111111111",
  42169=>"100000001",
  42170=>"001011111",
  42171=>"000011101",
  42172=>"111100100",
  42173=>"000011000",
  42174=>"000000000",
  42175=>"111111001",
  42176=>"111100100",
  42177=>"000000000",
  42178=>"111011010",
  42179=>"011111111",
  42180=>"000000000",
  42181=>"000010011",
  42182=>"011011000",
  42183=>"111111111",
  42184=>"111011011",
  42185=>"111111110",
  42186=>"111110110",
  42187=>"001000000",
  42188=>"111111111",
  42189=>"111111100",
  42190=>"000000011",
  42191=>"000000011",
  42192=>"101001000",
  42193=>"111011000",
  42194=>"000100100",
  42195=>"000000000",
  42196=>"000001111",
  42197=>"000000111",
  42198=>"011111111",
  42199=>"001000000",
  42200=>"000101000",
  42201=>"001011011",
  42202=>"111101100",
  42203=>"000000011",
  42204=>"000000011",
  42205=>"110110000",
  42206=>"100101101",
  42207=>"000000001",
  42208=>"000000000",
  42209=>"111111000",
  42210=>"000000000",
  42211=>"011000000",
  42212=>"111000100",
  42213=>"110111111",
  42214=>"000000000",
  42215=>"001000000",
  42216=>"000000000",
  42217=>"111111111",
  42218=>"011001111",
  42219=>"000000000",
  42220=>"000000000",
  42221=>"001001111",
  42222=>"110000100",
  42223=>"000001100",
  42224=>"111011011",
  42225=>"000000100",
  42226=>"001000110",
  42227=>"010110110",
  42228=>"000000000",
  42229=>"000000110",
  42230=>"111111110",
  42231=>"000000000",
  42232=>"101001000",
  42233=>"101100111",
  42234=>"111111111",
  42235=>"111111111",
  42236=>"111101101",
  42237=>"111111111",
  42238=>"111111110",
  42239=>"000111110",
  42240=>"000001001",
  42241=>"011011011",
  42242=>"000000000",
  42243=>"111111111",
  42244=>"000000000",
  42245=>"110011011",
  42246=>"000000000",
  42247=>"000000000",
  42248=>"100000000",
  42249=>"000001000",
  42250=>"111110100",
  42251=>"111111111",
  42252=>"100100111",
  42253=>"110000110",
  42254=>"000001111",
  42255=>"101101110",
  42256=>"101101111",
  42257=>"111100000",
  42258=>"100100111",
  42259=>"011011001",
  42260=>"000000000",
  42261=>"110111111",
  42262=>"111011011",
  42263=>"111111001",
  42264=>"111011011",
  42265=>"000100111",
  42266=>"000000000",
  42267=>"000000100",
  42268=>"000000000",
  42269=>"011000110",
  42270=>"111111111",
  42271=>"000000101",
  42272=>"111111111",
  42273=>"001000001",
  42274=>"111100100",
  42275=>"000100111",
  42276=>"011111110",
  42277=>"100000000",
  42278=>"000011011",
  42279=>"111111111",
  42280=>"011111100",
  42281=>"000000001",
  42282=>"111111100",
  42283=>"000001001",
  42284=>"001001111",
  42285=>"001011111",
  42286=>"000111111",
  42287=>"110111110",
  42288=>"011001001",
  42289=>"000000000",
  42290=>"001000000",
  42291=>"001001001",
  42292=>"111111111",
  42293=>"000000111",
  42294=>"000100000",
  42295=>"000000000",
  42296=>"000000000",
  42297=>"000111111",
  42298=>"011111110",
  42299=>"111000000",
  42300=>"100100100",
  42301=>"101011111",
  42302=>"000000000",
  42303=>"000000000",
  42304=>"000000001",
  42305=>"100110000",
  42306=>"000011100",
  42307=>"011111111",
  42308=>"000000000",
  42309=>"000000000",
  42310=>"000000000",
  42311=>"000000100",
  42312=>"111111111",
  42313=>"110001011",
  42314=>"000010010",
  42315=>"011111100",
  42316=>"111100100",
  42317=>"000001011",
  42318=>"111111111",
  42319=>"111111111",
  42320=>"001001000",
  42321=>"110111111",
  42322=>"111110010",
  42323=>"111111000",
  42324=>"001000000",
  42325=>"110100011",
  42326=>"100000111",
  42327=>"111111101",
  42328=>"111111010",
  42329=>"001000000",
  42330=>"000001011",
  42331=>"000000000",
  42332=>"111101000",
  42333=>"111111111",
  42334=>"111111111",
  42335=>"111111011",
  42336=>"111111011",
  42337=>"111000100",
  42338=>"110110000",
  42339=>"000000000",
  42340=>"111110110",
  42341=>"000110111",
  42342=>"111100000",
  42343=>"111111111",
  42344=>"011111110",
  42345=>"000000000",
  42346=>"111111011",
  42347=>"110010010",
  42348=>"111111011",
  42349=>"010000000",
  42350=>"111111111",
  42351=>"111111000",
  42352=>"000000000",
  42353=>"001001101",
  42354=>"000000100",
  42355=>"000000000",
  42356=>"100000000",
  42357=>"000010010",
  42358=>"000000000",
  42359=>"000110100",
  42360=>"111000010",
  42361=>"100000000",
  42362=>"000000100",
  42363=>"111111111",
  42364=>"111101000",
  42365=>"111000100",
  42366=>"100100000",
  42367=>"000000000",
  42368=>"110110110",
  42369=>"000000110",
  42370=>"101011011",
  42371=>"111111111",
  42372=>"000000101",
  42373=>"000000000",
  42374=>"110110001",
  42375=>"010110010",
  42376=>"111101111",
  42377=>"000110111",
  42378=>"110000111",
  42379=>"111001101",
  42380=>"100100100",
  42381=>"001001100",
  42382=>"000011111",
  42383=>"000000000",
  42384=>"111101111",
  42385=>"111111111",
  42386=>"111111111",
  42387=>"000000000",
  42388=>"011111111",
  42389=>"110110100",
  42390=>"011000011",
  42391=>"011011111",
  42392=>"100001111",
  42393=>"000110110",
  42394=>"100100111",
  42395=>"000000001",
  42396=>"000000000",
  42397=>"111111111",
  42398=>"000011011",
  42399=>"100100111",
  42400=>"000111111",
  42401=>"110010101",
  42402=>"010010110",
  42403=>"100100111",
  42404=>"000100100",
  42405=>"001111111",
  42406=>"001000111",
  42407=>"000000000",
  42408=>"000000000",
  42409=>"010111100",
  42410=>"111111111",
  42411=>"000011110",
  42412=>"111111000",
  42413=>"111000111",
  42414=>"000000000",
  42415=>"101111111",
  42416=>"000110001",
  42417=>"111111110",
  42418=>"011010000",
  42419=>"111111111",
  42420=>"001011011",
  42421=>"011110111",
  42422=>"111011001",
  42423=>"000000000",
  42424=>"110000001",
  42425=>"000000000",
  42426=>"000000000",
  42427=>"111111101",
  42428=>"000000000",
  42429=>"000000000",
  42430=>"101001001",
  42431=>"111011011",
  42432=>"111111111",
  42433=>"000001001",
  42434=>"000001001",
  42435=>"000000000",
  42436=>"110110110",
  42437=>"001011111",
  42438=>"000000000",
  42439=>"000000000",
  42440=>"000000100",
  42441=>"100000000",
  42442=>"000000000",
  42443=>"111110000",
  42444=>"001000111",
  42445=>"000001111",
  42446=>"001111101",
  42447=>"111111111",
  42448=>"100111111",
  42449=>"000000000",
  42450=>"011011000",
  42451=>"101001000",
  42452=>"001000000",
  42453=>"011111111",
  42454=>"110101111",
  42455=>"001101101",
  42456=>"000000000",
  42457=>"111110110",
  42458=>"011111111",
  42459=>"011111111",
  42460=>"111111001",
  42461=>"111010010",
  42462=>"101100000",
  42463=>"000000000",
  42464=>"111111111",
  42465=>"000111001",
  42466=>"011111111",
  42467=>"111111111",
  42468=>"010111111",
  42469=>"101001000",
  42470=>"000011011",
  42471=>"000000100",
  42472=>"000000000",
  42473=>"000000000",
  42474=>"111110000",
  42475=>"100000000",
  42476=>"001011111",
  42477=>"000000100",
  42478=>"011011011",
  42479=>"000000000",
  42480=>"000111111",
  42481=>"110011000",
  42482=>"000000100",
  42483=>"111111111",
  42484=>"111111101",
  42485=>"111111111",
  42486=>"001111111",
  42487=>"001001001",
  42488=>"011011000",
  42489=>"100110110",
  42490=>"111110100",
  42491=>"111111111",
  42492=>"111111111",
  42493=>"000001111",
  42494=>"111111011",
  42495=>"011111111",
  42496=>"110010000",
  42497=>"000001101",
  42498=>"000000111",
  42499=>"000000000",
  42500=>"100100100",
  42501=>"111000000",
  42502=>"111000000",
  42503=>"111111111",
  42504=>"111000000",
  42505=>"000111110",
  42506=>"100000000",
  42507=>"000111011",
  42508=>"000100110",
  42509=>"111000000",
  42510=>"011001001",
  42511=>"111111111",
  42512=>"111001011",
  42513=>"000000100",
  42514=>"000000000",
  42515=>"111111011",
  42516=>"000000111",
  42517=>"101100111",
  42518=>"101111101",
  42519=>"000000111",
  42520=>"000001001",
  42521=>"000000000",
  42522=>"011000111",
  42523=>"100100110",
  42524=>"110110111",
  42525=>"001011110",
  42526=>"101100001",
  42527=>"111111000",
  42528=>"000000010",
  42529=>"000001011",
  42530=>"010110000",
  42531=>"000000111",
  42532=>"111110000",
  42533=>"111111011",
  42534=>"101101000",
  42535=>"000111001",
  42536=>"000011111",
  42537=>"000000111",
  42538=>"111111000",
  42539=>"000000000",
  42540=>"101111101",
  42541=>"001111111",
  42542=>"000111111",
  42543=>"000111110",
  42544=>"111001001",
  42545=>"000000011",
  42546=>"111111111",
  42547=>"000001001",
  42548=>"110110000",
  42549=>"000110111",
  42550=>"111111111",
  42551=>"111000000",
  42552=>"110110000",
  42553=>"111111000",
  42554=>"000000000",
  42555=>"000111111",
  42556=>"111001000",
  42557=>"000101111",
  42558=>"000011011",
  42559=>"000000000",
  42560=>"000100000",
  42561=>"000000000",
  42562=>"010111111",
  42563=>"100100100",
  42564=>"110110000",
  42565=>"001011110",
  42566=>"000110111",
  42567=>"000000001",
  42568=>"111011000",
  42569=>"000000000",
  42570=>"011001000",
  42571=>"111111001",
  42572=>"100101000",
  42573=>"111111011",
  42574=>"000000010",
  42575=>"111111111",
  42576=>"111111001",
  42577=>"001001111",
  42578=>"110000000",
  42579=>"111011000",
  42580=>"111110000",
  42581=>"000000000",
  42582=>"000001101",
  42583=>"000000000",
  42584=>"011101000",
  42585=>"000000000",
  42586=>"001111111",
  42587=>"011001011",
  42588=>"000000001",
  42589=>"000000000",
  42590=>"111111111",
  42591=>"111110101",
  42592=>"000000000",
  42593=>"111111111",
  42594=>"100000001",
  42595=>"000000111",
  42596=>"000000000",
  42597=>"101000000",
  42598=>"111111111",
  42599=>"000000000",
  42600=>"000111111",
  42601=>"000000000",
  42602=>"010000111",
  42603=>"111001000",
  42604=>"010111110",
  42605=>"000000000",
  42606=>"111111111",
  42607=>"000000000",
  42608=>"111111111",
  42609=>"000000001",
  42610=>"000001001",
  42611=>"111111001",
  42612=>"111000000",
  42613=>"000000000",
  42614=>"110000000",
  42615=>"000100111",
  42616=>"000101001",
  42617=>"001000000",
  42618=>"000000000",
  42619=>"000000111",
  42620=>"110000001",
  42621=>"000111001",
  42622=>"000000000",
  42623=>"000000000",
  42624=>"000000111",
  42625=>"011111111",
  42626=>"110110111",
  42627=>"011111111",
  42628=>"111111111",
  42629=>"000000011",
  42630=>"101110100",
  42631=>"110010010",
  42632=>"000000111",
  42633=>"000000000",
  42634=>"001000000",
  42635=>"111000010",
  42636=>"000000000",
  42637=>"001000000",
  42638=>"111111011",
  42639=>"000000000",
  42640=>"000111111",
  42641=>"000000000",
  42642=>"000111111",
  42643=>"111011000",
  42644=>"000100000",
  42645=>"111111110",
  42646=>"111111000",
  42647=>"111111111",
  42648=>"000001100",
  42649=>"000000111",
  42650=>"000000110",
  42651=>"111101001",
  42652=>"111111101",
  42653=>"000110111",
  42654=>"111111111",
  42655=>"111111000",
  42656=>"000000000",
  42657=>"000000000",
  42658=>"110101000",
  42659=>"111001111",
  42660=>"000000101",
  42661=>"111111000",
  42662=>"111111111",
  42663=>"100111110",
  42664=>"001001111",
  42665=>"000000111",
  42666=>"111010000",
  42667=>"000000000",
  42668=>"110111111",
  42669=>"100001001",
  42670=>"000111111",
  42671=>"000111111",
  42672=>"111111111",
  42673=>"010001000",
  42674=>"111111111",
  42675=>"000000000",
  42676=>"100000000",
  42677=>"100000000",
  42678=>"000000000",
  42679=>"101111111",
  42680=>"111111000",
  42681=>"000000111",
  42682=>"000001111",
  42683=>"000111111",
  42684=>"000000110",
  42685=>"100000111",
  42686=>"000000010",
  42687=>"111111111",
  42688=>"100101111",
  42689=>"011100101",
  42690=>"010000011",
  42691=>"111111111",
  42692=>"111111100",
  42693=>"000111111",
  42694=>"000100000",
  42695=>"001000000",
  42696=>"101000000",
  42697=>"100000000",
  42698=>"011100000",
  42699=>"000000111",
  42700=>"000000000",
  42701=>"011111000",
  42702=>"111010000",
  42703=>"000000100",
  42704=>"000010111",
  42705=>"100000000",
  42706=>"111111111",
  42707=>"000000111",
  42708=>"000000000",
  42709=>"111011011",
  42710=>"001010000",
  42711=>"001111100",
  42712=>"001111111",
  42713=>"111111111",
  42714=>"000110010",
  42715=>"000000000",
  42716=>"011011111",
  42717=>"000000000",
  42718=>"000100111",
  42719=>"111111100",
  42720=>"111100100",
  42721=>"001001001",
  42722=>"111111111",
  42723=>"111101001",
  42724=>"000000000",
  42725=>"111110100",
  42726=>"000000011",
  42727=>"111111000",
  42728=>"111000111",
  42729=>"011111111",
  42730=>"111111111",
  42731=>"111110111",
  42732=>"000000000",
  42733=>"000000000",
  42734=>"111111101",
  42735=>"000000000",
  42736=>"110111111",
  42737=>"110111101",
  42738=>"111111111",
  42739=>"000000110",
  42740=>"100100000",
  42741=>"111111100",
  42742=>"110000000",
  42743=>"111111110",
  42744=>"000011111",
  42745=>"001001111",
  42746=>"111111110",
  42747=>"000000000",
  42748=>"000011001",
  42749=>"000000001",
  42750=>"000111111",
  42751=>"011000000",
  42752=>"110111111",
  42753=>"111110101",
  42754=>"000000101",
  42755=>"000000000",
  42756=>"111111111",
  42757=>"100000000",
  42758=>"001001101",
  42759=>"000101101",
  42760=>"101111111",
  42761=>"101111111",
  42762=>"111111111",
  42763=>"111111000",
  42764=>"111101111",
  42765=>"000001111",
  42766=>"110110011",
  42767=>"000000000",
  42768=>"111111000",
  42769=>"000000000",
  42770=>"000000000",
  42771=>"111111111",
  42772=>"110000000",
  42773=>"000000101",
  42774=>"001001001",
  42775=>"000011000",
  42776=>"000000111",
  42777=>"110000000",
  42778=>"111111111",
  42779=>"111011000",
  42780=>"111111111",
  42781=>"000000000",
  42782=>"111111111",
  42783=>"000000000",
  42784=>"111111000",
  42785=>"000001000",
  42786=>"000100000",
  42787=>"001001011",
  42788=>"000000111",
  42789=>"111111111",
  42790=>"111101000",
  42791=>"011100000",
  42792=>"011000000",
  42793=>"000000111",
  42794=>"000000110",
  42795=>"000000000",
  42796=>"001000000",
  42797=>"111111000",
  42798=>"111111101",
  42799=>"000000111",
  42800=>"011011001",
  42801=>"000000000",
  42802=>"001011110",
  42803=>"000111111",
  42804=>"000000000",
  42805=>"000111111",
  42806=>"111101100",
  42807=>"111100111",
  42808=>"110110000",
  42809=>"000011011",
  42810=>"000010010",
  42811=>"111111000",
  42812=>"100100000",
  42813=>"111100000",
  42814=>"000111111",
  42815=>"000101000",
  42816=>"111111000",
  42817=>"000111111",
  42818=>"000000001",
  42819=>"000000111",
  42820=>"101100111",
  42821=>"111000000",
  42822=>"000000001",
  42823=>"001000000",
  42824=>"111111111",
  42825=>"000000000",
  42826=>"000100100",
  42827=>"000000111",
  42828=>"011000000",
  42829=>"111000000",
  42830=>"000000000",
  42831=>"000000000",
  42832=>"111111111",
  42833=>"000000000",
  42834=>"000011111",
  42835=>"111111001",
  42836=>"111000000",
  42837=>"011001000",
  42838=>"100100001",
  42839=>"000000111",
  42840=>"111111000",
  42841=>"111111111",
  42842=>"111111110",
  42843=>"111111000",
  42844=>"000000000",
  42845=>"000111111",
  42846=>"000000000",
  42847=>"110010001",
  42848=>"011111111",
  42849=>"000000000",
  42850=>"011011011",
  42851=>"000001010",
  42852=>"111100000",
  42853=>"001111111",
  42854=>"111111111",
  42855=>"111111011",
  42856=>"000100100",
  42857=>"111010110",
  42858=>"000100000",
  42859=>"110110110",
  42860=>"111011001",
  42861=>"000011011",
  42862=>"000000000",
  42863=>"000000000",
  42864=>"001011101",
  42865=>"111001001",
  42866=>"111000000",
  42867=>"011011000",
  42868=>"000000000",
  42869=>"111111111",
  42870=>"111111111",
  42871=>"000000000",
  42872=>"000111111",
  42873=>"111100000",
  42874=>"000000111",
  42875=>"111000000",
  42876=>"000111111",
  42877=>"111111111",
  42878=>"000001111",
  42879=>"111111111",
  42880=>"110011111",
  42881=>"111111111",
  42882=>"110111011",
  42883=>"000000000",
  42884=>"010110010",
  42885=>"000001000",
  42886=>"000110111",
  42887=>"111111111",
  42888=>"010111111",
  42889=>"000110110",
  42890=>"111111001",
  42891=>"111111111",
  42892=>"111011111",
  42893=>"111000000",
  42894=>"101000101",
  42895=>"000000111",
  42896=>"111111111",
  42897=>"001000000",
  42898=>"111111000",
  42899=>"010011000",
  42900=>"111000000",
  42901=>"000000000",
  42902=>"000000001",
  42903=>"000000011",
  42904=>"111111111",
  42905=>"100110000",
  42906=>"000000001",
  42907=>"111111000",
  42908=>"110111000",
  42909=>"110000000",
  42910=>"000000011",
  42911=>"001111110",
  42912=>"111111111",
  42913=>"001001011",
  42914=>"000000000",
  42915=>"111010111",
  42916=>"000000000",
  42917=>"010000000",
  42918=>"000001111",
  42919=>"111000000",
  42920=>"111111111",
  42921=>"111001001",
  42922=>"001111111",
  42923=>"000000110",
  42924=>"000101101",
  42925=>"100000010",
  42926=>"000000101",
  42927=>"011000000",
  42928=>"000000000",
  42929=>"110110100",
  42930=>"000000000",
  42931=>"000111111",
  42932=>"000110111",
  42933=>"010110111",
  42934=>"110000000",
  42935=>"110111111",
  42936=>"001000000",
  42937=>"100000100",
  42938=>"110100110",
  42939=>"001001111",
  42940=>"111111000",
  42941=>"100111111",
  42942=>"111001000",
  42943=>"100110110",
  42944=>"000000010",
  42945=>"000000000",
  42946=>"111111000",
  42947=>"000000000",
  42948=>"110111111",
  42949=>"000010001",
  42950=>"001111101",
  42951=>"011000000",
  42952=>"000111111",
  42953=>"100000001",
  42954=>"111001001",
  42955=>"111110111",
  42956=>"000000000",
  42957=>"111000000",
  42958=>"010111111",
  42959=>"000111111",
  42960=>"000000000",
  42961=>"000000100",
  42962=>"011000000",
  42963=>"110110111",
  42964=>"001000000",
  42965=>"100111111",
  42966=>"110001000",
  42967=>"001001001",
  42968=>"000001000",
  42969=>"011011001",
  42970=>"111111111",
  42971=>"100100110",
  42972=>"111111111",
  42973=>"000100111",
  42974=>"111111111",
  42975=>"111111000",
  42976=>"111111111",
  42977=>"111001001",
  42978=>"100111111",
  42979=>"111111000",
  42980=>"000100100",
  42981=>"010011111",
  42982=>"000110000",
  42983=>"110101001",
  42984=>"111111000",
  42985=>"000010110",
  42986=>"011111111",
  42987=>"111111111",
  42988=>"000111111",
  42989=>"001000100",
  42990=>"100000000",
  42991=>"110000000",
  42992=>"000001111",
  42993=>"000000000",
  42994=>"000011111",
  42995=>"001101000",
  42996=>"110110000",
  42997=>"000000000",
  42998=>"000100111",
  42999=>"011010000",
  43000=>"111000000",
  43001=>"001011000",
  43002=>"110000000",
  43003=>"111111000",
  43004=>"110110000",
  43005=>"110111111",
  43006=>"000111111",
  43007=>"110111000",
  43008=>"111110000",
  43009=>"000000000",
  43010=>"000000100",
  43011=>"000001000",
  43012=>"011111111",
  43013=>"000000000",
  43014=>"000000100",
  43015=>"000000000",
  43016=>"000000000",
  43017=>"111111000",
  43018=>"111111011",
  43019=>"000110110",
  43020=>"000000111",
  43021=>"100000010",
  43022=>"100111111",
  43023=>"000000000",
  43024=>"100110111",
  43025=>"000111111",
  43026=>"011001111",
  43027=>"111101100",
  43028=>"000011111",
  43029=>"000000000",
  43030=>"111111111",
  43031=>"111111111",
  43032=>"111111010",
  43033=>"110111000",
  43034=>"000000000",
  43035=>"111000000",
  43036=>"000100100",
  43037=>"110100100",
  43038=>"111111111",
  43039=>"111000111",
  43040=>"000101111",
  43041=>"000000001",
  43042=>"111111000",
  43043=>"000000100",
  43044=>"000111000",
  43045=>"111100000",
  43046=>"111111111",
  43047=>"000000000",
  43048=>"001000000",
  43049=>"000000000",
  43050=>"000110010",
  43051=>"111111110",
  43052=>"000011111",
  43053=>"111111000",
  43054=>"100100100",
  43055=>"111100100",
  43056=>"111111111",
  43057=>"000100000",
  43058=>"111100100",
  43059=>"011010000",
  43060=>"000001101",
  43061=>"100111011",
  43062=>"101111111",
  43063=>"000010010",
  43064=>"000000000",
  43065=>"111000001",
  43066=>"001011111",
  43067=>"000000000",
  43068=>"111111111",
  43069=>"111111111",
  43070=>"011111111",
  43071=>"001000101",
  43072=>"111111111",
  43073=>"000111111",
  43074=>"111010000",
  43075=>"111000100",
  43076=>"000011011",
  43077=>"000010010",
  43078=>"000000000",
  43079=>"111111111",
  43080=>"000110110",
  43081=>"000000111",
  43082=>"111110000",
  43083=>"000000111",
  43084=>"010000111",
  43085=>"110100111",
  43086=>"000000000",
  43087=>"011111111",
  43088=>"111011111",
  43089=>"101111111",
  43090=>"000010010",
  43091=>"000000000",
  43092=>"000000000",
  43093=>"101111111",
  43094=>"001011011",
  43095=>"000110111",
  43096=>"000000000",
  43097=>"001000000",
  43098=>"100000000",
  43099=>"111111111",
  43100=>"000000000",
  43101=>"111111111",
  43102=>"110110000",
  43103=>"100110110",
  43104=>"001000000",
  43105=>"010000010",
  43106=>"100100000",
  43107=>"000000001",
  43108=>"001000111",
  43109=>"011111111",
  43110=>"000000111",
  43111=>"000000000",
  43112=>"001111011",
  43113=>"000000000",
  43114=>"111111111",
  43115=>"111000000",
  43116=>"110110100",
  43117=>"000000000",
  43118=>"111111111",
  43119=>"010111111",
  43120=>"000011111",
  43121=>"111111011",
  43122=>"111111101",
  43123=>"011000000",
  43124=>"000000111",
  43125=>"111110000",
  43126=>"000000000",
  43127=>"000000000",
  43128=>"000000000",
  43129=>"000000000",
  43130=>"000000000",
  43131=>"111111111",
  43132=>"100110110",
  43133=>"000010010",
  43134=>"000000000",
  43135=>"000000000",
  43136=>"000000000",
  43137=>"111100000",
  43138=>"110000111",
  43139=>"000000000",
  43140=>"000000000",
  43141=>"100000111",
  43142=>"000000001",
  43143=>"000000111",
  43144=>"111111111",
  43145=>"000000111",
  43146=>"000001001",
  43147=>"111100100",
  43148=>"000001000",
  43149=>"111000000",
  43150=>"011111111",
  43151=>"000110110",
  43152=>"111111111",
  43153=>"100101111",
  43154=>"000000011",
  43155=>"110000000",
  43156=>"000000111",
  43157=>"000110110",
  43158=>"000000000",
  43159=>"111100100",
  43160=>"000001001",
  43161=>"111111111",
  43162=>"011111111",
  43163=>"111111111",
  43164=>"010000000",
  43165=>"111011011",
  43166=>"110110111",
  43167=>"000000010",
  43168=>"111011101",
  43169=>"001000000",
  43170=>"111111111",
  43171=>"000000000",
  43172=>"000000000",
  43173=>"000000000",
  43174=>"111000011",
  43175=>"111001001",
  43176=>"111011111",
  43177=>"000000010",
  43178=>"100000000",
  43179=>"111111111",
  43180=>"110101001",
  43181=>"001011000",
  43182=>"111110100",
  43183=>"000000000",
  43184=>"110111111",
  43185=>"011010010",
  43186=>"111111110",
  43187=>"000000000",
  43188=>"001000000",
  43189=>"011001000",
  43190=>"111111111",
  43191=>"000000000",
  43192=>"111010110",
  43193=>"111111000",
  43194=>"000011011",
  43195=>"000000101",
  43196=>"111111111",
  43197=>"111111000",
  43198=>"100000000",
  43199=>"000111001",
  43200=>"111111111",
  43201=>"111111111",
  43202=>"111100000",
  43203=>"100000011",
  43204=>"001011111",
  43205=>"011111111",
  43206=>"111100010",
  43207=>"111111110",
  43208=>"000000000",
  43209=>"000010110",
  43210=>"000010000",
  43211=>"000110000",
  43212=>"111001011",
  43213=>"111111011",
  43214=>"111000000",
  43215=>"011000000",
  43216=>"001000000",
  43217=>"100000001",
  43218=>"000000000",
  43219=>"011111111",
  43220=>"111111111",
  43221=>"111110111",
  43222=>"111111111",
  43223=>"000000000",
  43224=>"101111010",
  43225=>"111001000",
  43226=>"111011010",
  43227=>"001000101",
  43228=>"000000000",
  43229=>"111111111",
  43230=>"111111111",
  43231=>"010111011",
  43232=>"111111100",
  43233=>"000110110",
  43234=>"000000000",
  43235=>"111000100",
  43236=>"111111100",
  43237=>"011010111",
  43238=>"111111111",
  43239=>"000000000",
  43240=>"000100000",
  43241=>"000000000",
  43242=>"001000000",
  43243=>"001011111",
  43244=>"011000011",
  43245=>"000000010",
  43246=>"111001001",
  43247=>"000000111",
  43248=>"100110000",
  43249=>"001000001",
  43250=>"111101000",
  43251=>"000000000",
  43252=>"000000111",
  43253=>"000000000",
  43254=>"111011010",
  43255=>"000110111",
  43256=>"111111111",
  43257=>"011111111",
  43258=>"111001000",
  43259=>"000010111",
  43260=>"110110110",
  43261=>"011111110",
  43262=>"011000000",
  43263=>"000000100",
  43264=>"000000000",
  43265=>"000000000",
  43266=>"000010000",
  43267=>"111001000",
  43268=>"100000000",
  43269=>"000111110",
  43270=>"000000111",
  43271=>"111010111",
  43272=>"111011011",
  43273=>"000110111",
  43274=>"000001111",
  43275=>"011000000",
  43276=>"111111110",
  43277=>"101110111",
  43278=>"000010000",
  43279=>"111111111",
  43280=>"000000000",
  43281=>"111111111",
  43282=>"101101111",
  43283=>"000111110",
  43284=>"000011001",
  43285=>"001000000",
  43286=>"110110011",
  43287=>"000000111",
  43288=>"001001010",
  43289=>"100100111",
  43290=>"111000111",
  43291=>"000000111",
  43292=>"111111011",
  43293=>"111111010",
  43294=>"001011111",
  43295=>"000011111",
  43296=>"100000000",
  43297=>"001001011",
  43298=>"000000010",
  43299=>"111111111",
  43300=>"000110010",
  43301=>"000000000",
  43302=>"011000111",
  43303=>"111111000",
  43304=>"000000000",
  43305=>"000011010",
  43306=>"110111111",
  43307=>"000000000",
  43308=>"110110111",
  43309=>"111111110",
  43310=>"000000000",
  43311=>"000111110",
  43312=>"110110111",
  43313=>"011111111",
  43314=>"110111111",
  43315=>"000111111",
  43316=>"000000000",
  43317=>"000000000",
  43318=>"001000011",
  43319=>"000001000",
  43320=>"000000000",
  43321=>"000000111",
  43322=>"000000000",
  43323=>"000001000",
  43324=>"111010110",
  43325=>"110000000",
  43326=>"111111111",
  43327=>"111111111",
  43328=>"101101101",
  43329=>"000000000",
  43330=>"000000100",
  43331=>"000111011",
  43332=>"111111010",
  43333=>"111111111",
  43334=>"010010000",
  43335=>"000001001",
  43336=>"000000010",
  43337=>"111000000",
  43338=>"000000000",
  43339=>"111011011",
  43340=>"000000000",
  43341=>"011000000",
  43342=>"101000110",
  43343=>"000000000",
  43344=>"111111111",
  43345=>"000000000",
  43346=>"001000111",
  43347=>"001111111",
  43348=>"111001011",
  43349=>"011011111",
  43350=>"000000000",
  43351=>"111111100",
  43352=>"000000110",
  43353=>"111001000",
  43354=>"111111000",
  43355=>"011010010",
  43356=>"000000101",
  43357=>"010111111",
  43358=>"001000000",
  43359=>"011111011",
  43360=>"000000000",
  43361=>"000000000",
  43362=>"111101110",
  43363=>"000000000",
  43364=>"011111001",
  43365=>"011001000",
  43366=>"010000000",
  43367=>"111111001",
  43368=>"111110000",
  43369=>"110000000",
  43370=>"000000000",
  43371=>"100000000",
  43372=>"111001001",
  43373=>"000000111",
  43374=>"001111111",
  43375=>"111111011",
  43376=>"111111111",
  43377=>"111000000",
  43378=>"001100010",
  43379=>"000001000",
  43380=>"111111000",
  43381=>"110110000",
  43382=>"111111110",
  43383=>"000000111",
  43384=>"000000000",
  43385=>"000000000",
  43386=>"000000000",
  43387=>"011000000",
  43388=>"000000000",
  43389=>"110100110",
  43390=>"111111111",
  43391=>"011111111",
  43392=>"011011111",
  43393=>"010011000",
  43394=>"110011011",
  43395=>"000000001",
  43396=>"010110100",
  43397=>"111000000",
  43398=>"110110010",
  43399=>"100000000",
  43400=>"010010110",
  43401=>"000000111",
  43402=>"111100000",
  43403=>"101111111",
  43404=>"111111111",
  43405=>"000001111",
  43406=>"100000000",
  43407=>"000000001",
  43408=>"000000100",
  43409=>"111011001",
  43410=>"000010000",
  43411=>"011011011",
  43412=>"001111111",
  43413=>"000000000",
  43414=>"000000000",
  43415=>"000100110",
  43416=>"111100111",
  43417=>"111011000",
  43418=>"101100000",
  43419=>"111111010",
  43420=>"000000000",
  43421=>"000010110",
  43422=>"000000000",
  43423=>"001000110",
  43424=>"000110111",
  43425=>"110110110",
  43426=>"011101111",
  43427=>"000110000",
  43428=>"001000000",
  43429=>"000000000",
  43430=>"000110000",
  43431=>"000000000",
  43432=>"110000011",
  43433=>"111111110",
  43434=>"000000000",
  43435=>"001011000",
  43436=>"000000000",
  43437=>"111111111",
  43438=>"000000101",
  43439=>"011000000",
  43440=>"110111110",
  43441=>"000000000",
  43442=>"001001111",
  43443=>"001000111",
  43444=>"000000000",
  43445=>"111111111",
  43446=>"000100000",
  43447=>"001111111",
  43448=>"000001111",
  43449=>"001111111",
  43450=>"111111010",
  43451=>"001000000",
  43452=>"000000000",
  43453=>"110110110",
  43454=>"001000000",
  43455=>"101100000",
  43456=>"111011011",
  43457=>"111111111",
  43458=>"000000000",
  43459=>"001000000",
  43460=>"111011111",
  43461=>"010110100",
  43462=>"110100101",
  43463=>"000001001",
  43464=>"000000100",
  43465=>"000000000",
  43466=>"111111111",
  43467=>"010000000",
  43468=>"011000000",
  43469=>"111111111",
  43470=>"100000000",
  43471=>"011110000",
  43472=>"111110110",
  43473=>"000110110",
  43474=>"001000001",
  43475=>"111111011",
  43476=>"011011111",
  43477=>"101100000",
  43478=>"110100111",
  43479=>"000100100",
  43480=>"111111110",
  43481=>"111000100",
  43482=>"000000000",
  43483=>"110000000",
  43484=>"001111111",
  43485=>"001000100",
  43486=>"000000000",
  43487=>"111111110",
  43488=>"000000000",
  43489=>"111111001",
  43490=>"000111111",
  43491=>"000000000",
  43492=>"111111111",
  43493=>"001000000",
  43494=>"111111111",
  43495=>"001001000",
  43496=>"111111100",
  43497=>"001001101",
  43498=>"000011011",
  43499=>"000111111",
  43500=>"011000000",
  43501=>"110111110",
  43502=>"111111111",
  43503=>"000000000",
  43504=>"000000000",
  43505=>"000000011",
  43506=>"000001000",
  43507=>"111111001",
  43508=>"011111010",
  43509=>"001001111",
  43510=>"111110000",
  43511=>"000001011",
  43512=>"000000100",
  43513=>"011011010",
  43514=>"000111110",
  43515=>"001000010",
  43516=>"111111111",
  43517=>"100000110",
  43518=>"111111110",
  43519=>"000000000",
  43520=>"111111111",
  43521=>"111001011",
  43522=>"100100111",
  43523=>"001001001",
  43524=>"111010010",
  43525=>"000000000",
  43526=>"000000010",
  43527=>"010010010",
  43528=>"111101100",
  43529=>"110101001",
  43530=>"101001001",
  43531=>"011011001",
  43532=>"000010100",
  43533=>"010010011",
  43534=>"011011011",
  43535=>"000010011",
  43536=>"111111111",
  43537=>"001111001",
  43538=>"000000010",
  43539=>"111011000",
  43540=>"101101101",
  43541=>"101000100",
  43542=>"100000010",
  43543=>"100100110",
  43544=>"111101001",
  43545=>"010010000",
  43546=>"000000000",
  43547=>"111100000",
  43548=>"110010000",
  43549=>"000001111",
  43550=>"001011011",
  43551=>"011011000",
  43552=>"100101001",
  43553=>"001011001",
  43554=>"000110110",
  43555=>"100100100",
  43556=>"101101100",
  43557=>"011111100",
  43558=>"101111000",
  43559=>"111010001",
  43560=>"110110011",
  43561=>"111111111",
  43562=>"011011111",
  43563=>"111111011",
  43564=>"101111000",
  43565=>"111100011",
  43566=>"010010010",
  43567=>"000000001",
  43568=>"000000000",
  43569=>"000000000",
  43570=>"100100110",
  43571=>"100111111",
  43572=>"010110010",
  43573=>"000110110",
  43574=>"000010010",
  43575=>"010000101",
  43576=>"000011101",
  43577=>"101111010",
  43578=>"011011011",
  43579=>"111111111",
  43580=>"011011111",
  43581=>"100110111",
  43582=>"010010010",
  43583=>"111111111",
  43584=>"000011011",
  43585=>"111111111",
  43586=>"111101100",
  43587=>"111100101",
  43588=>"001001000",
  43589=>"000010010",
  43590=>"111111100",
  43591=>"000000001",
  43592=>"110110110",
  43593=>"101101111",
  43594=>"011011011",
  43595=>"001000000",
  43596=>"111111111",
  43597=>"100111010",
  43598=>"101101111",
  43599=>"110110010",
  43600=>"111001011",
  43601=>"001001001",
  43602=>"110110000",
  43603=>"010110110",
  43604=>"010010000",
  43605=>"111111001",
  43606=>"111000000",
  43607=>"000000010",
  43608=>"100100110",
  43609=>"111111011",
  43610=>"100100111",
  43611=>"000111111",
  43612=>"000100111",
  43613=>"101101100",
  43614=>"111111111",
  43615=>"000000010",
  43616=>"001000000",
  43617=>"001101101",
  43618=>"001011011",
  43619=>"110010000",
  43620=>"010000000",
  43621=>"101101000",
  43622=>"000000101",
  43623=>"000101111",
  43624=>"000000000",
  43625=>"100001001",
  43626=>"111001001",
  43627=>"000000101",
  43628=>"111111111",
  43629=>"000000010",
  43630=>"011010000",
  43631=>"101101101",
  43632=>"001101101",
  43633=>"000000000",
  43634=>"000010010",
  43635=>"111101001",
  43636=>"111111011",
  43637=>"000001001",
  43638=>"110110110",
  43639=>"100101101",
  43640=>"100000000",
  43641=>"010001111",
  43642=>"000101111",
  43643=>"101111111",
  43644=>"011010011",
  43645=>"000011011",
  43646=>"000010010",
  43647=>"000000000",
  43648=>"111101000",
  43649=>"111111001",
  43650=>"010011001",
  43651=>"111111000",
  43652=>"010011010",
  43653=>"111110110",
  43654=>"001001111",
  43655=>"000000001",
  43656=>"000000001",
  43657=>"110110010",
  43658=>"111111111",
  43659=>"111011000",
  43660=>"111101101",
  43661=>"011011000",
  43662=>"000001001",
  43663=>"000010010",
  43664=>"111101111",
  43665=>"110111000",
  43666=>"111111111",
  43667=>"000000001",
  43668=>"111111011",
  43669=>"010110000",
  43670=>"111011111",
  43671=>"011111001",
  43672=>"111111111",
  43673=>"010010010",
  43674=>"000000000",
  43675=>"111111111",
  43676=>"000111111",
  43677=>"110000000",
  43678=>"010011011",
  43679=>"111111011",
  43680=>"110110110",
  43681=>"000000111",
  43682=>"010011011",
  43683=>"110110111",
  43684=>"100100100",
  43685=>"000000000",
  43686=>"000001001",
  43687=>"000110000",
  43688=>"000000000",
  43689=>"001001001",
  43690=>"000101101",
  43691=>"111011111",
  43692=>"100101111",
  43693=>"111111111",
  43694=>"001001111",
  43695=>"111111111",
  43696=>"111111111",
  43697=>"111111110",
  43698=>"000000001",
  43699=>"101111111",
  43700=>"110111110",
  43701=>"011011110",
  43702=>"001111111",
  43703=>"111111111",
  43704=>"000000000",
  43705=>"010010010",
  43706=>"000000110",
  43707=>"111111110",
  43708=>"100100101",
  43709=>"110000000",
  43710=>"000110000",
  43711=>"101000100",
  43712=>"111111011",
  43713=>"111111111",
  43714=>"000000000",
  43715=>"001000100",
  43716=>"001000001",
  43717=>"101001011",
  43718=>"101101101",
  43719=>"111111111",
  43720=>"111001101",
  43721=>"010010010",
  43722=>"111101001",
  43723=>"111111111",
  43724=>"000000011",
  43725=>"001001001",
  43726=>"000000111",
  43727=>"100000011",
  43728=>"000000101",
  43729=>"010010111",
  43730=>"000010000",
  43731=>"110110010",
  43732=>"001000000",
  43733=>"011100000",
  43734=>"110111111",
  43735=>"110101000",
  43736=>"010000111",
  43737=>"000100110",
  43738=>"100101101",
  43739=>"010000000",
  43740=>"100010010",
  43741=>"010010010",
  43742=>"100000101",
  43743=>"101111111",
  43744=>"100100001",
  43745=>"011010101",
  43746=>"111111111",
  43747=>"111110010",
  43748=>"011001000",
  43749=>"100111110",
  43750=>"101101101",
  43751=>"000010010",
  43752=>"001001000",
  43753=>"000111011",
  43754=>"000000000",
  43755=>"000000101",
  43756=>"111011011",
  43757=>"101101101",
  43758=>"000001111",
  43759=>"000000000",
  43760=>"101101101",
  43761=>"100100101",
  43762=>"010010010",
  43763=>"010110111",
  43764=>"101111111",
  43765=>"000000000",
  43766=>"111100111",
  43767=>"000010010",
  43768=>"101001000",
  43769=>"000000000",
  43770=>"010010011",
  43771=>"000000001",
  43772=>"101101000",
  43773=>"001001001",
  43774=>"100000101",
  43775=>"011011000",
  43776=>"010011000",
  43777=>"011011011",
  43778=>"000000001",
  43779=>"111011011",
  43780=>"000000000",
  43781=>"110110111",
  43782=>"000000001",
  43783=>"001000101",
  43784=>"000000101",
  43785=>"100000000",
  43786=>"010000000",
  43787=>"001001011",
  43788=>"101000000",
  43789=>"001000111",
  43790=>"101001101",
  43791=>"111111111",
  43792=>"010000010",
  43793=>"111111111",
  43794=>"101101000",
  43795=>"010010110",
  43796=>"000011001",
  43797=>"001101101",
  43798=>"011011011",
  43799=>"111111010",
  43800=>"110110001",
  43801=>"101100001",
  43802=>"001111011",
  43803=>"111100100",
  43804=>"001110110",
  43805=>"110000000",
  43806=>"010010010",
  43807=>"110101111",
  43808=>"111111101",
  43809=>"110010110",
  43810=>"101101101",
  43811=>"010000000",
  43812=>"111011001",
  43813=>"000000010",
  43814=>"001111111",
  43815=>"101101111",
  43816=>"010011000",
  43817=>"000000000",
  43818=>"110110111",
  43819=>"000110100",
  43820=>"011000000",
  43821=>"001001001",
  43822=>"111011010",
  43823=>"010010010",
  43824=>"011010011",
  43825=>"000000000",
  43826=>"101101101",
  43827=>"101101101",
  43828=>"111111111",
  43829=>"001001001",
  43830=>"001101101",
  43831=>"000000000",
  43832=>"001001000",
  43833=>"000011111",
  43834=>"100110110",
  43835=>"111111011",
  43836=>"101101101",
  43837=>"011010011",
  43838=>"100111111",
  43839=>"000000000",
  43840=>"101101101",
  43841=>"111111111",
  43842=>"000000000",
  43843=>"010010010",
  43844=>"111111000",
  43845=>"100101100",
  43846=>"010111010",
  43847=>"111010010",
  43848=>"100100000",
  43849=>"101100100",
  43850=>"111111000",
  43851=>"111100110",
  43852=>"010000001",
  43853=>"000000000",
  43854=>"011111000",
  43855=>"100110100",
  43856=>"100110000",
  43857=>"111111101",
  43858=>"100111111",
  43859=>"100000000",
  43860=>"000000000",
  43861=>"111111111",
  43862=>"000000010",
  43863=>"001000001",
  43864=>"010110010",
  43865=>"010000000",
  43866=>"001001000",
  43867=>"000000100",
  43868=>"111000110",
  43869=>"000000000",
  43870=>"000111100",
  43871=>"001001111",
  43872=>"111001101",
  43873=>"101101001",
  43874=>"111111110",
  43875=>"011011011",
  43876=>"111100100",
  43877=>"010000000",
  43878=>"000001001",
  43879=>"111010011",
  43880=>"001011011",
  43881=>"011000000",
  43882=>"110111110",
  43883=>"001000011",
  43884=>"101001001",
  43885=>"101101100",
  43886=>"000010011",
  43887=>"111011000",
  43888=>"101101101",
  43889=>"111001001",
  43890=>"111101000",
  43891=>"011001001",
  43892=>"101100100",
  43893=>"010010010",
  43894=>"000100110",
  43895=>"011101111",
  43896=>"010010011",
  43897=>"111000011",
  43898=>"100101111",
  43899=>"000000011",
  43900=>"000001001",
  43901=>"000010010",
  43902=>"111101101",
  43903=>"001001011",
  43904=>"110110000",
  43905=>"111011111",
  43906=>"000000100",
  43907=>"111111101",
  43908=>"011111101",
  43909=>"000000000",
  43910=>"001001101",
  43911=>"000000111",
  43912=>"001001001",
  43913=>"001001001",
  43914=>"001110010",
  43915=>"111111111",
  43916=>"110110111",
  43917=>"010011001",
  43918=>"111111010",
  43919=>"001101001",
  43920=>"101100100",
  43921=>"110110110",
  43922=>"111100111",
  43923=>"001001001",
  43924=>"001000001",
  43925=>"101101000",
  43926=>"111000000",
  43927=>"110010000",
  43928=>"111111111",
  43929=>"001000000",
  43930=>"111111111",
  43931=>"010011111",
  43932=>"000110111",
  43933=>"000110111",
  43934=>"000000100",
  43935=>"000000000",
  43936=>"101101101",
  43937=>"110010010",
  43938=>"111010000",
  43939=>"000100000",
  43940=>"011010000",
  43941=>"101101001",
  43942=>"111110100",
  43943=>"101111111",
  43944=>"111010110",
  43945=>"100100101",
  43946=>"000000010",
  43947=>"000100010",
  43948=>"000000000",
  43949=>"111001111",
  43950=>"101111111",
  43951=>"000100100",
  43952=>"101101111",
  43953=>"011000000",
  43954=>"111111111",
  43955=>"100100000",
  43956=>"111111111",
  43957=>"111111110",
  43958=>"000110010",
  43959=>"111111111",
  43960=>"100110111",
  43961=>"101101101",
  43962=>"000000000",
  43963=>"000110011",
  43964=>"001000000",
  43965=>"111011000",
  43966=>"100001001",
  43967=>"011001000",
  43968=>"110000111",
  43969=>"101101111",
  43970=>"000000000",
  43971=>"100100000",
  43972=>"101010110",
  43973=>"111110000",
  43974=>"111001101",
  43975=>"000000000",
  43976=>"001111111",
  43977=>"111101100",
  43978=>"000010010",
  43979=>"001011111",
  43980=>"001001001",
  43981=>"111111100",
  43982=>"111011111",
  43983=>"101101100",
  43984=>"001000101",
  43985=>"111011001",
  43986=>"010001001",
  43987=>"111111110",
  43988=>"000001111",
  43989=>"000011011",
  43990=>"111111111",
  43991=>"001001001",
  43992=>"111111111",
  43993=>"100111011",
  43994=>"101100100",
  43995=>"000011000",
  43996=>"000011001",
  43997=>"011010001",
  43998=>"100100100",
  43999=>"001011010",
  44000=>"011001101",
  44001=>"000000000",
  44002=>"100100010",
  44003=>"100000100",
  44004=>"000100100",
  44005=>"000100110",
  44006=>"110000000",
  44007=>"100100101",
  44008=>"010011011",
  44009=>"101111111",
  44010=>"110101101",
  44011=>"000001011",
  44012=>"111111111",
  44013=>"111011001",
  44014=>"110110111",
  44015=>"010111111",
  44016=>"000000011",
  44017=>"101111111",
  44018=>"000000010",
  44019=>"111100110",
  44020=>"110110111",
  44021=>"000000100",
  44022=>"001001000",
  44023=>"011011111",
  44024=>"111111111",
  44025=>"110111111",
  44026=>"000000000",
  44027=>"111101101",
  44028=>"001000000",
  44029=>"111011011",
  44030=>"110010010",
  44031=>"110110110",
  44032=>"111111111",
  44033=>"001000000",
  44034=>"000100000",
  44035=>"101111111",
  44036=>"011111111",
  44037=>"001000101",
  44038=>"111111111",
  44039=>"100000000",
  44040=>"100111110",
  44041=>"000000110",
  44042=>"000000000",
  44043=>"000000111",
  44044=>"100000000",
  44045=>"111001110",
  44046=>"000000000",
  44047=>"111111111",
  44048=>"111100111",
  44049=>"111111111",
  44050=>"010000000",
  44051=>"110110110",
  44052=>"111111111",
  44053=>"111111111",
  44054=>"110011111",
  44055=>"000010110",
  44056=>"110110111",
  44057=>"111110100",
  44058=>"111111111",
  44059=>"100100110",
  44060=>"000001000",
  44061=>"000110000",
  44062=>"000000000",
  44063=>"000000000",
  44064=>"111000000",
  44065=>"111001111",
  44066=>"111010000",
  44067=>"011011000",
  44068=>"000000000",
  44069=>"111000101",
  44070=>"010000011",
  44071=>"010111011",
  44072=>"000000111",
  44073=>"000001001",
  44074=>"100111111",
  44075=>"111111000",
  44076=>"111111111",
  44077=>"111000000",
  44078=>"011111011",
  44079=>"000111000",
  44080=>"000000110",
  44081=>"000000000",
  44082=>"111111111",
  44083=>"111111111",
  44084=>"111000000",
  44085=>"000100100",
  44086=>"111000000",
  44087=>"010110110",
  44088=>"111111111",
  44089=>"111011111",
  44090=>"000000111",
  44091=>"111111010",
  44092=>"111100000",
  44093=>"111011011",
  44094=>"001001001",
  44095=>"000000100",
  44096=>"111111111",
  44097=>"111111111",
  44098=>"001111111",
  44099=>"111111110",
  44100=>"110111111",
  44101=>"110110100",
  44102=>"000000111",
  44103=>"000000000",
  44104=>"000000000",
  44105=>"001001001",
  44106=>"010000000",
  44107=>"000000000",
  44108=>"001011111",
  44109=>"000000000",
  44110=>"000000000",
  44111=>"111111011",
  44112=>"111111111",
  44113=>"110000000",
  44114=>"000000100",
  44115=>"000000010",
  44116=>"111111111",
  44117=>"001001101",
  44118=>"111000001",
  44119=>"100000100",
  44120=>"000000000",
  44121=>"000111111",
  44122=>"000001011",
  44123=>"000100111",
  44124=>"111111111",
  44125=>"111100111",
  44126=>"100100100",
  44127=>"011111111",
  44128=>"011011011",
  44129=>"111100000",
  44130=>"111100111",
  44131=>"000001010",
  44132=>"001000000",
  44133=>"100000000",
  44134=>"001100111",
  44135=>"000000000",
  44136=>"111111100",
  44137=>"000000001",
  44138=>"000000100",
  44139=>"011000101",
  44140=>"000100110",
  44141=>"000100100",
  44142=>"000001111",
  44143=>"000101111",
  44144=>"111111111",
  44145=>"011111111",
  44146=>"000000010",
  44147=>"000000000",
  44148=>"111110000",
  44149=>"100110111",
  44150=>"000000000",
  44151=>"111111111",
  44152=>"111011011",
  44153=>"000000110",
  44154=>"000000011",
  44155=>"000000000",
  44156=>"000110110",
  44157=>"111111111",
  44158=>"000000000",
  44159=>"011011011",
  44160=>"000111111",
  44161=>"111100000",
  44162=>"111111111",
  44163=>"000000000",
  44164=>"000011000",
  44165=>"011000000",
  44166=>"011110100",
  44167=>"000110100",
  44168=>"101111000",
  44169=>"110000000",
  44170=>"011011111",
  44171=>"000000000",
  44172=>"111111111",
  44173=>"110110000",
  44174=>"000111110",
  44175=>"100110110",
  44176=>"000000000",
  44177=>"000111111",
  44178=>"111110100",
  44179=>"111011000",
  44180=>"000000000",
  44181=>"000000000",
  44182=>"111111111",
  44183=>"000000000",
  44184=>"110000110",
  44185=>"000001000",
  44186=>"111111111",
  44187=>"111100110",
  44188=>"100110111",
  44189=>"000000111",
  44190=>"111001000",
  44191=>"111111011",
  44192=>"000000011",
  44193=>"111010000",
  44194=>"111011000",
  44195=>"111111111",
  44196=>"000000000",
  44197=>"000100100",
  44198=>"001001011",
  44199=>"000000000",
  44200=>"000000000",
  44201=>"011000100",
  44202=>"011011000",
  44203=>"111011111",
  44204=>"111011001",
  44205=>"010011001",
  44206=>"010010000",
  44207=>"000000000",
  44208=>"000010111",
  44209=>"001001011",
  44210=>"011111111",
  44211=>"000000000",
  44212=>"100100111",
  44213=>"111110000",
  44214=>"110111111",
  44215=>"000000001",
  44216=>"000000000",
  44217=>"111000000",
  44218=>"000000000",
  44219=>"110100000",
  44220=>"000000111",
  44221=>"000001001",
  44222=>"010000000",
  44223=>"111111111",
  44224=>"000111100",
  44225=>"001000111",
  44226=>"000000000",
  44227=>"000000111",
  44228=>"000000000",
  44229=>"010110000",
  44230=>"000100111",
  44231=>"000000111",
  44232=>"111111111",
  44233=>"011111111",
  44234=>"111111111",
  44235=>"011011000",
  44236=>"111010000",
  44237=>"000000000",
  44238=>"000000000",
  44239=>"111111101",
  44240=>"111111111",
  44241=>"000000011",
  44242=>"111010000",
  44243=>"000000000",
  44244=>"010000000",
  44245=>"011001000",
  44246=>"111111111",
  44247=>"001000000",
  44248=>"000000110",
  44249=>"111111111",
  44250=>"000000000",
  44251=>"000000000",
  44252=>"111011000",
  44253=>"000100100",
  44254=>"000100100",
  44255=>"110010011",
  44256=>"111111101",
  44257=>"111111111",
  44258=>"111111000",
  44259=>"000000000",
  44260=>"101101101",
  44261=>"110111111",
  44262=>"001111111",
  44263=>"111111111",
  44264=>"111111111",
  44265=>"000000000",
  44266=>"110000111",
  44267=>"000000001",
  44268=>"110110010",
  44269=>"111111111",
  44270=>"011111000",
  44271=>"000000000",
  44272=>"011011011",
  44273=>"110111111",
  44274=>"000000000",
  44275=>"000000000",
  44276=>"111111000",
  44277=>"100111111",
  44278=>"000000000",
  44279=>"000000000",
  44280=>"000000000",
  44281=>"000000110",
  44282=>"000000000",
  44283=>"001000000",
  44284=>"000000111",
  44285=>"000000011",
  44286=>"000000000",
  44287=>"100110110",
  44288=>"000000000",
  44289=>"111111111",
  44290=>"010111111",
  44291=>"000100111",
  44292=>"110000111",
  44293=>"010010111",
  44294=>"000000000",
  44295=>"110111111",
  44296=>"111111111",
  44297=>"000000000",
  44298=>"000100100",
  44299=>"110111100",
  44300=>"111011011",
  44301=>"000000000",
  44302=>"000000000",
  44303=>"001000111",
  44304=>"110000001",
  44305=>"111111111",
  44306=>"000000001",
  44307=>"000010000",
  44308=>"001000000",
  44309=>"100000001",
  44310=>"111111000",
  44311=>"000111110",
  44312=>"110110111",
  44313=>"000000000",
  44314=>"111001001",
  44315=>"111101000",
  44316=>"100111111",
  44317=>"000000001",
  44318=>"111111000",
  44319=>"000100000",
  44320=>"110000000",
  44321=>"000000000",
  44322=>"000001000",
  44323=>"110011011",
  44324=>"111001000",
  44325=>"000001000",
  44326=>"101000000",
  44327=>"000000000",
  44328=>"111111111",
  44329=>"111111111",
  44330=>"010110110",
  44331=>"111111111",
  44332=>"000110100",
  44333=>"011011111",
  44334=>"111111111",
  44335=>"000010111",
  44336=>"000101111",
  44337=>"000000000",
  44338=>"110010000",
  44339=>"111110111",
  44340=>"111111000",
  44341=>"010110110",
  44342=>"000010000",
  44343=>"000110000",
  44344=>"000000000",
  44345=>"000000000",
  44346=>"010000000",
  44347=>"111111001",
  44348=>"111111111",
  44349=>"000000000",
  44350=>"000000001",
  44351=>"111011000",
  44352=>"000110100",
  44353=>"110111111",
  44354=>"000000010",
  44355=>"000000000",
  44356=>"111000001",
  44357=>"110000100",
  44358=>"000000000",
  44359=>"000000111",
  44360=>"011000000",
  44361=>"111111111",
  44362=>"000010111",
  44363=>"001001001",
  44364=>"000000000",
  44365=>"111111111",
  44366=>"110000110",
  44367=>"111111111",
  44368=>"000000000",
  44369=>"000000100",
  44370=>"111111110",
  44371=>"111111100",
  44372=>"000001111",
  44373=>"000011011",
  44374=>"000000111",
  44375=>"111111111",
  44376=>"010111111",
  44377=>"111111111",
  44378=>"111111111",
  44379=>"110111111",
  44380=>"000000011",
  44381=>"110111110",
  44382=>"110110111",
  44383=>"100110111",
  44384=>"111111111",
  44385=>"000000000",
  44386=>"000100000",
  44387=>"111100100",
  44388=>"000011000",
  44389=>"111111011",
  44390=>"111110100",
  44391=>"000000000",
  44392=>"000000000",
  44393=>"011100110",
  44394=>"000000000",
  44395=>"000110011",
  44396=>"000000000",
  44397=>"000000000",
  44398=>"100000000",
  44399=>"000011011",
  44400=>"000001111",
  44401=>"001001000",
  44402=>"010111110",
  44403=>"011011011",
  44404=>"000000000",
  44405=>"000000111",
  44406=>"000000000",
  44407=>"100100000",
  44408=>"001000001",
  44409=>"100000000",
  44410=>"011010000",
  44411=>"111111100",
  44412=>"111001111",
  44413=>"111110110",
  44414=>"110000000",
  44415=>"111111111",
  44416=>"000000100",
  44417=>"000000001",
  44418=>"111111011",
  44419=>"111111111",
  44420=>"000000000",
  44421=>"000000000",
  44422=>"111111111",
  44423=>"110011000",
  44424=>"000000101",
  44425=>"111010011",
  44426=>"001000100",
  44427=>"000100111",
  44428=>"000110111",
  44429=>"011011011",
  44430=>"111111111",
  44431=>"000000000",
  44432=>"111111111",
  44433=>"110001001",
  44434=>"000000000",
  44435=>"110111111",
  44436=>"000000111",
  44437=>"000100100",
  44438=>"111111111",
  44439=>"001000000",
  44440=>"010111111",
  44441=>"111001000",
  44442=>"111111111",
  44443=>"111111011",
  44444=>"111110111",
  44445=>"111011011",
  44446=>"001000000",
  44447=>"111111111",
  44448=>"101101111",
  44449=>"000000001",
  44450=>"000000000",
  44451=>"010111000",
  44452=>"000000100",
  44453=>"000000000",
  44454=>"111001111",
  44455=>"000000000",
  44456=>"000010000",
  44457=>"111111111",
  44458=>"000000000",
  44459=>"111110000",
  44460=>"000111111",
  44461=>"000000001",
  44462=>"011000000",
  44463=>"111111100",
  44464=>"111000000",
  44465=>"000000000",
  44466=>"111111110",
  44467=>"111111111",
  44468=>"000000000",
  44469=>"010000000",
  44470=>"000111111",
  44471=>"011111111",
  44472=>"000000000",
  44473=>"010010000",
  44474=>"111000100",
  44475=>"111111111",
  44476=>"100000000",
  44477=>"111010110",
  44478=>"000000000",
  44479=>"010011011",
  44480=>"000001111",
  44481=>"000011011",
  44482=>"111011111",
  44483=>"001001000",
  44484=>"000000110",
  44485=>"011000001",
  44486=>"000000000",
  44487=>"001001001",
  44488=>"000000000",
  44489=>"000000011",
  44490=>"111011011",
  44491=>"111001111",
  44492=>"000000000",
  44493=>"111111001",
  44494=>"111111100",
  44495=>"001111001",
  44496=>"001000000",
  44497=>"111011011",
  44498=>"001110111",
  44499=>"001101111",
  44500=>"000000000",
  44501=>"111111011",
  44502=>"000000110",
  44503=>"001000000",
  44504=>"000001011",
  44505=>"000000000",
  44506=>"000000000",
  44507=>"111000101",
  44508=>"100001011",
  44509=>"110110111",
  44510=>"111110111",
  44511=>"000000000",
  44512=>"111111000",
  44513=>"111111111",
  44514=>"001001000",
  44515=>"110000000",
  44516=>"000110000",
  44517=>"000000000",
  44518=>"000000000",
  44519=>"111111100",
  44520=>"001000001",
  44521=>"001111111",
  44522=>"111111101",
  44523=>"111111111",
  44524=>"111110111",
  44525=>"110110000",
  44526=>"111111111",
  44527=>"111111111",
  44528=>"000000000",
  44529=>"000000000",
  44530=>"111110111",
  44531=>"111111111",
  44532=>"000000000",
  44533=>"000111111",
  44534=>"000101000",
  44535=>"000000000",
  44536=>"000000000",
  44537=>"010110010",
  44538=>"111111111",
  44539=>"000000000",
  44540=>"000000111",
  44541=>"101100100",
  44542=>"000000000",
  44543=>"000000000",
  44544=>"111111111",
  44545=>"000101111",
  44546=>"111000000",
  44547=>"101000000",
  44548=>"111011000",
  44549=>"000000011",
  44550=>"000000000",
  44551=>"000000000",
  44552=>"000000000",
  44553=>"111011000",
  44554=>"100111011",
  44555=>"000110110",
  44556=>"111111110",
  44557=>"000000000",
  44558=>"010011000",
  44559=>"000000001",
  44560=>"111111111",
  44561=>"111111011",
  44562=>"000000001",
  44563=>"001000001",
  44564=>"111010000",
  44565=>"000000000",
  44566=>"010110000",
  44567=>"111111000",
  44568=>"001001111",
  44569=>"110000011",
  44570=>"010100000",
  44571=>"000000000",
  44572=>"000000000",
  44573=>"000000000",
  44574=>"100100111",
  44575=>"110110111",
  44576=>"000000000",
  44577=>"000001011",
  44578=>"000000110",
  44579=>"000000000",
  44580=>"111111111",
  44581=>"100111111",
  44582=>"111011011",
  44583=>"110110110",
  44584=>"000000011",
  44585=>"000000000",
  44586=>"111111111",
  44587=>"000011111",
  44588=>"111000000",
  44589=>"111000000",
  44590=>"111111111",
  44591=>"101100000",
  44592=>"000000100",
  44593=>"000000000",
  44594=>"000000000",
  44595=>"001000100",
  44596=>"000101111",
  44597=>"111111111",
  44598=>"001101111",
  44599=>"000000000",
  44600=>"110000000",
  44601=>"000000111",
  44602=>"011000000",
  44603=>"000000000",
  44604=>"001000001",
  44605=>"000000000",
  44606=>"110110110",
  44607=>"000000000",
  44608=>"000000000",
  44609=>"000101101",
  44610=>"000101100",
  44611=>"111111111",
  44612=>"110000000",
  44613=>"000000000",
  44614=>"101111111",
  44615=>"000000000",
  44616=>"001011010",
  44617=>"001000000",
  44618=>"000000000",
  44619=>"111010000",
  44620=>"000000000",
  44621=>"111111111",
  44622=>"110111010",
  44623=>"000000000",
  44624=>"000000000",
  44625=>"010110110",
  44626=>"111111111",
  44627=>"010011011",
  44628=>"111101111",
  44629=>"110110110",
  44630=>"111011000",
  44631=>"111111111",
  44632=>"000110110",
  44633=>"000000000",
  44634=>"111111111",
  44635=>"111111111",
  44636=>"010111111",
  44637=>"111111111",
  44638=>"000000000",
  44639=>"011011011",
  44640=>"100000000",
  44641=>"111111111",
  44642=>"111000000",
  44643=>"000000000",
  44644=>"000000000",
  44645=>"000100000",
  44646=>"000000000",
  44647=>"110110010",
  44648=>"111111111",
  44649=>"011111111",
  44650=>"011000100",
  44651=>"001111111",
  44652=>"111111111",
  44653=>"111011001",
  44654=>"000000111",
  44655=>"101111100",
  44656=>"000000000",
  44657=>"000000000",
  44658=>"111111111",
  44659=>"100110010",
  44660=>"001000000",
  44661=>"111110110",
  44662=>"000000000",
  44663=>"101000000",
  44664=>"000011000",
  44665=>"000000100",
  44666=>"000000000",
  44667=>"000000000",
  44668=>"011010010",
  44669=>"111111111",
  44670=>"111111000",
  44671=>"000000001",
  44672=>"000000000",
  44673=>"000000000",
  44674=>"111111111",
  44675=>"110110111",
  44676=>"011011110",
  44677=>"010000111",
  44678=>"000000000",
  44679=>"011010000",
  44680=>"000011111",
  44681=>"100000000",
  44682=>"111111111",
  44683=>"111111111",
  44684=>"000000000",
  44685=>"100100101",
  44686=>"000000110",
  44687=>"000000000",
  44688=>"111111111",
  44689=>"101111111",
  44690=>"000000000",
  44691=>"000100110",
  44692=>"000000000",
  44693=>"010000111",
  44694=>"111111111",
  44695=>"111111101",
  44696=>"111111111",
  44697=>"000000000",
  44698=>"111111000",
  44699=>"000000101",
  44700=>"101111011",
  44701=>"000000000",
  44702=>"000000000",
  44703=>"111111111",
  44704=>"000000000",
  44705=>"111110010",
  44706=>"110111111",
  44707=>"000111000",
  44708=>"111111111",
  44709=>"000000000",
  44710=>"000111111",
  44711=>"111111111",
  44712=>"001000000",
  44713=>"000000000",
  44714=>"000000000",
  44715=>"011010111",
  44716=>"000110111",
  44717=>"101110001",
  44718=>"101111111",
  44719=>"111111111",
  44720=>"011111111",
  44721=>"011011101",
  44722=>"111111111",
  44723=>"111111111",
  44724=>"100101001",
  44725=>"000000001",
  44726=>"111100111",
  44727=>"000000000",
  44728=>"000010110",
  44729=>"001011011",
  44730=>"111101000",
  44731=>"111111011",
  44732=>"000000000",
  44733=>"111111111",
  44734=>"111111111",
  44735=>"000110011",
  44736=>"111111111",
  44737=>"111001001",
  44738=>"100100000",
  44739=>"000100100",
  44740=>"000000000",
  44741=>"000000000",
  44742=>"000001000",
  44743=>"101111111",
  44744=>"101111111",
  44745=>"000000111",
  44746=>"000000000",
  44747=>"111111110",
  44748=>"111110111",
  44749=>"000000000",
  44750=>"000111100",
  44751=>"111111111",
  44752=>"000000111",
  44753=>"000000000",
  44754=>"111111111",
  44755=>"111101111",
  44756=>"111100000",
  44757=>"000001001",
  44758=>"000000000",
  44759=>"111111100",
  44760=>"110111111",
  44761=>"000000000",
  44762=>"111111000",
  44763=>"111111110",
  44764=>"111011111",
  44765=>"001000000",
  44766=>"000000000",
  44767=>"000001111",
  44768=>"011011001",
  44769=>"000000000",
  44770=>"000001100",
  44771=>"111111001",
  44772=>"011011111",
  44773=>"110111011",
  44774=>"111111000",
  44775=>"111111111",
  44776=>"111001000",
  44777=>"000000001",
  44778=>"111111100",
  44779=>"001011111",
  44780=>"100000000",
  44781=>"111000000",
  44782=>"000000000",
  44783=>"000000000",
  44784=>"100101111",
  44785=>"111100000",
  44786=>"000000011",
  44787=>"111111010",
  44788=>"100000111",
  44789=>"010010100",
  44790=>"000110111",
  44791=>"111000000",
  44792=>"000000000",
  44793=>"001101111",
  44794=>"010000000",
  44795=>"000100111",
  44796=>"111111111",
  44797=>"000000000",
  44798=>"000000000",
  44799=>"100000100",
  44800=>"011000010",
  44801=>"011011111",
  44802=>"111111111",
  44803=>"000000011",
  44804=>"011000000",
  44805=>"010010010",
  44806=>"111111110",
  44807=>"111111111",
  44808=>"111111111",
  44809=>"001000001",
  44810=>"111011000",
  44811=>"000000110",
  44812=>"110010111",
  44813=>"111001000",
  44814=>"111111100",
  44815=>"101100111",
  44816=>"111111111",
  44817=>"011101111",
  44818=>"001000001",
  44819=>"100000000",
  44820=>"100000000",
  44821=>"111111111",
  44822=>"111111101",
  44823=>"000111111",
  44824=>"111111111",
  44825=>"111100111",
  44826=>"111001011",
  44827=>"000000000",
  44828=>"111100000",
  44829=>"101000111",
  44830=>"111100000",
  44831=>"000000000",
  44832=>"100000000",
  44833=>"110010000",
  44834=>"011011111",
  44835=>"111111000",
  44836=>"000000000",
  44837=>"000000000",
  44838=>"000010111",
  44839=>"000000100",
  44840=>"111111111",
  44841=>"000000000",
  44842=>"000000110",
  44843=>"111001000",
  44844=>"111001111",
  44845=>"111111001",
  44846=>"111111111",
  44847=>"000011011",
  44848=>"000110110",
  44849=>"111111111",
  44850=>"000000110",
  44851=>"110111111",
  44852=>"111100101",
  44853=>"111111111",
  44854=>"111111111",
  44855=>"001110110",
  44856=>"111111010",
  44857=>"000000000",
  44858=>"110000000",
  44859=>"111101001",
  44860=>"000001000",
  44861=>"100110110",
  44862=>"000100000",
  44863=>"000001111",
  44864=>"000000110",
  44865=>"110110111",
  44866=>"000000111",
  44867=>"000000000",
  44868=>"100000000",
  44869=>"100000001",
  44870=>"000001111",
  44871=>"000000111",
  44872=>"000110101",
  44873=>"111000001",
  44874=>"011111110",
  44875=>"010010000",
  44876=>"111111111",
  44877=>"000100111",
  44878=>"001100100",
  44879=>"100110100",
  44880=>"000010110",
  44881=>"000000010",
  44882=>"001000000",
  44883=>"111111111",
  44884=>"000000000",
  44885=>"000000000",
  44886=>"000001111",
  44887=>"100111111",
  44888=>"000000000",
  44889=>"111111111",
  44890=>"000000000",
  44891=>"111111111",
  44892=>"000000011",
  44893=>"000110000",
  44894=>"000111111",
  44895=>"100111101",
  44896=>"001111111",
  44897=>"111111111",
  44898=>"110111110",
  44899=>"000000101",
  44900=>"000001111",
  44901=>"001110111",
  44902=>"001000001",
  44903=>"010010000",
  44904=>"100110000",
  44905=>"111111111",
  44906=>"000000000",
  44907=>"000001000",
  44908=>"000000000",
  44909=>"000001101",
  44910=>"000000001",
  44911=>"000111111",
  44912=>"011001101",
  44913=>"000000000",
  44914=>"000000001",
  44915=>"000000100",
  44916=>"001111111",
  44917=>"001000000",
  44918=>"000100110",
  44919=>"000000111",
  44920=>"100000000",
  44921=>"111000000",
  44922=>"000000110",
  44923=>"111111000",
  44924=>"111101111",
  44925=>"010000000",
  44926=>"001001000",
  44927=>"100001000",
  44928=>"010001001",
  44929=>"100010100",
  44930=>"100100100",
  44931=>"000010011",
  44932=>"000000111",
  44933=>"000000000",
  44934=>"111111000",
  44935=>"101111111",
  44936=>"001111001",
  44937=>"110100100",
  44938=>"000000000",
  44939=>"111111101",
  44940=>"001000000",
  44941=>"111111111",
  44942=>"010010000",
  44943=>"101000000",
  44944=>"011000000",
  44945=>"111110111",
  44946=>"111111111",
  44947=>"111110110",
  44948=>"001001001",
  44949=>"011001000",
  44950=>"110111111",
  44951=>"001011001",
  44952=>"000110111",
  44953=>"111111111",
  44954=>"111010000",
  44955=>"001000001",
  44956=>"111111100",
  44957=>"111010000",
  44958=>"111111111",
  44959=>"000110000",
  44960=>"111100100",
  44961=>"001001000",
  44962=>"000000000",
  44963=>"111110111",
  44964=>"011000000",
  44965=>"111000000",
  44966=>"111111111",
  44967=>"111110110",
  44968=>"111111011",
  44969=>"001011001",
  44970=>"111111111",
  44971=>"110110111",
  44972=>"001100000",
  44973=>"000001000",
  44974=>"101110100",
  44975=>"000100111",
  44976=>"111111111",
  44977=>"111111111",
  44978=>"100010000",
  44979=>"111111101",
  44980=>"000000000",
  44981=>"101000101",
  44982=>"111110110",
  44983=>"111001101",
  44984=>"010111111",
  44985=>"011000110",
  44986=>"111111010",
  44987=>"110111111",
  44988=>"110100110",
  44989=>"111111111",
  44990=>"000000000",
  44991=>"111110100",
  44992=>"000000000",
  44993=>"000000000",
  44994=>"111111000",
  44995=>"111111111",
  44996=>"111000000",
  44997=>"110100000",
  44998=>"010000000",
  44999=>"111111001",
  45000=>"011001000",
  45001=>"000000000",
  45002=>"111011011",
  45003=>"111111111",
  45004=>"000000000",
  45005=>"111110000",
  45006=>"101000111",
  45007=>"000101111",
  45008=>"100111110",
  45009=>"000110111",
  45010=>"001111111",
  45011=>"000000111",
  45012=>"001000000",
  45013=>"111111110",
  45014=>"000000000",
  45015=>"001001000",
  45016=>"000111111",
  45017=>"000000000",
  45018=>"000100000",
  45019=>"110100100",
  45020=>"000111011",
  45021=>"111010110",
  45022=>"110101111",
  45023=>"000011001",
  45024=>"111111011",
  45025=>"000000011",
  45026=>"000000111",
  45027=>"111011011",
  45028=>"110110111",
  45029=>"001000000",
  45030=>"101011011",
  45031=>"111111000",
  45032=>"000010111",
  45033=>"111111111",
  45034=>"000000111",
  45035=>"111011010",
  45036=>"111111110",
  45037=>"100110100",
  45038=>"000111110",
  45039=>"111001001",
  45040=>"000100111",
  45041=>"111111111",
  45042=>"001000010",
  45043=>"111111111",
  45044=>"000000111",
  45045=>"111000111",
  45046=>"000000001",
  45047=>"000000000",
  45048=>"100111111",
  45049=>"000000000",
  45050=>"111001111",
  45051=>"111110110",
  45052=>"000000000",
  45053=>"000000000",
  45054=>"101111111",
  45055=>"000000000",
  45056=>"001011010",
  45057=>"000111000",
  45058=>"111111000",
  45059=>"011010000",
  45060=>"111111111",
  45061=>"111111001",
  45062=>"000000100",
  45063=>"000000000",
  45064=>"111000000",
  45065=>"111111000",
  45066=>"110110000",
  45067=>"000000001",
  45068=>"101110111",
  45069=>"111010010",
  45070=>"000000000",
  45071=>"000000000",
  45072=>"110100100",
  45073=>"111000111",
  45074=>"111111110",
  45075=>"111101000",
  45076=>"000000000",
  45077=>"111110100",
  45078=>"000000000",
  45079=>"000000101",
  45080=>"111011000",
  45081=>"111111011",
  45082=>"111111011",
  45083=>"011001000",
  45084=>"111111100",
  45085=>"111111101",
  45086=>"110111110",
  45087=>"000000111",
  45088=>"000000010",
  45089=>"110111111",
  45090=>"000111111",
  45091=>"111100100",
  45092=>"000101000",
  45093=>"111111111",
  45094=>"111111110",
  45095=>"000110000",
  45096=>"000111111",
  45097=>"111111000",
  45098=>"000000000",
  45099=>"000000000",
  45100=>"001111111",
  45101=>"101000111",
  45102=>"000000111",
  45103=>"001001111",
  45104=>"000000111",
  45105=>"110100111",
  45106=>"100111111",
  45107=>"111111111",
  45108=>"000000011",
  45109=>"101001001",
  45110=>"111011011",
  45111=>"011011111",
  45112=>"000000000",
  45113=>"000000011",
  45114=>"111000000",
  45115=>"101001011",
  45116=>"111111111",
  45117=>"100000000",
  45118=>"110010000",
  45119=>"111010000",
  45120=>"001111111",
  45121=>"011000000",
  45122=>"010111011",
  45123=>"001001111",
  45124=>"000010110",
  45125=>"011011001",
  45126=>"111000000",
  45127=>"001000000",
  45128=>"111111100",
  45129=>"000000100",
  45130=>"001011001",
  45131=>"000011111",
  45132=>"000011111",
  45133=>"000000000",
  45134=>"000000000",
  45135=>"111111111",
  45136=>"000000000",
  45137=>"000000001",
  45138=>"011011000",
  45139=>"101110111",
  45140=>"111011011",
  45141=>"111111111",
  45142=>"111101000",
  45143=>"111111011",
  45144=>"000000000",
  45145=>"001000000",
  45146=>"011000111",
  45147=>"000000000",
  45148=>"000000101",
  45149=>"110111111",
  45150=>"000000000",
  45151=>"011001111",
  45152=>"100000000",
  45153=>"000001001",
  45154=>"000000000",
  45155=>"000000000",
  45156=>"100110011",
  45157=>"000001111",
  45158=>"110000000",
  45159=>"111111000",
  45160=>"101111111",
  45161=>"111101000",
  45162=>"000001000",
  45163=>"000000000",
  45164=>"001011101",
  45165=>"111101000",
  45166=>"000110110",
  45167=>"111111010",
  45168=>"000001101",
  45169=>"000000111",
  45170=>"000000001",
  45171=>"000000000",
  45172=>"000001111",
  45173=>"000110101",
  45174=>"100111111",
  45175=>"000000000",
  45176=>"000000111",
  45177=>"000010001",
  45178=>"000011011",
  45179=>"000100111",
  45180=>"111111110",
  45181=>"111111000",
  45182=>"000000001",
  45183=>"000000100",
  45184=>"111111000",
  45185=>"011011001",
  45186=>"111111111",
  45187=>"000011011",
  45188=>"000000000",
  45189=>"101000000",
  45190=>"001010000",
  45191=>"111000000",
  45192=>"111111111",
  45193=>"111111111",
  45194=>"000000010",
  45195=>"110110010",
  45196=>"010000000",
  45197=>"000000000",
  45198=>"000000001",
  45199=>"000000000",
  45200=>"100000000",
  45201=>"000000111",
  45202=>"000100111",
  45203=>"110110111",
  45204=>"010011011",
  45205=>"010000000",
  45206=>"111100101",
  45207=>"001000000",
  45208=>"111110000",
  45209=>"111101100",
  45210=>"100110000",
  45211=>"110111111",
  45212=>"111011011",
  45213=>"000000110",
  45214=>"111001011",
  45215=>"111111001",
  45216=>"111111000",
  45217=>"100100000",
  45218=>"000011111",
  45219=>"000000000",
  45220=>"101100100",
  45221=>"000000000",
  45222=>"111111000",
  45223=>"011000101",
  45224=>"111111000",
  45225=>"111111001",
  45226=>"111111010",
  45227=>"100111111",
  45228=>"110001101",
  45229=>"000000111",
  45230=>"111111111",
  45231=>"000000011",
  45232=>"000000111",
  45233=>"001001000",
  45234=>"000111111",
  45235=>"111011001",
  45236=>"000000000",
  45237=>"000010110",
  45238=>"000000000",
  45239=>"000000000",
  45240=>"110100111",
  45241=>"111111110",
  45242=>"100110110",
  45243=>"010011111",
  45244=>"111111111",
  45245=>"000000000",
  45246=>"111101101",
  45247=>"011001111",
  45248=>"010010000",
  45249=>"010111100",
  45250=>"000001100",
  45251=>"111111000",
  45252=>"100000010",
  45253=>"001001011",
  45254=>"000000000",
  45255=>"110111010",
  45256=>"110110111",
  45257=>"110111111",
  45258=>"001001111",
  45259=>"000000100",
  45260=>"000001111",
  45261=>"111111000",
  45262=>"000000110",
  45263=>"111111110",
  45264=>"000000000",
  45265=>"111111011",
  45266=>"001000000",
  45267=>"111111111",
  45268=>"100100111",
  45269=>"111011001",
  45270=>"111111000",
  45271=>"000110110",
  45272=>"011011001",
  45273=>"111111110",
  45274=>"000000000",
  45275=>"011111011",
  45276=>"111111011",
  45277=>"101000111",
  45278=>"000000010",
  45279=>"000000000",
  45280=>"111111001",
  45281=>"111111000",
  45282=>"001001011",
  45283=>"111100000",
  45284=>"111000011",
  45285=>"000000000",
  45286=>"111111000",
  45287=>"111111000",
  45288=>"011000000",
  45289=>"001001111",
  45290=>"000000110",
  45291=>"000000001",
  45292=>"000000111",
  45293=>"111111111",
  45294=>"010010000",
  45295=>"111111111",
  45296=>"000000000",
  45297=>"000101001",
  45298=>"000100111",
  45299=>"011111110",
  45300=>"011000000",
  45301=>"111000111",
  45302=>"111111101",
  45303=>"000000000",
  45304=>"000111111",
  45305=>"111001001",
  45306=>"001001001",
  45307=>"111111111",
  45308=>"001000010",
  45309=>"111111100",
  45310=>"000001000",
  45311=>"111111000",
  45312=>"010000000",
  45313=>"111111000",
  45314=>"111111000",
  45315=>"011000000",
  45316=>"000101101",
  45317=>"111111011",
  45318=>"000010000",
  45319=>"111011100",
  45320=>"110111010",
  45321=>"110010000",
  45322=>"011010000",
  45323=>"000000100",
  45324=>"010111111",
  45325=>"111111111",
  45326=>"110111011",
  45327=>"111010000",
  45328=>"010000111",
  45329=>"111000000",
  45330=>"011011101",
  45331=>"111111111",
  45332=>"000000000",
  45333=>"111111111",
  45334=>"111110111",
  45335=>"000000111",
  45336=>"001001001",
  45337=>"001000000",
  45338=>"001000111",
  45339=>"111000000",
  45340=>"111111001",
  45341=>"111111111",
  45342=>"111111111",
  45343=>"110111000",
  45344=>"100100000",
  45345=>"110111010",
  45346=>"011111111",
  45347=>"100000110",
  45348=>"100100100",
  45349=>"000000001",
  45350=>"111101111",
  45351=>"000000101",
  45352=>"110110000",
  45353=>"000000100",
  45354=>"101011011",
  45355=>"000100000",
  45356=>"111111011",
  45357=>"111011011",
  45358=>"000000000",
  45359=>"000111000",
  45360=>"111111111",
  45361=>"001001000",
  45362=>"011111111",
  45363=>"000110110",
  45364=>"000000000",
  45365=>"000111101",
  45366=>"000000001",
  45367=>"111111110",
  45368=>"111111111",
  45369=>"101000000",
  45370=>"000000000",
  45371=>"100111111",
  45372=>"000100100",
  45373=>"111111111",
  45374=>"111111101",
  45375=>"111111011",
  45376=>"101101100",
  45377=>"001001000",
  45378=>"011111000",
  45379=>"000000111",
  45380=>"011011011",
  45381=>"000111111",
  45382=>"000000000",
  45383=>"001000000",
  45384=>"000000111",
  45385=>"111001010",
  45386=>"000000011",
  45387=>"011001100",
  45388=>"010110100",
  45389=>"001000100",
  45390=>"000000000",
  45391=>"001101100",
  45392=>"011011111",
  45393=>"111111111",
  45394=>"010000111",
  45395=>"000000011",
  45396=>"000111011",
  45397=>"111011111",
  45398=>"000000000",
  45399=>"111111111",
  45400=>"000110000",
  45401=>"000000000",
  45402=>"001001111",
  45403=>"110010010",
  45404=>"111100100",
  45405=>"000000000",
  45406=>"011011001",
  45407=>"000101001",
  45408=>"000000000",
  45409=>"000000001",
  45410=>"011001111",
  45411=>"111111111",
  45412=>"000100000",
  45413=>"000000101",
  45414=>"111111000",
  45415=>"110000000",
  45416=>"000001001",
  45417=>"001011001",
  45418=>"000101001",
  45419=>"111111111",
  45420=>"000101111",
  45421=>"100100110",
  45422=>"111111111",
  45423=>"000000000",
  45424=>"111111111",
  45425=>"000000100",
  45426=>"001011000",
  45427=>"111111111",
  45428=>"010111000",
  45429=>"010010010",
  45430=>"010110111",
  45431=>"111111111",
  45432=>"110111000",
  45433=>"111001000",
  45434=>"010000011",
  45435=>"110110000",
  45436=>"111000100",
  45437=>"111011000",
  45438=>"110010000",
  45439=>"100000111",
  45440=>"000000111",
  45441=>"010011011",
  45442=>"100100110",
  45443=>"000000000",
  45444=>"000111111",
  45445=>"001000110",
  45446=>"000001101",
  45447=>"111111111",
  45448=>"000000000",
  45449=>"000000111",
  45450=>"011011000",
  45451=>"111111000",
  45452=>"101110111",
  45453=>"111111111",
  45454=>"000110111",
  45455=>"111111011",
  45456=>"011000010",
  45457=>"000000010",
  45458=>"101001111",
  45459=>"100100111",
  45460=>"000000100",
  45461=>"111011011",
  45462=>"111111101",
  45463=>"001001110",
  45464=>"111111111",
  45465=>"000000111",
  45466=>"111110000",
  45467=>"011111111",
  45468=>"000000110",
  45469=>"111111111",
  45470=>"111000111",
  45471=>"000000001",
  45472=>"111000000",
  45473=>"111111011",
  45474=>"000011111",
  45475=>"111111111",
  45476=>"111001110",
  45477=>"000100111",
  45478=>"000110110",
  45479=>"111000000",
  45480=>"000000000",
  45481=>"111011111",
  45482=>"110111111",
  45483=>"000000111",
  45484=>"000000000",
  45485=>"110111010",
  45486=>"000111111",
  45487=>"000000000",
  45488=>"100100000",
  45489=>"000000001",
  45490=>"111111100",
  45491=>"000000001",
  45492=>"011011011",
  45493=>"000000001",
  45494=>"110111000",
  45495=>"001000000",
  45496=>"111111000",
  45497=>"000100111",
  45498=>"011000000",
  45499=>"111111100",
  45500=>"001111111",
  45501=>"111010000",
  45502=>"101101101",
  45503=>"011001011",
  45504=>"111111011",
  45505=>"000110010",
  45506=>"000000111",
  45507=>"000000111",
  45508=>"100111111",
  45509=>"110111110",
  45510=>"111001011",
  45511=>"010110000",
  45512=>"111010110",
  45513=>"000000000",
  45514=>"111000111",
  45515=>"001000000",
  45516=>"011000000",
  45517=>"111000111",
  45518=>"100000011",
  45519=>"111000101",
  45520=>"111111111",
  45521=>"000000000",
  45522=>"100100001",
  45523=>"011001001",
  45524=>"111111111",
  45525=>"111101001",
  45526=>"001011000",
  45527=>"000000000",
  45528=>"000001000",
  45529=>"000000001",
  45530=>"000110100",
  45531=>"000000000",
  45532=>"001011011",
  45533=>"011000000",
  45534=>"100000011",
  45535=>"000001111",
  45536=>"111111000",
  45537=>"000000001",
  45538=>"000001111",
  45539=>"001001100",
  45540=>"000100111",
  45541=>"000001111",
  45542=>"000101111",
  45543=>"000010011",
  45544=>"110110110",
  45545=>"000110110",
  45546=>"111111101",
  45547=>"100100110",
  45548=>"101111111",
  45549=>"000001011",
  45550=>"101000000",
  45551=>"100000011",
  45552=>"000100111",
  45553=>"000000011",
  45554=>"111111010",
  45555=>"000000111",
  45556=>"000010000",
  45557=>"111011001",
  45558=>"000000001",
  45559=>"000001110",
  45560=>"111111111",
  45561=>"011001111",
  45562=>"000000101",
  45563=>"000000111",
  45564=>"111110000",
  45565=>"110111011",
  45566=>"110000000",
  45567=>"000000000",
  45568=>"110110111",
  45569=>"110110111",
  45570=>"101000000",
  45571=>"000000000",
  45572=>"111111111",
  45573=>"001000100",
  45574=>"000000000",
  45575=>"000000000",
  45576=>"111111101",
  45577=>"111000000",
  45578=>"000111111",
  45579=>"000111111",
  45580=>"000000001",
  45581=>"000000001",
  45582=>"111000001",
  45583=>"000000001",
  45584=>"111101001",
  45585=>"110110110",
  45586=>"100000000",
  45587=>"011001111",
  45588=>"111110111",
  45589=>"100000001",
  45590=>"000000001",
  45591=>"001011011",
  45592=>"000110111",
  45593=>"000000001",
  45594=>"111000101",
  45595=>"010001000",
  45596=>"111111111",
  45597=>"100110110",
  45598=>"000000100",
  45599=>"100110001",
  45600=>"111100001",
  45601=>"111111111",
  45602=>"111111011",
  45603=>"000100101",
  45604=>"000000101",
  45605=>"110100100",
  45606=>"111100100",
  45607=>"110111111",
  45608=>"110111000",
  45609=>"000000000",
  45610=>"000000000",
  45611=>"110100110",
  45612=>"111000000",
  45613=>"111111111",
  45614=>"010010010",
  45615=>"111001000",
  45616=>"000101111",
  45617=>"001001000",
  45618=>"010111111",
  45619=>"000000001",
  45620=>"010111111",
  45621=>"000000000",
  45622=>"000000000",
  45623=>"100100111",
  45624=>"000000010",
  45625=>"000000000",
  45626=>"000000000",
  45627=>"000111111",
  45628=>"000010111",
  45629=>"111100000",
  45630=>"001000100",
  45631=>"111000111",
  45632=>"111100000",
  45633=>"000000001",
  45634=>"110111011",
  45635=>"110010010",
  45636=>"111111110",
  45637=>"111001001",
  45638=>"111001001",
  45639=>"000000000",
  45640=>"001001001",
  45641=>"011000000",
  45642=>"110000100",
  45643=>"000000000",
  45644=>"111011000",
  45645=>"111111001",
  45646=>"000011011",
  45647=>"000001000",
  45648=>"000000000",
  45649=>"000000111",
  45650=>"000100111",
  45651=>"011011000",
  45652=>"111001001",
  45653=>"000100100",
  45654=>"001000000",
  45655=>"000000000",
  45656=>"000111111",
  45657=>"000000000",
  45658=>"111111000",
  45659=>"011011000",
  45660=>"100000000",
  45661=>"000000000",
  45662=>"000011010",
  45663=>"000000011",
  45664=>"000100111",
  45665=>"001000110",
  45666=>"111111110",
  45667=>"111001000",
  45668=>"111111111",
  45669=>"000000000",
  45670=>"110010111",
  45671=>"000010110",
  45672=>"110111110",
  45673=>"111111000",
  45674=>"011011100",
  45675=>"010000000",
  45676=>"000010000",
  45677=>"101101101",
  45678=>"011010000",
  45679=>"111111000",
  45680=>"110111111",
  45681=>"011001101",
  45682=>"011111000",
  45683=>"101001111",
  45684=>"100000001",
  45685=>"000000101",
  45686=>"000100111",
  45687=>"011000000",
  45688=>"001001001",
  45689=>"100100111",
  45690=>"000000101",
  45691=>"001001111",
  45692=>"100110100",
  45693=>"110111110",
  45694=>"000001000",
  45695=>"111111111",
  45696=>"000000000",
  45697=>"111111000",
  45698=>"111111110",
  45699=>"111101111",
  45700=>"111111111",
  45701=>"000000000",
  45702=>"000011111",
  45703=>"000111111",
  45704=>"000000111",
  45705=>"000000000",
  45706=>"010110000",
  45707=>"000001000",
  45708=>"010011101",
  45709=>"011000000",
  45710=>"000000111",
  45711=>"000000110",
  45712=>"011111011",
  45713=>"000000011",
  45714=>"000000000",
  45715=>"000000111",
  45716=>"000000100",
  45717=>"000000110",
  45718=>"000111111",
  45719=>"001000000",
  45720=>"000000111",
  45721=>"111011000",
  45722=>"111111111",
  45723=>"111111111",
  45724=>"001000000",
  45725=>"100000010",
  45726=>"000000000",
  45727=>"111011111",
  45728=>"111100110",
  45729=>"100100110",
  45730=>"110111111",
  45731=>"000100111",
  45732=>"000000111",
  45733=>"001000000",
  45734=>"000000001",
  45735=>"000000000",
  45736=>"111000000",
  45737=>"000000001",
  45738=>"100000101",
  45739=>"000000000",
  45740=>"011001000",
  45741=>"000000001",
  45742=>"000011011",
  45743=>"000000110",
  45744=>"111110111",
  45745=>"110100100",
  45746=>"110111110",
  45747=>"000000101",
  45748=>"110000001",
  45749=>"000000101",
  45750=>"101111010",
  45751=>"000000100",
  45752=>"111110111",
  45753=>"000000000",
  45754=>"000000000",
  45755=>"111111111",
  45756=>"001110111",
  45757=>"111111110",
  45758=>"111000110",
  45759=>"111111111",
  45760=>"100100000",
  45761=>"000010111",
  45762=>"110111111",
  45763=>"000000000",
  45764=>"000000010",
  45765=>"101001000",
  45766=>"000000000",
  45767=>"000111010",
  45768=>"000100100",
  45769=>"111111111",
  45770=>"000001000",
  45771=>"010011011",
  45772=>"000000111",
  45773=>"010000000",
  45774=>"011011111",
  45775=>"001001000",
  45776=>"001111111",
  45777=>"000100100",
  45778=>"011011011",
  45779=>"111111111",
  45780=>"000000000",
  45781=>"001011111",
  45782=>"101101101",
  45783=>"001010000",
  45784=>"111110110",
  45785=>"111011011",
  45786=>"111000001",
  45787=>"111100000",
  45788=>"000000000",
  45789=>"000110111",
  45790=>"000111111",
  45791=>"000000000",
  45792=>"000000111",
  45793=>"000000000",
  45794=>"111111111",
  45795=>"000000101",
  45796=>"000000001",
  45797=>"111110110",
  45798=>"000000000",
  45799=>"000100111",
  45800=>"000000000",
  45801=>"111001111",
  45802=>"111111111",
  45803=>"111111111",
  45804=>"110010111",
  45805=>"000000000",
  45806=>"110111111",
  45807=>"110111111",
  45808=>"000000000",
  45809=>"000000000",
  45810=>"111111111",
  45811=>"111011000",
  45812=>"110111110",
  45813=>"000000110",
  45814=>"111110011",
  45815=>"001000000",
  45816=>"000000000",
  45817=>"101000000",
  45818=>"001000111",
  45819=>"000000111",
  45820=>"011010000",
  45821=>"000111111",
  45822=>"000110000",
  45823=>"111111110",
  45824=>"000000000",
  45825=>"010111111",
  45826=>"011111111",
  45827=>"000100111",
  45828=>"000000101",
  45829=>"000000011",
  45830=>"110100110",
  45831=>"000000000",
  45832=>"000000000",
  45833=>"110111111",
  45834=>"111111111",
  45835=>"000000001",
  45836=>"100100100",
  45837=>"010000000",
  45838=>"000111001",
  45839=>"000100000",
  45840=>"000000011",
  45841=>"000000011",
  45842=>"001111111",
  45843=>"111111011",
  45844=>"000000000",
  45845=>"000001111",
  45846=>"011111011",
  45847=>"111111111",
  45848=>"110111010",
  45849=>"000011111",
  45850=>"101000111",
  45851=>"000000001",
  45852=>"110110100",
  45853=>"010000000",
  45854=>"000000000",
  45855=>"111111111",
  45856=>"000100111",
  45857=>"111001000",
  45858=>"000000000",
  45859=>"111011000",
  45860=>"111100000",
  45861=>"111111000",
  45862=>"000000000",
  45863=>"001001000",
  45864=>"000011111",
  45865=>"000000000",
  45866=>"001000110",
  45867=>"111111111",
  45868=>"011001000",
  45869=>"000111111",
  45870=>"110011000",
  45871=>"000011010",
  45872=>"001000000",
  45873=>"100000001",
  45874=>"111001101",
  45875=>"000011011",
  45876=>"000000000",
  45877=>"111100000",
  45878=>"000000000",
  45879=>"000000000",
  45880=>"111001000",
  45881=>"111100000",
  45882=>"110111111",
  45883=>"111111100",
  45884=>"101000000",
  45885=>"110111111",
  45886=>"000010010",
  45887=>"000101001",
  45888=>"000000111",
  45889=>"110010101",
  45890=>"001000000",
  45891=>"110000000",
  45892=>"000000111",
  45893=>"001000001",
  45894=>"101111111",
  45895=>"000000000",
  45896=>"001000000",
  45897=>"110000000",
  45898=>"000110110",
  45899=>"110000110",
  45900=>"000110000",
  45901=>"000010111",
  45902=>"111111001",
  45903=>"011000000",
  45904=>"011010110",
  45905=>"111111011",
  45906=>"100110000",
  45907=>"111111111",
  45908=>"001000000",
  45909=>"011011011",
  45910=>"000000000",
  45911=>"010011111",
  45912=>"001001000",
  45913=>"101111111",
  45914=>"000010000",
  45915=>"110000000",
  45916=>"111011101",
  45917=>"000110111",
  45918=>"011111111",
  45919=>"100010111",
  45920=>"111000000",
  45921=>"000000111",
  45922=>"100100000",
  45923=>"000000101",
  45924=>"110111110",
  45925=>"000001001",
  45926=>"000000000",
  45927=>"001101111",
  45928=>"110100100",
  45929=>"101101111",
  45930=>"001001000",
  45931=>"111111111",
  45932=>"001011001",
  45933=>"000010000",
  45934=>"000000111",
  45935=>"000000000",
  45936=>"111111110",
  45937=>"111111110",
  45938=>"000000000",
  45939=>"011011000",
  45940=>"111111111",
  45941=>"100111111",
  45942=>"111001100",
  45943=>"111011110",
  45944=>"000000000",
  45945=>"000000000",
  45946=>"000000000",
  45947=>"001000000",
  45948=>"100110001",
  45949=>"111000011",
  45950=>"000000000",
  45951=>"010011000",
  45952=>"000000000",
  45953=>"111011000",
  45954=>"010000000",
  45955=>"000000111",
  45956=>"101000101",
  45957=>"010000111",
  45958=>"000000100",
  45959=>"101111011",
  45960=>"001001001",
  45961=>"100000000",
  45962=>"111000000",
  45963=>"110111111",
  45964=>"000000111",
  45965=>"001001000",
  45966=>"000000000",
  45967=>"000010000",
  45968=>"101101001",
  45969=>"110000111",
  45970=>"111100111",
  45971=>"111001001",
  45972=>"000000000",
  45973=>"000001001",
  45974=>"111111111",
  45975=>"000000000",
  45976=>"000001011",
  45977=>"011011111",
  45978=>"100101111",
  45979=>"001111011",
  45980=>"101000100",
  45981=>"000000111",
  45982=>"111111000",
  45983=>"001001001",
  45984=>"111101111",
  45985=>"110110110",
  45986=>"110000000",
  45987=>"111101111",
  45988=>"000000000",
  45989=>"000000000",
  45990=>"101100000",
  45991=>"001001000",
  45992=>"000000000",
  45993=>"111001000",
  45994=>"000000111",
  45995=>"010000000",
  45996=>"000000101",
  45997=>"101111101",
  45998=>"010000000",
  45999=>"111111011",
  46000=>"000010111",
  46001=>"011000000",
  46002=>"101111111",
  46003=>"001000000",
  46004=>"110111010",
  46005=>"111000000",
  46006=>"111000000",
  46007=>"111110110",
  46008=>"001001000",
  46009=>"111101111",
  46010=>"111011011",
  46011=>"000101111",
  46012=>"011011000",
  46013=>"111111111",
  46014=>"000111111",
  46015=>"010110000",
  46016=>"001001101",
  46017=>"101111000",
  46018=>"110111011",
  46019=>"110110000",
  46020=>"111101000",
  46021=>"101000000",
  46022=>"000000000",
  46023=>"100100101",
  46024=>"000111111",
  46025=>"111000000",
  46026=>"101000001",
  46027=>"001000000",
  46028=>"000000000",
  46029=>"001001001",
  46030=>"000000000",
  46031=>"111101100",
  46032=>"000110111",
  46033=>"111111111",
  46034=>"000000000",
  46035=>"110111110",
  46036=>"111110100",
  46037=>"111111001",
  46038=>"001000001",
  46039=>"011000100",
  46040=>"111000100",
  46041=>"110110000",
  46042=>"010000010",
  46043=>"100000111",
  46044=>"000000000",
  46045=>"000000000",
  46046=>"100000000",
  46047=>"010000100",
  46048=>"000110000",
  46049=>"100111110",
  46050=>"111110011",
  46051=>"000000010",
  46052=>"001000000",
  46053=>"101101101",
  46054=>"111111111",
  46055=>"100000000",
  46056=>"000000111",
  46057=>"111111110",
  46058=>"111000000",
  46059=>"001000000",
  46060=>"110111110",
  46061=>"011000000",
  46062=>"111111111",
  46063=>"111111000",
  46064=>"111111010",
  46065=>"010111111",
  46066=>"100000000",
  46067=>"111000000",
  46068=>"111000000",
  46069=>"000000101",
  46070=>"000000101",
  46071=>"001001111",
  46072=>"111101100",
  46073=>"001001000",
  46074=>"000000011",
  46075=>"111000000",
  46076=>"001110110",
  46077=>"000000000",
  46078=>"000000000",
  46079=>"000000000",
  46080=>"111110110",
  46081=>"011000000",
  46082=>"000000100",
  46083=>"000000001",
  46084=>"000000000",
  46085=>"000000111",
  46086=>"000000000",
  46087=>"111101111",
  46088=>"100111110",
  46089=>"111101000",
  46090=>"111111111",
  46091=>"000010000",
  46092=>"100111111",
  46093=>"111110000",
  46094=>"000110101",
  46095=>"111111000",
  46096=>"000001000",
  46097=>"110111111",
  46098=>"000000011",
  46099=>"000000000",
  46100=>"111111000",
  46101=>"000000000",
  46102=>"000100000",
  46103=>"011101100",
  46104=>"000000000",
  46105=>"100000011",
  46106=>"000000000",
  46107=>"111011000",
  46108=>"111111111",
  46109=>"111110100",
  46110=>"111111111",
  46111=>"010111000",
  46112=>"111111101",
  46113=>"111111110",
  46114=>"000000000",
  46115=>"000000100",
  46116=>"001001001",
  46117=>"111111111",
  46118=>"111111111",
  46119=>"000011111",
  46120=>"111111110",
  46121=>"000000000",
  46122=>"111111111",
  46123=>"000000000",
  46124=>"000000000",
  46125=>"100011011",
  46126=>"000000111",
  46127=>"011000100",
  46128=>"000000000",
  46129=>"001000000",
  46130=>"000000000",
  46131=>"000111111",
  46132=>"100111111",
  46133=>"100100100",
  46134=>"000000001",
  46135=>"111111101",
  46136=>"111111111",
  46137=>"000001000",
  46138=>"111111111",
  46139=>"000111111",
  46140=>"100100000",
  46141=>"000000100",
  46142=>"111111010",
  46143=>"000000000",
  46144=>"111111000",
  46145=>"000000010",
  46146=>"000111011",
  46147=>"110100011",
  46148=>"000000000",
  46149=>"000000001",
  46150=>"111111111",
  46151=>"000000000",
  46152=>"110110011",
  46153=>"000000000",
  46154=>"110011111",
  46155=>"111111100",
  46156=>"000011010",
  46157=>"100111001",
  46158=>"000000000",
  46159=>"000000000",
  46160=>"000000000",
  46161=>"100110111",
  46162=>"111111000",
  46163=>"111111111",
  46164=>"001000000",
  46165=>"111111111",
  46166=>"111111000",
  46167=>"100000000",
  46168=>"111111111",
  46169=>"000000000",
  46170=>"000001011",
  46171=>"000100100",
  46172=>"000010110",
  46173=>"111111010",
  46174=>"111111111",
  46175=>"110111000",
  46176=>"110111111",
  46177=>"000111111",
  46178=>"000000000",
  46179=>"111111111",
  46180=>"111111111",
  46181=>"001101100",
  46182=>"111101111",
  46183=>"111110110",
  46184=>"111000000",
  46185=>"000000000",
  46186=>"000001001",
  46187=>"000010011",
  46188=>"111101111",
  46189=>"000001001",
  46190=>"111111100",
  46191=>"111111111",
  46192=>"111010000",
  46193=>"000000111",
  46194=>"110110111",
  46195=>"001000001",
  46196=>"001000101",
  46197=>"111101111",
  46198=>"000100101",
  46199=>"000000001",
  46200=>"000010011",
  46201=>"000000110",
  46202=>"000000000",
  46203=>"000100111",
  46204=>"100000100",
  46205=>"011111111",
  46206=>"000100100",
  46207=>"010010001",
  46208=>"101100100",
  46209=>"000000000",
  46210=>"000000000",
  46211=>"111111111",
  46212=>"111001001",
  46213=>"011001000",
  46214=>"101111111",
  46215=>"101111111",
  46216=>"000000111",
  46217=>"000101111",
  46218=>"000000000",
  46219=>"111000111",
  46220=>"111000000",
  46221=>"111111111",
  46222=>"000000011",
  46223=>"000000000",
  46224=>"111111111",
  46225=>"001011111",
  46226=>"111110000",
  46227=>"000000000",
  46228=>"000001111",
  46229=>"110111111",
  46230=>"111111111",
  46231=>"111100000",
  46232=>"000101001",
  46233=>"100000000",
  46234=>"000000101",
  46235=>"111111111",
  46236=>"000000000",
  46237=>"111111111",
  46238=>"000000000",
  46239=>"000000000",
  46240=>"000000000",
  46241=>"010010001",
  46242=>"001010100",
  46243=>"000000110",
  46244=>"000100110",
  46245=>"111000111",
  46246=>"000000100",
  46247=>"100000011",
  46248=>"111111111",
  46249=>"000000000",
  46250=>"000000000",
  46251=>"000000000",
  46252=>"000000000",
  46253=>"000000100",
  46254=>"000000001",
  46255=>"111111000",
  46256=>"111011000",
  46257=>"000111100",
  46258=>"000111110",
  46259=>"000000000",
  46260=>"111100110",
  46261=>"000000000",
  46262=>"011011011",
  46263=>"000000010",
  46264=>"000000000",
  46265=>"000000100",
  46266=>"000000000",
  46267=>"110100111",
  46268=>"111111011",
  46269=>"111111111",
  46270=>"111000111",
  46271=>"111111111",
  46272=>"001011100",
  46273=>"001000000",
  46274=>"001001001",
  46275=>"000000000",
  46276=>"000000000",
  46277=>"000000000",
  46278=>"001001001",
  46279=>"111111011",
  46280=>"000111111",
  46281=>"000000000",
  46282=>"001000000",
  46283=>"100000000",
  46284=>"000000000",
  46285=>"000100111",
  46286=>"111111111",
  46287=>"011111011",
  46288=>"111011001",
  46289=>"011111111",
  46290=>"001000111",
  46291=>"000000000",
  46292=>"000000001",
  46293=>"000000100",
  46294=>"000000000",
  46295=>"111000111",
  46296=>"111101011",
  46297=>"011111111",
  46298=>"111000000",
  46299=>"111111111",
  46300=>"000000100",
  46301=>"000100111",
  46302=>"000000000",
  46303=>"000000111",
  46304=>"000000000",
  46305=>"000111111",
  46306=>"110000000",
  46307=>"111111111",
  46308=>"111011001",
  46309=>"000000011",
  46310=>"111111111",
  46311=>"110111110",
  46312=>"000000000",
  46313=>"110100000",
  46314=>"001001000",
  46315=>"110001001",
  46316=>"101011000",
  46317=>"000000110",
  46318=>"000110111",
  46319=>"000000000",
  46320=>"000100101",
  46321=>"000000000",
  46322=>"000000000",
  46323=>"000000000",
  46324=>"000000111",
  46325=>"100100000",
  46326=>"110110100",
  46327=>"000000000",
  46328=>"111110010",
  46329=>"000000000",
  46330=>"000111111",
  46331=>"011111111",
  46332=>"000000000",
  46333=>"110011011",
  46334=>"000000000",
  46335=>"000000000",
  46336=>"110100100",
  46337=>"011011001",
  46338=>"011000000",
  46339=>"000000000",
  46340=>"100111101",
  46341=>"000000000",
  46342=>"111111111",
  46343=>"000000000",
  46344=>"111111111",
  46345=>"000000011",
  46346=>"111111111",
  46347=>"000000001",
  46348=>"000000000",
  46349=>"000000111",
  46350=>"111111111",
  46351=>"000000000",
  46352=>"000000000",
  46353=>"111000111",
  46354=>"101111111",
  46355=>"111111111",
  46356=>"001011000",
  46357=>"111111011",
  46358=>"111100000",
  46359=>"000011001",
  46360=>"110111111",
  46361=>"111111111",
  46362=>"000000001",
  46363=>"011100000",
  46364=>"000000000",
  46365=>"000000000",
  46366=>"111100111",
  46367=>"000000000",
  46368=>"000100111",
  46369=>"110111111",
  46370=>"101100111",
  46371=>"111001111",
  46372=>"111111111",
  46373=>"000000000",
  46374=>"000000011",
  46375=>"000100111",
  46376=>"000000000",
  46377=>"000000000",
  46378=>"111111001",
  46379=>"001110000",
  46380=>"110011111",
  46381=>"001001111",
  46382=>"000111000",
  46383=>"000000000",
  46384=>"000000001",
  46385=>"000000100",
  46386=>"110000101",
  46387=>"111100111",
  46388=>"111111110",
  46389=>"111111110",
  46390=>"111100000",
  46391=>"000000000",
  46392=>"111110000",
  46393=>"111111010",
  46394=>"010111000",
  46395=>"000000110",
  46396=>"000000111",
  46397=>"111000110",
  46398=>"111111011",
  46399=>"000000000",
  46400=>"111111000",
  46401=>"000000000",
  46402=>"111111111",
  46403=>"111000000",
  46404=>"000000000",
  46405=>"000000001",
  46406=>"000000000",
  46407=>"111111111",
  46408=>"000010010",
  46409=>"010110000",
  46410=>"000000010",
  46411=>"101000100",
  46412=>"111111111",
  46413=>"000000111",
  46414=>"000001011",
  46415=>"111111111",
  46416=>"000001001",
  46417=>"000000000",
  46418=>"000000011",
  46419=>"001000000",
  46420=>"000010111",
  46421=>"001011001",
  46422=>"000000000",
  46423=>"111111111",
  46424=>"111111110",
  46425=>"110110000",
  46426=>"000000000",
  46427=>"000000000",
  46428=>"000000100",
  46429=>"111111111",
  46430=>"111111111",
  46431=>"111111110",
  46432=>"000111111",
  46433=>"111111111",
  46434=>"110110110",
  46435=>"000000000",
  46436=>"000001101",
  46437=>"000000111",
  46438=>"000000000",
  46439=>"000111111",
  46440=>"111000000",
  46441=>"111011000",
  46442=>"111111111",
  46443=>"111111111",
  46444=>"000000000",
  46445=>"000000000",
  46446=>"110110000",
  46447=>"110011011",
  46448=>"000000000",
  46449=>"000000000",
  46450=>"011111101",
  46451=>"000000000",
  46452=>"111110001",
  46453=>"000000000",
  46454=>"000000000",
  46455=>"000000000",
  46456=>"011010010",
  46457=>"000000000",
  46458=>"000000000",
  46459=>"111111111",
  46460=>"111111111",
  46461=>"111010100",
  46462=>"000000000",
  46463=>"100000000",
  46464=>"110000101",
  46465=>"000110011",
  46466=>"000000000",
  46467=>"111111010",
  46468=>"001111111",
  46469=>"000111111",
  46470=>"001101111",
  46471=>"000000000",
  46472=>"100111111",
  46473=>"000001001",
  46474=>"110111010",
  46475=>"011111000",
  46476=>"111111111",
  46477=>"010000000",
  46478=>"111110100",
  46479=>"000000000",
  46480=>"000000000",
  46481=>"011000000",
  46482=>"111110100",
  46483=>"000000000",
  46484=>"111111000",
  46485=>"000000000",
  46486=>"000010011",
  46487=>"000100000",
  46488=>"000000000",
  46489=>"111110110",
  46490=>"111111111",
  46491=>"111111111",
  46492=>"000000111",
  46493=>"111111000",
  46494=>"000000010",
  46495=>"000000101",
  46496=>"111111111",
  46497=>"111011111",
  46498=>"010110111",
  46499=>"111111011",
  46500=>"000000000",
  46501=>"000011010",
  46502=>"101000000",
  46503=>"000100111",
  46504=>"111100000",
  46505=>"111011111",
  46506=>"010111111",
  46507=>"000110000",
  46508=>"110100101",
  46509=>"110011000",
  46510=>"111111010",
  46511=>"110111111",
  46512=>"000000000",
  46513=>"000000000",
  46514=>"001010000",
  46515=>"111111111",
  46516=>"111111110",
  46517=>"000000100",
  46518=>"000000000",
  46519=>"000000001",
  46520=>"111110000",
  46521=>"000000110",
  46522=>"111100000",
  46523=>"111000100",
  46524=>"111111010",
  46525=>"101111100",
  46526=>"111000110",
  46527=>"110110111",
  46528=>"000000111",
  46529=>"011111000",
  46530=>"111111111",
  46531=>"111111000",
  46532=>"011011011",
  46533=>"111011101",
  46534=>"111111000",
  46535=>"100000010",
  46536=>"000111101",
  46537=>"000001000",
  46538=>"000000000",
  46539=>"111111111",
  46540=>"110111000",
  46541=>"111111101",
  46542=>"111111100",
  46543=>"111111111",
  46544=>"010000000",
  46545=>"000000110",
  46546=>"111111111",
  46547=>"100000000",
  46548=>"011000000",
  46549=>"111010000",
  46550=>"000000000",
  46551=>"001011011",
  46552=>"000000000",
  46553=>"111111000",
  46554=>"000000000",
  46555=>"111100110",
  46556=>"000000000",
  46557=>"111111101",
  46558=>"111111111",
  46559=>"000000001",
  46560=>"000000011",
  46561=>"111111111",
  46562=>"111111111",
  46563=>"000110111",
  46564=>"111111111",
  46565=>"000101111",
  46566=>"010000001",
  46567=>"000000000",
  46568=>"111111000",
  46569=>"111111100",
  46570=>"110000000",
  46571=>"001001001",
  46572=>"111111111",
  46573=>"000001001",
  46574=>"000000000",
  46575=>"000000000",
  46576=>"000000011",
  46577=>"000101101",
  46578=>"111111111",
  46579=>"000000000",
  46580=>"000000000",
  46581=>"100001101",
  46582=>"000000000",
  46583=>"111001000",
  46584=>"111111000",
  46585=>"000000011",
  46586=>"111000000",
  46587=>"111001101",
  46588=>"010000001",
  46589=>"111111110",
  46590=>"111111111",
  46591=>"000000100",
  46592=>"111111111",
  46593=>"000010001",
  46594=>"100000000",
  46595=>"100111111",
  46596=>"101110111",
  46597=>"001011011",
  46598=>"110111111",
  46599=>"111111011",
  46600=>"000000000",
  46601=>"000001000",
  46602=>"011000000",
  46603=>"011000011",
  46604=>"000011000",
  46605=>"100000000",
  46606=>"011111111",
  46607=>"000000111",
  46608=>"000000000",
  46609=>"000000001",
  46610=>"100100000",
  46611=>"000010111",
  46612=>"111110000",
  46613=>"010011111",
  46614=>"110000101",
  46615=>"010011000",
  46616=>"000111111",
  46617=>"100100100",
  46618=>"000111000",
  46619=>"111100100",
  46620=>"111111000",
  46621=>"000010111",
  46622=>"100110100",
  46623=>"110110000",
  46624=>"111101000",
  46625=>"000011111",
  46626=>"001001000",
  46627=>"111111110",
  46628=>"000011111",
  46629=>"010011001",
  46630=>"000000000",
  46631=>"111110111",
  46632=>"100000111",
  46633=>"000000111",
  46634=>"111111111",
  46635=>"111100111",
  46636=>"000100111",
  46637=>"000000000",
  46638=>"100000000",
  46639=>"000000111",
  46640=>"000101111",
  46641=>"000000000",
  46642=>"000000000",
  46643=>"000000000",
  46644=>"000111111",
  46645=>"000011000",
  46646=>"111000000",
  46647=>"000000000",
  46648=>"000000111",
  46649=>"000000000",
  46650=>"000001000",
  46651=>"111111111",
  46652=>"000111111",
  46653=>"101000111",
  46654=>"001111110",
  46655=>"111111000",
  46656=>"111101000",
  46657=>"011000110",
  46658=>"111111111",
  46659=>"111000111",
  46660=>"000000000",
  46661=>"001001001",
  46662=>"101000000",
  46663=>"000010000",
  46664=>"001001011",
  46665=>"000000000",
  46666=>"111101101",
  46667=>"111111111",
  46668=>"111101001",
  46669=>"000011111",
  46670=>"111111111",
  46671=>"010000000",
  46672=>"111001111",
  46673=>"111111000",
  46674=>"110100000",
  46675=>"000000100",
  46676=>"000000110",
  46677=>"111111111",
  46678=>"101000101",
  46679=>"000000111",
  46680=>"000000100",
  46681=>"101000111",
  46682=>"111010000",
  46683=>"100001001",
  46684=>"111110100",
  46685=>"001101111",
  46686=>"111111011",
  46687=>"111000000",
  46688=>"010110110",
  46689=>"111111100",
  46690=>"000000000",
  46691=>"111111111",
  46692=>"000111100",
  46693=>"100100111",
  46694=>"111011000",
  46695=>"000000000",
  46696=>"000000000",
  46697=>"111111110",
  46698=>"001011000",
  46699=>"111111010",
  46700=>"111111000",
  46701=>"011111111",
  46702=>"000000010",
  46703=>"111100100",
  46704=>"000000111",
  46705=>"000000111",
  46706=>"000111111",
  46707=>"111100000",
  46708=>"000000111",
  46709=>"100100000",
  46710=>"000000010",
  46711=>"000000110",
  46712=>"100111111",
  46713=>"111111011",
  46714=>"000111111",
  46715=>"111000000",
  46716=>"011011100",
  46717=>"000010000",
  46718=>"101100111",
  46719=>"000000110",
  46720=>"111011000",
  46721=>"110000000",
  46722=>"111000000",
  46723=>"000111111",
  46724=>"000000111",
  46725=>"111111111",
  46726=>"110110111",
  46727=>"110111111",
  46728=>"111111000",
  46729=>"011000001",
  46730=>"000111111",
  46731=>"111111000",
  46732=>"111011011",
  46733=>"000000111",
  46734=>"001111111",
  46735=>"110100111",
  46736=>"111111110",
  46737=>"000000000",
  46738=>"111000100",
  46739=>"000110000",
  46740=>"110110100",
  46741=>"100100111",
  46742=>"111110111",
  46743=>"000011000",
  46744=>"110111000",
  46745=>"001111101",
  46746=>"111000000",
  46747=>"001000000",
  46748=>"001000100",
  46749=>"110111001",
  46750=>"101000011",
  46751=>"011111111",
  46752=>"000001011",
  46753=>"111110000",
  46754=>"111000010",
  46755=>"000000111",
  46756=>"000111111",
  46757=>"100110111",
  46758=>"111011000",
  46759=>"110111111",
  46760=>"111001111",
  46761=>"111111111",
  46762=>"111000000",
  46763=>"000011000",
  46764=>"011001001",
  46765=>"110000000",
  46766=>"111100000",
  46767=>"000001000",
  46768=>"111111111",
  46769=>"000000100",
  46770=>"011111000",
  46771=>"111110010",
  46772=>"000110111",
  46773=>"000101111",
  46774=>"000000001",
  46775=>"001001111",
  46776=>"001000110",
  46777=>"000000000",
  46778=>"000101111",
  46779=>"100001001",
  46780=>"111111100",
  46781=>"000000011",
  46782=>"111111111",
  46783=>"000101111",
  46784=>"000100101",
  46785=>"111101111",
  46786=>"000000111",
  46787=>"000000000",
  46788=>"111111111",
  46789=>"000000111",
  46790=>"111001111",
  46791=>"000100111",
  46792=>"000000111",
  46793=>"011001000",
  46794=>"111111001",
  46795=>"000111111",
  46796=>"111011000",
  46797=>"110011011",
  46798=>"000001111",
  46799=>"111101000",
  46800=>"000000110",
  46801=>"000000111",
  46802=>"000110000",
  46803=>"000000000",
  46804=>"110110111",
  46805=>"100000000",
  46806=>"001000000",
  46807=>"111111111",
  46808=>"111111101",
  46809=>"111000000",
  46810=>"111001000",
  46811=>"000110111",
  46812=>"111001010",
  46813=>"000000000",
  46814=>"000000110",
  46815=>"111101111",
  46816=>"000110111",
  46817=>"000011111",
  46818=>"111111110",
  46819=>"101000111",
  46820=>"000000111",
  46821=>"101111111",
  46822=>"000000000",
  46823=>"111111111",
  46824=>"001111111",
  46825=>"101100000",
  46826=>"011111101",
  46827=>"000000000",
  46828=>"111100000",
  46829=>"101101001",
  46830=>"101100110",
  46831=>"111111000",
  46832=>"000100000",
  46833=>"111110100",
  46834=>"001000001",
  46835=>"110000000",
  46836=>"010111110",
  46837=>"111111100",
  46838=>"000110110",
  46839=>"111000000",
  46840=>"101100111",
  46841=>"000000100",
  46842=>"111001111",
  46843=>"101100000",
  46844=>"000011111",
  46845=>"110010010",
  46846=>"111000000",
  46847=>"111000111",
  46848=>"000110000",
  46849=>"000100000",
  46850=>"111111000",
  46851=>"000000111",
  46852=>"001000000",
  46853=>"001001000",
  46854=>"100101001",
  46855=>"001000111",
  46856=>"000000000",
  46857=>"000110000",
  46858=>"111111111",
  46859=>"001111111",
  46860=>"111111011",
  46861=>"111011011",
  46862=>"001110111",
  46863=>"111111000",
  46864=>"111111100",
  46865=>"000000000",
  46866=>"101111111",
  46867=>"000000111",
  46868=>"001011000",
  46869=>"000001000",
  46870=>"110111110",
  46871=>"000100111",
  46872=>"111111111",
  46873=>"000100000",
  46874=>"111111110",
  46875=>"111101001",
  46876=>"100000000",
  46877=>"111110000",
  46878=>"101111111",
  46879=>"000000000",
  46880=>"000000000",
  46881=>"111111111",
  46882=>"111111001",
  46883=>"111000000",
  46884=>"111111111",
  46885=>"111111101",
  46886=>"111000000",
  46887=>"100000000",
  46888=>"110100000",
  46889=>"011111111",
  46890=>"111001000",
  46891=>"111100010",
  46892=>"111111111",
  46893=>"110100000",
  46894=>"111011011",
  46895=>"111100000",
  46896=>"011111010",
  46897=>"000000000",
  46898=>"111110000",
  46899=>"000000110",
  46900=>"111000001",
  46901=>"000010111",
  46902=>"001000000",
  46903=>"111111111",
  46904=>"000000000",
  46905=>"000000000",
  46906=>"111100100",
  46907=>"000001000",
  46908=>"001111111",
  46909=>"000000000",
  46910=>"000000000",
  46911=>"000000001",
  46912=>"111000100",
  46913=>"000100111",
  46914=>"100000000",
  46915=>"000000101",
  46916=>"111111111",
  46917=>"111111111",
  46918=>"001001101",
  46919=>"000000000",
  46920=>"111101100",
  46921=>"000000000",
  46922=>"101111111",
  46923=>"111011000",
  46924=>"000000000",
  46925=>"111111111",
  46926=>"100100111",
  46927=>"111111111",
  46928=>"000010111",
  46929=>"101111111",
  46930=>"111011000",
  46931=>"000111111",
  46932=>"010000000",
  46933=>"000000000",
  46934=>"001001001",
  46935=>"100000000",
  46936=>"000000100",
  46937=>"111100110",
  46938=>"000000111",
  46939=>"111110000",
  46940=>"110010111",
  46941=>"000000000",
  46942=>"111001000",
  46943=>"111000011",
  46944=>"000111111",
  46945=>"011111000",
  46946=>"011011000",
  46947=>"111001001",
  46948=>"000000000",
  46949=>"000000000",
  46950=>"000111111",
  46951=>"000000001",
  46952=>"111100000",
  46953=>"000000000",
  46954=>"000111111",
  46955=>"011010000",
  46956=>"010011001",
  46957=>"011001111",
  46958=>"111111000",
  46959=>"000000111",
  46960=>"111100000",
  46961=>"100111111",
  46962=>"000000010",
  46963=>"001111111",
  46964=>"111111111",
  46965=>"111100100",
  46966=>"001000110",
  46967=>"000000111",
  46968=>"111101111",
  46969=>"100110000",
  46970=>"000100000",
  46971=>"110000000",
  46972=>"011111111",
  46973=>"001000110",
  46974=>"111000000",
  46975=>"111001000",
  46976=>"001000111",
  46977=>"010111001",
  46978=>"000000110",
  46979=>"111101111",
  46980=>"000000111",
  46981=>"100000000",
  46982=>"111111111",
  46983=>"010010001",
  46984=>"111111111",
  46985=>"011000100",
  46986=>"101001001",
  46987=>"100100000",
  46988=>"111000011",
  46989=>"111111110",
  46990=>"001000000",
  46991=>"100111111",
  46992=>"001101001",
  46993=>"000000101",
  46994=>"111111111",
  46995=>"111100100",
  46996=>"111001000",
  46997=>"000110100",
  46998=>"111001011",
  46999=>"010011111",
  47000=>"000000111",
  47001=>"000000000",
  47002=>"000000001",
  47003=>"111110111",
  47004=>"000000000",
  47005=>"000000000",
  47006=>"000001011",
  47007=>"110000000",
  47008=>"000000000",
  47009=>"111100100",
  47010=>"011000100",
  47011=>"111111111",
  47012=>"111001011",
  47013=>"000010000",
  47014=>"111000000",
  47015=>"111111111",
  47016=>"000000000",
  47017=>"101001001",
  47018=>"101000001",
  47019=>"100000000",
  47020=>"000111111",
  47021=>"000000000",
  47022=>"111101000",
  47023=>"100000000",
  47024=>"111111111",
  47025=>"111111111",
  47026=>"111111011",
  47027=>"101000000",
  47028=>"111100000",
  47029=>"001001000",
  47030=>"111111100",
  47031=>"000011000",
  47032=>"000000000",
  47033=>"011011111",
  47034=>"000001000",
  47035=>"000000000",
  47036=>"000000010",
  47037=>"001000011",
  47038=>"000000000",
  47039=>"111011001",
  47040=>"001001000",
  47041=>"111111000",
  47042=>"111010000",
  47043=>"111111111",
  47044=>"001000111",
  47045=>"001001111",
  47046=>"000110111",
  47047=>"111111111",
  47048=>"111111010",
  47049=>"110100100",
  47050=>"101111011",
  47051=>"000111000",
  47052=>"000000000",
  47053=>"000101000",
  47054=>"100000011",
  47055=>"101100100",
  47056=>"111111111",
  47057=>"111000000",
  47058=>"001000111",
  47059=>"111111100",
  47060=>"110110110",
  47061=>"011000000",
  47062=>"000000011",
  47063=>"000000000",
  47064=>"111000000",
  47065=>"111011010",
  47066=>"000000000",
  47067=>"111000000",
  47068=>"111011011",
  47069=>"000101111",
  47070=>"000000000",
  47071=>"111111111",
  47072=>"000000000",
  47073=>"000111001",
  47074=>"111100100",
  47075=>"000000000",
  47076=>"111011001",
  47077=>"000000001",
  47078=>"010111000",
  47079=>"111001000",
  47080=>"110110111",
  47081=>"000000100",
  47082=>"001011000",
  47083=>"001111101",
  47084=>"111101000",
  47085=>"100100000",
  47086=>"000111111",
  47087=>"000011111",
  47088=>"111111111",
  47089=>"111000000",
  47090=>"011010011",
  47091=>"101000111",
  47092=>"000111111",
  47093=>"000000000",
  47094=>"110111000",
  47095=>"100010000",
  47096=>"000001001",
  47097=>"111100000",
  47098=>"000000000",
  47099=>"110000000",
  47100=>"000011010",
  47101=>"010000000",
  47102=>"000001000",
  47103=>"000000110",
  47104=>"111111111",
  47105=>"000000000",
  47106=>"000111111",
  47107=>"001000011",
  47108=>"001000000",
  47109=>"000000000",
  47110=>"110110000",
  47111=>"111111100",
  47112=>"000000000",
  47113=>"111111111",
  47114=>"111111111",
  47115=>"000000000",
  47116=>"001111100",
  47117=>"111000000",
  47118=>"101101101",
  47119=>"111111000",
  47120=>"111111111",
  47121=>"000000000",
  47122=>"000000100",
  47123=>"000000111",
  47124=>"000010110",
  47125=>"000000111",
  47126=>"000000111",
  47127=>"011011001",
  47128=>"001110110",
  47129=>"111111110",
  47130=>"000000101",
  47131=>"111110000",
  47132=>"000000000",
  47133=>"111111000",
  47134=>"111101111",
  47135=>"011011000",
  47136=>"000000000",
  47137=>"000000100",
  47138=>"001001000",
  47139=>"001000000",
  47140=>"111111111",
  47141=>"010111111",
  47142=>"000000000",
  47143=>"111111111",
  47144=>"001111100",
  47145=>"000000000",
  47146=>"000000000",
  47147=>"110000000",
  47148=>"111111111",
  47149=>"100000000",
  47150=>"011001000",
  47151=>"110110111",
  47152=>"111111111",
  47153=>"111101000",
  47154=>"000000000",
  47155=>"000000000",
  47156=>"000000111",
  47157=>"111100100",
  47158=>"110100100",
  47159=>"000010111",
  47160=>"101111111",
  47161=>"000000000",
  47162=>"101001000",
  47163=>"001000000",
  47164=>"111111111",
  47165=>"110100000",
  47166=>"100110100",
  47167=>"100111000",
  47168=>"000000000",
  47169=>"011001011",
  47170=>"000111111",
  47171=>"000000000",
  47172=>"010000000",
  47173=>"000000000",
  47174=>"110000001",
  47175=>"111111111",
  47176=>"111111111",
  47177=>"000000000",
  47178=>"111111000",
  47179=>"110111101",
  47180=>"000000000",
  47181=>"000000100",
  47182=>"111111111",
  47183=>"111111111",
  47184=>"000000000",
  47185=>"111111001",
  47186=>"000010111",
  47187=>"111001000",
  47188=>"100100100",
  47189=>"110111110",
  47190=>"000111111",
  47191=>"000000001",
  47192=>"000000000",
  47193=>"000000000",
  47194=>"000000111",
  47195=>"011111001",
  47196=>"000000001",
  47197=>"111111101",
  47198=>"001101000",
  47199=>"111111110",
  47200=>"000000000",
  47201=>"111111111",
  47202=>"000000000",
  47203=>"011000001",
  47204=>"001110000",
  47205=>"000000000",
  47206=>"000110000",
  47207=>"001111111",
  47208=>"000000000",
  47209=>"000000111",
  47210=>"100100111",
  47211=>"111111111",
  47212=>"011010110",
  47213=>"000100100",
  47214=>"100000000",
  47215=>"111111111",
  47216=>"000100101",
  47217=>"101111000",
  47218=>"101100101",
  47219=>"000001001",
  47220=>"000000000",
  47221=>"011111111",
  47222=>"100000111",
  47223=>"100000010",
  47224=>"100000000",
  47225=>"111111100",
  47226=>"101100110",
  47227=>"111111001",
  47228=>"001001000",
  47229=>"111111111",
  47230=>"000000000",
  47231=>"011011000",
  47232=>"010111010",
  47233=>"001000011",
  47234=>"111111111",
  47235=>"111000000",
  47236=>"000100101",
  47237=>"111111111",
  47238=>"000000000",
  47239=>"010100000",
  47240=>"111000100",
  47241=>"000000110",
  47242=>"110111011",
  47243=>"111111111",
  47244=>"111111111",
  47245=>"010110000",
  47246=>"111000000",
  47247=>"000001001",
  47248=>"100000101",
  47249=>"101111001",
  47250=>"001111101",
  47251=>"000000110",
  47252=>"100100000",
  47253=>"001101111",
  47254=>"111001000",
  47255=>"111100110",
  47256=>"000000000",
  47257=>"000000000",
  47258=>"111111111",
  47259=>"111111111",
  47260=>"000100100",
  47261=>"000001001",
  47262=>"100111111",
  47263=>"000000000",
  47264=>"000000000",
  47265=>"010000000",
  47266=>"000110001",
  47267=>"000010000",
  47268=>"001100100",
  47269=>"000000000",
  47270=>"110111111",
  47271=>"000000111",
  47272=>"011011000",
  47273=>"101100000",
  47274=>"000000000",
  47275=>"000111111",
  47276=>"111111111",
  47277=>"011001001",
  47278=>"111111000",
  47279=>"110100000",
  47280=>"000010000",
  47281=>"111011101",
  47282=>"111110110",
  47283=>"000000000",
  47284=>"110011000",
  47285=>"000000111",
  47286=>"111111111",
  47287=>"000000000",
  47288=>"111101000",
  47289=>"000000000",
  47290=>"000000100",
  47291=>"000110111",
  47292=>"000000000",
  47293=>"000000000",
  47294=>"111111111",
  47295=>"111111111",
  47296=>"000001011",
  47297=>"111111111",
  47298=>"001111111",
  47299=>"101101111",
  47300=>"111000111",
  47301=>"000000000",
  47302=>"000000010",
  47303=>"101000101",
  47304=>"000010000",
  47305=>"111111001",
  47306=>"001001000",
  47307=>"100101111",
  47308=>"000100000",
  47309=>"111111111",
  47310=>"000011010",
  47311=>"000000000",
  47312=>"111110000",
  47313=>"111111111",
  47314=>"010111000",
  47315=>"000010000",
  47316=>"111110111",
  47317=>"001001111",
  47318=>"000000111",
  47319=>"000001001",
  47320=>"111111111",
  47321=>"000111111",
  47322=>"000000000",
  47323=>"000110111",
  47324=>"000000000",
  47325=>"000000001",
  47326=>"111111111",
  47327=>"000000000",
  47328=>"001111000",
  47329=>"111111111",
  47330=>"110110000",
  47331=>"111110110",
  47332=>"000000000",
  47333=>"110111110",
  47334=>"101111101",
  47335=>"110100100",
  47336=>"100000000",
  47337=>"101111111",
  47338=>"110110101",
  47339=>"111111101",
  47340=>"011000000",
  47341=>"000000000",
  47342=>"000000111",
  47343=>"010111011",
  47344=>"111010110",
  47345=>"000110111",
  47346=>"001011111",
  47347=>"010010000",
  47348=>"111111111",
  47349=>"000001001",
  47350=>"111110000",
  47351=>"000000000",
  47352=>"000000100",
  47353=>"000000111",
  47354=>"000000000",
  47355=>"001000000",
  47356=>"000000001",
  47357=>"000001000",
  47358=>"000001111",
  47359=>"100111111",
  47360=>"110110110",
  47361=>"111101101",
  47362=>"111111011",
  47363=>"001111110",
  47364=>"111111111",
  47365=>"001011010",
  47366=>"111111000",
  47367=>"000111111",
  47368=>"111111010",
  47369=>"111000111",
  47370=>"010111011",
  47371=>"000101000",
  47372=>"110111100",
  47373=>"111111110",
  47374=>"001001111",
  47375=>"000000000",
  47376=>"001000000",
  47377=>"111111111",
  47378=>"001111011",
  47379=>"000111101",
  47380=>"000000000",
  47381=>"100100111",
  47382=>"011001001",
  47383=>"000000100",
  47384=>"111111111",
  47385=>"000000000",
  47386=>"001111111",
  47387=>"000010111",
  47388=>"001111100",
  47389=>"010000000",
  47390=>"010000000",
  47391=>"111111001",
  47392=>"100110100",
  47393=>"000000011",
  47394=>"000000110",
  47395=>"111111101",
  47396=>"111111100",
  47397=>"010010111",
  47398=>"111111111",
  47399=>"001111111",
  47400=>"111000000",
  47401=>"000000000",
  47402=>"000000010",
  47403=>"000000001",
  47404=>"000111111",
  47405=>"111111111",
  47406=>"000000000",
  47407=>"100000000",
  47408=>"000000000",
  47409=>"111011010",
  47410=>"100010111",
  47411=>"101111111",
  47412=>"110000000",
  47413=>"000000000",
  47414=>"000000000",
  47415=>"000011001",
  47416=>"000000000",
  47417=>"000101111",
  47418=>"000000101",
  47419=>"000000000",
  47420=>"000000000",
  47421=>"000000000",
  47422=>"100111111",
  47423=>"110111010",
  47424=>"101100111",
  47425=>"000000101",
  47426=>"000110000",
  47427=>"000000000",
  47428=>"110000000",
  47429=>"001011111",
  47430=>"000000000",
  47431=>"111111111",
  47432=>"011111111",
  47433=>"000000000",
  47434=>"100000000",
  47435=>"100000000",
  47436=>"000000000",
  47437=>"011111011",
  47438=>"000010110",
  47439=>"000000110",
  47440=>"000101111",
  47441=>"000111111",
  47442=>"001011111",
  47443=>"110010111",
  47444=>"111111111",
  47445=>"000000001",
  47446=>"110100111",
  47447=>"000000001",
  47448=>"111111111",
  47449=>"010000000",
  47450=>"011111000",
  47451=>"111111111",
  47452=>"000000000",
  47453=>"011011011",
  47454=>"110011011",
  47455=>"111001111",
  47456=>"111110111",
  47457=>"001001111",
  47458=>"111110111",
  47459=>"111100100",
  47460=>"001000100",
  47461=>"000000000",
  47462=>"001000001",
  47463=>"000000000",
  47464=>"110110100",
  47465=>"111101000",
  47466=>"000000000",
  47467=>"000000000",
  47468=>"000000000",
  47469=>"000000100",
  47470=>"000000000",
  47471=>"000000001",
  47472=>"011001000",
  47473=>"000011111",
  47474=>"010110000",
  47475=>"111111111",
  47476=>"100110110",
  47477=>"000000000",
  47478=>"000101001",
  47479=>"000000001",
  47480=>"000000000",
  47481=>"000000011",
  47482=>"001000000",
  47483=>"100000001",
  47484=>"001101000",
  47485=>"111111111",
  47486=>"000000100",
  47487=>"111111110",
  47488=>"000100101",
  47489=>"111111111",
  47490=>"000000000",
  47491=>"000000100",
  47492=>"000000000",
  47493=>"000000000",
  47494=>"110001011",
  47495=>"111111111",
  47496=>"111110000",
  47497=>"000001111",
  47498=>"111111011",
  47499=>"111001000",
  47500=>"101000000",
  47501=>"100000000",
  47502=>"000000110",
  47503=>"000011000",
  47504=>"011011010",
  47505=>"110111000",
  47506=>"110110000",
  47507=>"000000000",
  47508=>"000000000",
  47509=>"000000000",
  47510=>"111111111",
  47511=>"001001001",
  47512=>"100111111",
  47513=>"111111011",
  47514=>"010000110",
  47515=>"000000110",
  47516=>"011111111",
  47517=>"010111100",
  47518=>"111011011",
  47519=>"000000000",
  47520=>"001110111",
  47521=>"110111111",
  47522=>"111111111",
  47523=>"000000111",
  47524=>"000100000",
  47525=>"000000000",
  47526=>"000000000",
  47527=>"001001000",
  47528=>"000000000",
  47529=>"100000000",
  47530=>"000111111",
  47531=>"000000000",
  47532=>"000000000",
  47533=>"000011000",
  47534=>"000011111",
  47535=>"111000000",
  47536=>"011001000",
  47537=>"111000000",
  47538=>"000000011",
  47539=>"001000111",
  47540=>"111111000",
  47541=>"111101111",
  47542=>"110111111",
  47543=>"000001101",
  47544=>"000000111",
  47545=>"111110100",
  47546=>"111111111",
  47547=>"011111111",
  47548=>"111111111",
  47549=>"111111111",
  47550=>"111111111",
  47551=>"101110101",
  47552=>"011011010",
  47553=>"111000000",
  47554=>"000100000",
  47555=>"000000000",
  47556=>"000001001",
  47557=>"100000111",
  47558=>"000000000",
  47559=>"001101001",
  47560=>"000000001",
  47561=>"000000000",
  47562=>"000000000",
  47563=>"010000011",
  47564=>"010000001",
  47565=>"000000000",
  47566=>"100100000",
  47567=>"110110111",
  47568=>"000000011",
  47569=>"000000110",
  47570=>"000000111",
  47571=>"111111111",
  47572=>"000011000",
  47573=>"111101101",
  47574=>"001111000",
  47575=>"110100100",
  47576=>"111111110",
  47577=>"000000000",
  47578=>"001111001",
  47579=>"000011111",
  47580=>"000000000",
  47581=>"000010000",
  47582=>"111111111",
  47583=>"001000000",
  47584=>"001000100",
  47585=>"110000000",
  47586=>"000000010",
  47587=>"000100111",
  47588=>"000000001",
  47589=>"000111111",
  47590=>"000000000",
  47591=>"000000000",
  47592=>"000111111",
  47593=>"111111110",
  47594=>"111110111",
  47595=>"000000000",
  47596=>"000111011",
  47597=>"100100000",
  47598=>"111111111",
  47599=>"000010100",
  47600=>"000000000",
  47601=>"000001111",
  47602=>"000000000",
  47603=>"111010000",
  47604=>"110101100",
  47605=>"000000000",
  47606=>"000000111",
  47607=>"100110111",
  47608=>"111101111",
  47609=>"000000000",
  47610=>"100001000",
  47611=>"111111111",
  47612=>"001001110",
  47613=>"000000000",
  47614=>"000000011",
  47615=>"000000000",
  47616=>"111000000",
  47617=>"011011010",
  47618=>"000000000",
  47619=>"111111111",
  47620=>"000000100",
  47621=>"111111110",
  47622=>"111111111",
  47623=>"000000000",
  47624=>"001111111",
  47625=>"111111110",
  47626=>"000000111",
  47627=>"000000111",
  47628=>"000001111",
  47629=>"110110111",
  47630=>"011111111",
  47631=>"111111111",
  47632=>"000100000",
  47633=>"001011111",
  47634=>"111111111",
  47635=>"100100000",
  47636=>"111111101",
  47637=>"001000000",
  47638=>"111111100",
  47639=>"001000001",
  47640=>"000000000",
  47641=>"111111111",
  47642=>"111111101",
  47643=>"000010011",
  47644=>"100000000",
  47645=>"010110111",
  47646=>"110110111",
  47647=>"111111000",
  47648=>"000000000",
  47649=>"000000010",
  47650=>"111111111",
  47651=>"111010011",
  47652=>"001001111",
  47653=>"100000011",
  47654=>"111111111",
  47655=>"001000000",
  47656=>"111111110",
  47657=>"000000000",
  47658=>"000000001",
  47659=>"110000111",
  47660=>"000000000",
  47661=>"000000000",
  47662=>"000010000",
  47663=>"111111111",
  47664=>"111111110",
  47665=>"001000100",
  47666=>"000000000",
  47667=>"001000111",
  47668=>"000110000",
  47669=>"111111010",
  47670=>"000000000",
  47671=>"011111111",
  47672=>"000010000",
  47673=>"010000000",
  47674=>"001001000",
  47675=>"000000111",
  47676=>"111111111",
  47677=>"100000000",
  47678=>"111000000",
  47679=>"101111111",
  47680=>"000000010",
  47681=>"000000000",
  47682=>"111111111",
  47683=>"100100111",
  47684=>"001001100",
  47685=>"111111111",
  47686=>"101100100",
  47687=>"111111111",
  47688=>"111111111",
  47689=>"111101111",
  47690=>"000000100",
  47691=>"110110111",
  47692=>"100000111",
  47693=>"111111101",
  47694=>"011011000",
  47695=>"111111111",
  47696=>"111111111",
  47697=>"111111110",
  47698=>"100000000",
  47699=>"001001011",
  47700=>"000000000",
  47701=>"110110111",
  47702=>"001011111",
  47703=>"111111111",
  47704=>"111111111",
  47705=>"000000000",
  47706=>"100000000",
  47707=>"110111111",
  47708=>"111111111",
  47709=>"111111111",
  47710=>"111111111",
  47711=>"111101111",
  47712=>"111111111",
  47713=>"000010111",
  47714=>"110100000",
  47715=>"111000111",
  47716=>"011011011",
  47717=>"001111111",
  47718=>"110110000",
  47719=>"000111111",
  47720=>"111111100",
  47721=>"000000000",
  47722=>"111000000",
  47723=>"010111110",
  47724=>"100000000",
  47725=>"000000000",
  47726=>"111110111",
  47727=>"010110111",
  47728=>"111111010",
  47729=>"110110100",
  47730=>"000000000",
  47731=>"011001111",
  47732=>"000000000",
  47733=>"000000000",
  47734=>"000110111",
  47735=>"111110000",
  47736=>"111011000",
  47737=>"001000001",
  47738=>"000000000",
  47739=>"010111111",
  47740=>"010110110",
  47741=>"100111111",
  47742=>"111010000",
  47743=>"000000000",
  47744=>"111111111",
  47745=>"111111000",
  47746=>"111001001",
  47747=>"111000000",
  47748=>"111111111",
  47749=>"111111111",
  47750=>"000000000",
  47751=>"000000000",
  47752=>"001000001",
  47753=>"000000001",
  47754=>"111111111",
  47755=>"000100000",
  47756=>"111111111",
  47757=>"101111111",
  47758=>"000000000",
  47759=>"011000000",
  47760=>"000001011",
  47761=>"000011111",
  47762=>"111111000",
  47763=>"111111111",
  47764=>"000000000",
  47765=>"000000100",
  47766=>"001001001",
  47767=>"111111111",
  47768=>"000000100",
  47769=>"000000000",
  47770=>"111111111",
  47771=>"000011011",
  47772=>"111110100",
  47773=>"001000000",
  47774=>"000000001",
  47775=>"011111111",
  47776=>"100100000",
  47777=>"000000000",
  47778=>"010111111",
  47779=>"111111011",
  47780=>"000000000",
  47781=>"111111111",
  47782=>"000000000",
  47783=>"000000000",
  47784=>"111111111",
  47785=>"001110110",
  47786=>"000111111",
  47787=>"111000000",
  47788=>"000000000",
  47789=>"000000000",
  47790=>"111111111",
  47791=>"001001111",
  47792=>"000111100",
  47793=>"111111111",
  47794=>"111111000",
  47795=>"111111111",
  47796=>"111111011",
  47797=>"111111111",
  47798=>"111111111",
  47799=>"000000000",
  47800=>"101000100",
  47801=>"000000100",
  47802=>"000000000",
  47803=>"011011000",
  47804=>"011011111",
  47805=>"111111111",
  47806=>"111111111",
  47807=>"000100100",
  47808=>"111111111",
  47809=>"111110111",
  47810=>"110010000",
  47811=>"111111110",
  47812=>"111100111",
  47813=>"000000000",
  47814=>"110110110",
  47815=>"010000110",
  47816=>"100100111",
  47817=>"001000111",
  47818=>"000000000",
  47819=>"111111111",
  47820=>"000000000",
  47821=>"000010011",
  47822=>"111111111",
  47823=>"000000000",
  47824=>"111111111",
  47825=>"000000111",
  47826=>"001111110",
  47827=>"000000000",
  47828=>"000000000",
  47829=>"000000000",
  47830=>"000000000",
  47831=>"110111111",
  47832=>"011110000",
  47833=>"001100111",
  47834=>"111110110",
  47835=>"111101101",
  47836=>"111101111",
  47837=>"000011111",
  47838=>"011011001",
  47839=>"111001000",
  47840=>"000000000",
  47841=>"100111111",
  47842=>"011011000",
  47843=>"111111100",
  47844=>"111111111",
  47845=>"111111111",
  47846=>"011000011",
  47847=>"101000000",
  47848=>"000111100",
  47849=>"000000000",
  47850=>"111111100",
  47851=>"000000000",
  47852=>"000110111",
  47853=>"111010011",
  47854=>"001111111",
  47855=>"001111111",
  47856=>"111011000",
  47857=>"111011011",
  47858=>"000100000",
  47859=>"111011000",
  47860=>"111111000",
  47861=>"011011001",
  47862=>"001000000",
  47863=>"100000000",
  47864=>"111111011",
  47865=>"000000000",
  47866=>"100111111",
  47867=>"110110000",
  47868=>"111111111",
  47869=>"001011111",
  47870=>"100000000",
  47871=>"111111000",
  47872=>"000000000",
  47873=>"000000000",
  47874=>"000010000",
  47875=>"000011011",
  47876=>"111111110",
  47877=>"000000000",
  47878=>"010111110",
  47879=>"001001111",
  47880=>"111110110",
  47881=>"111011000",
  47882=>"111111111",
  47883=>"001000000",
  47884=>"000000010",
  47885=>"000000111",
  47886=>"000000000",
  47887=>"111110110",
  47888=>"001000000",
  47889=>"000100111",
  47890=>"000001000",
  47891=>"000000101",
  47892=>"000001001",
  47893=>"000110000",
  47894=>"001100100",
  47895=>"111111111",
  47896=>"000000000",
  47897=>"111111111",
  47898=>"100000000",
  47899=>"000000000",
  47900=>"011111111",
  47901=>"001111110",
  47902=>"111111111",
  47903=>"111000111",
  47904=>"000000000",
  47905=>"111111111",
  47906=>"111111111",
  47907=>"001000101",
  47908=>"111001001",
  47909=>"000100001",
  47910=>"000000100",
  47911=>"000000110",
  47912=>"000111111",
  47913=>"100000000",
  47914=>"001000110",
  47915=>"111010000",
  47916=>"011000000",
  47917=>"000000000",
  47918=>"101000011",
  47919=>"000000000",
  47920=>"000000000",
  47921=>"111111111",
  47922=>"000000000",
  47923=>"010011000",
  47924=>"111000000",
  47925=>"000110110",
  47926=>"111111110",
  47927=>"111101111",
  47928=>"111111000",
  47929=>"000111111",
  47930=>"000000000",
  47931=>"000000000",
  47932=>"111111111",
  47933=>"111111110",
  47934=>"000000000",
  47935=>"111111111",
  47936=>"000000000",
  47937=>"111111111",
  47938=>"001000100",
  47939=>"111111111",
  47940=>"001011000",
  47941=>"111111111",
  47942=>"101101101",
  47943=>"110111111",
  47944=>"111111000",
  47945=>"100111111",
  47946=>"111001111",
  47947=>"000000111",
  47948=>"000000000",
  47949=>"111111101",
  47950=>"000000000",
  47951=>"110000000",
  47952=>"000000000",
  47953=>"010000110",
  47954=>"111011011",
  47955=>"111111101",
  47956=>"000000000",
  47957=>"011011011",
  47958=>"111111111",
  47959=>"001000000",
  47960=>"111011111",
  47961=>"111111111",
  47962=>"000000000",
  47963=>"111001000",
  47964=>"000000000",
  47965=>"100110110",
  47966=>"000000101",
  47967=>"000000000",
  47968=>"111111111",
  47969=>"000000000",
  47970=>"001001001",
  47971=>"111111111",
  47972=>"000000001",
  47973=>"000000000",
  47974=>"111111111",
  47975=>"111111111",
  47976=>"100010011",
  47977=>"010000010",
  47978=>"111111111",
  47979=>"000000010",
  47980=>"000000000",
  47981=>"100111111",
  47982=>"000011111",
  47983=>"111111111",
  47984=>"000000000",
  47985=>"000000000",
  47986=>"000000111",
  47987=>"111111111",
  47988=>"111111011",
  47989=>"111111111",
  47990=>"011000000",
  47991=>"000000000",
  47992=>"111100111",
  47993=>"011111110",
  47994=>"111111111",
  47995=>"110110010",
  47996=>"001000000",
  47997=>"110110000",
  47998=>"111111111",
  47999=>"111111111",
  48000=>"110000001",
  48001=>"000000100",
  48002=>"111111111",
  48003=>"000000000",
  48004=>"111111111",
  48005=>"001001001",
  48006=>"001000000",
  48007=>"101100000",
  48008=>"000000000",
  48009=>"111001000",
  48010=>"000000000",
  48011=>"100111111",
  48012=>"111111111",
  48013=>"111011011",
  48014=>"000000000",
  48015=>"000000010",
  48016=>"010010000",
  48017=>"000001000",
  48018=>"000000000",
  48019=>"111111111",
  48020=>"000000000",
  48021=>"000000000",
  48022=>"111111111",
  48023=>"111111111",
  48024=>"111000000",
  48025=>"000000001",
  48026=>"000000000",
  48027=>"001001000",
  48028=>"000000000",
  48029=>"000110111",
  48030=>"100100000",
  48031=>"111111111",
  48032=>"000000000",
  48033=>"001001000",
  48034=>"100110111",
  48035=>"011111111",
  48036=>"001001111",
  48037=>"000110111",
  48038=>"111111110",
  48039=>"000000000",
  48040=>"000100111",
  48041=>"111111111",
  48042=>"000000101",
  48043=>"100010000",
  48044=>"111111111",
  48045=>"111010111",
  48046=>"010000000",
  48047=>"111111000",
  48048=>"111000001",
  48049=>"111111111",
  48050=>"111111111",
  48051=>"000000001",
  48052=>"000000000",
  48053=>"111111111",
  48054=>"110110000",
  48055=>"001001001",
  48056=>"111011000",
  48057=>"000000000",
  48058=>"111111111",
  48059=>"000000111",
  48060=>"111111111",
  48061=>"000000100",
  48062=>"111100000",
  48063=>"000000000",
  48064=>"000000000",
  48065=>"000000000",
  48066=>"001111111",
  48067=>"111111010",
  48068=>"100100000",
  48069=>"111000010",
  48070=>"000000000",
  48071=>"110100100",
  48072=>"111111111",
  48073=>"000000000",
  48074=>"000000000",
  48075=>"111111111",
  48076=>"111111000",
  48077=>"000000000",
  48078=>"001001000",
  48079=>"111111111",
  48080=>"011011000",
  48081=>"000011010",
  48082=>"001001111",
  48083=>"000000110",
  48084=>"000000000",
  48085=>"111111110",
  48086=>"000000000",
  48087=>"101101111",
  48088=>"111111111",
  48089=>"000000101",
  48090=>"000000000",
  48091=>"000000000",
  48092=>"000001000",
  48093=>"111111111",
  48094=>"111111111",
  48095=>"000000101",
  48096=>"111111111",
  48097=>"000000000",
  48098=>"010001000",
  48099=>"000001001",
  48100=>"101110111",
  48101=>"111111100",
  48102=>"000100111",
  48103=>"111111011",
  48104=>"111111110",
  48105=>"100000000",
  48106=>"000110000",
  48107=>"111100111",
  48108=>"111111111",
  48109=>"100000000",
  48110=>"000010000",
  48111=>"001001001",
  48112=>"001000001",
  48113=>"000000000",
  48114=>"000000000",
  48115=>"000000000",
  48116=>"000000000",
  48117=>"111111111",
  48118=>"000000000",
  48119=>"111111110",
  48120=>"011011111",
  48121=>"000000000",
  48122=>"111100100",
  48123=>"111111111",
  48124=>"111111111",
  48125=>"000000111",
  48126=>"000000000",
  48127=>"000000000",
  48128=>"011011111",
  48129=>"111111111",
  48130=>"111000011",
  48131=>"000000000",
  48132=>"011010100",
  48133=>"000000000",
  48134=>"111000000",
  48135=>"000000111",
  48136=>"001001111",
  48137=>"000000111",
  48138=>"000000100",
  48139=>"000000000",
  48140=>"110010001",
  48141=>"000000111",
  48142=>"100111111",
  48143=>"111111111",
  48144=>"000000000",
  48145=>"111111111",
  48146=>"111111111",
  48147=>"000000110",
  48148=>"110110100",
  48149=>"111111001",
  48150=>"111111111",
  48151=>"101000001",
  48152=>"001000100",
  48153=>"100111111",
  48154=>"111001010",
  48155=>"011011001",
  48156=>"111111111",
  48157=>"111111111",
  48158=>"110110000",
  48159=>"000000000",
  48160=>"111010000",
  48161=>"001001000",
  48162=>"110000100",
  48163=>"000000000",
  48164=>"000100000",
  48165=>"111111111",
  48166=>"111000011",
  48167=>"000001111",
  48168=>"100000101",
  48169=>"000000000",
  48170=>"101001111",
  48171=>"000000011",
  48172=>"101100000",
  48173=>"001001000",
  48174=>"000001000",
  48175=>"000000000",
  48176=>"001111110",
  48177=>"000000000",
  48178=>"110110111",
  48179=>"000000111",
  48180=>"111111000",
  48181=>"111111001",
  48182=>"000000000",
  48183=>"111100100",
  48184=>"000000010",
  48185=>"000110110",
  48186=>"000000000",
  48187=>"100000000",
  48188=>"000000000",
  48189=>"011000001",
  48190=>"111110110",
  48191=>"111000000",
  48192=>"010000000",
  48193=>"111101001",
  48194=>"000000000",
  48195=>"111111111",
  48196=>"000111100",
  48197=>"001111111",
  48198=>"011010000",
  48199=>"111111111",
  48200=>"000000000",
  48201=>"000000000",
  48202=>"011011111",
  48203=>"110111111",
  48204=>"000000000",
  48205=>"110000000",
  48206=>"111011111",
  48207=>"110111111",
  48208=>"000000000",
  48209=>"111111111",
  48210=>"000010111",
  48211=>"111111100",
  48212=>"000000000",
  48213=>"000000000",
  48214=>"011000000",
  48215=>"110110110",
  48216=>"000000000",
  48217=>"000000000",
  48218=>"111111111",
  48219=>"000000000",
  48220=>"111111111",
  48221=>"111010000",
  48222=>"111111110",
  48223=>"000000000",
  48224=>"000111111",
  48225=>"000000000",
  48226=>"100000000",
  48227=>"010011011",
  48228=>"001111001",
  48229=>"000000000",
  48230=>"000000000",
  48231=>"111111111",
  48232=>"111111001",
  48233=>"000000000",
  48234=>"111111000",
  48235=>"101111111",
  48236=>"011111111",
  48237=>"110111111",
  48238=>"000000000",
  48239=>"111111111",
  48240=>"100111010",
  48241=>"100111111",
  48242=>"000000000",
  48243=>"111101001",
  48244=>"000100111",
  48245=>"110110000",
  48246=>"000000000",
  48247=>"000000000",
  48248=>"000000000",
  48249=>"001000000",
  48250=>"000000000",
  48251=>"000000000",
  48252=>"111000000",
  48253=>"000011111",
  48254=>"000000000",
  48255=>"000000111",
  48256=>"011011111",
  48257=>"000000000",
  48258=>"000000000",
  48259=>"101100000",
  48260=>"000111111",
  48261=>"100100111",
  48262=>"011011011",
  48263=>"000000101",
  48264=>"111111111",
  48265=>"111111111",
  48266=>"111111111",
  48267=>"011111111",
  48268=>"011011111",
  48269=>"100100000",
  48270=>"111111011",
  48271=>"110111110",
  48272=>"110010010",
  48273=>"000110111",
  48274=>"000000110",
  48275=>"100000111",
  48276=>"000111111",
  48277=>"111011111",
  48278=>"000010111",
  48279=>"000000000",
  48280=>"111111111",
  48281=>"000100111",
  48282=>"110000100",
  48283=>"111111000",
  48284=>"111100100",
  48285=>"110101100",
  48286=>"110110111",
  48287=>"000000000",
  48288=>"111100110",
  48289=>"111111111",
  48290=>"000000000",
  48291=>"111000000",
  48292=>"110110111",
  48293=>"000000000",
  48294=>"111111111",
  48295=>"110110110",
  48296=>"111111111",
  48297=>"000000000",
  48298=>"111000000",
  48299=>"011111111",
  48300=>"000000110",
  48301=>"101101100",
  48302=>"111111001",
  48303=>"001111001",
  48304=>"011111111",
  48305=>"000000000",
  48306=>"111111111",
  48307=>"111110000",
  48308=>"000000000",
  48309=>"000000000",
  48310=>"000000011",
  48311=>"000111111",
  48312=>"100110110",
  48313=>"000000000",
  48314=>"111110111",
  48315=>"010000111",
  48316=>"110000000",
  48317=>"011000000",
  48318=>"111111000",
  48319=>"000000000",
  48320=>"000000000",
  48321=>"000001001",
  48322=>"111111110",
  48323=>"000000000",
  48324=>"010010000",
  48325=>"000000000",
  48326=>"101110110",
  48327=>"001011001",
  48328=>"000000000",
  48329=>"111101111",
  48330=>"000000000",
  48331=>"111110111",
  48332=>"111111110",
  48333=>"000100110",
  48334=>"000000101",
  48335=>"000000000",
  48336=>"000000000",
  48337=>"001011000",
  48338=>"000000000",
  48339=>"000000000",
  48340=>"110100110",
  48341=>"111111110",
  48342=>"011011000",
  48343=>"100100100",
  48344=>"000000100",
  48345=>"001111111",
  48346=>"100000000",
  48347=>"000000000",
  48348=>"110111000",
  48349=>"000001000",
  48350=>"000011000",
  48351=>"000000000",
  48352=>"000101111",
  48353=>"000000000",
  48354=>"111111000",
  48355=>"000000110",
  48356=>"000000111",
  48357=>"001000000",
  48358=>"010111111",
  48359=>"000000111",
  48360=>"111111111",
  48361=>"100000000",
  48362=>"111111111",
  48363=>"000000110",
  48364=>"111111111",
  48365=>"000101111",
  48366=>"000000011",
  48367=>"000000111",
  48368=>"000000000",
  48369=>"000100101",
  48370=>"111111001",
  48371=>"100101101",
  48372=>"010111111",
  48373=>"000000000",
  48374=>"110001000",
  48375=>"100000000",
  48376=>"000000111",
  48377=>"111110110",
  48378=>"000111111",
  48379=>"001000001",
  48380=>"111111010",
  48381=>"001111111",
  48382=>"111110110",
  48383=>"111111111",
  48384=>"000000000",
  48385=>"111111111",
  48386=>"111111111",
  48387=>"000011111",
  48388=>"000000100",
  48389=>"111111111",
  48390=>"111100111",
  48391=>"000111111",
  48392=>"111111111",
  48393=>"000000000",
  48394=>"111111010",
  48395=>"001111010",
  48396=>"111001001",
  48397=>"111111001",
  48398=>"000110110",
  48399=>"000110111",
  48400=>"111111110",
  48401=>"000100100",
  48402=>"000000000",
  48403=>"000000111",
  48404=>"111110000",
  48405=>"111111110",
  48406=>"011011110",
  48407=>"111111111",
  48408=>"111111011",
  48409=>"111111110",
  48410=>"000000000",
  48411=>"000000000",
  48412=>"000000000",
  48413=>"000000001",
  48414=>"111111101",
  48415=>"111111111",
  48416=>"110100010",
  48417=>"000001101",
  48418=>"011000001",
  48419=>"110110000",
  48420=>"000000000",
  48421=>"111111111",
  48422=>"000000000",
  48423=>"000000000",
  48424=>"000000011",
  48425=>"000010000",
  48426=>"111000000",
  48427=>"000111101",
  48428=>"000000000",
  48429=>"000000000",
  48430=>"111110111",
  48431=>"000000011",
  48432=>"010010000",
  48433=>"010001001",
  48434=>"111111111",
  48435=>"000110111",
  48436=>"000000000",
  48437=>"110111111",
  48438=>"101111111",
  48439=>"111111101",
  48440=>"000000000",
  48441=>"111001001",
  48442=>"111010010",
  48443=>"000000000",
  48444=>"101111111",
  48445=>"111001111",
  48446=>"000000000",
  48447=>"000110111",
  48448=>"000000000",
  48449=>"110000000",
  48450=>"111001001",
  48451=>"111111011",
  48452=>"011011010",
  48453=>"111001001",
  48454=>"000010111",
  48455=>"100000000",
  48456=>"000000000",
  48457=>"000111101",
  48458=>"111111111",
  48459=>"010000000",
  48460=>"011011011",
  48461=>"000000000",
  48462=>"110000000",
  48463=>"000100000",
  48464=>"111011011",
  48465=>"000110111",
  48466=>"000000000",
  48467=>"000011000",
  48468=>"000000000",
  48469=>"011011011",
  48470=>"000000000",
  48471=>"000100000",
  48472=>"111110100",
  48473=>"110111111",
  48474=>"000001001",
  48475=>"000000100",
  48476=>"000000000",
  48477=>"000000000",
  48478=>"000000000",
  48479=>"111111111",
  48480=>"010111000",
  48481=>"000000000",
  48482=>"111011000",
  48483=>"000000000",
  48484=>"100000000",
  48485=>"000000000",
  48486=>"111111111",
  48487=>"000000000",
  48488=>"001000000",
  48489=>"000001011",
  48490=>"000000000",
  48491=>"011101101",
  48492=>"000000010",
  48493=>"000100111",
  48494=>"000000000",
  48495=>"000000000",
  48496=>"000000000",
  48497=>"000000000",
  48498=>"000000111",
  48499=>"001001101",
  48500=>"000000000",
  48501=>"000000000",
  48502=>"100000001",
  48503=>"111111000",
  48504=>"111111000",
  48505=>"001000011",
  48506=>"111111111",
  48507=>"000000000",
  48508=>"000000000",
  48509=>"000000000",
  48510=>"111111111",
  48511=>"000000000",
  48512=>"110100110",
  48513=>"010010000",
  48514=>"110110111",
  48515=>"010000000",
  48516=>"111111111",
  48517=>"111111111",
  48518=>"000000000",
  48519=>"101000111",
  48520=>"111111111",
  48521=>"000000000",
  48522=>"000000011",
  48523=>"111011001",
  48524=>"110111111",
  48525=>"011001100",
  48526=>"100000000",
  48527=>"000000000",
  48528=>"000000000",
  48529=>"000000000",
  48530=>"110100000",
  48531=>"110110111",
  48532=>"111111111",
  48533=>"011010000",
  48534=>"110111111",
  48535=>"101101001",
  48536=>"111111000",
  48537=>"000000000",
  48538=>"010110111",
  48539=>"101101000",
  48540=>"000010000",
  48541=>"001001000",
  48542=>"111111000",
  48543=>"000000000",
  48544=>"010000000",
  48545=>"001111001",
  48546=>"111100100",
  48547=>"011111111",
  48548=>"100100000",
  48549=>"000000000",
  48550=>"000100111",
  48551=>"011011110",
  48552=>"000000000",
  48553=>"000000000",
  48554=>"111001111",
  48555=>"111111111",
  48556=>"110110110",
  48557=>"000000000",
  48558=>"111100110",
  48559=>"000000000",
  48560=>"111111111",
  48561=>"000110000",
  48562=>"000001111",
  48563=>"000100101",
  48564=>"111111100",
  48565=>"100000100",
  48566=>"111101111",
  48567=>"000000000",
  48568=>"000001000",
  48569=>"000001111",
  48570=>"110010001",
  48571=>"111111011",
  48572=>"001001001",
  48573=>"000000100",
  48574=>"001000000",
  48575=>"000000000",
  48576=>"000000000",
  48577=>"111111111",
  48578=>"010111111",
  48579=>"011111111",
  48580=>"111101100",
  48581=>"111111101",
  48582=>"100111100",
  48583=>"111101001",
  48584=>"111100111",
  48585=>"000001001",
  48586=>"000000000",
  48587=>"100111111",
  48588=>"101000000",
  48589=>"110111011",
  48590=>"101001000",
  48591=>"000000000",
  48592=>"001010000",
  48593=>"111111111",
  48594=>"100101000",
  48595=>"000000000",
  48596=>"010110000",
  48597=>"011001111",
  48598=>"000000000",
  48599=>"000111111",
  48600=>"000110011",
  48601=>"000000000",
  48602=>"000000100",
  48603=>"110000000",
  48604=>"100111111",
  48605=>"000100000",
  48606=>"000000000",
  48607=>"111110110",
  48608=>"111100000",
  48609=>"000100111",
  48610=>"111111111",
  48611=>"100100100",
  48612=>"111111001",
  48613=>"111111111",
  48614=>"110100000",
  48615=>"000000000",
  48616=>"111111101",
  48617=>"111111111",
  48618=>"000001111",
  48619=>"111111101",
  48620=>"110111111",
  48621=>"000000000",
  48622=>"111111111",
  48623=>"000000000",
  48624=>"000000000",
  48625=>"000000000",
  48626=>"111110100",
  48627=>"000000000",
  48628=>"111111111",
  48629=>"000000000",
  48630=>"111111111",
  48631=>"111111000",
  48632=>"001111111",
  48633=>"100101001",
  48634=>"001000100",
  48635=>"000000000",
  48636=>"111111111",
  48637=>"110111111",
  48638=>"000000000",
  48639=>"000000000",
  48640=>"001000001",
  48641=>"000000000",
  48642=>"111111000",
  48643=>"000000000",
  48644=>"100110100",
  48645=>"100100100",
  48646=>"111111111",
  48647=>"111111111",
  48648=>"010111011",
  48649=>"000000000",
  48650=>"000000001",
  48651=>"111000000",
  48652=>"000110110",
  48653=>"110111110",
  48654=>"000100111",
  48655=>"001001000",
  48656=>"111111111",
  48657=>"000000000",
  48658=>"000111111",
  48659=>"111111110",
  48660=>"000000000",
  48661=>"111000111",
  48662=>"000111111",
  48663=>"000101100",
  48664=>"010000000",
  48665=>"111111111",
  48666=>"101001110",
  48667=>"001101000",
  48668=>"000000111",
  48669=>"111111111",
  48670=>"111111000",
  48671=>"111111111",
  48672=>"000000000",
  48673=>"111110110",
  48674=>"111111111",
  48675=>"111111001",
  48676=>"111111110",
  48677=>"000111000",
  48678=>"101001111",
  48679=>"101000001",
  48680=>"000001111",
  48681=>"000000000",
  48682=>"000000000",
  48683=>"000000111",
  48684=>"000000000",
  48685=>"000000000",
  48686=>"000000000",
  48687=>"011111111",
  48688=>"000000110",
  48689=>"100111001",
  48690=>"001101110",
  48691=>"111111111",
  48692=>"000111111",
  48693=>"111110100",
  48694=>"000000000",
  48695=>"000000110",
  48696=>"011000000",
  48697=>"100000110",
  48698=>"000000000",
  48699=>"110000000",
  48700=>"111100111",
  48701=>"111011000",
  48702=>"111111001",
  48703=>"111111111",
  48704=>"000000100",
  48705=>"100100100",
  48706=>"000000000",
  48707=>"111111111",
  48708=>"111111000",
  48709=>"000001111",
  48710=>"000000000",
  48711=>"011111000",
  48712=>"000001111",
  48713=>"111100110",
  48714=>"010111000",
  48715=>"111010000",
  48716=>"111111100",
  48717=>"111111000",
  48718=>"011010010",
  48719=>"110000000",
  48720=>"000111010",
  48721=>"000000000",
  48722=>"111100000",
  48723=>"111110110",
  48724=>"000000000",
  48725=>"111111111",
  48726=>"111000100",
  48727=>"000101111",
  48728=>"001000100",
  48729=>"111101111",
  48730=>"000000100",
  48731=>"100100000",
  48732=>"111111000",
  48733=>"001001001",
  48734=>"111101111",
  48735=>"000000000",
  48736=>"100000000",
  48737=>"111110111",
  48738=>"111111111",
  48739=>"001000000",
  48740=>"000000000",
  48741=>"101000000",
  48742=>"000100000",
  48743=>"100111111",
  48744=>"000000000",
  48745=>"111011000",
  48746=>"111000000",
  48747=>"001000001",
  48748=>"111111100",
  48749=>"100001001",
  48750=>"111111111",
  48751=>"010111111",
  48752=>"000000000",
  48753=>"111111000",
  48754=>"000111111",
  48755=>"110100100",
  48756=>"000000001",
  48757=>"000000100",
  48758=>"000000000",
  48759=>"000100000",
  48760=>"000111111",
  48761=>"000111111",
  48762=>"011000000",
  48763=>"000000000",
  48764=>"100110110",
  48765=>"000111111",
  48766=>"000000000",
  48767=>"000000000",
  48768=>"000000000",
  48769=>"010000111",
  48770=>"000000000",
  48771=>"111011001",
  48772=>"111001111",
  48773=>"000000101",
  48774=>"111111100",
  48775=>"010011011",
  48776=>"011000000",
  48777=>"000111111",
  48778=>"111111010",
  48779=>"000000000",
  48780=>"000010111",
  48781=>"100101111",
  48782=>"111111000",
  48783=>"111111111",
  48784=>"000000000",
  48785=>"110110000",
  48786=>"111111111",
  48787=>"111111111",
  48788=>"001111111",
  48789=>"000001111",
  48790=>"000110111",
  48791=>"111111111",
  48792=>"000001001",
  48793=>"111111110",
  48794=>"111111001",
  48795=>"000011000",
  48796=>"111111111",
  48797=>"100110000",
  48798=>"110101001",
  48799=>"000101101",
  48800=>"111110111",
  48801=>"001000000",
  48802=>"000000000",
  48803=>"111111010",
  48804=>"000000000",
  48805=>"111111000",
  48806=>"011001011",
  48807=>"111110110",
  48808=>"001111111",
  48809=>"000001000",
  48810=>"000111111",
  48811=>"000000001",
  48812=>"111111111",
  48813=>"111111110",
  48814=>"000000000",
  48815=>"111111000",
  48816=>"000000000",
  48817=>"111111011",
  48818=>"111111010",
  48819=>"010111110",
  48820=>"000000101",
  48821=>"000000111",
  48822=>"111111111",
  48823=>"000000000",
  48824=>"001001000",
  48825=>"000000000",
  48826=>"100000000",
  48827=>"000001001",
  48828=>"111111101",
  48829=>"111111110",
  48830=>"111111111",
  48831=>"001011111",
  48832=>"000000000",
  48833=>"000000001",
  48834=>"111111100",
  48835=>"000000111",
  48836=>"111111111",
  48837=>"111111000",
  48838=>"111000000",
  48839=>"011111111",
  48840=>"000000010",
  48841=>"000000000",
  48842=>"101100000",
  48843=>"000000000",
  48844=>"111111000",
  48845=>"000000000",
  48846=>"000000101",
  48847=>"100000000",
  48848=>"000001011",
  48849=>"000000000",
  48850=>"000000000",
  48851=>"100000000",
  48852=>"000000111",
  48853=>"000000110",
  48854=>"000011111",
  48855=>"011111000",
  48856=>"111110000",
  48857=>"110110111",
  48858=>"111111111",
  48859=>"111111111",
  48860=>"101100111",
  48861=>"111000000",
  48862=>"000000000",
  48863=>"111001000",
  48864=>"000000000",
  48865=>"110110111",
  48866=>"000000111",
  48867=>"000010000",
  48868=>"001001111",
  48869=>"101001000",
  48870=>"111111111",
  48871=>"111111110",
  48872=>"111111010",
  48873=>"000001000",
  48874=>"111110000",
  48875=>"010000000",
  48876=>"010011001",
  48877=>"000001111",
  48878=>"100110110",
  48879=>"000000000",
  48880=>"000000100",
  48881=>"011110111",
  48882=>"001111111",
  48883=>"001000000",
  48884=>"000000000",
  48885=>"000110011",
  48886=>"011111110",
  48887=>"110111101",
  48888=>"110110111",
  48889=>"000000000",
  48890=>"001011000",
  48891=>"111001000",
  48892=>"000000111",
  48893=>"100000110",
  48894=>"111000000",
  48895=>"111000111",
  48896=>"100000000",
  48897=>"100100111",
  48898=>"111111111",
  48899=>"111111111",
  48900=>"111101000",
  48901=>"111111100",
  48902=>"101111101",
  48903=>"000000100",
  48904=>"000000000",
  48905=>"111111111",
  48906=>"000001011",
  48907=>"000000000",
  48908=>"001001001",
  48909=>"000000000",
  48910=>"111100000",
  48911=>"111110000",
  48912=>"000000000",
  48913=>"000111111",
  48914=>"000000111",
  48915=>"111111000",
  48916=>"000000000",
  48917=>"000000000",
  48918=>"000000100",
  48919=>"111111000",
  48920=>"001000000",
  48921=>"000000000",
  48922=>"000001001",
  48923=>"000000000",
  48924=>"000000100",
  48925=>"111100111",
  48926=>"000000000",
  48927=>"011111111",
  48928=>"000000111",
  48929=>"000010011",
  48930=>"000000000",
  48931=>"000000111",
  48932=>"111111010",
  48933=>"111111111",
  48934=>"000101101",
  48935=>"000110011",
  48936=>"001001001",
  48937=>"111111000",
  48938=>"111110000",
  48939=>"111110000",
  48940=>"111111101",
  48941=>"010101001",
  48942=>"000110000",
  48943=>"111000001",
  48944=>"011111000",
  48945=>"000000110",
  48946=>"111111110",
  48947=>"111111111",
  48948=>"111101000",
  48949=>"011011101",
  48950=>"011001000",
  48951=>"000111101",
  48952=>"000111010",
  48953=>"000000000",
  48954=>"111111000",
  48955=>"101111010",
  48956=>"111111111",
  48957=>"111111000",
  48958=>"000000000",
  48959=>"111000000",
  48960=>"000011010",
  48961=>"001001010",
  48962=>"101111110",
  48963=>"000000000",
  48964=>"001000100",
  48965=>"110111111",
  48966=>"000101111",
  48967=>"001011000",
  48968=>"111011000",
  48969=>"000000000",
  48970=>"001000101",
  48971=>"010100101",
  48972=>"000110111",
  48973=>"111111111",
  48974=>"101000001",
  48975=>"111111111",
  48976=>"011001001",
  48977=>"111101001",
  48978=>"110111111",
  48979=>"001101000",
  48980=>"111001000",
  48981=>"001011001",
  48982=>"111111111",
  48983=>"000110100",
  48984=>"000000000",
  48985=>"000000000",
  48986=>"001111000",
  48987=>"111110111",
  48988=>"000000000",
  48989=>"000000000",
  48990=>"000000000",
  48991=>"001001011",
  48992=>"010111110",
  48993=>"111111111",
  48994=>"111111000",
  48995=>"111101111",
  48996=>"000000110",
  48997=>"000000111",
  48998=>"000000000",
  48999=>"011111111",
  49000=>"000000110",
  49001=>"000000000",
  49002=>"111111100",
  49003=>"010111100",
  49004=>"000000000",
  49005=>"000000000",
  49006=>"111111111",
  49007=>"000000000",
  49008=>"000000000",
  49009=>"000000000",
  49010=>"111111011",
  49011=>"100111111",
  49012=>"000000010",
  49013=>"111111000",
  49014=>"000000000",
  49015=>"000000000",
  49016=>"111111111",
  49017=>"011001001",
  49018=>"000000111",
  49019=>"111111000",
  49020=>"000000000",
  49021=>"000000111",
  49022=>"001001111",
  49023=>"111111111",
  49024=>"110111111",
  49025=>"111111000",
  49026=>"000000111",
  49027=>"100000011",
  49028=>"111000111",
  49029=>"111111111",
  49030=>"100100000",
  49031=>"111111100",
  49032=>"000000100",
  49033=>"111000000",
  49034=>"110100000",
  49035=>"111111110",
  49036=>"110000000",
  49037=>"000000100",
  49038=>"001001000",
  49039=>"000000000",
  49040=>"000000000",
  49041=>"111001111",
  49042=>"000000100",
  49043=>"111111001",
  49044=>"111111000",
  49045=>"000010010",
  49046=>"111011000",
  49047=>"000000000",
  49048=>"111111001",
  49049=>"000000000",
  49050=>"000000100",
  49051=>"001111110",
  49052=>"001001001",
  49053=>"111111000",
  49054=>"100111001",
  49055=>"111000000",
  49056=>"000111111",
  49057=>"011011001",
  49058=>"111100000",
  49059=>"000000011",
  49060=>"111111111",
  49061=>"110111011",
  49062=>"000000000",
  49063=>"110111111",
  49064=>"111111111",
  49065=>"000001111",
  49066=>"111111010",
  49067=>"100000000",
  49068=>"000000111",
  49069=>"111111111",
  49070=>"000100110",
  49071=>"111111111",
  49072=>"110000000",
  49073=>"111111111",
  49074=>"000000000",
  49075=>"000000001",
  49076=>"000000001",
  49077=>"111011111",
  49078=>"001000000",
  49079=>"000000111",
  49080=>"111111111",
  49081=>"001111110",
  49082=>"111111001",
  49083=>"000000111",
  49084=>"000011011",
  49085=>"111111110",
  49086=>"000000000",
  49087=>"100100000",
  49088=>"111111000",
  49089=>"110000010",
  49090=>"111111011",
  49091=>"000000001",
  49092=>"000000000",
  49093=>"101000101",
  49094=>"111011000",
  49095=>"000001000",
  49096=>"000000000",
  49097=>"100000000",
  49098=>"100000100",
  49099=>"000000111",
  49100=>"111110000",
  49101=>"000000110",
  49102=>"000000000",
  49103=>"000000011",
  49104=>"111010000",
  49105=>"111111111",
  49106=>"000000000",
  49107=>"111110110",
  49108=>"111111000",
  49109=>"011000000",
  49110=>"101001111",
  49111=>"000001001",
  49112=>"001001000",
  49113=>"110101111",
  49114=>"111011000",
  49115=>"111111000",
  49116=>"000010000",
  49117=>"111111110",
  49118=>"111111000",
  49119=>"111111111",
  49120=>"000000010",
  49121=>"000000111",
  49122=>"110111100",
  49123=>"111111000",
  49124=>"000000111",
  49125=>"000111111",
  49126=>"111000111",
  49127=>"111010011",
  49128=>"001001000",
  49129=>"110110110",
  49130=>"000000000",
  49131=>"000000111",
  49132=>"111111000",
  49133=>"000000000",
  49134=>"111101100",
  49135=>"110111111",
  49136=>"000000000",
  49137=>"110000000",
  49138=>"011000000",
  49139=>"111110110",
  49140=>"101000100",
  49141=>"000111111",
  49142=>"000000000",
  49143=>"111111000",
  49144=>"000001000",
  49145=>"001001001",
  49146=>"000000110",
  49147=>"111111111",
  49148=>"100000000",
  49149=>"111001001",
  49150=>"111111010",
  49151=>"001001111",
  49152=>"111111010",
  49153=>"000100100",
  49154=>"111111000",
  49155=>"000000111",
  49156=>"111111101",
  49157=>"000000110",
  49158=>"011000000",
  49159=>"111100111",
  49160=>"000000000",
  49161=>"110000000",
  49162=>"000100100",
  49163=>"111111000",
  49164=>"110100000",
  49165=>"111100100",
  49166=>"111000001",
  49167=>"001011001",
  49168=>"111011111",
  49169=>"111000000",
  49170=>"001111111",
  49171=>"011000000",
  49172=>"111110110",
  49173=>"000000111",
  49174=>"111111111",
  49175=>"111111111",
  49176=>"111100000",
  49177=>"100000111",
  49178=>"111111111",
  49179=>"111111111",
  49180=>"100000100",
  49181=>"000011111",
  49182=>"000000011",
  49183=>"111000000",
  49184=>"000111011",
  49185=>"111111111",
  49186=>"000000111",
  49187=>"111111000",
  49188=>"111111010",
  49189=>"101000000",
  49190=>"110111110",
  49191=>"000000000",
  49192=>"000100101",
  49193=>"011111011",
  49194=>"000000000",
  49195=>"001110000",
  49196=>"111001111",
  49197=>"000000000",
  49198=>"100000000",
  49199=>"111111111",
  49200=>"100000000",
  49201=>"000000011",
  49202=>"100100000",
  49203=>"111101000",
  49204=>"100111011",
  49205=>"000000111",
  49206=>"001000111",
  49207=>"000000011",
  49208=>"100111111",
  49209=>"111010000",
  49210=>"001011111",
  49211=>"001000000",
  49212=>"111000000",
  49213=>"111110000",
  49214=>"110110000",
  49215=>"111111111",
  49216=>"111110110",
  49217=>"110000000",
  49218=>"000001000",
  49219=>"101000111",
  49220=>"000000111",
  49221=>"001111111",
  49222=>"000000000",
  49223=>"000000000",
  49224=>"000000110",
  49225=>"111111000",
  49226=>"001000111",
  49227=>"111111111",
  49228=>"111111110",
  49229=>"111000000",
  49230=>"000000100",
  49231=>"111111000",
  49232=>"000000000",
  49233=>"111000011",
  49234=>"111111000",
  49235=>"111011111",
  49236=>"000100111",
  49237=>"111100100",
  49238=>"111100000",
  49239=>"000111111",
  49240=>"110100110",
  49241=>"111111101",
  49242=>"111111101",
  49243=>"000110000",
  49244=>"000100000",
  49245=>"000000000",
  49246=>"001100100",
  49247=>"110111111",
  49248=>"000000010",
  49249=>"111111111",
  49250=>"111111000",
  49251=>"111000011",
  49252=>"110110000",
  49253=>"010111000",
  49254=>"000111111",
  49255=>"001001111",
  49256=>"111011101",
  49257=>"000000111",
  49258=>"011000111",
  49259=>"111111010",
  49260=>"111011000",
  49261=>"001000000",
  49262=>"001000000",
  49263=>"111001011",
  49264=>"111000000",
  49265=>"000111111",
  49266=>"000111011",
  49267=>"000000000",
  49268=>"000000000",
  49269=>"001011000",
  49270=>"000000100",
  49271=>"111101000",
  49272=>"110111110",
  49273=>"100100101",
  49274=>"000000000",
  49275=>"000000000",
  49276=>"111111011",
  49277=>"000111111",
  49278=>"000000110",
  49279=>"111111000",
  49280=>"110000000",
  49281=>"001000000",
  49282=>"000000111",
  49283=>"111100000",
  49284=>"000001001",
  49285=>"111111000",
  49286=>"111111111",
  49287=>"000101111",
  49288=>"101100111",
  49289=>"111000111",
  49290=>"000000000",
  49291=>"000000000",
  49292=>"111000000",
  49293=>"001111001",
  49294=>"001000000",
  49295=>"111010000",
  49296=>"100101111",
  49297=>"100000000",
  49298=>"000000100",
  49299=>"001000111",
  49300=>"100000000",
  49301=>"000000111",
  49302=>"000000100",
  49303=>"000000000",
  49304=>"100101100",
  49305=>"111100000",
  49306=>"111111000",
  49307=>"111001000",
  49308=>"111111111",
  49309=>"000000101",
  49310=>"001111111",
  49311=>"000111111",
  49312=>"111111111",
  49313=>"101111111",
  49314=>"000000111",
  49315=>"011000100",
  49316=>"111111000",
  49317=>"000010111",
  49318=>"100000010",
  49319=>"000111111",
  49320=>"000100110",
  49321=>"000101001",
  49322=>"000000111",
  49323=>"110000011",
  49324=>"111110010",
  49325=>"101111111",
  49326=>"110001101",
  49327=>"001000000",
  49328=>"101110111",
  49329=>"110000001",
  49330=>"110111111",
  49331=>"000000000",
  49332=>"001000111",
  49333=>"110110010",
  49334=>"000111111",
  49335=>"111111110",
  49336=>"000000000",
  49337=>"111111111",
  49338=>"110000000",
  49339=>"111111111",
  49340=>"000000011",
  49341=>"000000010",
  49342=>"000000100",
  49343=>"010000000",
  49344=>"111111000",
  49345=>"000000111",
  49346=>"100000000",
  49347=>"000000000",
  49348=>"001111111",
  49349=>"111111011",
  49350=>"111111000",
  49351=>"100011011",
  49352=>"000000000",
  49353=>"000000111",
  49354=>"111101001",
  49355=>"000000000",
  49356=>"010000000",
  49357=>"001001011",
  49358=>"111111000",
  49359=>"000000000",
  49360=>"111111111",
  49361=>"111011011",
  49362=>"000100000",
  49363=>"000000111",
  49364=>"001001111",
  49365=>"111110000",
  49366=>"111000000",
  49367=>"100000000",
  49368=>"100000111",
  49369=>"001000111",
  49370=>"111000001",
  49371=>"000000000",
  49372=>"111111111",
  49373=>"000000000",
  49374=>"000011111",
  49375=>"001111111",
  49376=>"000000000",
  49377=>"010000000",
  49378=>"000000111",
  49379=>"111110110",
  49380=>"000000000",
  49381=>"000000011",
  49382=>"111011000",
  49383=>"111000001",
  49384=>"000000111",
  49385=>"011111001",
  49386=>"111111001",
  49387=>"111000000",
  49388=>"111111111",
  49389=>"011111101",
  49390=>"111110110",
  49391=>"001100000",
  49392=>"011001000",
  49393=>"111110100",
  49394=>"011111111",
  49395=>"100111111",
  49396=>"000000111",
  49397=>"000100101",
  49398=>"000110100",
  49399=>"001000000",
  49400=>"000000000",
  49401=>"000111111",
  49402=>"111110000",
  49403=>"111111010",
  49404=>"110111111",
  49405=>"011001000",
  49406=>"000000111",
  49407=>"000000000",
  49408=>"111000000",
  49409=>"001000001",
  49410=>"000000000",
  49411=>"111110000",
  49412=>"000000111",
  49413=>"110100111",
  49414=>"111111111",
  49415=>"100000000",
  49416=>"111111000",
  49417=>"000000000",
  49418=>"001000100",
  49419=>"111111111",
  49420=>"100000000",
  49421=>"000001111",
  49422=>"100000000",
  49423=>"000000011",
  49424=>"000000000",
  49425=>"100111111",
  49426=>"000000000",
  49427=>"000000100",
  49428=>"001001111",
  49429=>"000000111",
  49430=>"000000001",
  49431=>"000000000",
  49432=>"111111000",
  49433=>"100110100",
  49434=>"000101111",
  49435=>"111000111",
  49436=>"111111000",
  49437=>"111000111",
  49438=>"000000001",
  49439=>"000111111",
  49440=>"111111000",
  49441=>"111111011",
  49442=>"111001000",
  49443=>"000000111",
  49444=>"111111000",
  49445=>"000000111",
  49446=>"101101111",
  49447=>"111111001",
  49448=>"111101111",
  49449=>"111000000",
  49450=>"000000000",
  49451=>"000111110",
  49452=>"111100000",
  49453=>"101001001",
  49454=>"000000000",
  49455=>"000000000",
  49456=>"000000000",
  49457=>"111110000",
  49458=>"111111000",
  49459=>"000000000",
  49460=>"001001000",
  49461=>"000000111",
  49462=>"000111101",
  49463=>"111000000",
  49464=>"111111011",
  49465=>"111100111",
  49466=>"000110000",
  49467=>"000000111",
  49468=>"000000111",
  49469=>"000000001",
  49470=>"100000000",
  49471=>"011111111",
  49472=>"111000100",
  49473=>"000000000",
  49474=>"111110000",
  49475=>"110111001",
  49476=>"001000000",
  49477=>"000000111",
  49478=>"111111111",
  49479=>"011000000",
  49480=>"111100000",
  49481=>"000000000",
  49482=>"001000111",
  49483=>"000011111",
  49484=>"001000011",
  49485=>"101001111",
  49486=>"001000110",
  49487=>"000111110",
  49488=>"000000111",
  49489=>"000000101",
  49490=>"111111000",
  49491=>"000000111",
  49492=>"010110111",
  49493=>"011011001",
  49494=>"000001011",
  49495=>"000100111",
  49496=>"000000111",
  49497=>"111110010",
  49498=>"100000000",
  49499=>"000000000",
  49500=>"010111000",
  49501=>"000100000",
  49502=>"100100101",
  49503=>"100000000",
  49504=>"111111000",
  49505=>"000000000",
  49506=>"000100111",
  49507=>"111111000",
  49508=>"111111111",
  49509=>"000000000",
  49510=>"000000000",
  49511=>"111110110",
  49512=>"000100111",
  49513=>"111111111",
  49514=>"111010000",
  49515=>"111111111",
  49516=>"000001001",
  49517=>"111111101",
  49518=>"010010000",
  49519=>"111111101",
  49520=>"100000000",
  49521=>"000110000",
  49522=>"000000001",
  49523=>"000001001",
  49524=>"010111111",
  49525=>"000000001",
  49526=>"100000000",
  49527=>"000000111",
  49528=>"101111011",
  49529=>"000000100",
  49530=>"000001101",
  49531=>"111111000",
  49532=>"111000000",
  49533=>"111111111",
  49534=>"000000001",
  49535=>"111001111",
  49536=>"111111111",
  49537=>"000000000",
  49538=>"110111111",
  49539=>"000000000",
  49540=>"000000111",
  49541=>"111100000",
  49542=>"111000000",
  49543=>"111111000",
  49544=>"000000111",
  49545=>"000000010",
  49546=>"111111011",
  49547=>"111111010",
  49548=>"111111100",
  49549=>"111111000",
  49550=>"110100000",
  49551=>"000011000",
  49552=>"000000000",
  49553=>"110111111",
  49554=>"110111001",
  49555=>"111111111",
  49556=>"011001101",
  49557=>"000000000",
  49558=>"111001001",
  49559=>"011001001",
  49560=>"000000011",
  49561=>"000010110",
  49562=>"000001111",
  49563=>"000111111",
  49564=>"011011000",
  49565=>"111111001",
  49566=>"001000001",
  49567=>"111111111",
  49568=>"011110000",
  49569=>"110111011",
  49570=>"111111000",
  49571=>"000001111",
  49572=>"101111101",
  49573=>"011000000",
  49574=>"111111110",
  49575=>"110000110",
  49576=>"000101111",
  49577=>"111111111",
  49578=>"011101111",
  49579=>"000000101",
  49580=>"000000000",
  49581=>"110000111",
  49582=>"010000000",
  49583=>"000000111",
  49584=>"011001000",
  49585=>"000000000",
  49586=>"000000000",
  49587=>"000000000",
  49588=>"100111110",
  49589=>"000001111",
  49590=>"000000000",
  49591=>"111001000",
  49592=>"101000000",
  49593=>"111111000",
  49594=>"000111111",
  49595=>"110111111",
  49596=>"011011111",
  49597=>"011000000",
  49598=>"011101001",
  49599=>"100000000",
  49600=>"000000111",
  49601=>"110000000",
  49602=>"111110110",
  49603=>"110110000",
  49604=>"111110000",
  49605=>"000000000",
  49606=>"111000000",
  49607=>"000000011",
  49608=>"001000000",
  49609=>"001000000",
  49610=>"000000000",
  49611=>"000000010",
  49612=>"111000000",
  49613=>"110111010",
  49614=>"111111011",
  49615=>"001000111",
  49616=>"101101001",
  49617=>"000001111",
  49618=>"011011000",
  49619=>"111111010",
  49620=>"000000111",
  49621=>"111000000",
  49622=>"101110100",
  49623=>"001001001",
  49624=>"100000000",
  49625=>"111101000",
  49626=>"110010010",
  49627=>"000000100",
  49628=>"111001011",
  49629=>"111111000",
  49630=>"111010000",
  49631=>"001001011",
  49632=>"110000001",
  49633=>"000000011",
  49634=>"000000010",
  49635=>"000000101",
  49636=>"111101000",
  49637=>"010111010",
  49638=>"000000000",
  49639=>"000000000",
  49640=>"111101001",
  49641=>"111111111",
  49642=>"100100111",
  49643=>"111111000",
  49644=>"111101111",
  49645=>"110100111",
  49646=>"000000000",
  49647=>"000000000",
  49648=>"100000000",
  49649=>"001001000",
  49650=>"100100100",
  49651=>"000001001",
  49652=>"111001000",
  49653=>"100101111",
  49654=>"001000100",
  49655=>"000111000",
  49656=>"111000000",
  49657=>"001001010",
  49658=>"000001000",
  49659=>"000000000",
  49660=>"110000000",
  49661=>"000000111",
  49662=>"111001111",
  49663=>"000000000",
  49664=>"111010011",
  49665=>"111011111",
  49666=>"101101111",
  49667=>"000000000",
  49668=>"001000111",
  49669=>"011011001",
  49670=>"000000000",
  49671=>"111111111",
  49672=>"000000000",
  49673=>"111111000",
  49674=>"100000000",
  49675=>"000000111",
  49676=>"000110111",
  49677=>"011000011",
  49678=>"000000000",
  49679=>"001000000",
  49680=>"111001100",
  49681=>"000000111",
  49682=>"000000011",
  49683=>"000000000",
  49684=>"000000000",
  49685=>"000000000",
  49686=>"001011001",
  49687=>"111111111",
  49688=>"000000000",
  49689=>"000110111",
  49690=>"111111111",
  49691=>"111111110",
  49692=>"110111110",
  49693=>"011111101",
  49694=>"000001111",
  49695=>"000000111",
  49696=>"000000000",
  49697=>"100111111",
  49698=>"111010100",
  49699=>"111111111",
  49700=>"111111111",
  49701=>"110110111",
  49702=>"001000000",
  49703=>"100100000",
  49704=>"110011111",
  49705=>"000111111",
  49706=>"111111111",
  49707=>"011001100",
  49708=>"111111001",
  49709=>"001111111",
  49710=>"000111111",
  49711=>"001111000",
  49712=>"000001111",
  49713=>"000000000",
  49714=>"110000000",
  49715=>"111000000",
  49716=>"100111111",
  49717=>"000000000",
  49718=>"001011111",
  49719=>"100100100",
  49720=>"111001000",
  49721=>"111111111",
  49722=>"000000000",
  49723=>"100110000",
  49724=>"111111110",
  49725=>"101100100",
  49726=>"010111000",
  49727=>"101000000",
  49728=>"111111111",
  49729=>"000000000",
  49730=>"000000100",
  49731=>"111111011",
  49732=>"000100110",
  49733=>"000000001",
  49734=>"000010000",
  49735=>"011000000",
  49736=>"100100111",
  49737=>"101101111",
  49738=>"011000000",
  49739=>"110000111",
  49740=>"111111111",
  49741=>"000000111",
  49742=>"100000000",
  49743=>"000000000",
  49744=>"011000000",
  49745=>"111110110",
  49746=>"100100000",
  49747=>"000000110",
  49748=>"000000100",
  49749=>"000000101",
  49750=>"000000000",
  49751=>"000111111",
  49752=>"000000000",
  49753=>"000000000",
  49754=>"000000001",
  49755=>"000000000",
  49756=>"111111111",
  49757=>"000011011",
  49758=>"100010011",
  49759=>"000000000",
  49760=>"101111011",
  49761=>"111111110",
  49762=>"111111111",
  49763=>"000000011",
  49764=>"001011111",
  49765=>"000000000",
  49766=>"111111000",
  49767=>"011011111",
  49768=>"110100000",
  49769=>"001001001",
  49770=>"110110111",
  49771=>"000000001",
  49772=>"011001000",
  49773=>"000000000",
  49774=>"111100110",
  49775=>"000001000",
  49776=>"000110111",
  49777=>"010000111",
  49778=>"000111111",
  49779=>"111111111",
  49780=>"000000000",
  49781=>"111111111",
  49782=>"101100100",
  49783=>"000000000",
  49784=>"111111111",
  49785=>"011001001",
  49786=>"100000000",
  49787=>"000000010",
  49788=>"110010000",
  49789=>"000000001",
  49790=>"100000000",
  49791=>"000000000",
  49792=>"100000100",
  49793=>"111111111",
  49794=>"111110000",
  49795=>"011111000",
  49796=>"001001000",
  49797=>"000000000",
  49798=>"000000000",
  49799=>"000000000",
  49800=>"111111000",
  49801=>"000000000",
  49802=>"000001000",
  49803=>"111111011",
  49804=>"111111101",
  49805=>"000000000",
  49806=>"111111111",
  49807=>"000111111",
  49808=>"111111011",
  49809=>"100110110",
  49810=>"000111100",
  49811=>"111111111",
  49812=>"111111001",
  49813=>"000100111",
  49814=>"111000000",
  49815=>"011111111",
  49816=>"111111110",
  49817=>"011000000",
  49818=>"001000110",
  49819=>"111111111",
  49820=>"000000000",
  49821=>"110111000",
  49822=>"111011001",
  49823=>"000000001",
  49824=>"111100000",
  49825=>"000011110",
  49826=>"000000000",
  49827=>"111100100",
  49828=>"000000000",
  49829=>"000000000",
  49830=>"111101110",
  49831=>"001111001",
  49832=>"111111111",
  49833=>"011111111",
  49834=>"000000000",
  49835=>"100100110",
  49836=>"111011000",
  49837=>"110110000",
  49838=>"000000000",
  49839=>"000011001",
  49840=>"000001000",
  49841=>"101011000",
  49842=>"001101110",
  49843=>"111101000",
  49844=>"000000000",
  49845=>"000000011",
  49846=>"000000000",
  49847=>"111111101",
  49848=>"001010010",
  49849=>"111111111",
  49850=>"000000000",
  49851=>"000000000",
  49852=>"000000011",
  49853=>"001001000",
  49854=>"100100110",
  49855=>"000110111",
  49856=>"000000110",
  49857=>"111111110",
  49858=>"100001001",
  49859=>"111111010",
  49860=>"000000000",
  49861=>"010011011",
  49862=>"000000000",
  49863=>"000000000",
  49864=>"111111111",
  49865=>"111111111",
  49866=>"000011111",
  49867=>"000011001",
  49868=>"000000110",
  49869=>"000100101",
  49870=>"000000000",
  49871=>"000000000",
  49872=>"001000000",
  49873=>"111111111",
  49874=>"001001010",
  49875=>"111111111",
  49876=>"000000000",
  49877=>"111000001",
  49878=>"000000000",
  49879=>"111110110",
  49880=>"000000111",
  49881=>"111000000",
  49882=>"000000000",
  49883=>"011011011",
  49884=>"111010000",
  49885=>"111111111",
  49886=>"000000000",
  49887=>"010000000",
  49888=>"000000000",
  49889=>"000000111",
  49890=>"000000000",
  49891=>"011000000",
  49892=>"111111011",
  49893=>"000000000",
  49894=>"000000000",
  49895=>"111111111",
  49896=>"111111000",
  49897=>"110000010",
  49898=>"111100000",
  49899=>"000000000",
  49900=>"001001000",
  49901=>"011011000",
  49902=>"111001000",
  49903=>"111000000",
  49904=>"111111111",
  49905=>"100000110",
  49906=>"111100000",
  49907=>"000000011",
  49908=>"000111011",
  49909=>"010000000",
  49910=>"111110110",
  49911=>"001001111",
  49912=>"111111110",
  49913=>"011111001",
  49914=>"001000111",
  49915=>"000000111",
  49916=>"110111110",
  49917=>"001000100",
  49918=>"011010111",
  49919=>"111000000",
  49920=>"000000000",
  49921=>"001011010",
  49922=>"111111111",
  49923=>"001111111",
  49924=>"110110100",
  49925=>"110100000",
  49926=>"111111100",
  49927=>"110110100",
  49928=>"001011111",
  49929=>"110000000",
  49930=>"111111111",
  49931=>"000000000",
  49932=>"111111000",
  49933=>"000000000",
  49934=>"111111111",
  49935=>"101111100",
  49936=>"000000010",
  49937=>"111111111",
  49938=>"100100111",
  49939=>"111111011",
  49940=>"000000000",
  49941=>"010111111",
  49942=>"000110000",
  49943=>"000000000",
  49944=>"111100111",
  49945=>"000001111",
  49946=>"000000111",
  49947=>"011000000",
  49948=>"001001011",
  49949=>"111000011",
  49950=>"111111111",
  49951=>"000000110",
  49952=>"111111011",
  49953=>"000000000",
  49954=>"001000010",
  49955=>"111111111",
  49956=>"001000000",
  49957=>"111111000",
  49958=>"000001000",
  49959=>"000011110",
  49960=>"011111000",
  49961=>"000001111",
  49962=>"100000001",
  49963=>"101001000",
  49964=>"000000000",
  49965=>"111111110",
  49966=>"000000000",
  49967=>"000000000",
  49968=>"111011111",
  49969=>"100000000",
  49970=>"000000000",
  49971=>"011111111",
  49972=>"000000000",
  49973=>"011111001",
  49974=>"100100000",
  49975=>"000000000",
  49976=>"101101000",
  49977=>"100101111",
  49978=>"111111001",
  49979=>"010000000",
  49980=>"111110110",
  49981=>"000000000",
  49982=>"111111111",
  49983=>"111110000",
  49984=>"111111111",
  49985=>"000011001",
  49986=>"000001101",
  49987=>"000111111",
  49988=>"000000110",
  49989=>"000011001",
  49990=>"001111111",
  49991=>"111111100",
  49992=>"111011001",
  49993=>"111111111",
  49994=>"111011000",
  49995=>"111111110",
  49996=>"001001000",
  49997=>"011000000",
  49998=>"000000000",
  49999=>"111111111",
  50000=>"000100111",
  50001=>"000000110",
  50002=>"110110000",
  50003=>"001101111",
  50004=>"101000111",
  50005=>"011011011",
  50006=>"111111010",
  50007=>"111110111",
  50008=>"111111110",
  50009=>"111000000",
  50010=>"001000110",
  50011=>"111011111",
  50012=>"010111000",
  50013=>"000111110",
  50014=>"111111011",
  50015=>"000000000",
  50016=>"000000000",
  50017=>"000101111",
  50018=>"000000111",
  50019=>"000011111",
  50020=>"111110110",
  50021=>"111111111",
  50022=>"000101111",
  50023=>"111110000",
  50024=>"011111011",
  50025=>"111011111",
  50026=>"111111100",
  50027=>"100101111",
  50028=>"001011000",
  50029=>"000101001",
  50030=>"000000000",
  50031=>"000000010",
  50032=>"111111111",
  50033=>"111001011",
  50034=>"111111011",
  50035=>"000000001",
  50036=>"111111100",
  50037=>"101111111",
  50038=>"000001001",
  50039=>"000000111",
  50040=>"111111000",
  50041=>"000100100",
  50042=>"000010010",
  50043=>"111111110",
  50044=>"000000000",
  50045=>"000000110",
  50046=>"000101111",
  50047=>"101111111",
  50048=>"100100111",
  50049=>"010010000",
  50050=>"000000000",
  50051=>"111111111",
  50052=>"000000000",
  50053=>"111111111",
  50054=>"111011000",
  50055=>"000000000",
  50056=>"000000000",
  50057=>"010111101",
  50058=>"011000000",
  50059=>"000100100",
  50060=>"101001101",
  50061=>"000100111",
  50062=>"000000000",
  50063=>"000011111",
  50064=>"000111111",
  50065=>"111111111",
  50066=>"111111111",
  50067=>"111111111",
  50068=>"100101000",
  50069=>"000000000",
  50070=>"000000000",
  50071=>"001000100",
  50072=>"111111111",
  50073=>"100000000",
  50074=>"000000110",
  50075=>"000000000",
  50076=>"000000000",
  50077=>"011111110",
  50078=>"000000000",
  50079=>"000000110",
  50080=>"001000000",
  50081=>"110111110",
  50082=>"000011110",
  50083=>"000000000",
  50084=>"111111111",
  50085=>"000000000",
  50086=>"101001001",
  50087=>"000000101",
  50088=>"001001000",
  50089=>"010111111",
  50090=>"001111001",
  50091=>"000000000",
  50092=>"000000000",
  50093=>"000010000",
  50094=>"011111100",
  50095=>"101111111",
  50096=>"111111111",
  50097=>"000100100",
  50098=>"100100000",
  50099=>"000000001",
  50100=>"000011111",
  50101=>"011011000",
  50102=>"111111111",
  50103=>"000111110",
  50104=>"001000000",
  50105=>"111011011",
  50106=>"000000111",
  50107=>"111111000",
  50108=>"100100000",
  50109=>"001110111",
  50110=>"000000000",
  50111=>"001111111",
  50112=>"011000000",
  50113=>"111111111",
  50114=>"000001011",
  50115=>"111111110",
  50116=>"111111100",
  50117=>"111111001",
  50118=>"111111111",
  50119=>"000000000",
  50120=>"010111110",
  50121=>"000000000",
  50122=>"111001001",
  50123=>"000000101",
  50124=>"000000000",
  50125=>"111111011",
  50126=>"011000000",
  50127=>"000000000",
  50128=>"101001000",
  50129=>"001011011",
  50130=>"011011111",
  50131=>"111111111",
  50132=>"111111111",
  50133=>"111111111",
  50134=>"000000001",
  50135=>"111111111",
  50136=>"000011001",
  50137=>"111101000",
  50138=>"111111110",
  50139=>"111111000",
  50140=>"100111111",
  50141=>"111111111",
  50142=>"000000011",
  50143=>"011111110",
  50144=>"000000011",
  50145=>"111111111",
  50146=>"000000000",
  50147=>"111111000",
  50148=>"101111111",
  50149=>"111000000",
  50150=>"010010000",
  50151=>"111000111",
  50152=>"001001000",
  50153=>"111111111",
  50154=>"000000000",
  50155=>"111011011",
  50156=>"000100000",
  50157=>"110111111",
  50158=>"011010010",
  50159=>"001111000",
  50160=>"000000000",
  50161=>"000000000",
  50162=>"100000111",
  50163=>"000001001",
  50164=>"000000000",
  50165=>"111111111",
  50166=>"000000100",
  50167=>"000100000",
  50168=>"000000000",
  50169=>"000000001",
  50170=>"000000000",
  50171=>"000000111",
  50172=>"111111000",
  50173=>"001111100",
  50174=>"000000011",
  50175=>"001111111",
  50176=>"010110110",
  50177=>"001000001",
  50178=>"000000010",
  50179=>"011011111",
  50180=>"111111111",
  50181=>"111001001",
  50182=>"100000000",
  50183=>"000000000",
  50184=>"111001011",
  50185=>"101001111",
  50186=>"111111111",
  50187=>"111111111",
  50188=>"001001001",
  50189=>"111000000",
  50190=>"111111111",
  50191=>"000000000",
  50192=>"111111111",
  50193=>"111000111",
  50194=>"111111111",
  50195=>"111000101",
  50196=>"000100111",
  50197=>"000000111",
  50198=>"000000000",
  50199=>"111011011",
  50200=>"111111111",
  50201=>"111111111",
  50202=>"000000000",
  50203=>"100100100",
  50204=>"000000000",
  50205=>"111111111",
  50206=>"001011100",
  50207=>"001011011",
  50208=>"001001000",
  50209=>"111111111",
  50210=>"000000000",
  50211=>"000011011",
  50212=>"111110100",
  50213=>"000000000",
  50214=>"011111111",
  50215=>"000001001",
  50216=>"111111101",
  50217=>"000111011",
  50218=>"111111111",
  50219=>"000000000",
  50220=>"111111011",
  50221=>"011001000",
  50222=>"111010000",
  50223=>"110111111",
  50224=>"111111110",
  50225=>"111111000",
  50226=>"000000000",
  50227=>"000000100",
  50228=>"000000000",
  50229=>"001001000",
  50230=>"000001001",
  50231=>"000000011",
  50232=>"000110110",
  50233=>"000110110",
  50234=>"000111111",
  50235=>"011000000",
  50236=>"001111111",
  50237=>"111111111",
  50238=>"111110111",
  50239=>"001000000",
  50240=>"001001000",
  50241=>"000000001",
  50242=>"001011111",
  50243=>"111111001",
  50244=>"110110110",
  50245=>"111111111",
  50246=>"110111010",
  50247=>"111111111",
  50248=>"011111011",
  50249=>"000000000",
  50250=>"110111111",
  50251=>"001011000",
  50252=>"110110000",
  50253=>"001001011",
  50254=>"111111111",
  50255=>"001111001",
  50256=>"001011001",
  50257=>"111110010",
  50258=>"010011000",
  50259=>"011011001",
  50260=>"101001001",
  50261=>"000000000",
  50262=>"000010111",
  50263=>"110111111",
  50264=>"000000000",
  50265=>"000000000",
  50266=>"000000010",
  50267=>"100110000",
  50268=>"000000000",
  50269=>"000000000",
  50270=>"011111111",
  50271=>"000000000",
  50272=>"000000110",
  50273=>"111111111",
  50274=>"101000000",
  50275=>"110000000",
  50276=>"010000000",
  50277=>"111111111",
  50278=>"000000000",
  50279=>"111111001",
  50280=>"011000000",
  50281=>"000100111",
  50282=>"111111111",
  50283=>"000000000",
  50284=>"010011011",
  50285=>"111111111",
  50286=>"111111111",
  50287=>"110110010",
  50288=>"000110000",
  50289=>"000001000",
  50290=>"001001101",
  50291=>"000100010",
  50292=>"110100000",
  50293=>"100000000",
  50294=>"010111111",
  50295=>"000000000",
  50296=>"111101000",
  50297=>"001011011",
  50298=>"111000000",
  50299=>"000000000",
  50300=>"010110110",
  50301=>"000000001",
  50302=>"100000000",
  50303=>"011000101",
  50304=>"111111111",
  50305=>"111111111",
  50306=>"011000000",
  50307=>"110111110",
  50308=>"111100111",
  50309=>"111111101",
  50310=>"000000000",
  50311=>"000000000",
  50312=>"000000011",
  50313=>"000000011",
  50314=>"111111000",
  50315=>"001111111",
  50316=>"000000011",
  50317=>"000010000",
  50318=>"111011000",
  50319=>"111001100",
  50320=>"000000000",
  50321=>"111110111",
  50322=>"010111010",
  50323=>"000001001",
  50324=>"101101110",
  50325=>"111111111",
  50326=>"000010011",
  50327=>"011000000",
  50328=>"001001001",
  50329=>"001001111",
  50330=>"101000100",
  50331=>"000000001",
  50332=>"111110000",
  50333=>"101101100",
  50334=>"111111111",
  50335=>"111111101",
  50336=>"000000000",
  50337=>"000000000",
  50338=>"000000000",
  50339=>"000000101",
  50340=>"001001000",
  50341=>"111111111",
  50342=>"000000000",
  50343=>"001100110",
  50344=>"000010011",
  50345=>"101001001",
  50346=>"111101111",
  50347=>"001111111",
  50348=>"000000000",
  50349=>"001011000",
  50350=>"000111111",
  50351=>"000000010",
  50352=>"110110000",
  50353=>"111111010",
  50354=>"000000000",
  50355=>"111000000",
  50356=>"110110111",
  50357=>"000000000",
  50358=>"011111011",
  50359=>"111111111",
  50360=>"000011000",
  50361=>"111011111",
  50362=>"101101001",
  50363=>"000000001",
  50364=>"000000000",
  50365=>"111111111",
  50366=>"000000010",
  50367=>"100110111",
  50368=>"000000000",
  50369=>"110111011",
  50370=>"111111111",
  50371=>"000000000",
  50372=>"111111111",
  50373=>"001000000",
  50374=>"111101111",
  50375=>"000101111",
  50376=>"110100000",
  50377=>"111111110",
  50378=>"001000001",
  50379=>"111111000",
  50380=>"000100100",
  50381=>"111111110",
  50382=>"111111001",
  50383=>"000000101",
  50384=>"100111111",
  50385=>"000000001",
  50386=>"000000011",
  50387=>"000000001",
  50388=>"000000000",
  50389=>"001101100",
  50390=>"000111111",
  50391=>"001000000",
  50392=>"001001000",
  50393=>"010110111",
  50394=>"000000000",
  50395=>"111000000",
  50396=>"000110111",
  50397=>"000000111",
  50398=>"001000111",
  50399=>"000000001",
  50400=>"000000000",
  50401=>"000000000",
  50402=>"111111111",
  50403=>"000011111",
  50404=>"000000111",
  50405=>"111011000",
  50406=>"111010000",
  50407=>"111111111",
  50408=>"000110111",
  50409=>"111111011",
  50410=>"111001001",
  50411=>"111111001",
  50412=>"011011000",
  50413=>"011011111",
  50414=>"011111111",
  50415=>"000000000",
  50416=>"110110111",
  50417=>"010111111",
  50418=>"110110111",
  50419=>"000000000",
  50420=>"110110000",
  50421=>"000011011",
  50422=>"101111111",
  50423=>"000000000",
  50424=>"000000111",
  50425=>"111111101",
  50426=>"000000000",
  50427=>"110010010",
  50428=>"111011111",
  50429=>"000000000",
  50430=>"001111111",
  50431=>"111110010",
  50432=>"000000000",
  50433=>"001011000",
  50434=>"111111111",
  50435=>"000000000",
  50436=>"100000000",
  50437=>"000100111",
  50438=>"110111011",
  50439=>"011011110",
  50440=>"111110110",
  50441=>"000100111",
  50442=>"111111001",
  50443=>"110111111",
  50444=>"000000000",
  50445=>"011111111",
  50446=>"111111111",
  50447=>"011111110",
  50448=>"110111101",
  50449=>"000001111",
  50450=>"000000111",
  50451=>"010110010",
  50452=>"111001111",
  50453=>"001000000",
  50454=>"000000001",
  50455=>"110111000",
  50456=>"111111111",
  50457=>"000000011",
  50458=>"000000000",
  50459=>"111000000",
  50460=>"110100000",
  50461=>"000000000",
  50462=>"000000000",
  50463=>"111111111",
  50464=>"111110000",
  50465=>"110111111",
  50466=>"111110010",
  50467=>"000100000",
  50468=>"101111111",
  50469=>"100110001",
  50470=>"000100110",
  50471=>"001000000",
  50472=>"111011111",
  50473=>"001001001",
  50474=>"001000000",
  50475=>"000011111",
  50476=>"111100000",
  50477=>"011001000",
  50478=>"110110110",
  50479=>"000000000",
  50480=>"001001001",
  50481=>"111111111",
  50482=>"100000001",
  50483=>"111111111",
  50484=>"010000110",
  50485=>"000001101",
  50486=>"000011000",
  50487=>"000101111",
  50488=>"001001011",
  50489=>"000001000",
  50490=>"000000011",
  50491=>"000000011",
  50492=>"000000000",
  50493=>"010000000",
  50494=>"001111101",
  50495=>"100100000",
  50496=>"000011111",
  50497=>"000111000",
  50498=>"001001000",
  50499=>"000000111",
  50500=>"111110000",
  50501=>"000010010",
  50502=>"111000000",
  50503=>"000000111",
  50504=>"111111000",
  50505=>"111000000",
  50506=>"001000000",
  50507=>"111110110",
  50508=>"000000001",
  50509=>"110000111",
  50510=>"111111000",
  50511=>"110010000",
  50512=>"110000100",
  50513=>"011111111",
  50514=>"010000000",
  50515=>"111111111",
  50516=>"111111000",
  50517=>"101111111",
  50518=>"111111111",
  50519=>"000000000",
  50520=>"000000100",
  50521=>"110000000",
  50522=>"000000000",
  50523=>"001111111",
  50524=>"000001001",
  50525=>"110010010",
  50526=>"011001011",
  50527=>"111111011",
  50528=>"000111011",
  50529=>"000000000",
  50530=>"111001001",
  50531=>"000001011",
  50532=>"000000110",
  50533=>"001001101",
  50534=>"001001001",
  50535=>"000000000",
  50536=>"111111111",
  50537=>"101000000",
  50538=>"001000001",
  50539=>"000000000",
  50540=>"000000001",
  50541=>"001111011",
  50542=>"000000111",
  50543=>"000000000",
  50544=>"110100100",
  50545=>"000110111",
  50546=>"101000111",
  50547=>"011111100",
  50548=>"110111000",
  50549=>"110110100",
  50550=>"000111111",
  50551=>"111111011",
  50552=>"101000001",
  50553=>"111111111",
  50554=>"000000000",
  50555=>"001011000",
  50556=>"111111111",
  50557=>"000111111",
  50558=>"101001001",
  50559=>"101111111",
  50560=>"000000011",
  50561=>"101101011",
  50562=>"001011111",
  50563=>"110100000",
  50564=>"101000000",
  50565=>"111111110",
  50566=>"000000100",
  50567=>"101101111",
  50568=>"111011111",
  50569=>"100000000",
  50570=>"011001001",
  50571=>"100000000",
  50572=>"001001101",
  50573=>"000000000",
  50574=>"011111111",
  50575=>"110110111",
  50576=>"101100100",
  50577=>"000110111",
  50578=>"001000001",
  50579=>"000000000",
  50580=>"111111011",
  50581=>"001110100",
  50582=>"001111111",
  50583=>"000011011",
  50584=>"111111111",
  50585=>"101110111",
  50586=>"000000000",
  50587=>"001011111",
  50588=>"000000000",
  50589=>"111000000",
  50590=>"110000000",
  50591=>"001001001",
  50592=>"011000100",
  50593=>"011111011",
  50594=>"000010000",
  50595=>"000010010",
  50596=>"011111111",
  50597=>"111011000",
  50598=>"111111100",
  50599=>"000110111",
  50600=>"000000000",
  50601=>"000101000",
  50602=>"000111111",
  50603=>"111111011",
  50604=>"111101000",
  50605=>"111111110",
  50606=>"001111000",
  50607=>"111111111",
  50608=>"011011010",
  50609=>"001001001",
  50610=>"000000000",
  50611=>"000000000",
  50612=>"000000000",
  50613=>"000000101",
  50614=>"111110111",
  50615=>"000000001",
  50616=>"000001111",
  50617=>"000010110",
  50618=>"111101000",
  50619=>"100000001",
  50620=>"011111111",
  50621=>"000001111",
  50622=>"001000000",
  50623=>"000010000",
  50624=>"000000000",
  50625=>"110110000",
  50626=>"000000000",
  50627=>"011011000",
  50628=>"000000000",
  50629=>"001011111",
  50630=>"000000000",
  50631=>"000000110",
  50632=>"100000000",
  50633=>"111010000",
  50634=>"000000000",
  50635=>"000000000",
  50636=>"011011000",
  50637=>"000001111",
  50638=>"000110111",
  50639=>"111110111",
  50640=>"111111111",
  50641=>"010110100",
  50642=>"100100100",
  50643=>"111110100",
  50644=>"001000101",
  50645=>"010010000",
  50646=>"111101001",
  50647=>"100100101",
  50648=>"011111111",
  50649=>"001001000",
  50650=>"000001111",
  50651=>"000000111",
  50652=>"110111111",
  50653=>"000000000",
  50654=>"000100111",
  50655=>"001011111",
  50656=>"110000000",
  50657=>"111101111",
  50658=>"000000001",
  50659=>"111111111",
  50660=>"111111111",
  50661=>"111010011",
  50662=>"111111111",
  50663=>"010111111",
  50664=>"111111111",
  50665=>"111001001",
  50666=>"001000000",
  50667=>"000000000",
  50668=>"000000000",
  50669=>"101101001",
  50670=>"111111101",
  50671=>"111101111",
  50672=>"000000000",
  50673=>"111000111",
  50674=>"111111111",
  50675=>"000000000",
  50676=>"110110001",
  50677=>"111111111",
  50678=>"000000000",
  50679=>"011011111",
  50680=>"010010000",
  50681=>"111110000",
  50682=>"111100111",
  50683=>"111111000",
  50684=>"000111000",
  50685=>"001001010",
  50686=>"000001001",
  50687=>"000000000",
  50688=>"000010000",
  50689=>"000000001",
  50690=>"000000000",
  50691=>"111111111",
  50692=>"000000100",
  50693=>"111111111",
  50694=>"000111111",
  50695=>"011001000",
  50696=>"110110111",
  50697=>"000100111",
  50698=>"111110100",
  50699=>"011000000",
  50700=>"110000000",
  50701=>"111111111",
  50702=>"001001011",
  50703=>"000000000",
  50704=>"000000110",
  50705=>"000111011",
  50706=>"111111111",
  50707=>"111111111",
  50708=>"111111000",
  50709=>"000000111",
  50710=>"000000111",
  50711=>"100000000",
  50712=>"111111001",
  50713=>"000000011",
  50714=>"100000010",
  50715=>"110000000",
  50716=>"000000111",
  50717=>"000000000",
  50718=>"010000000",
  50719=>"111111011",
  50720=>"000110111",
  50721=>"111001000",
  50722=>"111111111",
  50723=>"111011111",
  50724=>"001000000",
  50725=>"011111111",
  50726=>"100111111",
  50727=>"000000000",
  50728=>"111111000",
  50729=>"000000111",
  50730=>"000000010",
  50731=>"001110110",
  50732=>"111000011",
  50733=>"110111000",
  50734=>"001111111",
  50735=>"111111111",
  50736=>"011011010",
  50737=>"000000110",
  50738=>"111011001",
  50739=>"000000100",
  50740=>"000000000",
  50741=>"000111111",
  50742=>"000011000",
  50743=>"111111111",
  50744=>"111111111",
  50745=>"111111000",
  50746=>"111100000",
  50747=>"100110010",
  50748=>"000000000",
  50749=>"100000000",
  50750=>"000111011",
  50751=>"000000111",
  50752=>"111111110",
  50753=>"111111110",
  50754=>"111111100",
  50755=>"111111000",
  50756=>"000110111",
  50757=>"100100110",
  50758=>"111111111",
  50759=>"101000000",
  50760=>"011111111",
  50761=>"001101100",
  50762=>"111111110",
  50763=>"110111111",
  50764=>"000000101",
  50765=>"110110100",
  50766=>"111000000",
  50767=>"111010000",
  50768=>"000000000",
  50769=>"011000011",
  50770=>"010010111",
  50771=>"000000100",
  50772=>"000000101",
  50773=>"101100100",
  50774=>"110101000",
  50775=>"111000000",
  50776=>"111110111",
  50777=>"000001111",
  50778=>"011111101",
  50779=>"001111110",
  50780=>"000000111",
  50781=>"111000000",
  50782=>"111011000",
  50783=>"111111110",
  50784=>"111000001",
  50785=>"111001000",
  50786=>"000000000",
  50787=>"111001000",
  50788=>"000000001",
  50789=>"000100111",
  50790=>"000000011",
  50791=>"000111111",
  50792=>"000111111",
  50793=>"000000000",
  50794=>"110000001",
  50795=>"000000000",
  50796=>"111110110",
  50797=>"000111111",
  50798=>"000000010",
  50799=>"110000000",
  50800=>"000011111",
  50801=>"111111111",
  50802=>"000000110",
  50803=>"001000000",
  50804=>"110111111",
  50805=>"011111000",
  50806=>"000011111",
  50807=>"000111111",
  50808=>"000000000",
  50809=>"110111101",
  50810=>"001000000",
  50811=>"001000000",
  50812=>"110111111",
  50813=>"111110100",
  50814=>"000100110",
  50815=>"110111111",
  50816=>"111100111",
  50817=>"000000000",
  50818=>"111111111",
  50819=>"000111111",
  50820=>"010101111",
  50821=>"000100111",
  50822=>"011100110",
  50823=>"110010011",
  50824=>"000000000",
  50825=>"000000111",
  50826=>"000000110",
  50827=>"110111100",
  50828=>"111001111",
  50829=>"110111000",
  50830=>"111011111",
  50831=>"111000000",
  50832=>"000000001",
  50833=>"000111011",
  50834=>"001110000",
  50835=>"111111000",
  50836=>"000000110",
  50837=>"100111111",
  50838=>"000100100",
  50839=>"011000000",
  50840=>"000110110",
  50841=>"101111000",
  50842=>"001000000",
  50843=>"001011111",
  50844=>"101111000",
  50845=>"000111111",
  50846=>"001001001",
  50847=>"101111100",
  50848=>"001011001",
  50849=>"111111111",
  50850=>"111111111",
  50851=>"000000110",
  50852=>"000000000",
  50853=>"000001011",
  50854=>"011111011",
  50855=>"000111111",
  50856=>"000000111",
  50857=>"010000010",
  50858=>"000000000",
  50859=>"111000000",
  50860=>"111111000",
  50861=>"000000011",
  50862=>"111100111",
  50863=>"000000111",
  50864=>"000000010",
  50865=>"000000111",
  50866=>"111111111",
  50867=>"000100101",
  50868=>"111111010",
  50869=>"111000000",
  50870=>"110000000",
  50871=>"111111110",
  50872=>"000000000",
  50873=>"000000000",
  50874=>"000000000",
  50875=>"000000001",
  50876=>"010110000",
  50877=>"010110000",
  50878=>"110111111",
  50879=>"111111110",
  50880=>"111101111",
  50881=>"000001111",
  50882=>"010110111",
  50883=>"110011010",
  50884=>"000000000",
  50885=>"111101111",
  50886=>"110111111",
  50887=>"110000000",
  50888=>"111111010",
  50889=>"001000000",
  50890=>"000000100",
  50891=>"000000100",
  50892=>"001001001",
  50893=>"110111111",
  50894=>"110111111",
  50895=>"000000101",
  50896=>"100000000",
  50897=>"000000000",
  50898=>"011111111",
  50899=>"000010110",
  50900=>"001100000",
  50901=>"011011101",
  50902=>"011101001",
  50903=>"010000000",
  50904=>"000000000",
  50905=>"100000000",
  50906=>"111111000",
  50907=>"000000111",
  50908=>"111111000",
  50909=>"111101111",
  50910=>"000000111",
  50911=>"000000000",
  50912=>"110111111",
  50913=>"000010000",
  50914=>"111111111",
  50915=>"111110000",
  50916=>"101101111",
  50917=>"110111111",
  50918=>"111111000",
  50919=>"111000000",
  50920=>"000000110",
  50921=>"111111110",
  50922=>"000010111",
  50923=>"110011011",
  50924=>"100000000",
  50925=>"000000111",
  50926=>"111111000",
  50927=>"010000000",
  50928=>"100100111",
  50929=>"000001111",
  50930=>"111111111",
  50931=>"000000011",
  50932=>"110110100",
  50933=>"111111000",
  50934=>"000001011",
  50935=>"111000110",
  50936=>"000000000",
  50937=>"100100000",
  50938=>"111111111",
  50939=>"110000000",
  50940=>"111000000",
  50941=>"001001111",
  50942=>"000000000",
  50943=>"011000000",
  50944=>"000110111",
  50945=>"000000001",
  50946=>"010000111",
  50947=>"000000000",
  50948=>"000110000",
  50949=>"111111111",
  50950=>"111110000",
  50951=>"111101000",
  50952=>"111111000",
  50953=>"111100110",
  50954=>"010111110",
  50955=>"110110111",
  50956=>"111000000",
  50957=>"000000101",
  50958=>"000000000",
  50959=>"000000000",
  50960=>"110100001",
  50961=>"111101111",
  50962=>"001000101",
  50963=>"100111011",
  50964=>"111111110",
  50965=>"100010000",
  50966=>"001001000",
  50967=>"111111000",
  50968=>"000001111",
  50969=>"111000000",
  50970=>"111111101",
  50971=>"000000000",
  50972=>"000000001",
  50973=>"000000000",
  50974=>"000000000",
  50975=>"111011000",
  50976=>"000111111",
  50977=>"111111111",
  50978=>"000000001",
  50979=>"111111101",
  50980=>"000000110",
  50981=>"110111111",
  50982=>"001000000",
  50983=>"000000111",
  50984=>"000000000",
  50985=>"000111111",
  50986=>"111100000",
  50987=>"100000100",
  50988=>"000001111",
  50989=>"000001011",
  50990=>"111111111",
  50991=>"000111110",
  50992=>"111111111",
  50993=>"110110110",
  50994=>"111111111",
  50995=>"111111111",
  50996=>"111000100",
  50997=>"000000001",
  50998=>"000000000",
  50999=>"111111110",
  51000=>"111000000",
  51001=>"000000111",
  51002=>"000000001",
  51003=>"110000000",
  51004=>"000000000",
  51005=>"000000000",
  51006=>"000000000",
  51007=>"110111000",
  51008=>"010000000",
  51009=>"111000110",
  51010=>"111111110",
  51011=>"111000111",
  51012=>"111111100",
  51013=>"111000001",
  51014=>"000001000",
  51015=>"011010000",
  51016=>"111111000",
  51017=>"100000000",
  51018=>"000001000",
  51019=>"111111000",
  51020=>"111111111",
  51021=>"100100111",
  51022=>"110111111",
  51023=>"000000110",
  51024=>"110110110",
  51025=>"000110111",
  51026=>"111000000",
  51027=>"000000001",
  51028=>"000000111",
  51029=>"011011011",
  51030=>"000000111",
  51031=>"101001001",
  51032=>"111111010",
  51033=>"000011001",
  51034=>"111110110",
  51035=>"000000000",
  51036=>"000000111",
  51037=>"000000000",
  51038=>"101000011",
  51039=>"111111111",
  51040=>"000000000",
  51041=>"000001011",
  51042=>"111001001",
  51043=>"010111000",
  51044=>"111111000",
  51045=>"001000001",
  51046=>"100111001",
  51047=>"110100100",
  51048=>"111111000",
  51049=>"000000000",
  51050=>"000000001",
  51051=>"110111110",
  51052=>"000000100",
  51053=>"000000000",
  51054=>"111111111",
  51055=>"000000110",
  51056=>"011001000",
  51057=>"000000000",
  51058=>"000110100",
  51059=>"111110111",
  51060=>"000000000",
  51061=>"000000111",
  51062=>"101111111",
  51063=>"111111111",
  51064=>"000011111",
  51065=>"111010000",
  51066=>"111011000",
  51067=>"111110111",
  51068=>"110110100",
  51069=>"010011000",
  51070=>"000000000",
  51071=>"000111111",
  51072=>"000000100",
  51073=>"011011011",
  51074=>"000011011",
  51075=>"101000000",
  51076=>"110111111",
  51077=>"000111110",
  51078=>"010111111",
  51079=>"111001000",
  51080=>"001000000",
  51081=>"000000111",
  51082=>"000000000",
  51083=>"111111111",
  51084=>"100001111",
  51085=>"000000011",
  51086=>"000000000",
  51087=>"000111000",
  51088=>"000001000",
  51089=>"111111000",
  51090=>"000000000",
  51091=>"000000000",
  51092=>"110111111",
  51093=>"010010000",
  51094=>"001000101",
  51095=>"000000000",
  51096=>"000110110",
  51097=>"000000000",
  51098=>"111110110",
  51099=>"111001011",
  51100=>"110110000",
  51101=>"000000110",
  51102=>"000000000",
  51103=>"000000111",
  51104=>"001000000",
  51105=>"000010111",
  51106=>"000000000",
  51107=>"111101001",
  51108=>"001001111",
  51109=>"110000000",
  51110=>"111000001",
  51111=>"111111000",
  51112=>"111111110",
  51113=>"001000001",
  51114=>"000000000",
  51115=>"100100111",
  51116=>"011011000",
  51117=>"000000011",
  51118=>"111110010",
  51119=>"111111000",
  51120=>"000000000",
  51121=>"000100111",
  51122=>"000000111",
  51123=>"010000111",
  51124=>"000000001",
  51125=>"101111111",
  51126=>"001001100",
  51127=>"000000101",
  51128=>"000000111",
  51129=>"000000111",
  51130=>"100000000",
  51131=>"111100100",
  51132=>"010110110",
  51133=>"111000111",
  51134=>"000000111",
  51135=>"101000000",
  51136=>"000000111",
  51137=>"111001011",
  51138=>"111111111",
  51139=>"000111000",
  51140=>"000000100",
  51141=>"011001111",
  51142=>"011011010",
  51143=>"110000000",
  51144=>"001000000",
  51145=>"000000000",
  51146=>"111000000",
  51147=>"111000111",
  51148=>"000000000",
  51149=>"111111000",
  51150=>"011001000",
  51151=>"100100111",
  51152=>"000000000",
  51153=>"111111000",
  51154=>"000000000",
  51155=>"111101111",
  51156=>"000001001",
  51157=>"111111000",
  51158=>"001001000",
  51159=>"101011010",
  51160=>"000000110",
  51161=>"000000001",
  51162=>"011111111",
  51163=>"111111011",
  51164=>"111101111",
  51165=>"111010111",
  51166=>"111110001",
  51167=>"000000001",
  51168=>"010111011",
  51169=>"111111110",
  51170=>"111111011",
  51171=>"000111111",
  51172=>"000000110",
  51173=>"100000100",
  51174=>"111111110",
  51175=>"111100100",
  51176=>"111110111",
  51177=>"111111111",
  51178=>"000000110",
  51179=>"001000111",
  51180=>"101111111",
  51181=>"000000000",
  51182=>"000000110",
  51183=>"000000000",
  51184=>"000000000",
  51185=>"000000000",
  51186=>"000000101",
  51187=>"000000101",
  51188=>"000000000",
  51189=>"000000000",
  51190=>"000111111",
  51191=>"001110111",
  51192=>"000010010",
  51193=>"100000000",
  51194=>"111111001",
  51195=>"010111001",
  51196=>"111111110",
  51197=>"111111000",
  51198=>"001011111",
  51199=>"000000000",
  51200=>"111110110",
  51201=>"100110010",
  51202=>"111111011",
  51203=>"001101000",
  51204=>"000001011",
  51205=>"000011111",
  51206=>"111101000",
  51207=>"000000000",
  51208=>"000001000",
  51209=>"100111111",
  51210=>"000011011",
  51211=>"111011000",
  51212=>"111101111",
  51213=>"010010000",
  51214=>"011000000",
  51215=>"011011001",
  51216=>"111110111",
  51217=>"101101111",
  51218=>"111111100",
  51219=>"111111010",
  51220=>"111111001",
  51221=>"000000000",
  51222=>"010010000",
  51223=>"111111101",
  51224=>"110111000",
  51225=>"111110111",
  51226=>"111000000",
  51227=>"101111001",
  51228=>"000000001",
  51229=>"110110000",
  51230=>"000000000",
  51231=>"111011111",
  51232=>"000000000",
  51233=>"001001000",
  51234=>"000011000",
  51235=>"111111011",
  51236=>"111110110",
  51237=>"000100100",
  51238=>"011111111",
  51239=>"011111111",
  51240=>"000010000",
  51241=>"000111111",
  51242=>"111110111",
  51243=>"110110000",
  51244=>"011011001",
  51245=>"110110000",
  51246=>"111101101",
  51247=>"100111011",
  51248=>"000000000",
  51249=>"101000000",
  51250=>"001000001",
  51251=>"000000111",
  51252=>"100000000",
  51253=>"001001001",
  51254=>"000001000",
  51255=>"001011111",
  51256=>"111111000",
  51257=>"000000010",
  51258=>"001011000",
  51259=>"111011001",
  51260=>"111111111",
  51261=>"001011001",
  51262=>"111111111",
  51263=>"000000000",
  51264=>"001001001",
  51265=>"000100110",
  51266=>"000100101",
  51267=>"000000111",
  51268=>"100100000",
  51269=>"101111111",
  51270=>"111110000",
  51271=>"111111111",
  51272=>"011001001",
  51273=>"111001001",
  51274=>"111111111",
  51275=>"011001001",
  51276=>"110110000",
  51277=>"000000101",
  51278=>"001001000",
  51279=>"111111111",
  51280=>"011011010",
  51281=>"000110000",
  51282=>"001011011",
  51283=>"111001001",
  51284=>"100100110",
  51285=>"111111111",
  51286=>"000001101",
  51287=>"000001001",
  51288=>"111111110",
  51289=>"000001010",
  51290=>"000010011",
  51291=>"011001001",
  51292=>"000000000",
  51293=>"111111001",
  51294=>"011011000",
  51295=>"101111001",
  51296=>"000000000",
  51297=>"000000000",
  51298=>"000000000",
  51299=>"000110100",
  51300=>"100000000",
  51301=>"111111111",
  51302=>"000000001",
  51303=>"000011111",
  51304=>"000011111",
  51305=>"110100111",
  51306=>"000010000",
  51307=>"000101111",
  51308=>"000000000",
  51309=>"001111111",
  51310=>"111111001",
  51311=>"000000001",
  51312=>"110110000",
  51313=>"011111111",
  51314=>"001001000",
  51315=>"111111011",
  51316=>"011011010",
  51317=>"111111111",
  51318=>"000011011",
  51319=>"000001001",
  51320=>"100100100",
  51321=>"111111111",
  51322=>"111001111",
  51323=>"000000000",
  51324=>"111111011",
  51325=>"111111111",
  51326=>"111111111",
  51327=>"111111111",
  51328=>"000000000",
  51329=>"000000111",
  51330=>"111111111",
  51331=>"110111111",
  51332=>"000000000",
  51333=>"111111111",
  51334=>"110111010",
  51335=>"010010000",
  51336=>"010000000",
  51337=>"101111110",
  51338=>"111101101",
  51339=>"001001011",
  51340=>"000010010",
  51341=>"111111111",
  51342=>"000000000",
  51343=>"000001001",
  51344=>"111111111",
  51345=>"101100100",
  51346=>"110011111",
  51347=>"000000000",
  51348=>"100100000",
  51349=>"011111000",
  51350=>"111111111",
  51351=>"110111010",
  51352=>"110110000",
  51353=>"011111111",
  51354=>"011110000",
  51355=>"110111010",
  51356=>"011111110",
  51357=>"000110111",
  51358=>"011011111",
  51359=>"011111011",
  51360=>"000000000",
  51361=>"001111001",
  51362=>"000000000",
  51363=>"111111011",
  51364=>"011001011",
  51365=>"111101111",
  51366=>"111111111",
  51367=>"010010000",
  51368=>"111011001",
  51369=>"111111111",
  51370=>"000100101",
  51371=>"000000000",
  51372=>"111111111",
  51373=>"111111000",
  51374=>"100101111",
  51375=>"111111111",
  51376=>"010111011",
  51377=>"001010110",
  51378=>"000000000",
  51379=>"000000000",
  51380=>"000000111",
  51381=>"000000000",
  51382=>"000000000",
  51383=>"000000000",
  51384=>"110100000",
  51385=>"000000000",
  51386=>"101000000",
  51387=>"110111111",
  51388=>"111111111",
  51389=>"100110111",
  51390=>"111111111",
  51391=>"000000111",
  51392=>"111111111",
  51393=>"000000000",
  51394=>"100111111",
  51395=>"111111000",
  51396=>"000000000",
  51397=>"010000000",
  51398=>"110010110",
  51399=>"000001111",
  51400=>"110111110",
  51401=>"101111111",
  51402=>"000000001",
  51403=>"111111111",
  51404=>"111110000",
  51405=>"111111111",
  51406=>"000000001",
  51407=>"111100111",
  51408=>"111111011",
  51409=>"111111011",
  51410=>"111010000",
  51411=>"001101111",
  51412=>"100100000",
  51413=>"000011011",
  51414=>"110110010",
  51415=>"000000110",
  51416=>"011000000",
  51417=>"000100000",
  51418=>"011011010",
  51419=>"000000000",
  51420=>"011011001",
  51421=>"111111111",
  51422=>"100000000",
  51423=>"111111000",
  51424=>"111111010",
  51425=>"110110000",
  51426=>"100111001",
  51427=>"101000000",
  51428=>"111100111",
  51429=>"000110110",
  51430=>"111111111",
  51431=>"111111000",
  51432=>"110110100",
  51433=>"110110111",
  51434=>"000000000",
  51435=>"111101111",
  51436=>"110111111",
  51437=>"011111010",
  51438=>"100000111",
  51439=>"011111001",
  51440=>"111110100",
  51441=>"011011011",
  51442=>"111011100",
  51443=>"110101100",
  51444=>"111111111",
  51445=>"110110100",
  51446=>"111111111",
  51447=>"010011011",
  51448=>"111111111",
  51449=>"000000000",
  51450=>"111111111",
  51451=>"000000000",
  51452=>"001000100",
  51453=>"011111111",
  51454=>"001000111",
  51455=>"011111000",
  51456=>"000000000",
  51457=>"000000000",
  51458=>"111111111",
  51459=>"000000000",
  51460=>"000111011",
  51461=>"000000000",
  51462=>"000000000",
  51463=>"101111111",
  51464=>"000000000",
  51465=>"011000100",
  51466=>"110110111",
  51467=>"111111111",
  51468=>"110110000",
  51469=>"001000000",
  51470=>"011000000",
  51471=>"100100111",
  51472=>"111111111",
  51473=>"110111111",
  51474=>"011001001",
  51475=>"110111101",
  51476=>"111111011",
  51477=>"000000000",
  51478=>"011011001",
  51479=>"110010110",
  51480=>"110111000",
  51481=>"111111111",
  51482=>"011001111",
  51483=>"000000010",
  51484=>"100100100",
  51485=>"000000000",
  51486=>"011011000",
  51487=>"111111011",
  51488=>"111100000",
  51489=>"000000001",
  51490=>"111111000",
  51491=>"111011111",
  51492=>"011000000",
  51493=>"111111111",
  51494=>"111111111",
  51495=>"001101001",
  51496=>"111000100",
  51497=>"011011111",
  51498=>"011111011",
  51499=>"010000000",
  51500=>"111111111",
  51501=>"010001011",
  51502=>"111000000",
  51503=>"000000000",
  51504=>"000000000",
  51505=>"101111111",
  51506=>"000001000",
  51507=>"000000000",
  51508=>"000000000",
  51509=>"000000000",
  51510=>"000000000",
  51511=>"000110000",
  51512=>"010111111",
  51513=>"011011011",
  51514=>"111111111",
  51515=>"000000000",
  51516=>"111111111",
  51517=>"000000000",
  51518=>"000100111",
  51519=>"001001001",
  51520=>"000000000",
  51521=>"111111111",
  51522=>"000000000",
  51523=>"111111111",
  51524=>"011111000",
  51525=>"111111110",
  51526=>"001000000",
  51527=>"111010010",
  51528=>"000110000",
  51529=>"000011001",
  51530=>"111111011",
  51531=>"110010011",
  51532=>"111111110",
  51533=>"011011001",
  51534=>"111111011",
  51535=>"010111111",
  51536=>"111111000",
  51537=>"001001001",
  51538=>"000000110",
  51539=>"011001001",
  51540=>"001000000",
  51541=>"111101111",
  51542=>"000000000",
  51543=>"101111100",
  51544=>"111111111",
  51545=>"111111111",
  51546=>"111111111",
  51547=>"000001001",
  51548=>"000000000",
  51549=>"000000000",
  51550=>"000000000",
  51551=>"011011111",
  51552=>"000000000",
  51553=>"111111111",
  51554=>"000000000",
  51555=>"111111111",
  51556=>"011000001",
  51557=>"000000011",
  51558=>"010010110",
  51559=>"110010000",
  51560=>"110111111",
  51561=>"010000111",
  51562=>"100000111",
  51563=>"000000000",
  51564=>"110110100",
  51565=>"000000000",
  51566=>"000000100",
  51567=>"000000111",
  51568=>"000000000",
  51569=>"111111111",
  51570=>"001111001",
  51571=>"111111110",
  51572=>"101111000",
  51573=>"000000000",
  51574=>"000100111",
  51575=>"000000000",
  51576=>"000000000",
  51577=>"000010000",
  51578=>"111111000",
  51579=>"011111111",
  51580=>"111111111",
  51581=>"111111010",
  51582=>"111111111",
  51583=>"100111101",
  51584=>"111111111",
  51585=>"000101111",
  51586=>"001001111",
  51587=>"000000111",
  51588=>"000001001",
  51589=>"011111010",
  51590=>"000000000",
  51591=>"100100111",
  51592=>"011001000",
  51593=>"001101000",
  51594=>"111111111",
  51595=>"111111010",
  51596=>"111111111",
  51597=>"110111110",
  51598=>"010010000",
  51599=>"000010000",
  51600=>"111111111",
  51601=>"001111001",
  51602=>"000000000",
  51603=>"111111111",
  51604=>"111111011",
  51605=>"011101111",
  51606=>"111101111",
  51607=>"111111111",
  51608=>"000000001",
  51609=>"111010110",
  51610=>"011001000",
  51611=>"111111111",
  51612=>"111111111",
  51613=>"000000000",
  51614=>"001000000",
  51615=>"000000111",
  51616=>"111111111",
  51617=>"111111111",
  51618=>"000000000",
  51619=>"000111111",
  51620=>"010000100",
  51621=>"000100101",
  51622=>"111111000",
  51623=>"111000000",
  51624=>"000110000",
  51625=>"011001011",
  51626=>"000000001",
  51627=>"100100000",
  51628=>"111111111",
  51629=>"111111110",
  51630=>"000110110",
  51631=>"001001000",
  51632=>"000000100",
  51633=>"110101101",
  51634=>"000110000",
  51635=>"111111111",
  51636=>"100000000",
  51637=>"001001001",
  51638=>"111001001",
  51639=>"001001000",
  51640=>"111001011",
  51641=>"110110101",
  51642=>"000101111",
  51643=>"000101011",
  51644=>"100100110",
  51645=>"011001001",
  51646=>"111111000",
  51647=>"011011001",
  51648=>"000000000",
  51649=>"111111111",
  51650=>"000000000",
  51651=>"011011001",
  51652=>"000000000",
  51653=>"000000100",
  51654=>"100000000",
  51655=>"000000100",
  51656=>"110110010",
  51657=>"111000110",
  51658=>"000000111",
  51659=>"111111111",
  51660=>"100100111",
  51661=>"001000000",
  51662=>"000000000",
  51663=>"110000000",
  51664=>"110000000",
  51665=>"000111110",
  51666=>"011001001",
  51667=>"111111111",
  51668=>"000000110",
  51669=>"000010000",
  51670=>"000000000",
  51671=>"110011001",
  51672=>"000100101",
  51673=>"100110100",
  51674=>"000000000",
  51675=>"000111111",
  51676=>"000000000",
  51677=>"111111111",
  51678=>"101001000",
  51679=>"010011110",
  51680=>"000000000",
  51681=>"001101110",
  51682=>"000000000",
  51683=>"000000000",
  51684=>"100110011",
  51685=>"100100101",
  51686=>"111011011",
  51687=>"001111001",
  51688=>"000111111",
  51689=>"001001111",
  51690=>"000000111",
  51691=>"111111111",
  51692=>"011111011",
  51693=>"111110110",
  51694=>"000111000",
  51695=>"000000000",
  51696=>"101101111",
  51697=>"000000101",
  51698=>"001001001",
  51699=>"010010000",
  51700=>"111111000",
  51701=>"000000000",
  51702=>"010011000",
  51703=>"001101101",
  51704=>"000000011",
  51705=>"100110100",
  51706=>"010011010",
  51707=>"111000000",
  51708=>"010000000",
  51709=>"000010110",
  51710=>"111111111",
  51711=>"001001101",
  51712=>"000000110",
  51713=>"000000000",
  51714=>"000000000",
  51715=>"000000110",
  51716=>"000000000",
  51717=>"111111111",
  51718=>"111111111",
  51719=>"100000000",
  51720=>"000000000",
  51721=>"111111111",
  51722=>"110010000",
  51723=>"000000000",
  51724=>"111111000",
  51725=>"111111111",
  51726=>"111011000",
  51727=>"111111111",
  51728=>"001111001",
  51729=>"111000000",
  51730=>"000001111",
  51731=>"111111001",
  51732=>"011000000",
  51733=>"111000000",
  51734=>"000011011",
  51735=>"011000001",
  51736=>"111111111",
  51737=>"101000001",
  51738=>"000000000",
  51739=>"111011001",
  51740=>"000000000",
  51741=>"111000001",
  51742=>"001111111",
  51743=>"000000000",
  51744=>"011111111",
  51745=>"111011000",
  51746=>"000000000",
  51747=>"111111111",
  51748=>"111111111",
  51749=>"111111111",
  51750=>"000100111",
  51751=>"111000001",
  51752=>"101000000",
  51753=>"110111010",
  51754=>"000000000",
  51755=>"111000000",
  51756=>"111001111",
  51757=>"001111111",
  51758=>"000000000",
  51759=>"110110111",
  51760=>"101011011",
  51761=>"000000000",
  51762=>"000111111",
  51763=>"111110100",
  51764=>"000000111",
  51765=>"111111111",
  51766=>"000111101",
  51767=>"011011111",
  51768=>"000000000",
  51769=>"111000100",
  51770=>"000000000",
  51771=>"110110010",
  51772=>"000000000",
  51773=>"000010000",
  51774=>"111111011",
  51775=>"100100000",
  51776=>"000000000",
  51777=>"000000010",
  51778=>"011011000",
  51779=>"111111001",
  51780=>"110000001",
  51781=>"000000000",
  51782=>"110010000",
  51783=>"111111111",
  51784=>"100100000",
  51785=>"000000111",
  51786=>"100100100",
  51787=>"000000001",
  51788=>"111110111",
  51789=>"110000110",
  51790=>"011000000",
  51791=>"111011001",
  51792=>"000100000",
  51793=>"000000110",
  51794=>"000111111",
  51795=>"000000111",
  51796=>"000000000",
  51797=>"111100101",
  51798=>"001111111",
  51799=>"000000111",
  51800=>"000000000",
  51801=>"100100100",
  51802=>"000000110",
  51803=>"111111111",
  51804=>"111111011",
  51805=>"111111111",
  51806=>"110111011",
  51807=>"000000000",
  51808=>"001000001",
  51809=>"111011010",
  51810=>"000000000",
  51811=>"110000000",
  51812=>"000000000",
  51813=>"001111111",
  51814=>"110111111",
  51815=>"000000101",
  51816=>"000000000",
  51817=>"000111111",
  51818=>"110100101",
  51819=>"111111000",
  51820=>"010010000",
  51821=>"111111111",
  51822=>"111111000",
  51823=>"110110110",
  51824=>"111111000",
  51825=>"100111110",
  51826=>"100000000",
  51827=>"111000000",
  51828=>"000000100",
  51829=>"111111111",
  51830=>"000011010",
  51831=>"001001011",
  51832=>"000000000",
  51833=>"111111111",
  51834=>"011000000",
  51835=>"011011000",
  51836=>"110110000",
  51837=>"100100111",
  51838=>"000000000",
  51839=>"000000000",
  51840=>"111000000",
  51841=>"111011011",
  51842=>"100000000",
  51843=>"110000100",
  51844=>"000000000",
  51845=>"000000000",
  51846=>"110011000",
  51847=>"000000000",
  51848=>"010110111",
  51849=>"000000000",
  51850=>"011111000",
  51851=>"000000000",
  51852=>"000000000",
  51853=>"111111111",
  51854=>"000111111",
  51855=>"111000111",
  51856=>"000100110",
  51857=>"000000000",
  51858=>"100110111",
  51859=>"111111010",
  51860=>"011001001",
  51861=>"000000000",
  51862=>"000000000",
  51863=>"000000000",
  51864=>"000000000",
  51865=>"001101000",
  51866=>"011111111",
  51867=>"000000000",
  51868=>"111111111",
  51869=>"000000000",
  51870=>"111101111",
  51871=>"111100100",
  51872=>"111000111",
  51873=>"111101000",
  51874=>"110111110",
  51875=>"010110100",
  51876=>"001111000",
  51877=>"110111111",
  51878=>"000000111",
  51879=>"001001101",
  51880=>"111011001",
  51881=>"001011001",
  51882=>"000000000",
  51883=>"000000000",
  51884=>"000000111",
  51885=>"100010110",
  51886=>"000111001",
  51887=>"000001101",
  51888=>"111111111",
  51889=>"011011101",
  51890=>"111111111",
  51891=>"000000000",
  51892=>"111111111",
  51893=>"000001000",
  51894=>"111111111",
  51895=>"100000000",
  51896=>"100111001",
  51897=>"101001111",
  51898=>"000000000",
  51899=>"001001000",
  51900=>"001000000",
  51901=>"011001111",
  51902=>"111111001",
  51903=>"000000000",
  51904=>"111111000",
  51905=>"000101111",
  51906=>"000011001",
  51907=>"000000000",
  51908=>"000111111",
  51909=>"100111111",
  51910=>"111110111",
  51911=>"000000000",
  51912=>"000111111",
  51913=>"111111000",
  51914=>"000110110",
  51915=>"011111111",
  51916=>"111100110",
  51917=>"111111111",
  51918=>"111111111",
  51919=>"001000000",
  51920=>"110111000",
  51921=>"001011001",
  51922=>"001010100",
  51923=>"111111111",
  51924=>"111100111",
  51925=>"111101100",
  51926=>"000000000",
  51927=>"111111000",
  51928=>"001111111",
  51929=>"111110000",
  51930=>"111111111",
  51931=>"100100111",
  51932=>"000000100",
  51933=>"000000110",
  51934=>"000000000",
  51935=>"100111111",
  51936=>"000000000",
  51937=>"000000000",
  51938=>"111011011",
  51939=>"000000100",
  51940=>"000000111",
  51941=>"001101111",
  51942=>"001000110",
  51943=>"000000000",
  51944=>"001000000",
  51945=>"111001000",
  51946=>"111111100",
  51947=>"001000000",
  51948=>"111111111",
  51949=>"111000110",
  51950=>"000001111",
  51951=>"000111011",
  51952=>"111101111",
  51953=>"110011000",
  51954=>"000110000",
  51955=>"000000110",
  51956=>"101011111",
  51957=>"000000000",
  51958=>"000001111",
  51959=>"000000110",
  51960=>"000000001",
  51961=>"111111001",
  51962=>"000010111",
  51963=>"101101111",
  51964=>"111011000",
  51965=>"000000000",
  51966=>"000000000",
  51967=>"001000111",
  51968=>"111111111",
  51969=>"000000000",
  51970=>"111111110",
  51971=>"101001111",
  51972=>"110111111",
  51973=>"111111100",
  51974=>"000111111",
  51975=>"011011010",
  51976=>"110110000",
  51977=>"000000000",
  51978=>"000000000",
  51979=>"101111111",
  51980=>"011001000",
  51981=>"100111111",
  51982=>"001001000",
  51983=>"011001001",
  51984=>"000011110",
  51985=>"000000000",
  51986=>"011000111",
  51987=>"000001111",
  51988=>"111110100",
  51989=>"111111011",
  51990=>"100101111",
  51991=>"111111001",
  51992=>"110000000",
  51993=>"111111111",
  51994=>"000000010",
  51995=>"001011111",
  51996=>"111111111",
  51997=>"110110110",
  51998=>"000000001",
  51999=>"111111111",
  52000=>"111110110",
  52001=>"111110000",
  52002=>"001001111",
  52003=>"111111111",
  52004=>"100001000",
  52005=>"111011000",
  52006=>"110110111",
  52007=>"111111000",
  52008=>"000000100",
  52009=>"000000011",
  52010=>"000000000",
  52011=>"010110000",
  52012=>"000000000",
  52013=>"111001000",
  52014=>"111111000",
  52015=>"000000001",
  52016=>"000000001",
  52017=>"111111111",
  52018=>"111111111",
  52019=>"100100100",
  52020=>"000000000",
  52021=>"111011101",
  52022=>"000011001",
  52023=>"000000000",
  52024=>"111000000",
  52025=>"110111111",
  52026=>"111111111",
  52027=>"111111011",
  52028=>"001000000",
  52029=>"011111111",
  52030=>"111111011",
  52031=>"111111000",
  52032=>"111111000",
  52033=>"000100110",
  52034=>"000000011",
  52035=>"000000001",
  52036=>"000000000",
  52037=>"110000000",
  52038=>"001000000",
  52039=>"000000111",
  52040=>"000001001",
  52041=>"000011000",
  52042=>"111000000",
  52043=>"111110000",
  52044=>"110110111",
  52045=>"111111111",
  52046=>"001001000",
  52047=>"000001001",
  52048=>"000001011",
  52049=>"000000111",
  52050=>"010011001",
  52051=>"111110011",
  52052=>"000000000",
  52053=>"000010011",
  52054=>"111111000",
  52055=>"000000001",
  52056=>"111111111",
  52057=>"101111100",
  52058=>"111110000",
  52059=>"111001001",
  52060=>"000000000",
  52061=>"111111111",
  52062=>"000000000",
  52063=>"111111001",
  52064=>"000000000",
  52065=>"000001101",
  52066=>"111111111",
  52067=>"000000000",
  52068=>"001001111",
  52069=>"000111111",
  52070=>"111101111",
  52071=>"000001001",
  52072=>"110000000",
  52073=>"101100000",
  52074=>"001000000",
  52075=>"000100000",
  52076=>"000000000",
  52077=>"000000000",
  52078=>"111101101",
  52079=>"000000000",
  52080=>"000000000",
  52081=>"001001111",
  52082=>"000110111",
  52083=>"111110111",
  52084=>"011010000",
  52085=>"110100001",
  52086=>"100110110",
  52087=>"000000000",
  52088=>"111111111",
  52089=>"110000111",
  52090=>"111111111",
  52091=>"000001001",
  52092=>"000000000",
  52093=>"111111111",
  52094=>"000000000",
  52095=>"100100000",
  52096=>"111101100",
  52097=>"011011111",
  52098=>"110100110",
  52099=>"000101000",
  52100=>"110010010",
  52101=>"110010000",
  52102=>"000011111",
  52103=>"011010000",
  52104=>"111111011",
  52105=>"000000000",
  52106=>"000001000",
  52107=>"000001111",
  52108=>"110111000",
  52109=>"111000000",
  52110=>"110101111",
  52111=>"100000000",
  52112=>"000000000",
  52113=>"111011000",
  52114=>"000000111",
  52115=>"110000000",
  52116=>"000111111",
  52117=>"000000011",
  52118=>"000000000",
  52119=>"110110110",
  52120=>"101101000",
  52121=>"111111110",
  52122=>"100000000",
  52123=>"000000001",
  52124=>"100001111",
  52125=>"111111111",
  52126=>"111011111",
  52127=>"000000000",
  52128=>"001011001",
  52129=>"001011111",
  52130=>"000100001",
  52131=>"010000000",
  52132=>"000000000",
  52133=>"111111111",
  52134=>"000000000",
  52135=>"000000000",
  52136=>"111010000",
  52137=>"000110000",
  52138=>"100100000",
  52139=>"001000000",
  52140=>"000000000",
  52141=>"111111111",
  52142=>"000000000",
  52143=>"011011011",
  52144=>"110010110",
  52145=>"000100000",
  52146=>"111111111",
  52147=>"000000000",
  52148=>"011000000",
  52149=>"000000000",
  52150=>"111111111",
  52151=>"000010000",
  52152=>"000000111",
  52153=>"000111000",
  52154=>"100101111",
  52155=>"000000100",
  52156=>"111111100",
  52157=>"100111111",
  52158=>"011111111",
  52159=>"100000000",
  52160=>"111010111",
  52161=>"000100000",
  52162=>"000000000",
  52163=>"000000000",
  52164=>"111111000",
  52165=>"000111111",
  52166=>"110001011",
  52167=>"000000000",
  52168=>"000100000",
  52169=>"111111111",
  52170=>"000000000",
  52171=>"111111011",
  52172=>"111111111",
  52173=>"000000000",
  52174=>"000000111",
  52175=>"111010111",
  52176=>"110110000",
  52177=>"111011001",
  52178=>"011000100",
  52179=>"111011000",
  52180=>"001000000",
  52181=>"000000000",
  52182=>"000000000",
  52183=>"110000000",
  52184=>"111111111",
  52185=>"000000000",
  52186=>"000110000",
  52187=>"000000011",
  52188=>"110111001",
  52189=>"000000100",
  52190=>"011010000",
  52191=>"110100111",
  52192=>"111000111",
  52193=>"111110001",
  52194=>"111110100",
  52195=>"000000001",
  52196=>"000000100",
  52197=>"111111111",
  52198=>"000000000",
  52199=>"111111000",
  52200=>"101111111",
  52201=>"000000000",
  52202=>"000000111",
  52203=>"110110011",
  52204=>"100110000",
  52205=>"011011011",
  52206=>"100100000",
  52207=>"000000000",
  52208=>"001001001",
  52209=>"111111111",
  52210=>"111111000",
  52211=>"111001001",
  52212=>"001001000",
  52213=>"000000000",
  52214=>"110110111",
  52215=>"000000110",
  52216=>"000000000",
  52217=>"001001111",
  52218=>"111111111",
  52219=>"111101111",
  52220=>"000000100",
  52221=>"000000000",
  52222=>"000000011",
  52223=>"001001111",
  52224=>"111111110",
  52225=>"000000000",
  52226=>"111111111",
  52227=>"000000100",
  52228=>"100000100",
  52229=>"100100111",
  52230=>"100000000",
  52231=>"000000000",
  52232=>"111100101",
  52233=>"100111101",
  52234=>"111001111",
  52235=>"001000000",
  52236=>"111111110",
  52237=>"110000000",
  52238=>"111111000",
  52239=>"000000110",
  52240=>"100001001",
  52241=>"000000000",
  52242=>"111111111",
  52243=>"000000111",
  52244=>"111111111",
  52245=>"000100100",
  52246=>"101000000",
  52247=>"111111110",
  52248=>"100000000",
  52249=>"111001000",
  52250=>"111111111",
  52251=>"000000010",
  52252=>"111101111",
  52253=>"111111000",
  52254=>"011011000",
  52255=>"000000000",
  52256=>"000000000",
  52257=>"000001100",
  52258=>"111001001",
  52259=>"110000111",
  52260=>"110000000",
  52261=>"000000010",
  52262=>"000000000",
  52263=>"001000000",
  52264=>"111101100",
  52265=>"000000101",
  52266=>"000000000",
  52267=>"000000001",
  52268=>"000000011",
  52269=>"111111110",
  52270=>"111111001",
  52271=>"000110111",
  52272=>"000000000",
  52273=>"111011001",
  52274=>"000000001",
  52275=>"000000000",
  52276=>"011011010",
  52277=>"000001001",
  52278=>"110100111",
  52279=>"111101000",
  52280=>"001000000",
  52281=>"111000000",
  52282=>"111000100",
  52283=>"000010000",
  52284=>"111111111",
  52285=>"111111100",
  52286=>"001001001",
  52287=>"111100100",
  52288=>"000000000",
  52289=>"000000001",
  52290=>"111110110",
  52291=>"111111111",
  52292=>"111100110",
  52293=>"111111111",
  52294=>"000011010",
  52295=>"111111111",
  52296=>"111111111",
  52297=>"001000111",
  52298=>"101100111",
  52299=>"111100101",
  52300=>"111111111",
  52301=>"111111001",
  52302=>"000110111",
  52303=>"000000000",
  52304=>"000000010",
  52305=>"111000000",
  52306=>"000000111",
  52307=>"101000000",
  52308=>"000000000",
  52309=>"011111111",
  52310=>"000000111",
  52311=>"011111111",
  52312=>"111110111",
  52313=>"111111101",
  52314=>"111111011",
  52315=>"100100100",
  52316=>"000000000",
  52317=>"000000000",
  52318=>"111111111",
  52319=>"000000000",
  52320=>"110000000",
  52321=>"000000000",
  52322=>"000111101",
  52323=>"001000000",
  52324=>"111111111",
  52325=>"010000000",
  52326=>"111000000",
  52327=>"011011110",
  52328=>"000100111",
  52329=>"111111111",
  52330=>"101100100",
  52331=>"111111111",
  52332=>"001001001",
  52333=>"000111111",
  52334=>"000000001",
  52335=>"100000001",
  52336=>"000111111",
  52337=>"111111000",
  52338=>"011011011",
  52339=>"100000000",
  52340=>"000000000",
  52341=>"111110000",
  52342=>"000001001",
  52343=>"111101000",
  52344=>"111111111",
  52345=>"011000000",
  52346=>"111111111",
  52347=>"111011010",
  52348=>"110000001",
  52349=>"111111111",
  52350=>"111010000",
  52351=>"000000000",
  52352=>"000000000",
  52353=>"010000000",
  52354=>"000100111",
  52355=>"000000000",
  52356=>"000000000",
  52357=>"000000001",
  52358=>"000000000",
  52359=>"000000110",
  52360=>"100110111",
  52361=>"000000000",
  52362=>"000001101",
  52363=>"111111111",
  52364=>"111100000",
  52365=>"110111000",
  52366=>"111000110",
  52367=>"000000000",
  52368=>"000000000",
  52369=>"000000000",
  52370=>"000111111",
  52371=>"000000001",
  52372=>"111111110",
  52373=>"000000000",
  52374=>"111111000",
  52375=>"001000000",
  52376=>"110111111",
  52377=>"111101111",
  52378=>"000000000",
  52379=>"011011000",
  52380=>"000000000",
  52381=>"000000000",
  52382=>"000000000",
  52383=>"111111111",
  52384=>"000101100",
  52385=>"111001100",
  52386=>"001001000",
  52387=>"111111111",
  52388=>"111100111",
  52389=>"000000000",
  52390=>"111111111",
  52391=>"100100000",
  52392=>"111001011",
  52393=>"111111111",
  52394=>"111101001",
  52395=>"100000000",
  52396=>"000000000",
  52397=>"000000000",
  52398=>"111100110",
  52399=>"110001000",
  52400=>"111111111",
  52401=>"000000000",
  52402=>"000000000",
  52403=>"111111011",
  52404=>"000000000",
  52405=>"000001001",
  52406=>"111111111",
  52407=>"000000101",
  52408=>"111111111",
  52409=>"000000000",
  52410=>"111100100",
  52411=>"100100111",
  52412=>"111111001",
  52413=>"001000111",
  52414=>"000000001",
  52415=>"000001111",
  52416=>"000000000",
  52417=>"001111111",
  52418=>"111111110",
  52419=>"001111111",
  52420=>"000000000",
  52421=>"000011011",
  52422=>"000000000",
  52423=>"111001100",
  52424=>"010111111",
  52425=>"111111111",
  52426=>"000000100",
  52427=>"111011111",
  52428=>"111011011",
  52429=>"111000000",
  52430=>"100000001",
  52431=>"110000111",
  52432=>"101111111",
  52433=>"000000000",
  52434=>"111111000",
  52435=>"000000000",
  52436=>"111111010",
  52437=>"111111011",
  52438=>"111111111",
  52439=>"000000111",
  52440=>"110111111",
  52441=>"111000000",
  52442=>"000000000",
  52443=>"111100000",
  52444=>"110101111",
  52445=>"111111111",
  52446=>"000001001",
  52447=>"000000011",
  52448=>"000000000",
  52449=>"111111111",
  52450=>"011111111",
  52451=>"000000000",
  52452=>"000000110",
  52453=>"001001001",
  52454=>"100000000",
  52455=>"111000000",
  52456=>"011000000",
  52457=>"101111001",
  52458=>"111000000",
  52459=>"000000001",
  52460=>"111111000",
  52461=>"111111111",
  52462=>"110110110",
  52463=>"111111011",
  52464=>"010000000",
  52465=>"000000111",
  52466=>"000011111",
  52467=>"000000000",
  52468=>"111111000",
  52469=>"000000000",
  52470=>"001101111",
  52471=>"111111000",
  52472=>"110000000",
  52473=>"000011000",
  52474=>"000101111",
  52475=>"000000000",
  52476=>"110111111",
  52477=>"001001011",
  52478=>"100000000",
  52479=>"000000000",
  52480=>"000000000",
  52481=>"000000001",
  52482=>"000000000",
  52483=>"111111111",
  52484=>"001101001",
  52485=>"000000000",
  52486=>"000000000",
  52487=>"111111111",
  52488=>"000010000",
  52489=>"011001000",
  52490=>"011011011",
  52491=>"111111110",
  52492=>"000000000",
  52493=>"001000000",
  52494=>"101010001",
  52495=>"011010010",
  52496=>"111111000",
  52497=>"100110111",
  52498=>"111001100",
  52499=>"111111111",
  52500=>"110111000",
  52501=>"111111000",
  52502=>"111100010",
  52503=>"100111111",
  52504=>"111111111",
  52505=>"100000000",
  52506=>"000100010",
  52507=>"110100000",
  52508=>"111000010",
  52509=>"110111111",
  52510=>"110110111",
  52511=>"000000000",
  52512=>"001100000",
  52513=>"000010000",
  52514=>"111111111",
  52515=>"110100110",
  52516=>"000100111",
  52517=>"000000001",
  52518=>"110100000",
  52519=>"100100000",
  52520=>"110111000",
  52521=>"111111111",
  52522=>"100100100",
  52523=>"000000001",
  52524=>"000000000",
  52525=>"111111110",
  52526=>"110110111",
  52527=>"110111111",
  52528=>"111111111",
  52529=>"101111110",
  52530=>"110110110",
  52531=>"000111111",
  52532=>"111101011",
  52533=>"001011111",
  52534=>"001000111",
  52535=>"000000000",
  52536=>"010110000",
  52537=>"111111111",
  52538=>"111111111",
  52539=>"011000001",
  52540=>"000111111",
  52541=>"111111000",
  52542=>"111100100",
  52543=>"111111011",
  52544=>"000000000",
  52545=>"101101111",
  52546=>"100000000",
  52547=>"111111010",
  52548=>"100000000",
  52549=>"111111111",
  52550=>"000000000",
  52551=>"111100110",
  52552=>"011000001",
  52553=>"001111111",
  52554=>"111110111",
  52555=>"000000000",
  52556=>"011000000",
  52557=>"000000111",
  52558=>"100110010",
  52559=>"110111111",
  52560=>"000011000",
  52561=>"001100100",
  52562=>"110000110",
  52563=>"111000000",
  52564=>"000000000",
  52565=>"011001111",
  52566=>"000110000",
  52567=>"000000000",
  52568=>"111110011",
  52569=>"111111111",
  52570=>"010000000",
  52571=>"111010111",
  52572=>"000111111",
  52573=>"111111111",
  52574=>"111111100",
  52575=>"001000000",
  52576=>"111111111",
  52577=>"001100000",
  52578=>"111001000",
  52579=>"111011011",
  52580=>"000000000",
  52581=>"000000000",
  52582=>"111111111",
  52583=>"011111111",
  52584=>"010000011",
  52585=>"111111010",
  52586=>"111110100",
  52587=>"111111111",
  52588=>"000000111",
  52589=>"111110111",
  52590=>"000000000",
  52591=>"000101001",
  52592=>"010000000",
  52593=>"011111111",
  52594=>"100100101",
  52595=>"111111111",
  52596=>"000000001",
  52597=>"111110111",
  52598=>"000111111",
  52599=>"000000000",
  52600=>"111111111",
  52601=>"000100000",
  52602=>"000000001",
  52603=>"000100111",
  52604=>"111111111",
  52605=>"111111111",
  52606=>"111111111",
  52607=>"000001111",
  52608=>"111011001",
  52609=>"111101101",
  52610=>"111111111",
  52611=>"000000000",
  52612=>"111011110",
  52613=>"010110110",
  52614=>"000000110",
  52615=>"000110111",
  52616=>"000000111",
  52617=>"111111011",
  52618=>"000000111",
  52619=>"011011000",
  52620=>"100100111",
  52621=>"110110110",
  52622=>"111111010",
  52623=>"000000001",
  52624=>"001000000",
  52625=>"100000000",
  52626=>"111011000",
  52627=>"111111111",
  52628=>"000000000",
  52629=>"000000000",
  52630=>"111000111",
  52631=>"100000110",
  52632=>"011000000",
  52633=>"000000000",
  52634=>"110010101",
  52635=>"111111111",
  52636=>"000010010",
  52637=>"111111101",
  52638=>"000000000",
  52639=>"111111111",
  52640=>"100101111",
  52641=>"101111011",
  52642=>"000000111",
  52643=>"111111111",
  52644=>"100000000",
  52645=>"100000000",
  52646=>"111111111",
  52647=>"000000100",
  52648=>"011011011",
  52649=>"000100111",
  52650=>"000111111",
  52651=>"000000000",
  52652=>"110111111",
  52653=>"111111100",
  52654=>"111111111",
  52655=>"111111111",
  52656=>"111111000",
  52657=>"000000000",
  52658=>"000000000",
  52659=>"111111111",
  52660=>"111110000",
  52661=>"111101111",
  52662=>"000100111",
  52663=>"000000000",
  52664=>"111111111",
  52665=>"011111011",
  52666=>"100001111",
  52667=>"000000111",
  52668=>"111111001",
  52669=>"111111101",
  52670=>"000000000",
  52671=>"001011001",
  52672=>"000000000",
  52673=>"111000000",
  52674=>"000010010",
  52675=>"010111111",
  52676=>"111110110",
  52677=>"101000000",
  52678=>"001000100",
  52679=>"111111011",
  52680=>"000000000",
  52681=>"111000111",
  52682=>"000010000",
  52683=>"000000000",
  52684=>"010111111",
  52685=>"100001001",
  52686=>"111011011",
  52687=>"100000111",
  52688=>"000000111",
  52689=>"101000000",
  52690=>"111111000",
  52691=>"000000000",
  52692=>"111111111",
  52693=>"101111111",
  52694=>"101101000",
  52695=>"000000000",
  52696=>"000000000",
  52697=>"110011000",
  52698=>"111000111",
  52699=>"000000011",
  52700=>"111111111",
  52701=>"000000100",
  52702=>"000000000",
  52703=>"100100000",
  52704=>"001011111",
  52705=>"000000110",
  52706=>"111111000",
  52707=>"110100110",
  52708=>"111111111",
  52709=>"111111111",
  52710=>"111100101",
  52711=>"110111111",
  52712=>"000000000",
  52713=>"000001011",
  52714=>"000000000",
  52715=>"000101011",
  52716=>"110000000",
  52717=>"001011001",
  52718=>"011111111",
  52719=>"110110111",
  52720=>"001000101",
  52721=>"000010000",
  52722=>"111111111",
  52723=>"000001000",
  52724=>"111111111",
  52725=>"111111111",
  52726=>"010000000",
  52727=>"001011011",
  52728=>"001011000",
  52729=>"111111111",
  52730=>"000000000",
  52731=>"000001001",
  52732=>"001101000",
  52733=>"000000000",
  52734=>"000000000",
  52735=>"111111111",
  52736=>"111000110",
  52737=>"000000000",
  52738=>"001111111",
  52739=>"100000101",
  52740=>"000110111",
  52741=>"101000001",
  52742=>"111101101",
  52743=>"111111111",
  52744=>"100110111",
  52745=>"000101110",
  52746=>"110110111",
  52747=>"111000000",
  52748=>"011010000",
  52749=>"111111000",
  52750=>"000111111",
  52751=>"111111111",
  52752=>"111111010",
  52753=>"111111111",
  52754=>"110110100",
  52755=>"000111111",
  52756=>"001001111",
  52757=>"011000001",
  52758=>"011000000",
  52759=>"111000000",
  52760=>"111111111",
  52761=>"111011000",
  52762=>"101111000",
  52763=>"000000111",
  52764=>"111000000",
  52765=>"000000010",
  52766=>"111110110",
  52767=>"111110000",
  52768=>"000000111",
  52769=>"111000000",
  52770=>"110000000",
  52771=>"011111011",
  52772=>"000000011",
  52773=>"000000000",
  52774=>"110001001",
  52775=>"111000111",
  52776=>"111111001",
  52777=>"000000000",
  52778=>"111111111",
  52779=>"111011111",
  52780=>"111001010",
  52781=>"000000111",
  52782=>"010000000",
  52783=>"000000001",
  52784=>"011000000",
  52785=>"011111110",
  52786=>"101001000",
  52787=>"000000000",
  52788=>"111100000",
  52789=>"110111010",
  52790=>"111111101",
  52791=>"111111011",
  52792=>"110110111",
  52793=>"000000000",
  52794=>"000000111",
  52795=>"100000111",
  52796=>"001111011",
  52797=>"101100100",
  52798=>"000100100",
  52799=>"111100111",
  52800=>"000001111",
  52801=>"010000111",
  52802=>"111101000",
  52803=>"000000000",
  52804=>"010000010",
  52805=>"000000111",
  52806=>"000000001",
  52807=>"111111111",
  52808=>"111110111",
  52809=>"000000011",
  52810=>"011011110",
  52811=>"111111000",
  52812=>"111101001",
  52813=>"000000111",
  52814=>"111111111",
  52815=>"111111011",
  52816=>"011001111",
  52817=>"000011111",
  52818=>"000000001",
  52819=>"111011000",
  52820=>"000000001",
  52821=>"000100000",
  52822=>"111011001",
  52823=>"000000000",
  52824=>"110000001",
  52825=>"111101111",
  52826=>"111111111",
  52827=>"100000000",
  52828=>"111111100",
  52829=>"111111011",
  52830=>"011110000",
  52831=>"111001011",
  52832=>"110100111",
  52833=>"111111010",
  52834=>"000000000",
  52835=>"010000111",
  52836=>"000000000",
  52837=>"000000000",
  52838=>"111111010",
  52839=>"111111111",
  52840=>"111110110",
  52841=>"001000000",
  52842=>"000000000",
  52843=>"001000000",
  52844=>"000000101",
  52845=>"000000000",
  52846=>"111111111",
  52847=>"111111111",
  52848=>"000111111",
  52849=>"111111000",
  52850=>"100110111",
  52851=>"111111111",
  52852=>"000000111",
  52853=>"111110000",
  52854=>"011000001",
  52855=>"101100101",
  52856=>"010111000",
  52857=>"111110111",
  52858=>"111001001",
  52859=>"111111111",
  52860=>"110110000",
  52861=>"101001001",
  52862=>"000000000",
  52863=>"000001001",
  52864=>"001101111",
  52865=>"111000000",
  52866=>"010011111",
  52867=>"111100100",
  52868=>"000100111",
  52869=>"111111111",
  52870=>"001001101",
  52871=>"000000000",
  52872=>"111101000",
  52873=>"111111111",
  52874=>"000111111",
  52875=>"111110110",
  52876=>"000000110",
  52877=>"111000000",
  52878=>"111101100",
  52879=>"001001001",
  52880=>"011001011",
  52881=>"000000000",
  52882=>"000010111",
  52883=>"111100000",
  52884=>"000000100",
  52885=>"001011111",
  52886=>"111111111",
  52887=>"011111011",
  52888=>"111011000",
  52889=>"111111000",
  52890=>"110001001",
  52891=>"110110000",
  52892=>"000000000",
  52893=>"000000000",
  52894=>"111111111",
  52895=>"111010000",
  52896=>"111001000",
  52897=>"000000001",
  52898=>"000000111",
  52899=>"000001111",
  52900=>"000000010",
  52901=>"000000110",
  52902=>"001001000",
  52903=>"010010010",
  52904=>"111000111",
  52905=>"110111111",
  52906=>"111111111",
  52907=>"000000111",
  52908=>"000000000",
  52909=>"011100110",
  52910=>"000000000",
  52911=>"111111001",
  52912=>"011001111",
  52913=>"111000000",
  52914=>"111111111",
  52915=>"111000001",
  52916=>"111000000",
  52917=>"111000000",
  52918=>"000000000",
  52919=>"111111110",
  52920=>"111111111",
  52921=>"111111011",
  52922=>"111111000",
  52923=>"011001000",
  52924=>"000000011",
  52925=>"000001011",
  52926=>"000000001",
  52927=>"000000101",
  52928=>"000000111",
  52929=>"111111110",
  52930=>"001101011",
  52931=>"011111111",
  52932=>"100000000",
  52933=>"111000001",
  52934=>"111111111",
  52935=>"100000100",
  52936=>"000000000",
  52937=>"000000000",
  52938=>"000000001",
  52939=>"000111111",
  52940=>"111111100",
  52941=>"110110100",
  52942=>"111101101",
  52943=>"000000000",
  52944=>"110011111",
  52945=>"000000001",
  52946=>"011000111",
  52947=>"110000000",
  52948=>"000000000",
  52949=>"110111000",
  52950=>"100101000",
  52951=>"111000000",
  52952=>"111111111",
  52953=>"001000000",
  52954=>"101000000",
  52955=>"101111111",
  52956=>"100000000",
  52957=>"100000110",
  52958=>"000000000",
  52959=>"100111011",
  52960=>"000111111",
  52961=>"111111110",
  52962=>"110010011",
  52963=>"111111111",
  52964=>"101101100",
  52965=>"111000000",
  52966=>"111110000",
  52967=>"000000000",
  52968=>"000000100",
  52969=>"000001111",
  52970=>"000000101",
  52971=>"110111111",
  52972=>"001011000",
  52973=>"110110011",
  52974=>"111111111",
  52975=>"011111111",
  52976=>"111111111",
  52977=>"000000001",
  52978=>"000000000",
  52979=>"000000001",
  52980=>"000000001",
  52981=>"111100110",
  52982=>"111000000",
  52983=>"000000000",
  52984=>"111111111",
  52985=>"111001000",
  52986=>"001111111",
  52987=>"000000111",
  52988=>"101001000",
  52989=>"001001111",
  52990=>"111100100",
  52991=>"000111111",
  52992=>"111111000",
  52993=>"011000110",
  52994=>"000110111",
  52995=>"000001111",
  52996=>"000000000",
  52997=>"101111111",
  52998=>"000000000",
  52999=>"000000101",
  53000=>"000000110",
  53001=>"001000000",
  53002=>"111011000",
  53003=>"111111111",
  53004=>"000000001",
  53005=>"000100111",
  53006=>"000000001",
  53007=>"111111001",
  53008=>"111111100",
  53009=>"000000000",
  53010=>"101101100",
  53011=>"000000000",
  53012=>"111000110",
  53013=>"001011011",
  53014=>"111000000",
  53015=>"111000000",
  53016=>"001111000",
  53017=>"111111111",
  53018=>"000000000",
  53019=>"111000001",
  53020=>"111000000",
  53021=>"011010010",
  53022=>"000011001",
  53023=>"000111111",
  53024=>"000100100",
  53025=>"000111110",
  53026=>"100000111",
  53027=>"001011101",
  53028=>"011011111",
  53029=>"100101001",
  53030=>"110100100",
  53031=>"011000000",
  53032=>"100000000",
  53033=>"000000011",
  53034=>"111111011",
  53035=>"100111111",
  53036=>"011000000",
  53037=>"000101000",
  53038=>"100101100",
  53039=>"111111010",
  53040=>"111101111",
  53041=>"001011000",
  53042=>"110110100",
  53043=>"011111011",
  53044=>"100101001",
  53045=>"111110111",
  53046=>"001111000",
  53047=>"111011000",
  53048=>"000000000",
  53049=>"000000111",
  53050=>"001101001",
  53051=>"000000100",
  53052=>"110110110",
  53053=>"000000000",
  53054=>"111111011",
  53055=>"111111110",
  53056=>"011111111",
  53057=>"000000001",
  53058=>"111000001",
  53059=>"111000000",
  53060=>"011011011",
  53061=>"111111111",
  53062=>"100100000",
  53063=>"000000001",
  53064=>"000000000",
  53065=>"101000001",
  53066=>"011000000",
  53067=>"001000001",
  53068=>"111111111",
  53069=>"100100111",
  53070=>"000000001",
  53071=>"000000001",
  53072=>"111001000",
  53073=>"000000111",
  53074=>"000000110",
  53075=>"010000000",
  53076=>"100110000",
  53077=>"011011011",
  53078=>"011011111",
  53079=>"111100000",
  53080=>"111111000",
  53081=>"111111111",
  53082=>"001111111",
  53083=>"000100111",
  53084=>"001000001",
  53085=>"000000011",
  53086=>"101101111",
  53087=>"000001000",
  53088=>"000000000",
  53089=>"111111110",
  53090=>"111011001",
  53091=>"111111011",
  53092=>"000001011",
  53093=>"000000000",
  53094=>"000011111",
  53095=>"000000100",
  53096=>"111000100",
  53097=>"111011011",
  53098=>"001000000",
  53099=>"001001000",
  53100=>"100110000",
  53101=>"011111111",
  53102=>"000000000",
  53103=>"000001101",
  53104=>"011000000",
  53105=>"111011000",
  53106=>"000000101",
  53107=>"100100111",
  53108=>"001000000",
  53109=>"011111111",
  53110=>"000000111",
  53111=>"011001011",
  53112=>"111111111",
  53113=>"000000001",
  53114=>"111111111",
  53115=>"000111110",
  53116=>"011001011",
  53117=>"111111111",
  53118=>"100111111",
  53119=>"000100111",
  53120=>"111111010",
  53121=>"111111111",
  53122=>"000000000",
  53123=>"000000010",
  53124=>"110000001",
  53125=>"010111011",
  53126=>"111111000",
  53127=>"000000000",
  53128=>"111111111",
  53129=>"111000000",
  53130=>"000000100",
  53131=>"111111000",
  53132=>"001001111",
  53133=>"111101000",
  53134=>"111000000",
  53135=>"111111111",
  53136=>"000111000",
  53137=>"111011011",
  53138=>"111001111",
  53139=>"011111111",
  53140=>"111111111",
  53141=>"000010000",
  53142=>"000010111",
  53143=>"000000000",
  53144=>"001000000",
  53145=>"111111111",
  53146=>"000001111",
  53147=>"000000111",
  53148=>"111000000",
  53149=>"000000001",
  53150=>"000000000",
  53151=>"000000111",
  53152=>"001000000",
  53153=>"101111000",
  53154=>"100000000",
  53155=>"000001111",
  53156=>"000001111",
  53157=>"000111111",
  53158=>"111111111",
  53159=>"000000111",
  53160=>"010000000",
  53161=>"001111001",
  53162=>"111111111",
  53163=>"000000000",
  53164=>"000111111",
  53165=>"111111111",
  53166=>"000000111",
  53167=>"100011111",
  53168=>"101101110",
  53169=>"111000000",
  53170=>"000000001",
  53171=>"011011111",
  53172=>"000000000",
  53173=>"000001001",
  53174=>"111101111",
  53175=>"001001000",
  53176=>"000111001",
  53177=>"000100100",
  53178=>"011000000",
  53179=>"111111111",
  53180=>"100000011",
  53181=>"111111001",
  53182=>"110000011",
  53183=>"111000000",
  53184=>"100101000",
  53185=>"000011000",
  53186=>"000001001",
  53187=>"000111111",
  53188=>"000000100",
  53189=>"110001001",
  53190=>"000000000",
  53191=>"111110000",
  53192=>"111000000",
  53193=>"110110011",
  53194=>"101000000",
  53195=>"111111000",
  53196=>"000100000",
  53197=>"000000001",
  53198=>"000000111",
  53199=>"111000011",
  53200=>"110110111",
  53201=>"000000001",
  53202=>"100000000",
  53203=>"011011011",
  53204=>"101111100",
  53205=>"000001101",
  53206=>"000000000",
  53207=>"000000000",
  53208=>"101111101",
  53209=>"000101101",
  53210=>"011001000",
  53211=>"011111111",
  53212=>"111111011",
  53213=>"001000000",
  53214=>"111100000",
  53215=>"000100111",
  53216=>"011000000",
  53217=>"000000000",
  53218=>"011001000",
  53219=>"001000001",
  53220=>"111010110",
  53221=>"000111111",
  53222=>"000000000",
  53223=>"000000000",
  53224=>"000000000",
  53225=>"000000100",
  53226=>"000000000",
  53227=>"100110100",
  53228=>"001000000",
  53229=>"100000000",
  53230=>"000000101",
  53231=>"111011111",
  53232=>"000000000",
  53233=>"111111111",
  53234=>"000100100",
  53235=>"000000111",
  53236=>"011001000",
  53237=>"000000000",
  53238=>"000000000",
  53239=>"111111001",
  53240=>"011111010",
  53241=>"101001000",
  53242=>"000100111",
  53243=>"110000001",
  53244=>"110110111",
  53245=>"000000000",
  53246=>"111111111",
  53247=>"111111111",
  53248=>"010000010",
  53249=>"000000110",
  53250=>"111111111",
  53251=>"000000000",
  53252=>"101001000",
  53253=>"000000000",
  53254=>"001011001",
  53255=>"110000111",
  53256=>"000000011",
  53257=>"111111000",
  53258=>"011001101",
  53259=>"000111101",
  53260=>"000000000",
  53261=>"111111111",
  53262=>"000010000",
  53263=>"000011011",
  53264=>"000000100",
  53265=>"010011001",
  53266=>"000011111",
  53267=>"100000000",
  53268=>"111111111",
  53269=>"000000001",
  53270=>"001011011",
  53271=>"000000000",
  53272=>"111111111",
  53273=>"000011111",
  53274=>"000000000",
  53275=>"000111111",
  53276=>"000000111",
  53277=>"111111111",
  53278=>"100110000",
  53279=>"010000000",
  53280=>"111111111",
  53281=>"111111101",
  53282=>"110110110",
  53283=>"010010110",
  53284=>"111111000",
  53285=>"000000111",
  53286=>"111110100",
  53287=>"111000000",
  53288=>"101101011",
  53289=>"111111111",
  53290=>"111111111",
  53291=>"111111110",
  53292=>"000000000",
  53293=>"000000000",
  53294=>"000000000",
  53295=>"100111000",
  53296=>"111100110",
  53297=>"000011000",
  53298=>"000000000",
  53299=>"111001000",
  53300=>"111101000",
  53301=>"111011011",
  53302=>"011000000",
  53303=>"111111111",
  53304=>"000000010",
  53305=>"010000000",
  53306=>"111111111",
  53307=>"111111111",
  53308=>"111001000",
  53309=>"111111111",
  53310=>"000100100",
  53311=>"111000000",
  53312=>"000000000",
  53313=>"101111000",
  53314=>"111111111",
  53315=>"111101001",
  53316=>"000000011",
  53317=>"000011011",
  53318=>"000000000",
  53319=>"001001001",
  53320=>"111111111",
  53321=>"001000000",
  53322=>"000000000",
  53323=>"111111000",
  53324=>"000000000",
  53325=>"000000000",
  53326=>"101101001",
  53327=>"000000000",
  53328=>"000011111",
  53329=>"000000000",
  53330=>"111111000",
  53331=>"001001111",
  53332=>"001000000",
  53333=>"111111011",
  53334=>"100001111",
  53335=>"000000000",
  53336=>"111111111",
  53337=>"001000000",
  53338=>"111111111",
  53339=>"000000000",
  53340=>"000101100",
  53341=>"000111001",
  53342=>"111111001",
  53343=>"111010000",
  53344=>"100000000",
  53345=>"111100000",
  53346=>"111000000",
  53347=>"000000000",
  53348=>"000010000",
  53349=>"011001001",
  53350=>"011000000",
  53351=>"000000000",
  53352=>"111111111",
  53353=>"110111110",
  53354=>"001000000",
  53355=>"110111000",
  53356=>"001000010",
  53357=>"000000000",
  53358=>"000000111",
  53359=>"000000111",
  53360=>"000000000",
  53361=>"111000111",
  53362=>"000100100",
  53363=>"111110000",
  53364=>"000000000",
  53365=>"011011000",
  53366=>"101111111",
  53367=>"001001111",
  53368=>"000111111",
  53369=>"000110100",
  53370=>"000000110",
  53371=>"000000000",
  53372=>"110100110",
  53373=>"011011000",
  53374=>"000001111",
  53375=>"000000000",
  53376=>"000000000",
  53377=>"111110000",
  53378=>"111111011",
  53379=>"100000001",
  53380=>"000100100",
  53381=>"101000000",
  53382=>"000000000",
  53383=>"000000000",
  53384=>"000110011",
  53385=>"000000000",
  53386=>"101101101",
  53387=>"011111011",
  53388=>"111100111",
  53389=>"001010000",
  53390=>"111111111",
  53391=>"000000000",
  53392=>"000000100",
  53393=>"111100000",
  53394=>"000000000",
  53395=>"110110110",
  53396=>"110000000",
  53397=>"000110111",
  53398=>"000011111",
  53399=>"111100110",
  53400=>"000000000",
  53401=>"000000000",
  53402=>"110111111",
  53403=>"111111101",
  53404=>"110111111",
  53405=>"000000110",
  53406=>"111111111",
  53407=>"000000111",
  53408=>"111111111",
  53409=>"011011011",
  53410=>"111111111",
  53411=>"111111111",
  53412=>"000000001",
  53413=>"111111111",
  53414=>"100100000",
  53415=>"110010010",
  53416=>"011011011",
  53417=>"000011000",
  53418=>"111010000",
  53419=>"010010000",
  53420=>"111111000",
  53421=>"110111101",
  53422=>"110111111",
  53423=>"011000100",
  53424=>"111111111",
  53425=>"111011000",
  53426=>"111111111",
  53427=>"111111111",
  53428=>"011111111",
  53429=>"010011000",
  53430=>"010000000",
  53431=>"111111100",
  53432=>"111111111",
  53433=>"111111111",
  53434=>"010000000",
  53435=>"010000000",
  53436=>"000111111",
  53437=>"001011001",
  53438=>"000000000",
  53439=>"001111011",
  53440=>"111111111",
  53441=>"001101111",
  53442=>"000000001",
  53443=>"000000000",
  53444=>"000110000",
  53445=>"000000000",
  53446=>"110000000",
  53447=>"111100100",
  53448=>"000111111",
  53449=>"000000000",
  53450=>"000000000",
  53451=>"111100100",
  53452=>"111111110",
  53453=>"111111111",
  53454=>"111001111",
  53455=>"111001000",
  53456=>"010011111",
  53457=>"000000100",
  53458=>"110010111",
  53459=>"000000000",
  53460=>"111101101",
  53461=>"111110100",
  53462=>"000111111",
  53463=>"111111111",
  53464=>"110000000",
  53465=>"000000000",
  53466=>"000000000",
  53467=>"011111001",
  53468=>"111111110",
  53469=>"111111111",
  53470=>"111111111",
  53471=>"000000000",
  53472=>"111111111",
  53473=>"110111011",
  53474=>"000000000",
  53475=>"111111111",
  53476=>"000110000",
  53477=>"000000000",
  53478=>"011011011",
  53479=>"110110111",
  53480=>"110111000",
  53481=>"111111111",
  53482=>"001000111",
  53483=>"111111111",
  53484=>"000000000",
  53485=>"000000000",
  53486=>"100000000",
  53487=>"000000000",
  53488=>"101001011",
  53489=>"000001001",
  53490=>"000000000",
  53491=>"100100000",
  53492=>"011011000",
  53493=>"000000000",
  53494=>"110111001",
  53495=>"111111111",
  53496=>"000001000",
  53497=>"011111111",
  53498=>"111111011",
  53499=>"000000011",
  53500=>"000000000",
  53501=>"000000000",
  53502=>"111001001",
  53503=>"000000000",
  53504=>"111111000",
  53505=>"011011010",
  53506=>"100000101",
  53507=>"111111111",
  53508=>"001111000",
  53509=>"111110111",
  53510=>"110100000",
  53511=>"111011100",
  53512=>"111111000",
  53513=>"100111111",
  53514=>"011111111",
  53515=>"100101111",
  53516=>"001001001",
  53517=>"101111111",
  53518=>"100000110",
  53519=>"111011000",
  53520=>"000011000",
  53521=>"000000001",
  53522=>"111111111",
  53523=>"110111111",
  53524=>"000001010",
  53525=>"011010011",
  53526=>"110110100",
  53527=>"000000000",
  53528=>"111011111",
  53529=>"111001101",
  53530=>"111011101",
  53531=>"000000000",
  53532=>"100100100",
  53533=>"000001111",
  53534=>"001111111",
  53535=>"101100111",
  53536=>"000100100",
  53537=>"011111111",
  53538=>"111100111",
  53539=>"111001111",
  53540=>"000010111",
  53541=>"111111111",
  53542=>"000000000",
  53543=>"000000011",
  53544=>"000000111",
  53545=>"000001001",
  53546=>"111000111",
  53547=>"100111001",
  53548=>"011011000",
  53549=>"000000000",
  53550=>"111111111",
  53551=>"011011000",
  53552=>"011111011",
  53553=>"111111110",
  53554=>"000000000",
  53555=>"010011111",
  53556=>"001011010",
  53557=>"000000001",
  53558=>"000000000",
  53559=>"011000000",
  53560=>"010010010",
  53561=>"111101111",
  53562=>"000101100",
  53563=>"001111111",
  53564=>"111110100",
  53565=>"111111111",
  53566=>"000000000",
  53567=>"111000000",
  53568=>"000000000",
  53569=>"101111111",
  53570=>"111111001",
  53571=>"000000100",
  53572=>"110110110",
  53573=>"111011010",
  53574=>"000010000",
  53575=>"010000000",
  53576=>"100000000",
  53577=>"111011011",
  53578=>"000000111",
  53579=>"000000000",
  53580=>"000011000",
  53581=>"001001001",
  53582=>"111111111",
  53583=>"000000000",
  53584=>"011010100",
  53585=>"111111111",
  53586=>"111111100",
  53587=>"111111111",
  53588=>"000111111",
  53589=>"011011011",
  53590=>"000000000",
  53591=>"111011000",
  53592=>"011111111",
  53593=>"000000001",
  53594=>"111100000",
  53595=>"000101100",
  53596=>"000111111",
  53597=>"111111100",
  53598=>"111010110",
  53599=>"000001111",
  53600=>"000000000",
  53601=>"000000000",
  53602=>"011000000",
  53603=>"001101111",
  53604=>"000010010",
  53605=>"000000000",
  53606=>"000000000",
  53607=>"111111111",
  53608=>"100110100",
  53609=>"000000000",
  53610=>"110100100",
  53611=>"000000000",
  53612=>"000001001",
  53613=>"011011111",
  53614=>"000001000",
  53615=>"000010000",
  53616=>"111001000",
  53617=>"000000000",
  53618=>"000001101",
  53619=>"111100101",
  53620=>"011011000",
  53621=>"111111111",
  53622=>"111000000",
  53623=>"000010000",
  53624=>"000000000",
  53625=>"000000000",
  53626=>"000000000",
  53627=>"000110111",
  53628=>"000000010",
  53629=>"000000110",
  53630=>"000010000",
  53631=>"111000111",
  53632=>"111111111",
  53633=>"000100111",
  53634=>"000011011",
  53635=>"000000000",
  53636=>"111000000",
  53637=>"111111111",
  53638=>"000000000",
  53639=>"110110111",
  53640=>"111110110",
  53641=>"111000000",
  53642=>"000000000",
  53643=>"111111110",
  53644=>"111111111",
  53645=>"000100000",
  53646=>"101111111",
  53647=>"000000000",
  53648=>"000000000",
  53649=>"111111111",
  53650=>"111111111",
  53651=>"000010111",
  53652=>"000000000",
  53653=>"000000000",
  53654=>"000000000",
  53655=>"000000000",
  53656=>"011111111",
  53657=>"110110110",
  53658=>"000000000",
  53659=>"111111111",
  53660=>"111111000",
  53661=>"111110011",
  53662=>"000000000",
  53663=>"000000000",
  53664=>"000011011",
  53665=>"010010111",
  53666=>"100101111",
  53667=>"000000000",
  53668=>"111001111",
  53669=>"111111110",
  53670=>"111111111",
  53671=>"110111111",
  53672=>"010110111",
  53673=>"000000110",
  53674=>"000000000",
  53675=>"110101101",
  53676=>"000011111",
  53677=>"110111111",
  53678=>"010010110",
  53679=>"000000100",
  53680=>"111111000",
  53681=>"100101100",
  53682=>"000111111",
  53683=>"001001011",
  53684=>"111111111",
  53685=>"000000000",
  53686=>"111111111",
  53687=>"000000000",
  53688=>"000011111",
  53689=>"000000100",
  53690=>"000000000",
  53691=>"001001011",
  53692=>"000111111",
  53693=>"000000100",
  53694=>"100000000",
  53695=>"110011111",
  53696=>"100000000",
  53697=>"000000000",
  53698=>"111011011",
  53699=>"111000000",
  53700=>"111111011",
  53701=>"111110110",
  53702=>"000000000",
  53703=>"000000111",
  53704=>"001000000",
  53705=>"111110000",
  53706=>"000000001",
  53707=>"000000011",
  53708=>"000000000",
  53709=>"000100000",
  53710=>"000000000",
  53711=>"100110111",
  53712=>"000011111",
  53713=>"001001101",
  53714=>"011111111",
  53715=>"100000000",
  53716=>"011000010",
  53717=>"011111111",
  53718=>"000100000",
  53719=>"000000000",
  53720=>"111000000",
  53721=>"000111111",
  53722=>"001011011",
  53723=>"111010000",
  53724=>"000001001",
  53725=>"111111111",
  53726=>"111011111",
  53727=>"011011000",
  53728=>"010000110",
  53729=>"111111111",
  53730=>"000000001",
  53731=>"110100111",
  53732=>"000000000",
  53733=>"000000000",
  53734=>"111111000",
  53735=>"111111111",
  53736=>"100111111",
  53737=>"000000000",
  53738=>"111100100",
  53739=>"000000000",
  53740=>"000001111",
  53741=>"000000000",
  53742=>"100101111",
  53743=>"011111100",
  53744=>"011011000",
  53745=>"111111111",
  53746=>"111111111",
  53747=>"100110110",
  53748=>"011001111",
  53749=>"111001001",
  53750=>"000000000",
  53751=>"000000000",
  53752=>"000000000",
  53753=>"001001001",
  53754=>"001011000",
  53755=>"111111111",
  53756=>"111000000",
  53757=>"111111110",
  53758=>"011110000",
  53759=>"000000000",
  53760=>"000000110",
  53761=>"000000000",
  53762=>"111111111",
  53763=>"111110000",
  53764=>"111111111",
  53765=>"000000000",
  53766=>"111000000",
  53767=>"111111111",
  53768=>"000000111",
  53769=>"000011111",
  53770=>"101111011",
  53771=>"111110000",
  53772=>"000000000",
  53773=>"111110110",
  53774=>"111011000",
  53775=>"000000110",
  53776=>"111100000",
  53777=>"110111110",
  53778=>"001000110",
  53779=>"000000100",
  53780=>"000000111",
  53781=>"111101111",
  53782=>"000000111",
  53783=>"100110100",
  53784=>"111100101",
  53785=>"111111111",
  53786=>"001111111",
  53787=>"111111011",
  53788=>"000000000",
  53789=>"000000000",
  53790=>"000000000",
  53791=>"111001001",
  53792=>"010010000",
  53793=>"000100100",
  53794=>"001001111",
  53795=>"111110010",
  53796=>"111011000",
  53797=>"111111111",
  53798=>"000000000",
  53799=>"001111111",
  53800=>"100000001",
  53801=>"000111101",
  53802=>"101101111",
  53803=>"111111111",
  53804=>"000100111",
  53805=>"010111011",
  53806=>"001000111",
  53807=>"100000111",
  53808=>"111110100",
  53809=>"010000000",
  53810=>"000000000",
  53811=>"101101111",
  53812=>"001111001",
  53813=>"000010000",
  53814=>"100000000",
  53815=>"111111000",
  53816=>"000011011",
  53817=>"100000100",
  53818=>"101000000",
  53819=>"100100100",
  53820=>"111100000",
  53821=>"101000001",
  53822=>"011011011",
  53823=>"000000101",
  53824=>"111101001",
  53825=>"010111111",
  53826=>"111111100",
  53827=>"000000111",
  53828=>"000000000",
  53829=>"111111110",
  53830=>"111101101",
  53831=>"101111111",
  53832=>"000000000",
  53833=>"111001000",
  53834=>"000000101",
  53835=>"100100000",
  53836=>"001000111",
  53837=>"111100000",
  53838=>"000000000",
  53839=>"110111010",
  53840=>"100100110",
  53841=>"001100000",
  53842=>"110101111",
  53843=>"110110000",
  53844=>"000000000",
  53845=>"111111111",
  53846=>"100000111",
  53847=>"100110111",
  53848=>"111111111",
  53849=>"110000000",
  53850=>"000000000",
  53851=>"110100110",
  53852=>"000000000",
  53853=>"111111101",
  53854=>"110100111",
  53855=>"000001001",
  53856=>"000000000",
  53857=>"111111000",
  53858=>"000000000",
  53859=>"000100100",
  53860=>"110110100",
  53861=>"101100011",
  53862=>"000000001",
  53863=>"101101011",
  53864=>"111001000",
  53865=>"111111000",
  53866=>"111000110",
  53867=>"000000000",
  53868=>"110110000",
  53869=>"111001000",
  53870=>"000000000",
  53871=>"111111001",
  53872=>"100000111",
  53873=>"111111111",
  53874=>"011111101",
  53875=>"100000010",
  53876=>"111111111",
  53877=>"111111000",
  53878=>"100000100",
  53879=>"000011000",
  53880=>"000000000",
  53881=>"000110111",
  53882=>"100000000",
  53883=>"111111000",
  53884=>"000000100",
  53885=>"111111101",
  53886=>"000000000",
  53887=>"111111000",
  53888=>"001001111",
  53889=>"010011111",
  53890=>"111111101",
  53891=>"111010010",
  53892=>"111111111",
  53893=>"100000101",
  53894=>"000000000",
  53895=>"000000100",
  53896=>"000001111",
  53897=>"100000111",
  53898=>"110110000",
  53899=>"000011001",
  53900=>"100001111",
  53901=>"111111001",
  53902=>"011111111",
  53903=>"111111000",
  53904=>"100100000",
  53905=>"111111111",
  53906=>"111111000",
  53907=>"001111000",
  53908=>"110110110",
  53909=>"111111000",
  53910=>"001011111",
  53911=>"001000000",
  53912=>"111101000",
  53913=>"100111000",
  53914=>"100110111",
  53915=>"000000000",
  53916=>"111111111",
  53917=>"000000010",
  53918=>"001000000",
  53919=>"100000000",
  53920=>"111111111",
  53921=>"001001000",
  53922=>"111001101",
  53923=>"110100000",
  53924=>"000000000",
  53925=>"111110000",
  53926=>"111111100",
  53927=>"000000001",
  53928=>"111111111",
  53929=>"000110110",
  53930=>"000010000",
  53931=>"111010000",
  53932=>"001110110",
  53933=>"000001001",
  53934=>"111110110",
  53935=>"000000111",
  53936=>"000111010",
  53937=>"110010111",
  53938=>"111111100",
  53939=>"111101000",
  53940=>"110000000",
  53941=>"010110111",
  53942=>"000001011",
  53943=>"111111111",
  53944=>"000000010",
  53945=>"001000110",
  53946=>"100110111",
  53947=>"010110111",
  53948=>"100000100",
  53949=>"011000100",
  53950=>"111101111",
  53951=>"111110111",
  53952=>"000000000",
  53953=>"001000000",
  53954=>"010010000",
  53955=>"000000110",
  53956=>"101100110",
  53957=>"001000000",
  53958=>"010111111",
  53959=>"011011011",
  53960=>"100100111",
  53961=>"000000010",
  53962=>"011000000",
  53963=>"000000000",
  53964=>"100100110",
  53965=>"100100000",
  53966=>"111110110",
  53967=>"110000110",
  53968=>"001000000",
  53969=>"000011111",
  53970=>"000000000",
  53971=>"100000000",
  53972=>"111101000",
  53973=>"111111111",
  53974=>"000000001",
  53975=>"111111000",
  53976=>"001011010",
  53977=>"000000110",
  53978=>"111111111",
  53979=>"111111111",
  53980=>"000000100",
  53981=>"111101000",
  53982=>"000111111",
  53983=>"111011011",
  53984=>"000000000",
  53985=>"000110111",
  53986=>"111111000",
  53987=>"111111111",
  53988=>"110111001",
  53989=>"111001011",
  53990=>"110100100",
  53991=>"101001111",
  53992=>"000000110",
  53993=>"000100111",
  53994=>"101101111",
  53995=>"000011011",
  53996=>"000000001",
  53997=>"011111111",
  53998=>"000000110",
  53999=>"000000000",
  54000=>"000100111",
  54001=>"101101001",
  54002=>"000000000",
  54003=>"001001011",
  54004=>"111111110",
  54005=>"100010000",
  54006=>"111101000",
  54007=>"111111000",
  54008=>"111111000",
  54009=>"111111111",
  54010=>"000000111",
  54011=>"100101101",
  54012=>"001101111",
  54013=>"110110000",
  54014=>"100110101",
  54015=>"111100001",
  54016=>"001000100",
  54017=>"000000011",
  54018=>"111111010",
  54019=>"110111111",
  54020=>"001000101",
  54021=>"011010000",
  54022=>"110110110",
  54023=>"010011010",
  54024=>"000000110",
  54025=>"011011010",
  54026=>"000000001",
  54027=>"111111000",
  54028=>"110110110",
  54029=>"101001001",
  54030=>"111111111",
  54031=>"111110110",
  54032=>"111111100",
  54033=>"000000000",
  54034=>"101100100",
  54035=>"001000001",
  54036=>"100110111",
  54037=>"000110000",
  54038=>"011110111",
  54039=>"000100111",
  54040=>"000010110",
  54041=>"011011000",
  54042=>"101101111",
  54043=>"000000100",
  54044=>"000011001",
  54045=>"111111100",
  54046=>"000000000",
  54047=>"000000000",
  54048=>"000000000",
  54049=>"000000000",
  54050=>"111111011",
  54051=>"011001000",
  54052=>"000100110",
  54053=>"000000000",
  54054=>"010110000",
  54055=>"111111111",
  54056=>"111111110",
  54057=>"111111111",
  54058=>"111011111",
  54059=>"101101111",
  54060=>"111110111",
  54061=>"011011111",
  54062=>"111000000",
  54063=>"111111111",
  54064=>"111001111",
  54065=>"111001000",
  54066=>"111111010",
  54067=>"000000111",
  54068=>"011101001",
  54069=>"000001001",
  54070=>"000000110",
  54071=>"100101111",
  54072=>"000111111",
  54073=>"111101000",
  54074=>"000000000",
  54075=>"000101111",
  54076=>"111110000",
  54077=>"111001000",
  54078=>"000000000",
  54079=>"111111110",
  54080=>"001000000",
  54081=>"111111000",
  54082=>"001000100",
  54083=>"001000101",
  54084=>"000000000",
  54085=>"001001111",
  54086=>"000000111",
  54087=>"101101111",
  54088=>"110111000",
  54089=>"000000000",
  54090=>"111111001",
  54091=>"000000000",
  54092=>"111111011",
  54093=>"000000110",
  54094=>"000000010",
  54095=>"000110110",
  54096=>"011011011",
  54097=>"111110001",
  54098=>"111100001",
  54099=>"111111111",
  54100=>"101101111",
  54101=>"011011001",
  54102=>"010010011",
  54103=>"111001001",
  54104=>"000000111",
  54105=>"010000000",
  54106=>"111111111",
  54107=>"111110000",
  54108=>"000000000",
  54109=>"000000101",
  54110=>"000010010",
  54111=>"000001001",
  54112=>"111011001",
  54113=>"000000111",
  54114=>"000010001",
  54115=>"111111111",
  54116=>"000111111",
  54117=>"000000000",
  54118=>"000010000",
  54119=>"001000100",
  54120=>"001000010",
  54121=>"000000101",
  54122=>"000000000",
  54123=>"100001011",
  54124=>"111111110",
  54125=>"100100101",
  54126=>"000100000",
  54127=>"000000000",
  54128=>"000000000",
  54129=>"000000000",
  54130=>"010010011",
  54131=>"000000011",
  54132=>"000000000",
  54133=>"111011111",
  54134=>"100000000",
  54135=>"000000111",
  54136=>"000001001",
  54137=>"100110110",
  54138=>"001111110",
  54139=>"111111110",
  54140=>"000000000",
  54141=>"111111010",
  54142=>"111110110",
  54143=>"000000000",
  54144=>"111111111",
  54145=>"100000000",
  54146=>"100100100",
  54147=>"000101001",
  54148=>"111110100",
  54149=>"110111111",
  54150=>"100111100",
  54151=>"111111111",
  54152=>"101101110",
  54153=>"101000001",
  54154=>"110000000",
  54155=>"000000011",
  54156=>"111100100",
  54157=>"000001001",
  54158=>"000000000",
  54159=>"100100110",
  54160=>"000001001",
  54161=>"111111101",
  54162=>"100110111",
  54163=>"001011001",
  54164=>"000000000",
  54165=>"000000000",
  54166=>"100000000",
  54167=>"000001001",
  54168=>"111011000",
  54169=>"100100100",
  54170=>"000001001",
  54171=>"111011001",
  54172=>"111011111",
  54173=>"110111101",
  54174=>"110111110",
  54175=>"000100111",
  54176=>"000001000",
  54177=>"000011101",
  54178=>"111011011",
  54179=>"100100100",
  54180=>"111111000",
  54181=>"000000000",
  54182=>"010000111",
  54183=>"000000000",
  54184=>"110100110",
  54185=>"000000100",
  54186=>"111110000",
  54187=>"000000000",
  54188=>"111111010",
  54189=>"101111011",
  54190=>"111111111",
  54191=>"111110100",
  54192=>"101100100",
  54193=>"111000000",
  54194=>"000010110",
  54195=>"101111101",
  54196=>"100111111",
  54197=>"100000111",
  54198=>"000000111",
  54199=>"011011111",
  54200=>"000000101",
  54201=>"101101100",
  54202=>"000000001",
  54203=>"101000000",
  54204=>"100101101",
  54205=>"111111110",
  54206=>"000000000",
  54207=>"000000000",
  54208=>"000000000",
  54209=>"111111111",
  54210=>"000000000",
  54211=>"000000000",
  54212=>"000000111",
  54213=>"100000111",
  54214=>"000010110",
  54215=>"000111011",
  54216=>"111111110",
  54217=>"111111100",
  54218=>"101000101",
  54219=>"001011111",
  54220=>"011010010",
  54221=>"000000000",
  54222=>"100001011",
  54223=>"111111111",
  54224=>"100111000",
  54225=>"111000110",
  54226=>"000011101",
  54227=>"111111111",
  54228=>"000000000",
  54229=>"000001100",
  54230=>"000000001",
  54231=>"100100000",
  54232=>"110111111",
  54233=>"000010111",
  54234=>"111110100",
  54235=>"000000001",
  54236=>"111101010",
  54237=>"111110110",
  54238=>"000000101",
  54239=>"100000000",
  54240=>"000000001",
  54241=>"110111111",
  54242=>"100111000",
  54243=>"010011010",
  54244=>"110110011",
  54245=>"000010110",
  54246=>"000000001",
  54247=>"001101111",
  54248=>"011001000",
  54249=>"000000000",
  54250=>"000000011",
  54251=>"111111000",
  54252=>"100000000",
  54253=>"100110111",
  54254=>"001000101",
  54255=>"010010000",
  54256=>"000100000",
  54257=>"000111111",
  54258=>"111111000",
  54259=>"110111111",
  54260=>"000000111",
  54261=>"001000000",
  54262=>"000001101",
  54263=>"000000111",
  54264=>"011111000",
  54265=>"000000100",
  54266=>"001001011",
  54267=>"000100000",
  54268=>"001011110",
  54269=>"101010111",
  54270=>"101001000",
  54271=>"100100111",
  54272=>"111011111",
  54273=>"000111111",
  54274=>"001000000",
  54275=>"111000000",
  54276=>"000000111",
  54277=>"111100000",
  54278=>"111000000",
  54279=>"000000111",
  54280=>"100100100",
  54281=>"001001000",
  54282=>"110110000",
  54283=>"000000000",
  54284=>"111111000",
  54285=>"111001000",
  54286=>"000000000",
  54287=>"000000000",
  54288=>"001001000",
  54289=>"000110111",
  54290=>"100100010",
  54291=>"000011111",
  54292=>"000111111",
  54293=>"111111100",
  54294=>"111000000",
  54295=>"011011011",
  54296=>"000000000",
  54297=>"110000000",
  54298=>"000111111",
  54299=>"110111111",
  54300=>"100100000",
  54301=>"001011001",
  54302=>"011000100",
  54303=>"110110111",
  54304=>"100000000",
  54305=>"110000000",
  54306=>"111111111",
  54307=>"111111111",
  54308=>"010011011",
  54309=>"000111111",
  54310=>"000110110",
  54311=>"100000101",
  54312=>"101000000",
  54313=>"111111111",
  54314=>"010111111",
  54315=>"111111111",
  54316=>"111111011",
  54317=>"111111000",
  54318=>"101111111",
  54319=>"000111100",
  54320=>"001000000",
  54321=>"000011000",
  54322=>"110100000",
  54323=>"000000000",
  54324=>"011111111",
  54325=>"111001011",
  54326=>"100010010",
  54327=>"101101001",
  54328=>"100110111",
  54329=>"111111111",
  54330=>"111111111",
  54331=>"110111111",
  54332=>"000000000",
  54333=>"001101101",
  54334=>"000000000",
  54335=>"100101111",
  54336=>"111011000",
  54337=>"011011010",
  54338=>"000000000",
  54339=>"001001000",
  54340=>"001000000",
  54341=>"100110110",
  54342=>"001001011",
  54343=>"000000110",
  54344=>"000000000",
  54345=>"000000111",
  54346=>"000000000",
  54347=>"000000100",
  54348=>"011011011",
  54349=>"111111100",
  54350=>"000000000",
  54351=>"100111111",
  54352=>"100110111",
  54353=>"001111011",
  54354=>"000111111",
  54355=>"000000000",
  54356=>"000000000",
  54357=>"100111100",
  54358=>"000000000",
  54359=>"110000000",
  54360=>"001101111",
  54361=>"000101111",
  54362=>"111101100",
  54363=>"111011111",
  54364=>"111111011",
  54365=>"100000000",
  54366=>"100111111",
  54367=>"000000000",
  54368=>"111111111",
  54369=>"111111111",
  54370=>"110100100",
  54371=>"111111000",
  54372=>"000000000",
  54373=>"101000010",
  54374=>"000111111",
  54375=>"000000100",
  54376=>"111111111",
  54377=>"111100111",
  54378=>"111111111",
  54379=>"000000000",
  54380=>"000000001",
  54381=>"000111111",
  54382=>"000001001",
  54383=>"111111011",
  54384=>"000010000",
  54385=>"000000000",
  54386=>"011111110",
  54387=>"000000000",
  54388=>"000000100",
  54389=>"101101101",
  54390=>"000000101",
  54391=>"011111111",
  54392=>"100000000",
  54393=>"010111110",
  54394=>"110110011",
  54395=>"010000000",
  54396=>"100000000",
  54397=>"000000000",
  54398=>"011111111",
  54399=>"110010010",
  54400=>"100000000",
  54401=>"111001001",
  54402=>"111011011",
  54403=>"000000000",
  54404=>"111111111",
  54405=>"011111100",
  54406=>"000111001",
  54407=>"110000000",
  54408=>"111111000",
  54409=>"110000000",
  54410=>"101001000",
  54411=>"000111111",
  54412=>"100111100",
  54413=>"000000000",
  54414=>"111111000",
  54415=>"010111111",
  54416=>"000000000",
  54417=>"010000000",
  54418=>"000000000",
  54419=>"010000000",
  54420=>"000000000",
  54421=>"111001001",
  54422=>"111111110",
  54423=>"000000011",
  54424=>"101100111",
  54425=>"000010000",
  54426=>"000000000",
  54427=>"100001000",
  54428=>"000000001",
  54429=>"110110000",
  54430=>"111010010",
  54431=>"111111000",
  54432=>"111000000",
  54433=>"110111010",
  54434=>"110100000",
  54435=>"001000101",
  54436=>"111101111",
  54437=>"000100101",
  54438=>"111001000",
  54439=>"101101100",
  54440=>"010000111",
  54441=>"011000000",
  54442=>"000000000",
  54443=>"000001000",
  54444=>"111100101",
  54445=>"100101000",
  54446=>"000000111",
  54447=>"110010011",
  54448=>"000111111",
  54449=>"100100100",
  54450=>"010111010",
  54451=>"111001000",
  54452=>"110110000",
  54453=>"100111110",
  54454=>"111000010",
  54455=>"000000000",
  54456=>"111111111",
  54457=>"111111011",
  54458=>"111100110",
  54459=>"011111111",
  54460=>"000110000",
  54461=>"000111001",
  54462=>"000000101",
  54463=>"111111111",
  54464=>"111100000",
  54465=>"111111111",
  54466=>"011011001",
  54467=>"010011111",
  54468=>"000010111",
  54469=>"111111111",
  54470=>"111111111",
  54471=>"100000100",
  54472=>"111010000",
  54473=>"011011001",
  54474=>"001000000",
  54475=>"011000101",
  54476=>"111111111",
  54477=>"000000100",
  54478=>"100110111",
  54479=>"011111110",
  54480=>"100110110",
  54481=>"000000000",
  54482=>"000000000",
  54483=>"000000110",
  54484=>"101100000",
  54485=>"111111111",
  54486=>"100111111",
  54487=>"000111011",
  54488=>"111101111",
  54489=>"000000011",
  54490=>"111111111",
  54491=>"111111111",
  54492=>"000000100",
  54493=>"100100111",
  54494=>"111111111",
  54495=>"101111111",
  54496=>"110100000",
  54497=>"000111111",
  54498=>"011000000",
  54499=>"100000111",
  54500=>"000110100",
  54501=>"111100111",
  54502=>"011000111",
  54503=>"111111111",
  54504=>"001011001",
  54505=>"111000000",
  54506=>"000000000",
  54507=>"000000011",
  54508=>"000000000",
  54509=>"110111111",
  54510=>"001111111",
  54511=>"111011111",
  54512=>"110000000",
  54513=>"111001001",
  54514=>"000000000",
  54515=>"100000000",
  54516=>"111111111",
  54517=>"011001001",
  54518=>"111001000",
  54519=>"000000000",
  54520=>"111111000",
  54521=>"111111001",
  54522=>"000101111",
  54523=>"101111111",
  54524=>"110100100",
  54525=>"010111011",
  54526=>"000000100",
  54527=>"110111111",
  54528=>"111110111",
  54529=>"000000110",
  54530=>"000000000",
  54531=>"100111011",
  54532=>"111111111",
  54533=>"001001111",
  54534=>"111101111",
  54535=>"000011111",
  54536=>"111111111",
  54537=>"000000111",
  54538=>"100000000",
  54539=>"000000111",
  54540=>"111111111",
  54541=>"001000001",
  54542=>"000100111",
  54543=>"001000000",
  54544=>"000000000",
  54545=>"111110000",
  54546=>"000011000",
  54547=>"000000000",
  54548=>"000000011",
  54549=>"000000000",
  54550=>"111111111",
  54551=>"111111111",
  54552=>"111111011",
  54553=>"100010000",
  54554=>"111111111",
  54555=>"111111111",
  54556=>"000000000",
  54557=>"100101111",
  54558=>"000111111",
  54559=>"100010011",
  54560=>"111001100",
  54561=>"111111111",
  54562=>"000000000",
  54563=>"111110000",
  54564=>"001110110",
  54565=>"000000001",
  54566=>"000110111",
  54567=>"000001011",
  54568=>"000000011",
  54569=>"111111111",
  54570=>"100111111",
  54571=>"000001011",
  54572=>"010000100",
  54573=>"000100000",
  54574=>"010000111",
  54575=>"000000110",
  54576=>"000001001",
  54577=>"000000111",
  54578=>"011000111",
  54579=>"000111111",
  54580=>"111111110",
  54581=>"000000011",
  54582=>"111001111",
  54583=>"000000000",
  54584=>"111110000",
  54585=>"000001011",
  54586=>"111011111",
  54587=>"111000000",
  54588=>"000000000",
  54589=>"100111001",
  54590=>"111001001",
  54591=>"010110110",
  54592=>"000000000",
  54593=>"110100000",
  54594=>"100111111",
  54595=>"000001001",
  54596=>"111111111",
  54597=>"111111100",
  54598=>"101111011",
  54599=>"111000000",
  54600=>"011010111",
  54601=>"000000000",
  54602=>"110111111",
  54603=>"110000001",
  54604=>"110100011",
  54605=>"000000000",
  54606=>"111100110",
  54607=>"000111111",
  54608=>"111011000",
  54609=>"000101111",
  54610=>"000001001",
  54611=>"111111110",
  54612=>"111111010",
  54613=>"000000000",
  54614=>"111111111",
  54615=>"111011000",
  54616=>"000000111",
  54617=>"111111000",
  54618=>"101101000",
  54619=>"111001111",
  54620=>"111111000",
  54621=>"110111100",
  54622=>"010011011",
  54623=>"111111001",
  54624=>"010110001",
  54625=>"000001000",
  54626=>"111100000",
  54627=>"111110000",
  54628=>"001001111",
  54629=>"000000000",
  54630=>"101001001",
  54631=>"001111111",
  54632=>"011010111",
  54633=>"111011001",
  54634=>"000010000",
  54635=>"000000000",
  54636=>"000000001",
  54637=>"000100110",
  54638=>"111011010",
  54639=>"111011011",
  54640=>"110110110",
  54641=>"110000000",
  54642=>"000111111",
  54643=>"111111111",
  54644=>"111111111",
  54645=>"000000000",
  54646=>"000000000",
  54647=>"110111111",
  54648=>"111011000",
  54649=>"000000001",
  54650=>"011000000",
  54651=>"111111111",
  54652=>"111011101",
  54653=>"111111001",
  54654=>"110110010",
  54655=>"111000000",
  54656=>"101001000",
  54657=>"100111101",
  54658=>"100100111",
  54659=>"110111111",
  54660=>"110000000",
  54661=>"001011011",
  54662=>"000000111",
  54663=>"000000001",
  54664=>"000001001",
  54665=>"011100111",
  54666=>"000000000",
  54667=>"011011001",
  54668=>"011000001",
  54669=>"111111111",
  54670=>"000000000",
  54671=>"000000000",
  54672=>"000011011",
  54673=>"000000011",
  54674=>"101011000",
  54675=>"110100001",
  54676=>"110110000",
  54677=>"111100110",
  54678=>"000000000",
  54679=>"100000110",
  54680=>"111111111",
  54681=>"000000010",
  54682=>"101000111",
  54683=>"111111111",
  54684=>"000000000",
  54685=>"000110110",
  54686=>"110100110",
  54687=>"000111111",
  54688=>"100110111",
  54689=>"110110111",
  54690=>"100000111",
  54691=>"110000000",
  54692=>"011011011",
  54693=>"101110110",
  54694=>"000000000",
  54695=>"011000001",
  54696=>"000000010",
  54697=>"000000111",
  54698=>"011000000",
  54699=>"011010111",
  54700=>"000111111",
  54701=>"000000001",
  54702=>"111100000",
  54703=>"000000000",
  54704=>"000000000",
  54705=>"011111111",
  54706=>"111000000",
  54707=>"000000110",
  54708=>"111000000",
  54709=>"011010111",
  54710=>"000111111",
  54711=>"000000011",
  54712=>"000000000",
  54713=>"000011000",
  54714=>"100001111",
  54715=>"001000000",
  54716=>"000110111",
  54717=>"000000000",
  54718=>"111111100",
  54719=>"111111111",
  54720=>"000000001",
  54721=>"000000000",
  54722=>"111111111",
  54723=>"000001001",
  54724=>"000000000",
  54725=>"111010001",
  54726=>"000001101",
  54727=>"100000000",
  54728=>"111011111",
  54729=>"001000000",
  54730=>"000000000",
  54731=>"000000000",
  54732=>"001001000",
  54733=>"000110011",
  54734=>"000001001",
  54735=>"110000000",
  54736=>"001000000",
  54737=>"111110111",
  54738=>"111010000",
  54739=>"000010111",
  54740=>"100000000",
  54741=>"111111111",
  54742=>"000110001",
  54743=>"000100100",
  54744=>"111000000",
  54745=>"111000000",
  54746=>"000000000",
  54747=>"110111111",
  54748=>"010000000",
  54749=>"111000000",
  54750=>"111110000",
  54751=>"100100100",
  54752=>"000000000",
  54753=>"111111111",
  54754=>"000000000",
  54755=>"000001111",
  54756=>"000000000",
  54757=>"010010110",
  54758=>"001000001",
  54759=>"000000110",
  54760=>"100111111",
  54761=>"100000000",
  54762=>"111110001",
  54763=>"111000100",
  54764=>"000110111",
  54765=>"001000000",
  54766=>"000001000",
  54767=>"101100000",
  54768=>"000100111",
  54769=>"000000011",
  54770=>"110010010",
  54771=>"000000000",
  54772=>"111111110",
  54773=>"000000000",
  54774=>"111110010",
  54775=>"000000000",
  54776=>"110110000",
  54777=>"111101101",
  54778=>"111111010",
  54779=>"011111111",
  54780=>"000000000",
  54781=>"101001000",
  54782=>"000000000",
  54783=>"111111011",
  54784=>"000000000",
  54785=>"010000000",
  54786=>"000000101",
  54787=>"010110110",
  54788=>"001011011",
  54789=>"000010110",
  54790=>"001000000",
  54791=>"111111111",
  54792=>"011011111",
  54793=>"001001001",
  54794=>"001000000",
  54795=>"000000000",
  54796=>"100100000",
  54797=>"000000101",
  54798=>"010000001",
  54799=>"111111100",
  54800=>"000100100",
  54801=>"110010001",
  54802=>"111111111",
  54803=>"111111110",
  54804=>"001101001",
  54805=>"000001001",
  54806=>"000010110",
  54807=>"000000000",
  54808=>"010110110",
  54809=>"100001000",
  54810=>"100101111",
  54811=>"000110100",
  54812=>"000000000",
  54813=>"011110000",
  54814=>"000000000",
  54815=>"000110110",
  54816=>"111100100",
  54817=>"111110000",
  54818=>"111110110",
  54819=>"111111111",
  54820=>"001001001",
  54821=>"110110110",
  54822=>"001001001",
  54823=>"000000011",
  54824=>"000000000",
  54825=>"111111111",
  54826=>"010000001",
  54827=>"000011111",
  54828=>"111111111",
  54829=>"111111000",
  54830=>"010110110",
  54831=>"000000001",
  54832=>"110100110",
  54833=>"101111001",
  54834=>"000000100",
  54835=>"111111111",
  54836=>"111111000",
  54837=>"110110110",
  54838=>"011001001",
  54839=>"000110110",
  54840=>"110111111",
  54841=>"000111111",
  54842=>"110111111",
  54843=>"111100111",
  54844=>"001001001",
  54845=>"111111111",
  54846=>"001011111",
  54847=>"111111111",
  54848=>"001001000",
  54849=>"001011001",
  54850=>"111001000",
  54851=>"000000000",
  54852=>"100100100",
  54853=>"011000100",
  54854=>"110000000",
  54855=>"000000000",
  54856=>"111111001",
  54857=>"101101101",
  54858=>"110110111",
  54859=>"000000000",
  54860=>"010010000",
  54861=>"000011111",
  54862=>"010010111",
  54863=>"000000001",
  54864=>"000000111",
  54865=>"111111100",
  54866=>"001000001",
  54867=>"110110110",
  54868=>"110111110",
  54869=>"110111011",
  54870=>"000000001",
  54871=>"111111111",
  54872=>"000100111",
  54873=>"101101101",
  54874=>"110111111",
  54875=>"100100100",
  54876=>"001001001",
  54877=>"011011111",
  54878=>"100000000",
  54879=>"111111001",
  54880=>"000001111",
  54881=>"111111110",
  54882=>"000100111",
  54883=>"000000000",
  54884=>"101001000",
  54885=>"111110111",
  54886=>"000110110",
  54887=>"011000000",
  54888=>"000111111",
  54889=>"001010011",
  54890=>"000110010",
  54891=>"110111111",
  54892=>"001000000",
  54893=>"000000000",
  54894=>"000010000",
  54895=>"000000000",
  54896=>"110011111",
  54897=>"110110000",
  54898=>"111111011",
  54899=>"000000110",
  54900=>"000000000",
  54901=>"111000000",
  54902=>"000000001",
  54903=>"111000000",
  54904=>"100100100",
  54905=>"000000000",
  54906=>"111000000",
  54907=>"000000000",
  54908=>"100110100",
  54909=>"110110100",
  54910=>"100100111",
  54911=>"001011001",
  54912=>"101111100",
  54913=>"010110111",
  54914=>"000000000",
  54915=>"111111110",
  54916=>"001001001",
  54917=>"111111111",
  54918=>"000000000",
  54919=>"010000000",
  54920=>"000000000",
  54921=>"011111111",
  54922=>"001001001",
  54923=>"000000000",
  54924=>"000101111",
  54925=>"111111111",
  54926=>"010010111",
  54927=>"000000000",
  54928=>"010110110",
  54929=>"100000000",
  54930=>"010010111",
  54931=>"111011001",
  54932=>"111100111",
  54933=>"001000000",
  54934=>"000000001",
  54935=>"110100100",
  54936=>"001000001",
  54937=>"111111001",
  54938=>"111110000",
  54939=>"000000000",
  54940=>"110111111",
  54941=>"000000000",
  54942=>"100110000",
  54943=>"000000000",
  54944=>"000011111",
  54945=>"110111111",
  54946=>"111111111",
  54947=>"001001101",
  54948=>"111111011",
  54949=>"110010010",
  54950=>"000000000",
  54951=>"111111111",
  54952=>"000000001",
  54953=>"001001001",
  54954=>"101001111",
  54955=>"010000010",
  54956=>"111111101",
  54957=>"000000000",
  54958=>"111100110",
  54959=>"000000101",
  54960=>"010010010",
  54961=>"011110000",
  54962=>"010111010",
  54963=>"110110010",
  54964=>"000000000",
  54965=>"111000000",
  54966=>"000000000",
  54967=>"010110110",
  54968=>"000000100",
  54969=>"111111001",
  54970=>"111001000",
  54971=>"011110110",
  54972=>"001001101",
  54973=>"000000001",
  54974=>"111111111",
  54975=>"101101111",
  54976=>"000000000",
  54977=>"111110110",
  54978=>"111111111",
  54979=>"111010000",
  54980=>"011100111",
  54981=>"000001101",
  54982=>"100000100",
  54983=>"000000001",
  54984=>"000000110",
  54985=>"000111111",
  54986=>"000000001",
  54987=>"101000000",
  54988=>"010011110",
  54989=>"111111111",
  54990=>"000000000",
  54991=>"111000000",
  54992=>"000000000",
  54993=>"001000000",
  54994=>"111101111",
  54995=>"001000000",
  54996=>"000000100",
  54997=>"001000100",
  54998=>"000000000",
  54999=>"001001001",
  55000=>"111111000",
  55001=>"111111111",
  55002=>"001000000",
  55003=>"100101111",
  55004=>"000000000",
  55005=>"000111111",
  55006=>"000001101",
  55007=>"001000000",
  55008=>"000001001",
  55009=>"000011011",
  55010=>"000000000",
  55011=>"111111111",
  55012=>"101111110",
  55013=>"001001011",
  55014=>"111000000",
  55015=>"010010110",
  55016=>"110111111",
  55017=>"000001001",
  55018=>"001011001",
  55019=>"000000000",
  55020=>"011011001",
  55021=>"000000000",
  55022=>"000000001",
  55023=>"001000001",
  55024=>"001100000",
  55025=>"010010111",
  55026=>"110100010",
  55027=>"000010111",
  55028=>"011110010",
  55029=>"111000000",
  55030=>"000111111",
  55031=>"110111010",
  55032=>"111111100",
  55033=>"000000000",
  55034=>"000001000",
  55035=>"100100100",
  55036=>"001001011",
  55037=>"010010110",
  55038=>"000000011",
  55039=>"000000110",
  55040=>"000000000",
  55041=>"000000001",
  55042=>"111001000",
  55043=>"000000111",
  55044=>"000000000",
  55045=>"111000000",
  55046=>"110110111",
  55047=>"000000001",
  55048=>"000000000",
  55049=>"111111111",
  55050=>"011110111",
  55051=>"001101111",
  55052=>"000000000",
  55053=>"111111010",
  55054=>"100110011",
  55055=>"110100000",
  55056=>"000010011",
  55057=>"000011111",
  55058=>"000000000",
  55059=>"010110111",
  55060=>"000000000",
  55061=>"111111111",
  55062=>"111111111",
  55063=>"000100110",
  55064=>"110110110",
  55065=>"111111110",
  55066=>"000000000",
  55067=>"111110111",
  55068=>"000000000",
  55069=>"000100111",
  55070=>"001001001",
  55071=>"111111111",
  55072=>"000000000",
  55073=>"000000000",
  55074=>"110111010",
  55075=>"000000000",
  55076=>"001001000",
  55077=>"000011111",
  55078=>"000000000",
  55079=>"010010000",
  55080=>"001000000",
  55081=>"011111110",
  55082=>"010110110",
  55083=>"000000001",
  55084=>"111111111",
  55085=>"000110110",
  55086=>"011010000",
  55087=>"111111111",
  55088=>"010110110",
  55089=>"111001001",
  55090=>"111111110",
  55091=>"000000010",
  55092=>"000101111",
  55093=>"111101111",
  55094=>"000001111",
  55095=>"000100111",
  55096=>"111101110",
  55097=>"101000000",
  55098=>"111000000",
  55099=>"110011011",
  55100=>"001000100",
  55101=>"000110110",
  55102=>"011000000",
  55103=>"111110101",
  55104=>"000000000",
  55105=>"010110000",
  55106=>"000101000",
  55107=>"001001001",
  55108=>"000001110",
  55109=>"000111111",
  55110=>"001001001",
  55111=>"111111001",
  55112=>"000000000",
  55113=>"001000001",
  55114=>"000000000",
  55115=>"001000001",
  55116=>"000000000",
  55117=>"000001000",
  55118=>"011111100",
  55119=>"100100100",
  55120=>"110000100",
  55121=>"000000000",
  55122=>"111111111",
  55123=>"000001101",
  55124=>"001000000",
  55125=>"001011011",
  55126=>"000000111",
  55127=>"101111111",
  55128=>"011000000",
  55129=>"001000000",
  55130=>"001000000",
  55131=>"000010011",
  55132=>"000000000",
  55133=>"111011010",
  55134=>"110110110",
  55135=>"000000000",
  55136=>"101001001",
  55137=>"000000000",
  55138=>"110000000",
  55139=>"101001001",
  55140=>"000000001",
  55141=>"010011110",
  55142=>"100100111",
  55143=>"000000000",
  55144=>"000000000",
  55145=>"000010010",
  55146=>"001000000",
  55147=>"000110100",
  55148=>"111110100",
  55149=>"001111100",
  55150=>"001001001",
  55151=>"000000000",
  55152=>"000000000",
  55153=>"000000010",
  55154=>"011101111",
  55155=>"010011000",
  55156=>"000000000",
  55157=>"111110111",
  55158=>"111111111",
  55159=>"001011000",
  55160=>"101000001",
  55161=>"000000001",
  55162=>"000101111",
  55163=>"000000000",
  55164=>"000111110",
  55165=>"000000010",
  55166=>"001001000",
  55167=>"001000000",
  55168=>"000001011",
  55169=>"011000001",
  55170=>"111011011",
  55171=>"000000001",
  55172=>"101101101",
  55173=>"110111111",
  55174=>"100000001",
  55175=>"001000000",
  55176=>"000110110",
  55177=>"111111111",
  55178=>"000000001",
  55179=>"000000000",
  55180=>"000000111",
  55181=>"110000000",
  55182=>"100100110",
  55183=>"000000000",
  55184=>"000000000",
  55185=>"111111111",
  55186=>"000011111",
  55187=>"001001001",
  55188=>"000000000",
  55189=>"110000000",
  55190=>"000000000",
  55191=>"101111011",
  55192=>"000000000",
  55193=>"111000111",
  55194=>"111111111",
  55195=>"110110111",
  55196=>"111101001",
  55197=>"000001111",
  55198=>"100100000",
  55199=>"000000000",
  55200=>"000000000",
  55201=>"011011011",
  55202=>"001000001",
  55203=>"110111110",
  55204=>"010000000",
  55205=>"010111001",
  55206=>"001100000",
  55207=>"000111111",
  55208=>"101001001",
  55209=>"000000001",
  55210=>"000000111",
  55211=>"001111000",
  55212=>"000000100",
  55213=>"000000000",
  55214=>"000000001",
  55215=>"000110010",
  55216=>"000111100",
  55217=>"011111100",
  55218=>"000001111",
  55219=>"000011111",
  55220=>"000010000",
  55221=>"111100000",
  55222=>"000000111",
  55223=>"001001111",
  55224=>"000011011",
  55225=>"000000010",
  55226=>"000000011",
  55227=>"111111011",
  55228=>"000000000",
  55229=>"111010000",
  55230=>"000000000",
  55231=>"101000101",
  55232=>"111010010",
  55233=>"110110000",
  55234=>"011011011",
  55235=>"111111000",
  55236=>"110110110",
  55237=>"000000000",
  55238=>"000000000",
  55239=>"111111111",
  55240=>"000001000",
  55241=>"000001000",
  55242=>"000000001",
  55243=>"110111011",
  55244=>"011111010",
  55245=>"000000000",
  55246=>"000000001",
  55247=>"110110111",
  55248=>"111111010",
  55249=>"000000000",
  55250=>"111110110",
  55251=>"000000000",
  55252=>"101000000",
  55253=>"000000101",
  55254=>"000000000",
  55255=>"100000000",
  55256=>"110111111",
  55257=>"000110111",
  55258=>"111101000",
  55259=>"000000101",
  55260=>"111111011",
  55261=>"000000101",
  55262=>"100001101",
  55263=>"100000001",
  55264=>"100000000",
  55265=>"111001000",
  55266=>"010111111",
  55267=>"111110001",
  55268=>"000000000",
  55269=>"000000000",
  55270=>"101111010",
  55271=>"010010000",
  55272=>"111010011",
  55273=>"000000000",
  55274=>"001111000",
  55275=>"010001010",
  55276=>"111011111",
  55277=>"100100111",
  55278=>"111111111",
  55279=>"111001111",
  55280=>"111101000",
  55281=>"111000000",
  55282=>"011111111",
  55283=>"001001001",
  55284=>"000010011",
  55285=>"100100000",
  55286=>"000111011",
  55287=>"000010000",
  55288=>"111111011",
  55289=>"000000000",
  55290=>"011001111",
  55291=>"000001111",
  55292=>"110000011",
  55293=>"000000100",
  55294=>"001011000",
  55295=>"000000000",
  55296=>"000000111",
  55297=>"000000011",
  55298=>"111111111",
  55299=>"010000000",
  55300=>"110111110",
  55301=>"000000000",
  55302=>"111111111",
  55303=>"001001011",
  55304=>"111000100",
  55305=>"111111001",
  55306=>"000000101",
  55307=>"010010000",
  55308=>"000000000",
  55309=>"011111111",
  55310=>"111110111",
  55311=>"000000000",
  55312=>"000000001",
  55313=>"111111011",
  55314=>"111111000",
  55315=>"111000001",
  55316=>"000000000",
  55317=>"000000000",
  55318=>"111111111",
  55319=>"111111111",
  55320=>"111111111",
  55321=>"101100000",
  55322=>"000101111",
  55323=>"011000111",
  55324=>"000000000",
  55325=>"000110110",
  55326=>"111010001",
  55327=>"111000000",
  55328=>"111111011",
  55329=>"111111111",
  55330=>"111110000",
  55331=>"010111110",
  55332=>"110110101",
  55333=>"010000000",
  55334=>"000001011",
  55335=>"100000000",
  55336=>"110000000",
  55337=>"000000111",
  55338=>"111111111",
  55339=>"100000111",
  55340=>"000000100",
  55341=>"000001001",
  55342=>"111111111",
  55343=>"111010000",
  55344=>"000000000",
  55345=>"000000001",
  55346=>"111111110",
  55347=>"111111000",
  55348=>"111011001",
  55349=>"000000000",
  55350=>"111111000",
  55351=>"000000110",
  55352=>"111111001",
  55353=>"111010000",
  55354=>"101100111",
  55355=>"111011000",
  55356=>"100000000",
  55357=>"110110111",
  55358=>"000000000",
  55359=>"000000000",
  55360=>"000100111",
  55361=>"000110010",
  55362=>"000111111",
  55363=>"111111000",
  55364=>"000110000",
  55365=>"000000100",
  55366=>"000000001",
  55367=>"111111111",
  55368=>"000000001",
  55369=>"111100100",
  55370=>"111100111",
  55371=>"110111111",
  55372=>"001000111",
  55373=>"011000110",
  55374=>"111001000",
  55375=>"111101111",
  55376=>"111000000",
  55377=>"111000000",
  55378=>"111111111",
  55379=>"000011111",
  55380=>"000000011",
  55381=>"000100111",
  55382=>"000110000",
  55383=>"001000000",
  55384=>"010110110",
  55385=>"111101101",
  55386=>"011111111",
  55387=>"100111110",
  55388=>"000010111",
  55389=>"000000000",
  55390=>"111111111",
  55391=>"110110110",
  55392=>"110010000",
  55393=>"111111001",
  55394=>"111111100",
  55395=>"110000000",
  55396=>"000000101",
  55397=>"000111111",
  55398=>"000000111",
  55399=>"111001000",
  55400=>"001111111",
  55401=>"000111111",
  55402=>"111000110",
  55403=>"000000000",
  55404=>"000000111",
  55405=>"111111111",
  55406=>"111111111",
  55407=>"111111000",
  55408=>"000111011",
  55409=>"001000000",
  55410=>"000000101",
  55411=>"000100000",
  55412=>"111111111",
  55413=>"110000100",
  55414=>"000000111",
  55415=>"110111101",
  55416=>"100111000",
  55417=>"111111111",
  55418=>"001000000",
  55419=>"111011011",
  55420=>"110110111",
  55421=>"001000111",
  55422=>"110111000",
  55423=>"000000000",
  55424=>"111011000",
  55425=>"000000011",
  55426=>"111101100",
  55427=>"000000111",
  55428=>"111100101",
  55429=>"110111111",
  55430=>"111001111",
  55431=>"111000000",
  55432=>"000000111",
  55433=>"000000000",
  55434=>"100110100",
  55435=>"100000111",
  55436=>"001000000",
  55437=>"000000000",
  55438=>"000000011",
  55439=>"111011000",
  55440=>"111111111",
  55441=>"000000111",
  55442=>"111101000",
  55443=>"000000000",
  55444=>"110100111",
  55445=>"000000000",
  55446=>"001111111",
  55447=>"111111111",
  55448=>"000000000",
  55449=>"000000000",
  55450=>"111111000",
  55451=>"000000110",
  55452=>"001000111",
  55453=>"111111111",
  55454=>"111011010",
  55455=>"000000101",
  55456=>"000000000",
  55457=>"001000111",
  55458=>"110111111",
  55459=>"000011110",
  55460=>"110111000",
  55461=>"000000000",
  55462=>"111111111",
  55463=>"111111111",
  55464=>"001001000",
  55465=>"000000000",
  55466=>"000000000",
  55467=>"101000000",
  55468=>"111111111",
  55469=>"111111111",
  55470=>"000000111",
  55471=>"111111111",
  55472=>"110000000",
  55473=>"111000000",
  55474=>"111011010",
  55475=>"111111000",
  55476=>"111000111",
  55477=>"111111101",
  55478=>"001000111",
  55479=>"111111111",
  55480=>"111111111",
  55481=>"011111111",
  55482=>"000110100",
  55483=>"010000001",
  55484=>"001000000",
  55485=>"001000111",
  55486=>"000000111",
  55487=>"000000000",
  55488=>"111111111",
  55489=>"111101111",
  55490=>"000010111",
  55491=>"111111001",
  55492=>"111000000",
  55493=>"000000000",
  55494=>"111011000",
  55495=>"111111001",
  55496=>"000111111",
  55497=>"000000111",
  55498=>"000000000",
  55499=>"011000000",
  55500=>"000000000",
  55501=>"000000001",
  55502=>"111111111",
  55503=>"111111101",
  55504=>"111111110",
  55505=>"000000000",
  55506=>"000000000",
  55507=>"111101000",
  55508=>"110110000",
  55509=>"000000000",
  55510=>"111111011",
  55511=>"000000000",
  55512=>"000000111",
  55513=>"110111111",
  55514=>"110111111",
  55515=>"110111111",
  55516=>"111111111",
  55517=>"101111111",
  55518=>"000000111",
  55519=>"001101111",
  55520=>"111111111",
  55521=>"001011011",
  55522=>"001000000",
  55523=>"111111111",
  55524=>"111111111",
  55525=>"111111011",
  55526=>"111111111",
  55527=>"000000111",
  55528=>"001111111",
  55529=>"001001001",
  55530=>"100100111",
  55531=>"110100111",
  55532=>"000000000",
  55533=>"010010000",
  55534=>"000000000",
  55535=>"000000000",
  55536=>"000000000",
  55537=>"011000000",
  55538=>"000110111",
  55539=>"000000111",
  55540=>"011000000",
  55541=>"111111111",
  55542=>"011010011",
  55543=>"111111111",
  55544=>"000001001",
  55545=>"100000111",
  55546=>"000000000",
  55547=>"101000000",
  55548=>"011011000",
  55549=>"000000111",
  55550=>"000000000",
  55551=>"111110111",
  55552=>"111100000",
  55553=>"000010000",
  55554=>"011011011",
  55555=>"001001000",
  55556=>"111111111",
  55557=>"001000110",
  55558=>"111101110",
  55559=>"111101111",
  55560=>"111111000",
  55561=>"000001001",
  55562=>"111111101",
  55563=>"111111000",
  55564=>"110100000",
  55565=>"000000101",
  55566=>"110111001",
  55567=>"111111111",
  55568=>"000110000",
  55569=>"011000000",
  55570=>"000000000",
  55571=>"100000100",
  55572=>"101111111",
  55573=>"111111100",
  55574=>"111111001",
  55575=>"000000001",
  55576=>"000000111",
  55577=>"111101101",
  55578=>"110000000",
  55579=>"000110111",
  55580=>"011111100",
  55581=>"111001111",
  55582=>"100111111",
  55583=>"000000000",
  55584=>"000100111",
  55585=>"101111111",
  55586=>"000000110",
  55587=>"111111111",
  55588=>"000000000",
  55589=>"100100100",
  55590=>"001000000",
  55591=>"111101111",
  55592=>"111111111",
  55593=>"111111000",
  55594=>"011111111",
  55595=>"000000000",
  55596=>"000000000",
  55597=>"110110100",
  55598=>"111000010",
  55599=>"101000000",
  55600=>"000000101",
  55601=>"111111011",
  55602=>"000100000",
  55603=>"100100000",
  55604=>"111011111",
  55605=>"000000111",
  55606=>"111000000",
  55607=>"000000000",
  55608=>"111011111",
  55609=>"111111111",
  55610=>"000000111",
  55611=>"000000111",
  55612=>"000000000",
  55613=>"010000000",
  55614=>"000000000",
  55615=>"000000111",
  55616=>"111111000",
  55617=>"111111111",
  55618=>"000000011",
  55619=>"000000000",
  55620=>"000001000",
  55621=>"000000001",
  55622=>"111111111",
  55623=>"001111111",
  55624=>"000000000",
  55625=>"111011000",
  55626=>"000001111",
  55627=>"000000011",
  55628=>"000000000",
  55629=>"000010111",
  55630=>"000011111",
  55631=>"001000000",
  55632=>"001000000",
  55633=>"001000000",
  55634=>"000111111",
  55635=>"000000000",
  55636=>"001001000",
  55637=>"111111011",
  55638=>"000000101",
  55639=>"111111001",
  55640=>"101111111",
  55641=>"001111111",
  55642=>"111100111",
  55643=>"000000111",
  55644=>"000000100",
  55645=>"000000000",
  55646=>"111001001",
  55647=>"000000110",
  55648=>"111111111",
  55649=>"111111111",
  55650=>"001001000",
  55651=>"110000000",
  55652=>"101100100",
  55653=>"101100111",
  55654=>"111111111",
  55655=>"001000000",
  55656=>"000100111",
  55657=>"000000110",
  55658=>"001000000",
  55659=>"000001011",
  55660=>"111111111",
  55661=>"111111000",
  55662=>"111011111",
  55663=>"111101101",
  55664=>"111000000",
  55665=>"000000000",
  55666=>"000000111",
  55667=>"001000000",
  55668=>"000000111",
  55669=>"111101111",
  55670=>"111111001",
  55671=>"111111111",
  55672=>"000000111",
  55673=>"000000111",
  55674=>"001000000",
  55675=>"010010000",
  55676=>"000100100",
  55677=>"100110110",
  55678=>"111011000",
  55679=>"001001001",
  55680=>"110000000",
  55681=>"000011011",
  55682=>"000000001",
  55683=>"000000000",
  55684=>"111000000",
  55685=>"110110000",
  55686=>"000000000",
  55687=>"101001001",
  55688=>"001111111",
  55689=>"111000100",
  55690=>"000000000",
  55691=>"111111111",
  55692=>"111101000",
  55693=>"111000000",
  55694=>"000000000",
  55695=>"111111111",
  55696=>"111111011",
  55697=>"001000100",
  55698=>"000111111",
  55699=>"000001001",
  55700=>"000000110",
  55701=>"000000000",
  55702=>"110110100",
  55703=>"000000100",
  55704=>"110010000",
  55705=>"000010111",
  55706=>"111111000",
  55707=>"000000001",
  55708=>"000000111",
  55709=>"000000000",
  55710=>"111000000",
  55711=>"111111111",
  55712=>"000000111",
  55713=>"011011111",
  55714=>"000000000",
  55715=>"101000011",
  55716=>"111000000",
  55717=>"111111101",
  55718=>"111111111",
  55719=>"000000000",
  55720=>"000000000",
  55721=>"111110000",
  55722=>"000010000",
  55723=>"001000110",
  55724=>"000000000",
  55725=>"111111111",
  55726=>"000110101",
  55727=>"000000001",
  55728=>"010000000",
  55729=>"111111110",
  55730=>"111111111",
  55731=>"000100110",
  55732=>"011111111",
  55733=>"111111111",
  55734=>"110111100",
  55735=>"000000000",
  55736=>"010000110",
  55737=>"111100110",
  55738=>"111000001",
  55739=>"000000101",
  55740=>"000000000",
  55741=>"110000100",
  55742=>"111111111",
  55743=>"011011111",
  55744=>"001101100",
  55745=>"001000111",
  55746=>"111111111",
  55747=>"000111111",
  55748=>"111000111",
  55749=>"101110000",
  55750=>"001000111",
  55751=>"000111111",
  55752=>"000000111",
  55753=>"100111101",
  55754=>"111111111",
  55755=>"111111111",
  55756=>"010000000",
  55757=>"111111111",
  55758=>"110111111",
  55759=>"000000000",
  55760=>"000110000",
  55761=>"011111111",
  55762=>"000100100",
  55763=>"111111111",
  55764=>"000000001",
  55765=>"111111110",
  55766=>"011011000",
  55767=>"000000000",
  55768=>"000000111",
  55769=>"001001111",
  55770=>"100000000",
  55771=>"111110111",
  55772=>"001000001",
  55773=>"001000001",
  55774=>"111111101",
  55775=>"000000000",
  55776=>"000000000",
  55777=>"111111111",
  55778=>"111011001",
  55779=>"001000111",
  55780=>"110000000",
  55781=>"000000000",
  55782=>"000000000",
  55783=>"001000001",
  55784=>"000000001",
  55785=>"001111001",
  55786=>"110110100",
  55787=>"101000101",
  55788=>"000110111",
  55789=>"111011011",
  55790=>"001000000",
  55791=>"000000000",
  55792=>"111101100",
  55793=>"000000000",
  55794=>"101111111",
  55795=>"000110111",
  55796=>"000000001",
  55797=>"111111111",
  55798=>"010111011",
  55799=>"000100111",
  55800=>"111111010",
  55801=>"000000000",
  55802=>"101100111",
  55803=>"110110111",
  55804=>"111111111",
  55805=>"011000000",
  55806=>"111001111",
  55807=>"111111111",
  55808=>"111000000",
  55809=>"110100111",
  55810=>"111000001",
  55811=>"111111111",
  55812=>"111111111",
  55813=>"000000111",
  55814=>"111111100",
  55815=>"000000000",
  55816=>"100111011",
  55817=>"111011011",
  55818=>"011111111",
  55819=>"001000000",
  55820=>"011111111",
  55821=>"100000111",
  55822=>"000100111",
  55823=>"111111111",
  55824=>"000010000",
  55825=>"011111101",
  55826=>"000000000",
  55827=>"111111111",
  55828=>"000000000",
  55829=>"111000000",
  55830=>"000110110",
  55831=>"111100111",
  55832=>"000000001",
  55833=>"001011110",
  55834=>"111111111",
  55835=>"000000101",
  55836=>"011001001",
  55837=>"000110110",
  55838=>"011111111",
  55839=>"000000001",
  55840=>"000000011",
  55841=>"000001011",
  55842=>"111111111",
  55843=>"100101111",
  55844=>"111000110",
  55845=>"000000000",
  55846=>"000010111",
  55847=>"111111111",
  55848=>"000111011",
  55849=>"000100111",
  55850=>"111111111",
  55851=>"100000000",
  55852=>"110000000",
  55853=>"111010010",
  55854=>"000000000",
  55855=>"011011000",
  55856=>"011010001",
  55857=>"111111111",
  55858=>"111111100",
  55859=>"111111111",
  55860=>"000000111",
  55861=>"000100111",
  55862=>"011001000",
  55863=>"001010111",
  55864=>"111111010",
  55865=>"000000111",
  55866=>"000101111",
  55867=>"000000000",
  55868=>"000000000",
  55869=>"001100111",
  55870=>"110111000",
  55871=>"000000000",
  55872=>"110011000",
  55873=>"110000000",
  55874=>"000000011",
  55875=>"000000001",
  55876=>"011001001",
  55877=>"101111100",
  55878=>"111111110",
  55879=>"011111110",
  55880=>"000000000",
  55881=>"111111111",
  55882=>"111111000",
  55883=>"110110000",
  55884=>"000000000",
  55885=>"111111000",
  55886=>"000000100",
  55887=>"000111111",
  55888=>"010111111",
  55889=>"101000000",
  55890=>"111100111",
  55891=>"000001000",
  55892=>"000000000",
  55893=>"000000000",
  55894=>"000000111",
  55895=>"001000000",
  55896=>"111000111",
  55897=>"111100000",
  55898=>"111111000",
  55899=>"000000000",
  55900=>"111000001",
  55901=>"100111000",
  55902=>"111111001",
  55903=>"111111100",
  55904=>"000000100",
  55905=>"101000000",
  55906=>"000000001",
  55907=>"100111111",
  55908=>"111000011",
  55909=>"111011001",
  55910=>"001000000",
  55911=>"111110111",
  55912=>"000111111",
  55913=>"010000000",
  55914=>"111110000",
  55915=>"111000010",
  55916=>"111111111",
  55917=>"000000001",
  55918=>"000001001",
  55919=>"000111111",
  55920=>"000000000",
  55921=>"110110110",
  55922=>"000000001",
  55923=>"111001000",
  55924=>"101101000",
  55925=>"001001100",
  55926=>"111011001",
  55927=>"001000011",
  55928=>"010010000",
  55929=>"111000110",
  55930=>"000000000",
  55931=>"001000000",
  55932=>"011001001",
  55933=>"110011010",
  55934=>"111110000",
  55935=>"000111111",
  55936=>"111111011",
  55937=>"000000000",
  55938=>"000100100",
  55939=>"000100000",
  55940=>"111111111",
  55941=>"000000000",
  55942=>"000111000",
  55943=>"000000111",
  55944=>"111111111",
  55945=>"000001000",
  55946=>"111100000",
  55947=>"111010000",
  55948=>"110000001",
  55949=>"111111111",
  55950=>"110110110",
  55951=>"111011010",
  55952=>"000000000",
  55953=>"000001000",
  55954=>"111011000",
  55955=>"100001111",
  55956=>"010110111",
  55957=>"001001001",
  55958=>"111111111",
  55959=>"000000000",
  55960=>"111000001",
  55961=>"000000000",
  55962=>"111000000",
  55963=>"101101000",
  55964=>"001000110",
  55965=>"101000000",
  55966=>"110111111",
  55967=>"111000100",
  55968=>"011000000",
  55969=>"111100101",
  55970=>"110101101",
  55971=>"111000000",
  55972=>"001111000",
  55973=>"111111111",
  55974=>"111011111",
  55975=>"000000000",
  55976=>"000000000",
  55977=>"000000000",
  55978=>"111001111",
  55979=>"100110000",
  55980=>"000000010",
  55981=>"110110110",
  55982=>"010000110",
  55983=>"010101100",
  55984=>"111111000",
  55985=>"100101011",
  55986=>"010111010",
  55987=>"111101101",
  55988=>"011000000",
  55989=>"000000001",
  55990=>"000000000",
  55991=>"001000111",
  55992=>"100100000",
  55993=>"000111111",
  55994=>"000000000",
  55995=>"000010001",
  55996=>"100111111",
  55997=>"000000111",
  55998=>"111000000",
  55999=>"000000111",
  56000=>"011111111",
  56001=>"000111111",
  56002=>"011111111",
  56003=>"000111111",
  56004=>"111111111",
  56005=>"111000000",
  56006=>"000000110",
  56007=>"000001000",
  56008=>"000000000",
  56009=>"101000100",
  56010=>"000000111",
  56011=>"000000111",
  56012=>"000000000",
  56013=>"000110000",
  56014=>"000000000",
  56015=>"000000000",
  56016=>"101111111",
  56017=>"000111111",
  56018=>"100001111",
  56019=>"000000000",
  56020=>"000001000",
  56021=>"011111111",
  56022=>"011011011",
  56023=>"110110111",
  56024=>"111001111",
  56025=>"111111110",
  56026=>"111111111",
  56027=>"011011011",
  56028=>"011000110",
  56029=>"111000001",
  56030=>"100000000",
  56031=>"000000000",
  56032=>"111101000",
  56033=>"100101000",
  56034=>"111111111",
  56035=>"100111111",
  56036=>"000000000",
  56037=>"010100000",
  56038=>"011111111",
  56039=>"000000000",
  56040=>"111000000",
  56041=>"110111111",
  56042=>"000000111",
  56043=>"111111110",
  56044=>"110111010",
  56045=>"000000000",
  56046=>"111111111",
  56047=>"101000100",
  56048=>"111110000",
  56049=>"100000111",
  56050=>"111101001",
  56051=>"111001000",
  56052=>"111111000",
  56053=>"111110111",
  56054=>"000100100",
  56055=>"111010000",
  56056=>"000111111",
  56057=>"000110111",
  56058=>"001000000",
  56059=>"000000111",
  56060=>"000110000",
  56061=>"011000000",
  56062=>"000000000",
  56063=>"000001000",
  56064=>"001000000",
  56065=>"001001000",
  56066=>"100000000",
  56067=>"000000000",
  56068=>"111111000",
  56069=>"000000000",
  56070=>"000000000",
  56071=>"010000111",
  56072=>"111111111",
  56073=>"000000000",
  56074=>"000000101",
  56075=>"111110110",
  56076=>"000000000",
  56077=>"110010011",
  56078=>"000000001",
  56079=>"000111010",
  56080=>"001001101",
  56081=>"000000100",
  56082=>"000000000",
  56083=>"000010000",
  56084=>"111100110",
  56085=>"001000100",
  56086=>"000000000",
  56087=>"101000000",
  56088=>"000000000",
  56089=>"000111111",
  56090=>"111111111",
  56091=>"000000110",
  56092=>"011111111",
  56093=>"000000111",
  56094=>"011011000",
  56095=>"111100100",
  56096=>"100110011",
  56097=>"010010111",
  56098=>"001000000",
  56099=>"000000110",
  56100=>"101000001",
  56101=>"001100100",
  56102=>"100100100",
  56103=>"111001000",
  56104=>"000001111",
  56105=>"000000111",
  56106=>"111001100",
  56107=>"111010000",
  56108=>"111111111",
  56109=>"000000100",
  56110=>"101100000",
  56111=>"111000000",
  56112=>"111001111",
  56113=>"011111111",
  56114=>"111111111",
  56115=>"000111011",
  56116=>"000010010",
  56117=>"111111101",
  56118=>"111001000",
  56119=>"001110110",
  56120=>"011010000",
  56121=>"111000000",
  56122=>"110011001",
  56123=>"010011111",
  56124=>"001000000",
  56125=>"011111000",
  56126=>"100111001",
  56127=>"111111001",
  56128=>"111111100",
  56129=>"111011000",
  56130=>"001001001",
  56131=>"000000000",
  56132=>"000111111",
  56133=>"000000000",
  56134=>"000011011",
  56135=>"111111111",
  56136=>"100000000",
  56137=>"010111111",
  56138=>"101000100",
  56139=>"001111111",
  56140=>"000111111",
  56141=>"000001001",
  56142=>"011111111",
  56143=>"000100111",
  56144=>"000001000",
  56145=>"000000000",
  56146=>"000111111",
  56147=>"111111111",
  56148=>"011111111",
  56149=>"001111011",
  56150=>"110010011",
  56151=>"011111101",
  56152=>"111111110",
  56153=>"111111111",
  56154=>"000000111",
  56155=>"000100111",
  56156=>"011010111",
  56157=>"000000111",
  56158=>"001001001",
  56159=>"111111100",
  56160=>"010110110",
  56161=>"110010000",
  56162=>"000111111",
  56163=>"110000000",
  56164=>"000000100",
  56165=>"111111001",
  56166=>"111011011",
  56167=>"000001111",
  56168=>"000110110",
  56169=>"000100000",
  56170=>"011111001",
  56171=>"110110000",
  56172=>"011111111",
  56173=>"111101000",
  56174=>"000000000",
  56175=>"000000000",
  56176=>"111111111",
  56177=>"111111110",
  56178=>"000010111",
  56179=>"000000000",
  56180=>"100000001",
  56181=>"001111101",
  56182=>"111101000",
  56183=>"111111000",
  56184=>"111000000",
  56185=>"000111111",
  56186=>"000111111",
  56187=>"100101000",
  56188=>"101101111",
  56189=>"011111111",
  56190=>"000010000",
  56191=>"000000000",
  56192=>"000000000",
  56193=>"000000000",
  56194=>"000111011",
  56195=>"100100100",
  56196=>"000000111",
  56197=>"110000000",
  56198=>"000000110",
  56199=>"101000000",
  56200=>"110000000",
  56201=>"111011000",
  56202=>"000000001",
  56203=>"111111111",
  56204=>"001001111",
  56205=>"100100110",
  56206=>"111111110",
  56207=>"000000111",
  56208=>"000111111",
  56209=>"011111111",
  56210=>"110000000",
  56211=>"110111111",
  56212=>"000000111",
  56213=>"000111000",
  56214=>"001000000",
  56215=>"000011111",
  56216=>"111000001",
  56217=>"101011011",
  56218=>"111111110",
  56219=>"000111010",
  56220=>"011010010",
  56221=>"110110100",
  56222=>"111000000",
  56223=>"000111000",
  56224=>"001000000",
  56225=>"000011001",
  56226=>"110111111",
  56227=>"111010000",
  56228=>"010000111",
  56229=>"111111111",
  56230=>"111111000",
  56231=>"000000011",
  56232=>"000011011",
  56233=>"110111111",
  56234=>"111000000",
  56235=>"011111000",
  56236=>"011011111",
  56237=>"011000000",
  56238=>"000000111",
  56239=>"000000100",
  56240=>"111000000",
  56241=>"111111001",
  56242=>"000000110",
  56243=>"011111011",
  56244=>"111000111",
  56245=>"110111111",
  56246=>"110110110",
  56247=>"001000000",
  56248=>"111111101",
  56249=>"111010111",
  56250=>"000111111",
  56251=>"000000000",
  56252=>"000000000",
  56253=>"110111111",
  56254=>"011000000",
  56255=>"000000000",
  56256=>"111111100",
  56257=>"011011111",
  56258=>"110000010",
  56259=>"110110110",
  56260=>"001000000",
  56261=>"100100100",
  56262=>"111000000",
  56263=>"110010000",
  56264=>"100000000",
  56265=>"111111000",
  56266=>"010000000",
  56267=>"000000110",
  56268=>"101111000",
  56269=>"111000000",
  56270=>"010001111",
  56271=>"111000000",
  56272=>"000000111",
  56273=>"110011010",
  56274=>"000100110",
  56275=>"000000001",
  56276=>"000010011",
  56277=>"000111111",
  56278=>"000001111",
  56279=>"000111111",
  56280=>"111111111",
  56281=>"011011010",
  56282=>"001101110",
  56283=>"111110000",
  56284=>"111111111",
  56285=>"010000000",
  56286=>"000000111",
  56287=>"000000000",
  56288=>"111111000",
  56289=>"100100101",
  56290=>"111111000",
  56291=>"000000111",
  56292=>"111111111",
  56293=>"111100000",
  56294=>"001000000",
  56295=>"111001001",
  56296=>"110000000",
  56297=>"111001000",
  56298=>"000000000",
  56299=>"010111000",
  56300=>"100000111",
  56301=>"011101100",
  56302=>"001001001",
  56303=>"100000110",
  56304=>"111111111",
  56305=>"111000110",
  56306=>"000000001",
  56307=>"010000001",
  56308=>"010001000",
  56309=>"000000000",
  56310=>"110111111",
  56311=>"110000000",
  56312=>"000000000",
  56313=>"101001000",
  56314=>"000111111",
  56315=>"000011111",
  56316=>"000000001",
  56317=>"001101111",
  56318=>"000101110",
  56319=>"000110000",
  56320=>"111111110",
  56321=>"111111111",
  56322=>"000000000",
  56323=>"100100000",
  56324=>"101001001",
  56325=>"000000000",
  56326=>"110110110",
  56327=>"111101111",
  56328=>"111100100",
  56329=>"000000000",
  56330=>"010110000",
  56331=>"000110111",
  56332=>"000000000",
  56333=>"111111101",
  56334=>"111111111",
  56335=>"100000000",
  56336=>"111001000",
  56337=>"111111111",
  56338=>"011111111",
  56339=>"111111011",
  56340=>"000100101",
  56341=>"000000000",
  56342=>"000111111",
  56343=>"101000000",
  56344=>"111111111",
  56345=>"110111110",
  56346=>"000011111",
  56347=>"000000000",
  56348=>"111000100",
  56349=>"111000000",
  56350=>"110110111",
  56351=>"000000000",
  56352=>"000000111",
  56353=>"111111111",
  56354=>"000110010",
  56355=>"110110111",
  56356=>"000000000",
  56357=>"001000111",
  56358=>"000000000",
  56359=>"100111111",
  56360=>"111100100",
  56361=>"000000000",
  56362=>"000000000",
  56363=>"000000000",
  56364=>"111111111",
  56365=>"000000011",
  56366=>"111011000",
  56367=>"001000011",
  56368=>"000000000",
  56369=>"111110010",
  56370=>"101111111",
  56371=>"111111111",
  56372=>"000010000",
  56373=>"101100101",
  56374=>"000010000",
  56375=>"000001001",
  56376=>"000111111",
  56377=>"111111111",
  56378=>"000000001",
  56379=>"000111111",
  56380=>"111100111",
  56381=>"000000011",
  56382=>"111111111",
  56383=>"000000000",
  56384=>"000000000",
  56385=>"000000000",
  56386=>"111111111",
  56387=>"111111000",
  56388=>"000110110",
  56389=>"000000000",
  56390=>"111101000",
  56391=>"111111000",
  56392=>"000000100",
  56393=>"000000001",
  56394=>"000111010",
  56395=>"000111111",
  56396=>"000010111",
  56397=>"000000000",
  56398=>"010000000",
  56399=>"001000000",
  56400=>"000000000",
  56401=>"000000000",
  56402=>"000000110",
  56403=>"001111001",
  56404=>"111111111",
  56405=>"000000000",
  56406=>"100101111",
  56407=>"111010010",
  56408=>"111000001",
  56409=>"111101101",
  56410=>"000011111",
  56411=>"000000000",
  56412=>"110100100",
  56413=>"111111111",
  56414=>"001000000",
  56415=>"000000000",
  56416=>"111100101",
  56417=>"000000000",
  56418=>"111110100",
  56419=>"111111111",
  56420=>"111101101",
  56421=>"000000000",
  56422=>"000000000",
  56423=>"000011000",
  56424=>"000100111",
  56425=>"000110110",
  56426=>"110111110",
  56427=>"111111111",
  56428=>"101111111",
  56429=>"111111110",
  56430=>"111110111",
  56431=>"111110110",
  56432=>"011111111",
  56433=>"001101100",
  56434=>"111010110",
  56435=>"000000000",
  56436=>"100111000",
  56437=>"110110110",
  56438=>"001011111",
  56439=>"000000000",
  56440=>"000000000",
  56441=>"000000000",
  56442=>"110010010",
  56443=>"111000000",
  56444=>"000111111",
  56445=>"000011111",
  56446=>"110000000",
  56447=>"000000011",
  56448=>"000000000",
  56449=>"011011011",
  56450=>"111111110",
  56451=>"111110110",
  56452=>"000000001",
  56453=>"000000000",
  56454=>"111111111",
  56455=>"000000000",
  56456=>"111111111",
  56457=>"010111111",
  56458=>"000000110",
  56459=>"111000000",
  56460=>"111000010",
  56461=>"000000001",
  56462=>"000000000",
  56463=>"000000111",
  56464=>"111111111",
  56465=>"111111111",
  56466=>"001111111",
  56467=>"111100111",
  56468=>"111111111",
  56469=>"110110110",
  56470=>"000000100",
  56471=>"000000001",
  56472=>"111111111",
  56473=>"000000110",
  56474=>"111111111",
  56475=>"000000111",
  56476=>"101001001",
  56477=>"111111111",
  56478=>"111101101",
  56479=>"000000000",
  56480=>"100111010",
  56481=>"001000100",
  56482=>"000000000",
  56483=>"111111111",
  56484=>"100000001",
  56485=>"100000000",
  56486=>"011111100",
  56487=>"111111110",
  56488=>"000111011",
  56489=>"111000000",
  56490=>"111111111",
  56491=>"111111111",
  56492=>"000000100",
  56493=>"111111110",
  56494=>"111111111",
  56495=>"111111010",
  56496=>"000111111",
  56497=>"000000000",
  56498=>"110111110",
  56499=>"111111111",
  56500=>"000000000",
  56501=>"001000000",
  56502=>"111110000",
  56503=>"111111111",
  56504=>"111111111",
  56505=>"000000100",
  56506=>"111111111",
  56507=>"000000000",
  56508=>"110000000",
  56509=>"001000000",
  56510=>"111111111",
  56511=>"000111111",
  56512=>"111111111",
  56513=>"000101111",
  56514=>"000000000",
  56515=>"101111111",
  56516=>"111111000",
  56517=>"000000000",
  56518=>"101000000",
  56519=>"110000111",
  56520=>"000000001",
  56521=>"100111000",
  56522=>"111111110",
  56523=>"000000010",
  56524=>"001011011",
  56525=>"101000000",
  56526=>"000000010",
  56527=>"100111000",
  56528=>"000000000",
  56529=>"111110110",
  56530=>"111111111",
  56531=>"011111010",
  56532=>"110110000",
  56533=>"100111001",
  56534=>"000010111",
  56535=>"010110110",
  56536=>"000000000",
  56537=>"011111001",
  56538=>"000000000",
  56539=>"000000000",
  56540=>"000010111",
  56541=>"111111111",
  56542=>"000111111",
  56543=>"000000001",
  56544=>"011001111",
  56545=>"000000000",
  56546=>"111111011",
  56547=>"000000001",
  56548=>"000010010",
  56549=>"000000000",
  56550=>"110100000",
  56551=>"111100100",
  56552=>"110000001",
  56553=>"000001011",
  56554=>"111011001",
  56555=>"100000111",
  56556=>"110111000",
  56557=>"111111111",
  56558=>"111111111",
  56559=>"000000000",
  56560=>"101001000",
  56561=>"100111110",
  56562=>"111111111",
  56563=>"000000000",
  56564=>"000000000",
  56565=>"000000000",
  56566=>"110111111",
  56567=>"000000000",
  56568=>"010000000",
  56569=>"000000111",
  56570=>"000000000",
  56571=>"001001001",
  56572=>"100100111",
  56573=>"000000000",
  56574=>"110001001",
  56575=>"111110011",
  56576=>"000000000",
  56577=>"111101111",
  56578=>"111111111",
  56579=>"000101111",
  56580=>"111110111",
  56581=>"101001101",
  56582=>"111111111",
  56583=>"001111111",
  56584=>"000111111",
  56585=>"111110001",
  56586=>"011001011",
  56587=>"111111111",
  56588=>"111111111",
  56589=>"001111001",
  56590=>"100111111",
  56591=>"000000000",
  56592=>"110010000",
  56593=>"111111111",
  56594=>"000000000",
  56595=>"000110111",
  56596=>"000000000",
  56597=>"000000100",
  56598=>"111111111",
  56599=>"000000000",
  56600=>"000000000",
  56601=>"101111000",
  56602=>"000000110",
  56603=>"000000000",
  56604=>"110110111",
  56605=>"000000101",
  56606=>"010111111",
  56607=>"110111111",
  56608=>"111111110",
  56609=>"010000110",
  56610=>"111111110",
  56611=>"111011000",
  56612=>"111111111",
  56613=>"000000011",
  56614=>"110110110",
  56615=>"000100000",
  56616=>"111101101",
  56617=>"000000010",
  56618=>"001001100",
  56619=>"000000101",
  56620=>"000000000",
  56621=>"001111111",
  56622=>"111010111",
  56623=>"100000000",
  56624=>"111111110",
  56625=>"000000001",
  56626=>"111011111",
  56627=>"000000000",
  56628=>"111111111",
  56629=>"100110110",
  56630=>"111111111",
  56631=>"111011111",
  56632=>"000000000",
  56633=>"000000101",
  56634=>"110000000",
  56635=>"000001011",
  56636=>"111111111",
  56637=>"110000100",
  56638=>"101101100",
  56639=>"001101111",
  56640=>"001001000",
  56641=>"111011011",
  56642=>"100000100",
  56643=>"000000000",
  56644=>"111111111",
  56645=>"111110100",
  56646=>"000000000",
  56647=>"011011011",
  56648=>"110000000",
  56649=>"000000000",
  56650=>"100000100",
  56651=>"111111111",
  56652=>"110000000",
  56653=>"001000000",
  56654=>"111111110",
  56655=>"100100100",
  56656=>"111111000",
  56657=>"100111000",
  56658=>"111001001",
  56659=>"100011000",
  56660=>"110000000",
  56661=>"001001001",
  56662=>"000000010",
  56663=>"010000000",
  56664=>"111111111",
  56665=>"110000010",
  56666=>"100001111",
  56667=>"000000000",
  56668=>"000100110",
  56669=>"110000000",
  56670=>"000100110",
  56671=>"111111111",
  56672=>"000000100",
  56673=>"111111111",
  56674=>"110111111",
  56675=>"111101011",
  56676=>"111111111",
  56677=>"000000000",
  56678=>"000011000",
  56679=>"000111011",
  56680=>"111111111",
  56681=>"101101001",
  56682=>"111111111",
  56683=>"000011001",
  56684=>"011000000",
  56685=>"101011011",
  56686=>"000000000",
  56687=>"110100100",
  56688=>"111100100",
  56689=>"111111111",
  56690=>"011000101",
  56691=>"100000000",
  56692=>"111111111",
  56693=>"011111111",
  56694=>"111111000",
  56695=>"110000000",
  56696=>"111001000",
  56697=>"111111111",
  56698=>"000000000",
  56699=>"101101111",
  56700=>"000100110",
  56701=>"001000011",
  56702=>"111111111",
  56703=>"111101111",
  56704=>"111111111",
  56705=>"001000001",
  56706=>"000000001",
  56707=>"111110100",
  56708=>"111111111",
  56709=>"010010000",
  56710=>"000000000",
  56711=>"000000110",
  56712=>"000000000",
  56713=>"111111111",
  56714=>"000000000",
  56715=>"001001000",
  56716=>"111111111",
  56717=>"000100100",
  56718=>"000001011",
  56719=>"111111000",
  56720=>"111000000",
  56721=>"011000000",
  56722=>"111011010",
  56723=>"111111111",
  56724=>"001111111",
  56725=>"010010010",
  56726=>"111111111",
  56727=>"001001001",
  56728=>"000111111",
  56729=>"000000000",
  56730=>"000010000",
  56731=>"001100000",
  56732=>"000000000",
  56733=>"111000100",
  56734=>"001111001",
  56735=>"001000111",
  56736=>"010000000",
  56737=>"000000000",
  56738=>"000111111",
  56739=>"101111000",
  56740=>"000001111",
  56741=>"001000001",
  56742=>"000001111",
  56743=>"010000000",
  56744=>"110000000",
  56745=>"000000000",
  56746=>"100000000",
  56747=>"011011111",
  56748=>"110000000",
  56749=>"111001111",
  56750=>"111111111",
  56751=>"100111111",
  56752=>"110111111",
  56753=>"111000011",
  56754=>"111111110",
  56755=>"000010111",
  56756=>"000000100",
  56757=>"010001001",
  56758=>"110110111",
  56759=>"001000001",
  56760=>"111111111",
  56761=>"011011111",
  56762=>"000000100",
  56763=>"000000000",
  56764=>"011001011",
  56765=>"111110110",
  56766=>"000001000",
  56767=>"110111100",
  56768=>"111011001",
  56769=>"010011110",
  56770=>"111111111",
  56771=>"111001011",
  56772=>"111111000",
  56773=>"001011111",
  56774=>"111111111",
  56775=>"001001111",
  56776=>"000010011",
  56777=>"000000000",
  56778=>"010111110",
  56779=>"111111111",
  56780=>"000010110",
  56781=>"010011011",
  56782=>"011000110",
  56783=>"000111100",
  56784=>"001111111",
  56785=>"111111001",
  56786=>"011011111",
  56787=>"000000100",
  56788=>"011111100",
  56789=>"000000000",
  56790=>"011000000",
  56791=>"001000000",
  56792=>"100110000",
  56793=>"111111111",
  56794=>"101100111",
  56795=>"100111110",
  56796=>"001001011",
  56797=>"011111001",
  56798=>"111101111",
  56799=>"111111110",
  56800=>"000000000",
  56801=>"001011001",
  56802=>"111111111",
  56803=>"110100000",
  56804=>"111111111",
  56805=>"110000000",
  56806=>"001001101",
  56807=>"000100111",
  56808=>"000000000",
  56809=>"111111000",
  56810=>"100100101",
  56811=>"000000001",
  56812=>"000000101",
  56813=>"111111011",
  56814=>"111111111",
  56815=>"000000000",
  56816=>"110110111",
  56817=>"111111101",
  56818=>"111111100",
  56819=>"000001001",
  56820=>"011011000",
  56821=>"111000000",
  56822=>"111111000",
  56823=>"010000000",
  56824=>"000000000",
  56825=>"101111011",
  56826=>"110000000",
  56827=>"000000110",
  56828=>"000000000",
  56829=>"101001001",
  56830=>"001110000",
  56831=>"000100111",
  56832=>"010000000",
  56833=>"111101000",
  56834=>"101001011",
  56835=>"000000001",
  56836=>"111111111",
  56837=>"000000000",
  56838=>"000010111",
  56839=>"111111111",
  56840=>"000111001",
  56841=>"000000111",
  56842=>"111110110",
  56843=>"000011011",
  56844=>"111000100",
  56845=>"000011111",
  56846=>"101111111",
  56847=>"100101111",
  56848=>"111111110",
  56849=>"111111111",
  56850=>"111111011",
  56851=>"111111000",
  56852=>"111111111",
  56853=>"111111101",
  56854=>"110000000",
  56855=>"101111001",
  56856=>"000100100",
  56857=>"000000010",
  56858=>"001001100",
  56859=>"100110100",
  56860=>"111101111",
  56861=>"111111111",
  56862=>"111111111",
  56863=>"010010111",
  56864=>"111111111",
  56865=>"111111000",
  56866=>"100100111",
  56867=>"111111111",
  56868=>"000100001",
  56869=>"000000000",
  56870=>"000000000",
  56871=>"111111110",
  56872=>"111111111",
  56873=>"000101111",
  56874=>"111111111",
  56875=>"111110000",
  56876=>"111110100",
  56877=>"000111100",
  56878=>"111000100",
  56879=>"110100100",
  56880=>"011011010",
  56881=>"000000001",
  56882=>"101111111",
  56883=>"111111001",
  56884=>"111111111",
  56885=>"000110100",
  56886=>"111111110",
  56887=>"111111111",
  56888=>"000000001",
  56889=>"111000010",
  56890=>"111101001",
  56891=>"110000000",
  56892=>"111111111",
  56893=>"111011000",
  56894=>"111111111",
  56895=>"111100100",
  56896=>"111111111",
  56897=>"111000000",
  56898=>"000000000",
  56899=>"111111111",
  56900=>"001101100",
  56901=>"000000000",
  56902=>"000000000",
  56903=>"111000000",
  56904=>"000000010",
  56905=>"000000000",
  56906=>"111111111",
  56907=>"000000011",
  56908=>"110110111",
  56909=>"111000110",
  56910=>"000000000",
  56911=>"111110000",
  56912=>"111000000",
  56913=>"111111000",
  56914=>"111011000",
  56915=>"000000000",
  56916=>"000001011",
  56917=>"000000000",
  56918=>"000100111",
  56919=>"110000000",
  56920=>"001011110",
  56921=>"000000000",
  56922=>"110110110",
  56923=>"100000000",
  56924=>"000000000",
  56925=>"111000000",
  56926=>"010000000",
  56927=>"111000000",
  56928=>"000000000",
  56929=>"000000000",
  56930=>"111111011",
  56931=>"000000000",
  56932=>"000000000",
  56933=>"111000000",
  56934=>"000000010",
  56935=>"111111111",
  56936=>"000000000",
  56937=>"000000001",
  56938=>"001011011",
  56939=>"111111111",
  56940=>"111111001",
  56941=>"111011011",
  56942=>"000000000",
  56943=>"110111110",
  56944=>"111110110",
  56945=>"000000000",
  56946=>"100111111",
  56947=>"101111111",
  56948=>"000000000",
  56949=>"000000111",
  56950=>"111111111",
  56951=>"000011011",
  56952=>"000100000",
  56953=>"000000110",
  56954=>"000000000",
  56955=>"001001000",
  56956=>"110110110",
  56957=>"111110000",
  56958=>"000000000",
  56959=>"000001001",
  56960=>"111000111",
  56961=>"111000111",
  56962=>"000111111",
  56963=>"100111111",
  56964=>"110100100",
  56965=>"101111111",
  56966=>"111111110",
  56967=>"111111110",
  56968=>"111111011",
  56969=>"101100100",
  56970=>"001101111",
  56971=>"111100000",
  56972=>"111000000",
  56973=>"111110000",
  56974=>"110100000",
  56975=>"001000000",
  56976=>"000000000",
  56977=>"001001000",
  56978=>"111110111",
  56979=>"001000000",
  56980=>"110110100",
  56981=>"000000111",
  56982=>"111101100",
  56983=>"111010000",
  56984=>"011000000",
  56985=>"111111011",
  56986=>"100111111",
  56987=>"001001101",
  56988=>"110010000",
  56989=>"000111111",
  56990=>"000000000",
  56991=>"111111111",
  56992=>"111111100",
  56993=>"111000000",
  56994=>"111111111",
  56995=>"010110111",
  56996=>"000000000",
  56997=>"000000101",
  56998=>"000111111",
  56999=>"001000000",
  57000=>"000000000",
  57001=>"010111111",
  57002=>"111111111",
  57003=>"010000000",
  57004=>"111111111",
  57005=>"000000000",
  57006=>"001111111",
  57007=>"000110110",
  57008=>"111111000",
  57009=>"000011110",
  57010=>"000111111",
  57011=>"000000000",
  57012=>"111111000",
  57013=>"000000110",
  57014=>"000000000",
  57015=>"110000000",
  57016=>"100110100",
  57017=>"111101000",
  57018=>"000000000",
  57019=>"111110000",
  57020=>"000000000",
  57021=>"000000000",
  57022=>"000000000",
  57023=>"000001111",
  57024=>"111111111",
  57025=>"000000111",
  57026=>"111000000",
  57027=>"100111000",
  57028=>"100001001",
  57029=>"000000000",
  57030=>"000111111",
  57031=>"111111010",
  57032=>"111111111",
  57033=>"101111111",
  57034=>"000000100",
  57035=>"111111111",
  57036=>"000000000",
  57037=>"000010000",
  57038=>"111111111",
  57039=>"000001011",
  57040=>"010000000",
  57041=>"101000100",
  57042=>"111111110",
  57043=>"111010111",
  57044=>"100000000",
  57045=>"111111101",
  57046=>"010011011",
  57047=>"000001101",
  57048=>"000000011",
  57049=>"111111000",
  57050=>"111111111",
  57051=>"110110101",
  57052=>"000000000",
  57053=>"111111000",
  57054=>"111111011",
  57055=>"110000000",
  57056=>"111100100",
  57057=>"111111001",
  57058=>"110111101",
  57059=>"000110111",
  57060=>"000000000",
  57061=>"011011001",
  57062=>"110000000",
  57063=>"000000000",
  57064=>"000011000",
  57065=>"010010000",
  57066=>"000000111",
  57067=>"101100100",
  57068=>"000000111",
  57069=>"000000000",
  57070=>"100000000",
  57071=>"000111000",
  57072=>"000000000",
  57073=>"000111111",
  57074=>"111111111",
  57075=>"000000111",
  57076=>"000000000",
  57077=>"111100000",
  57078=>"000010000",
  57079=>"111111111",
  57080=>"111111111",
  57081=>"010100000",
  57082=>"000001111",
  57083=>"111111000",
  57084=>"111110000",
  57085=>"100000000",
  57086=>"010000000",
  57087=>"111010011",
  57088=>"000000001",
  57089=>"110110111",
  57090=>"111111111",
  57091=>"110110111",
  57092=>"111000000",
  57093=>"001100111",
  57094=>"111000000",
  57095=>"001001000",
  57096=>"001100101",
  57097=>"000000000",
  57098=>"111111111",
  57099=>"000000111",
  57100=>"000000000",
  57101=>"010011011",
  57102=>"111111011",
  57103=>"111011000",
  57104=>"110000000",
  57105=>"000000000",
  57106=>"111011000",
  57107=>"100001000",
  57108=>"111110000",
  57109=>"111111111",
  57110=>"110110100",
  57111=>"111111110",
  57112=>"000000100",
  57113=>"101000000",
  57114=>"000000000",
  57115=>"000110110",
  57116=>"111111000",
  57117=>"111000001",
  57118=>"111101001",
  57119=>"111000100",
  57120=>"011111111",
  57121=>"000001001",
  57122=>"000000111",
  57123=>"110000000",
  57124=>"000000110",
  57125=>"100100000",
  57126=>"111111111",
  57127=>"111101111",
  57128=>"100110111",
  57129=>"001001001",
  57130=>"001000000",
  57131=>"001001111",
  57132=>"000000000",
  57133=>"111000000",
  57134=>"111000000",
  57135=>"000000111",
  57136=>"110000000",
  57137=>"010111011",
  57138=>"110110111",
  57139=>"000000011",
  57140=>"000011000",
  57141=>"000101100",
  57142=>"111110000",
  57143=>"001000000",
  57144=>"111110111",
  57145=>"111010000",
  57146=>"000010011",
  57147=>"000000011",
  57148=>"000000000",
  57149=>"110010000",
  57150=>"001000000",
  57151=>"100110000",
  57152=>"111100101",
  57153=>"111000000",
  57154=>"000100110",
  57155=>"000000000",
  57156=>"011001000",
  57157=>"111111111",
  57158=>"001000000",
  57159=>"010000000",
  57160=>"111011111",
  57161=>"101000000",
  57162=>"100000000",
  57163=>"111111001",
  57164=>"110010000",
  57165=>"000000011",
  57166=>"110110011",
  57167=>"011111111",
  57168=>"000000001",
  57169=>"111011000",
  57170=>"111010000",
  57171=>"000111111",
  57172=>"010111111",
  57173=>"011011011",
  57174=>"010111111",
  57175=>"001000000",
  57176=>"000000000",
  57177=>"000010000",
  57178=>"001110110",
  57179=>"010000000",
  57180=>"000000000",
  57181=>"001001100",
  57182=>"110000000",
  57183=>"000001100",
  57184=>"000000000",
  57185=>"111111101",
  57186=>"100111111",
  57187=>"101111010",
  57188=>"111111111",
  57189=>"111111111",
  57190=>"011111111",
  57191=>"111010110",
  57192=>"111111110",
  57193=>"111101100",
  57194=>"111111111",
  57195=>"111111111",
  57196=>"110111000",
  57197=>"000000000",
  57198=>"111111111",
  57199=>"001000000",
  57200=>"001111011",
  57201=>"111101100",
  57202=>"000111111",
  57203=>"000000100",
  57204=>"111111101",
  57205=>"110000000",
  57206=>"000111111",
  57207=>"111111111",
  57208=>"000111111",
  57209=>"111111111",
  57210=>"101001000",
  57211=>"110110111",
  57212=>"111111111",
  57213=>"000001010",
  57214=>"000010011",
  57215=>"110000100",
  57216=>"001001001",
  57217=>"000000111",
  57218=>"000000011",
  57219=>"111011001",
  57220=>"000011011",
  57221=>"011010000",
  57222=>"001111111",
  57223=>"100000000",
  57224=>"000000000",
  57225=>"011111101",
  57226=>"000000000",
  57227=>"111110000",
  57228=>"101101111",
  57229=>"000100111",
  57230=>"111111100",
  57231=>"111111111",
  57232=>"111111000",
  57233=>"111000000",
  57234=>"111001001",
  57235=>"000000000",
  57236=>"111011001",
  57237=>"100111101",
  57238=>"111111111",
  57239=>"001000001",
  57240=>"111111111",
  57241=>"100100110",
  57242=>"000001010",
  57243=>"111111011",
  57244=>"000000000",
  57245=>"010000000",
  57246=>"000010010",
  57247=>"000011011",
  57248=>"111111110",
  57249=>"000000010",
  57250=>"000000000",
  57251=>"001001111",
  57252=>"110111101",
  57253=>"111001000",
  57254=>"110011000",
  57255=>"111111000",
  57256=>"111111111",
  57257=>"000100000",
  57258=>"000100111",
  57259=>"000000000",
  57260=>"001001001",
  57261=>"111001000",
  57262=>"001111111",
  57263=>"000000000",
  57264=>"111111100",
  57265=>"000000010",
  57266=>"101111111",
  57267=>"110110111",
  57268=>"100000000",
  57269=>"011111111",
  57270=>"000011111",
  57271=>"000111111",
  57272=>"111111100",
  57273=>"111010000",
  57274=>"011010111",
  57275=>"000000000",
  57276=>"111111000",
  57277=>"011011011",
  57278=>"000001111",
  57279=>"100100100",
  57280=>"000001011",
  57281=>"000101000",
  57282=>"111111111",
  57283=>"000000000",
  57284=>"111110000",
  57285=>"000000000",
  57286=>"111111000",
  57287=>"000100111",
  57288=>"011001100",
  57289=>"110110001",
  57290=>"011001000",
  57291=>"111111111",
  57292=>"101000000",
  57293=>"011011110",
  57294=>"100111111",
  57295=>"100011001",
  57296=>"000000000",
  57297=>"110100110",
  57298=>"000000010",
  57299=>"000001000",
  57300=>"000010111",
  57301=>"100000000",
  57302=>"010000000",
  57303=>"100100111",
  57304=>"111000101",
  57305=>"100100100",
  57306=>"100000000",
  57307=>"000110000",
  57308=>"000010111",
  57309=>"011011101",
  57310=>"000000000",
  57311=>"000111111",
  57312=>"011001111",
  57313=>"000000111",
  57314=>"110101000",
  57315=>"111000011",
  57316=>"111111110",
  57317=>"000000011",
  57318=>"001000000",
  57319=>"000000000",
  57320=>"111000001",
  57321=>"111110000",
  57322=>"111111000",
  57323=>"000000000",
  57324=>"111111111",
  57325=>"000000000",
  57326=>"111111001",
  57327=>"000000100",
  57328=>"000000000",
  57329=>"000111000",
  57330=>"111011100",
  57331=>"000101111",
  57332=>"110110000",
  57333=>"000010000",
  57334=>"000011010",
  57335=>"111111100",
  57336=>"010010111",
  57337=>"010000000",
  57338=>"111111111",
  57339=>"111111000",
  57340=>"110110000",
  57341=>"111111111",
  57342=>"111111111",
  57343=>"111001000",
  57344=>"100100000",
  57345=>"100100000",
  57346=>"000000000",
  57347=>"111111111",
  57348=>"001101111",
  57349=>"100000000",
  57350=>"000000000",
  57351=>"111111111",
  57352=>"010000000",
  57353=>"000000000",
  57354=>"001111111",
  57355=>"011111111",
  57356=>"000000000",
  57357=>"001001000",
  57358=>"000001001",
  57359=>"000000000",
  57360=>"000000001",
  57361=>"111111000",
  57362=>"000000000",
  57363=>"101000000",
  57364=>"000000000",
  57365=>"010111110",
  57366=>"111111111",
  57367=>"000101001",
  57368=>"000101111",
  57369=>"111111111",
  57370=>"111111011",
  57371=>"000010110",
  57372=>"111111111",
  57373=>"001001001",
  57374=>"011011001",
  57375=>"000000110",
  57376=>"111000000",
  57377=>"110110111",
  57378=>"101101111",
  57379=>"111011001",
  57380=>"111111111",
  57381=>"000000000",
  57382=>"000000000",
  57383=>"000000000",
  57384=>"111111000",
  57385=>"111110010",
  57386=>"000000000",
  57387=>"000110000",
  57388=>"010111111",
  57389=>"110101000",
  57390=>"010010000",
  57391=>"011011111",
  57392=>"111111111",
  57393=>"000000000",
  57394=>"000000000",
  57395=>"000000000",
  57396=>"000110110",
  57397=>"110111111",
  57398=>"001011000",
  57399=>"111111111",
  57400=>"000000010",
  57401=>"010000000",
  57402=>"111111111",
  57403=>"000000000",
  57404=>"111111110",
  57405=>"000000000",
  57406=>"000011011",
  57407=>"000000000",
  57408=>"000000000",
  57409=>"000000000",
  57410=>"111111111",
  57411=>"000000111",
  57412=>"001111011",
  57413=>"011011001",
  57414=>"011001111",
  57415=>"000000000",
  57416=>"000111011",
  57417=>"000000001",
  57418=>"111011000",
  57419=>"000100110",
  57420=>"101000000",
  57421=>"111000000",
  57422=>"000000000",
  57423=>"111111111",
  57424=>"000000000",
  57425=>"011001000",
  57426=>"000000000",
  57427=>"111111111",
  57428=>"000000000",
  57429=>"111111111",
  57430=>"001011000",
  57431=>"111111110",
  57432=>"000000000",
  57433=>"101001000",
  57434=>"111111111",
  57435=>"000000000",
  57436=>"111111111",
  57437=>"000101111",
  57438=>"000111100",
  57439=>"001111111",
  57440=>"100100111",
  57441=>"001111111",
  57442=>"011001000",
  57443=>"111111111",
  57444=>"000001001",
  57445=>"111110000",
  57446=>"011110000",
  57447=>"000100000",
  57448=>"010111111",
  57449=>"111000000",
  57450=>"000000010",
  57451=>"110111111",
  57452=>"110111011",
  57453=>"111111111",
  57454=>"111111111",
  57455=>"010110010",
  57456=>"000000000",
  57457=>"000000000",
  57458=>"011111011",
  57459=>"010010000",
  57460=>"000000000",
  57461=>"000000000",
  57462=>"000000000",
  57463=>"111111111",
  57464=>"000011111",
  57465=>"111101000",
  57466=>"000000111",
  57467=>"000000000",
  57468=>"000111111",
  57469=>"000000000",
  57470=>"000000000",
  57471=>"000000000",
  57472=>"000000000",
  57473=>"000110111",
  57474=>"111110100",
  57475=>"011011001",
  57476=>"000100111",
  57477=>"000000000",
  57478=>"001111001",
  57479=>"000000000",
  57480=>"010000000",
  57481=>"000000111",
  57482=>"100100111",
  57483=>"111111111",
  57484=>"000000000",
  57485=>"000000001",
  57486=>"000000100",
  57487=>"000100111",
  57488=>"111111111",
  57489=>"011011000",
  57490=>"000100101",
  57491=>"111111111",
  57492=>"111111111",
  57493=>"110111111",
  57494=>"010000000",
  57495=>"000001111",
  57496=>"111111111",
  57497=>"110111110",
  57498=>"000000000",
  57499=>"100000000",
  57500=>"000100000",
  57501=>"100101000",
  57502=>"011010110",
  57503=>"111111101",
  57504=>"000000000",
  57505=>"111101011",
  57506=>"000000000",
  57507=>"110000010",
  57508=>"010000000",
  57509=>"000101111",
  57510=>"000000000",
  57511=>"001001001",
  57512=>"000000100",
  57513=>"111111111",
  57514=>"000000000",
  57515=>"111111111",
  57516=>"010111111",
  57517=>"000001001",
  57518=>"111111011",
  57519=>"000010001",
  57520=>"000000000",
  57521=>"111111011",
  57522=>"111111110",
  57523=>"010111011",
  57524=>"011111111",
  57525=>"111111111",
  57526=>"011000000",
  57527=>"001000000",
  57528=>"111111111",
  57529=>"000000000",
  57530=>"101001001",
  57531=>"110110000",
  57532=>"000000000",
  57533=>"110110100",
  57534=>"111111111",
  57535=>"111110110",
  57536=>"111111111",
  57537=>"000000000",
  57538=>"110000000",
  57539=>"000000001",
  57540=>"000100011",
  57541=>"000111111",
  57542=>"111001000",
  57543=>"000000000",
  57544=>"111111111",
  57545=>"000000000",
  57546=>"111111111",
  57547=>"000000011",
  57548=>"100111111",
  57549=>"101111111",
  57550=>"001000111",
  57551=>"111011001",
  57552=>"000000000",
  57553=>"111111111",
  57554=>"000000001",
  57555=>"010010000",
  57556=>"111001111",
  57557=>"000000000",
  57558=>"000000000",
  57559=>"111111111",
  57560=>"111111111",
  57561=>"111101111",
  57562=>"000000111",
  57563=>"111000111",
  57564=>"000001001",
  57565=>"000100111",
  57566=>"000000000",
  57567=>"001011000",
  57568=>"001000011",
  57569=>"100110000",
  57570=>"111000000",
  57571=>"011011001",
  57572=>"010000111",
  57573=>"000000000",
  57574=>"000010111",
  57575=>"000010000",
  57576=>"000000000",
  57577=>"001001000",
  57578=>"000011001",
  57579=>"000000001",
  57580=>"111110000",
  57581=>"011001000",
  57582=>"111000000",
  57583=>"111111111",
  57584=>"000100111",
  57585=>"011011111",
  57586=>"111001000",
  57587=>"000000000",
  57588=>"000001011",
  57589=>"011001100",
  57590=>"001111011",
  57591=>"010000100",
  57592=>"111111111",
  57593=>"110000000",
  57594=>"000000000",
  57595=>"011001000",
  57596=>"110110111",
  57597=>"001001111",
  57598=>"010000001",
  57599=>"111111111",
  57600=>"000010000",
  57601=>"000111111",
  57602=>"111000000",
  57603=>"001111111",
  57604=>"110111101",
  57605=>"000000001",
  57606=>"111111000",
  57607=>"111111111",
  57608=>"111100000",
  57609=>"000000000",
  57610=>"000101111",
  57611=>"111111111",
  57612=>"101100000",
  57613=>"111111111",
  57614=>"101111111",
  57615=>"000000000",
  57616=>"000111111",
  57617=>"000000111",
  57618=>"000000011",
  57619=>"000000100",
  57620=>"001000000",
  57621=>"000000000",
  57622=>"011011000",
  57623=>"010000000",
  57624=>"001001001",
  57625=>"011011111",
  57626=>"111111011",
  57627=>"111111111",
  57628=>"000000000",
  57629=>"011000000",
  57630=>"000111110",
  57631=>"111111000",
  57632=>"101001000",
  57633=>"000000000",
  57634=>"000000000",
  57635=>"111111110",
  57636=>"100100100",
  57637=>"000011111",
  57638=>"000000000",
  57639=>"011011011",
  57640=>"000000000",
  57641=>"000000000",
  57642=>"100100011",
  57643=>"111111011",
  57644=>"000000000",
  57645=>"111001000",
  57646=>"111000111",
  57647=>"000011111",
  57648=>"000000000",
  57649=>"000111111",
  57650=>"111111111",
  57651=>"001000000",
  57652=>"111110111",
  57653=>"100111111",
  57654=>"000000000",
  57655=>"101011111",
  57656=>"000000010",
  57657=>"000000111",
  57658=>"000110110",
  57659=>"110011001",
  57660=>"111001001",
  57661=>"000000101",
  57662=>"111111111",
  57663=>"111011000",
  57664=>"111010011",
  57665=>"111001101",
  57666=>"110110111",
  57667=>"000000000",
  57668=>"000000000",
  57669=>"000000001",
  57670=>"111000000",
  57671=>"111111101",
  57672=>"000111011",
  57673=>"000000000",
  57674=>"111111111",
  57675=>"000000000",
  57676=>"000000000",
  57677=>"111011011",
  57678=>"000000000",
  57679=>"100111111",
  57680=>"001001001",
  57681=>"111111111",
  57682=>"000000100",
  57683=>"000000000",
  57684=>"000000000",
  57685=>"001000000",
  57686=>"111111111",
  57687=>"011000000",
  57688=>"111111111",
  57689=>"111010000",
  57690=>"111111111",
  57691=>"100111111",
  57692=>"001111110",
  57693=>"000000101",
  57694=>"000000011",
  57695=>"100000001",
  57696=>"111111111",
  57697=>"100000000",
  57698=>"100100111",
  57699=>"111111111",
  57700=>"111101100",
  57701=>"111111001",
  57702=>"000000111",
  57703=>"000000000",
  57704=>"000000000",
  57705=>"000000000",
  57706=>"000000001",
  57707=>"101001000",
  57708=>"010001000",
  57709=>"111100111",
  57710=>"000000000",
  57711=>"110000000",
  57712=>"110111110",
  57713=>"010110111",
  57714=>"001000000",
  57715=>"111111111",
  57716=>"000000000",
  57717=>"000000000",
  57718=>"000000101",
  57719=>"011011000",
  57720=>"111111111",
  57721=>"111110111",
  57722=>"011001011",
  57723=>"110111111",
  57724=>"000000000",
  57725=>"001001001",
  57726=>"000000000",
  57727=>"000000111",
  57728=>"100100100",
  57729=>"000000011",
  57730=>"110110100",
  57731=>"000001111",
  57732=>"111111111",
  57733=>"000000000",
  57734=>"011001000",
  57735=>"111111111",
  57736=>"000000000",
  57737=>"111111111",
  57738=>"001001011",
  57739=>"010111111",
  57740=>"111111111",
  57741=>"110111110",
  57742=>"000000000",
  57743=>"000000000",
  57744=>"110000000",
  57745=>"001001000",
  57746=>"100000000",
  57747=>"110100000",
  57748=>"100110111",
  57749=>"011011011",
  57750=>"011001001",
  57751=>"100000010",
  57752=>"100100100",
  57753=>"000000000",
  57754=>"101101101",
  57755=>"000000000",
  57756=>"001111110",
  57757=>"000001111",
  57758=>"100100110",
  57759=>"100110000",
  57760=>"111110100",
  57761=>"111111111",
  57762=>"001011011",
  57763=>"011011111",
  57764=>"000101101",
  57765=>"111111111",
  57766=>"000001001",
  57767=>"111001001",
  57768=>"000110000",
  57769=>"111111111",
  57770=>"000000001",
  57771=>"111001111",
  57772=>"000000000",
  57773=>"000000000",
  57774=>"111111100",
  57775=>"000000000",
  57776=>"110000000",
  57777=>"000101111",
  57778=>"000010001",
  57779=>"000101111",
  57780=>"000000000",
  57781=>"011111111",
  57782=>"111111111",
  57783=>"010111111",
  57784=>"000000010",
  57785=>"100000101",
  57786=>"111111111",
  57787=>"100100101",
  57788=>"111100000",
  57789=>"000111001",
  57790=>"001000000",
  57791=>"100000100",
  57792=>"111111111",
  57793=>"110111111",
  57794=>"000000000",
  57795=>"111111110",
  57796=>"001011001",
  57797=>"111001111",
  57798=>"111111111",
  57799=>"111111100",
  57800=>"000000000",
  57801=>"000001110",
  57802=>"000000110",
  57803=>"000000000",
  57804=>"111110000",
  57805=>"000000000",
  57806=>"111111011",
  57807=>"000011111",
  57808=>"000001111",
  57809=>"111111111",
  57810=>"111111111",
  57811=>"000000000",
  57812=>"111111110",
  57813=>"111100100",
  57814=>"000000000",
  57815=>"000000000",
  57816=>"011011011",
  57817=>"011011000",
  57818=>"000000000",
  57819=>"000000000",
  57820=>"000000011",
  57821=>"000011000",
  57822=>"111111111",
  57823=>"110110011",
  57824=>"111111111",
  57825=>"001011111",
  57826=>"010000000",
  57827=>"000000000",
  57828=>"100000000",
  57829=>"000100100",
  57830=>"100000000",
  57831=>"111111111",
  57832=>"001001011",
  57833=>"111111110",
  57834=>"000000000",
  57835=>"111111111",
  57836=>"101001001",
  57837=>"001000011",
  57838=>"111111111",
  57839=>"000000000",
  57840=>"000000001",
  57841=>"111111111",
  57842=>"111111111",
  57843=>"100111111",
  57844=>"001101111",
  57845=>"111111111",
  57846=>"000000000",
  57847=>"011011001",
  57848=>"000001111",
  57849=>"001111111",
  57850=>"010000110",
  57851=>"001000100",
  57852=>"000010111",
  57853=>"000000000",
  57854=>"000000000",
  57855=>"001001000",
  57856=>"110110111",
  57857=>"000000000",
  57858=>"000000111",
  57859=>"001000010",
  57860=>"000000000",
  57861=>"000000001",
  57862=>"111011000",
  57863=>"111111111",
  57864=>"111110011",
  57865=>"100100110",
  57866=>"010000000",
  57867=>"110100010",
  57868=>"111111111",
  57869=>"011001100",
  57870=>"000000000",
  57871=>"111000111",
  57872=>"000000000",
  57873=>"000000010",
  57874=>"000100100",
  57875=>"101001011",
  57876=>"111000111",
  57877=>"000000000",
  57878=>"000000001",
  57879=>"000100100",
  57880=>"110110110",
  57881=>"001011110",
  57882=>"000100111",
  57883=>"111111001",
  57884=>"000000000",
  57885=>"111111111",
  57886=>"000000000",
  57887=>"000000001",
  57888=>"000111111",
  57889=>"111000000",
  57890=>"000000111",
  57891=>"100000000",
  57892=>"111111111",
  57893=>"111111111",
  57894=>"000000000",
  57895=>"101111100",
  57896=>"110111111",
  57897=>"000110111",
  57898=>"110111010",
  57899=>"100000000",
  57900=>"000001111",
  57901=>"000111111",
  57902=>"001011111",
  57903=>"000101111",
  57904=>"001110000",
  57905=>"111111001",
  57906=>"000000100",
  57907=>"001000000",
  57908=>"000001001",
  57909=>"001001001",
  57910=>"110111111",
  57911=>"101111111",
  57912=>"011011000",
  57913=>"000000000",
  57914=>"111111111",
  57915=>"000000000",
  57916=>"000110111",
  57917=>"000000100",
  57918=>"001001000",
  57919=>"001000101",
  57920=>"111010110",
  57921=>"000101000",
  57922=>"000100111",
  57923=>"111111111",
  57924=>"010110110",
  57925=>"001000100",
  57926=>"000000000",
  57927=>"111111111",
  57928=>"001000111",
  57929=>"011011011",
  57930=>"111111111",
  57931=>"000000101",
  57932=>"101001111",
  57933=>"110000001",
  57934=>"000000100",
  57935=>"110111000",
  57936=>"111001000",
  57937=>"000000011",
  57938=>"000000110",
  57939=>"000111111",
  57940=>"000000000",
  57941=>"000000000",
  57942=>"000000000",
  57943=>"000000000",
  57944=>"111110000",
  57945=>"100100100",
  57946=>"000111111",
  57947=>"100110101",
  57948=>"000101101",
  57949=>"110111111",
  57950=>"110110010",
  57951=>"000111111",
  57952=>"001000000",
  57953=>"100110110",
  57954=>"001000000",
  57955=>"110111110",
  57956=>"100000001",
  57957=>"000000001",
  57958=>"000000111",
  57959=>"100100100",
  57960=>"100100000",
  57961=>"111000000",
  57962=>"000000000",
  57963=>"110110000",
  57964=>"100110111",
  57965=>"101000101",
  57966=>"111101100",
  57967=>"110110110",
  57968=>"111100000",
  57969=>"000001111",
  57970=>"111111011",
  57971=>"111110000",
  57972=>"010010000",
  57973=>"001000000",
  57974=>"000001111",
  57975=>"001011111",
  57976=>"000000000",
  57977=>"000001001",
  57978=>"000011011",
  57979=>"000000001",
  57980=>"110110110",
  57981=>"000100000",
  57982=>"000000000",
  57983=>"000100101",
  57984=>"001111111",
  57985=>"000000111",
  57986=>"000010111",
  57987=>"000000000",
  57988=>"001001001",
  57989=>"111111010",
  57990=>"000000001",
  57991=>"000000011",
  57992=>"000000011",
  57993=>"010010011",
  57994=>"111011111",
  57995=>"000110000",
  57996=>"100001101",
  57997=>"000010010",
  57998=>"001000111",
  57999=>"101111001",
  58000=>"000000001",
  58001=>"000000000",
  58002=>"010010000",
  58003=>"111110110",
  58004=>"001000000",
  58005=>"111111010",
  58006=>"111000000",
  58007=>"000001001",
  58008=>"001000001",
  58009=>"111000001",
  58010=>"000000001",
  58011=>"000011011",
  58012=>"010000100",
  58013=>"111110000",
  58014=>"000111111",
  58015=>"101110110",
  58016=>"100000100",
  58017=>"111000000",
  58018=>"000000001",
  58019=>"111111111",
  58020=>"001001001",
  58021=>"011001000",
  58022=>"111111111",
  58023=>"000000001",
  58024=>"001011111",
  58025=>"000000111",
  58026=>"000000000",
  58027=>"000000101",
  58028=>"111111001",
  58029=>"111111101",
  58030=>"111111101",
  58031=>"111111111",
  58032=>"001111111",
  58033=>"110110000",
  58034=>"111111111",
  58035=>"101101001",
  58036=>"000001101",
  58037=>"011000001",
  58038=>"111111111",
  58039=>"001000000",
  58040=>"111101000",
  58041=>"111111110",
  58042=>"001001111",
  58043=>"110000000",
  58044=>"000110010",
  58045=>"000100110",
  58046=>"111101001",
  58047=>"001001001",
  58048=>"000110111",
  58049=>"000110000",
  58050=>"000000000",
  58051=>"000000111",
  58052=>"111111101",
  58053=>"111000000",
  58054=>"000000000",
  58055=>"001111000",
  58056=>"000110110",
  58057=>"111110011",
  58058=>"110111010",
  58059=>"011011000",
  58060=>"111000000",
  58061=>"010111110",
  58062=>"000000101",
  58063=>"011011000",
  58064=>"011111111",
  58065=>"110110110",
  58066=>"000000000",
  58067=>"000000001",
  58068=>"000000100",
  58069=>"100110110",
  58070=>"111111111",
  58071=>"000111111",
  58072=>"000000101",
  58073=>"000000000",
  58074=>"011111111",
  58075=>"000000000",
  58076=>"110000000",
  58077=>"000011001",
  58078=>"000100111",
  58079=>"000000000",
  58080=>"111111000",
  58081=>"000000000",
  58082=>"111000000",
  58083=>"111111111",
  58084=>"111111111",
  58085=>"011111011",
  58086=>"000110101",
  58087=>"000001001",
  58088=>"111000000",
  58089=>"101101000",
  58090=>"111111111",
  58091=>"000000101",
  58092=>"011111111",
  58093=>"001001111",
  58094=>"010000000",
  58095=>"000000111",
  58096=>"110111111",
  58097=>"111001011",
  58098=>"111111111",
  58099=>"000000001",
  58100=>"111000000",
  58101=>"000000111",
  58102=>"100111000",
  58103=>"110111011",
  58104=>"100111111",
  58105=>"000000000",
  58106=>"000001001",
  58107=>"000010111",
  58108=>"000000001",
  58109=>"110110110",
  58110=>"000000000",
  58111=>"111011001",
  58112=>"111101101",
  58113=>"001001001",
  58114=>"000111111",
  58115=>"111111000",
  58116=>"101000000",
  58117=>"000010110",
  58118=>"000000111",
  58119=>"001001001",
  58120=>"000111001",
  58121=>"000000000",
  58122=>"000000000",
  58123=>"000000000",
  58124=>"001000000",
  58125=>"110001111",
  58126=>"111110000",
  58127=>"010011111",
  58128=>"000110111",
  58129=>"000000000",
  58130=>"001000101",
  58131=>"000000000",
  58132=>"110111111",
  58133=>"010111111",
  58134=>"101101100",
  58135=>"000001001",
  58136=>"001001001",
  58137=>"000000000",
  58138=>"000010000",
  58139=>"111110111",
  58140=>"010111010",
  58141=>"000000000",
  58142=>"111001000",
  58143=>"000000110",
  58144=>"000111110",
  58145=>"010110110",
  58146=>"111111010",
  58147=>"111111111",
  58148=>"111100100",
  58149=>"011000100",
  58150=>"111111110",
  58151=>"000100111",
  58152=>"011001001",
  58153=>"111111010",
  58154=>"001001111",
  58155=>"110000110",
  58156=>"011001000",
  58157=>"000001001",
  58158=>"100100001",
  58159=>"000000000",
  58160=>"000000001",
  58161=>"000000000",
  58162=>"000000010",
  58163=>"000101110",
  58164=>"000000000",
  58165=>"010011000",
  58166=>"000000000",
  58167=>"111110111",
  58168=>"001111000",
  58169=>"000000000",
  58170=>"111111001",
  58171=>"111111111",
  58172=>"000000101",
  58173=>"000111100",
  58174=>"000000000",
  58175=>"010010111",
  58176=>"000000000",
  58177=>"000000000",
  58178=>"001000000",
  58179=>"111111101",
  58180=>"000000111",
  58181=>"000111111",
  58182=>"001011111",
  58183=>"011000000",
  58184=>"111001001",
  58185=>"111110000",
  58186=>"001001001",
  58187=>"000000110",
  58188=>"000000110",
  58189=>"000000000",
  58190=>"100001111",
  58191=>"000000000",
  58192=>"000000000",
  58193=>"110111111",
  58194=>"000000000",
  58195=>"000000000",
  58196=>"001001101",
  58197=>"011011001",
  58198=>"111000000",
  58199=>"111001000",
  58200=>"111110011",
  58201=>"101110111",
  58202=>"111110010",
  58203=>"110100111",
  58204=>"000000001",
  58205=>"000000101",
  58206=>"001001011",
  58207=>"111111111",
  58208=>"111111101",
  58209=>"111111000",
  58210=>"100100101",
  58211=>"111111111",
  58212=>"011011111",
  58213=>"000000001",
  58214=>"000000000",
  58215=>"111111111",
  58216=>"000000001",
  58217=>"000000000",
  58218=>"011110110",
  58219=>"111111110",
  58220=>"100110111",
  58221=>"100111111",
  58222=>"010110000",
  58223=>"111010000",
  58224=>"100000000",
  58225=>"011001000",
  58226=>"000000010",
  58227=>"111111000",
  58228=>"111111111",
  58229=>"000000000",
  58230=>"000000000",
  58231=>"000010010",
  58232=>"111111101",
  58233=>"010011001",
  58234=>"110110010",
  58235=>"011011111",
  58236=>"000111111",
  58237=>"001001101",
  58238=>"000000111",
  58239=>"111111111",
  58240=>"010110110",
  58241=>"000000000",
  58242=>"100000001",
  58243=>"111110010",
  58244=>"000000000",
  58245=>"010000000",
  58246=>"000110111",
  58247=>"000001101",
  58248=>"100110111",
  58249=>"000000000",
  58250=>"000000000",
  58251=>"111111001",
  58252=>"101101101",
  58253=>"000001111",
  58254=>"110111010",
  58255=>"100000000",
  58256=>"000000000",
  58257=>"000000000",
  58258=>"000000101",
  58259=>"000000001",
  58260=>"000000010",
  58261=>"000000000",
  58262=>"000000000",
  58263=>"001011011",
  58264=>"000000000",
  58265=>"000010010",
  58266=>"010000000",
  58267=>"001000000",
  58268=>"000101110",
  58269=>"110000011",
  58270=>"000001000",
  58271=>"100100110",
  58272=>"000000000",
  58273=>"010111111",
  58274=>"000000001",
  58275=>"111111000",
  58276=>"101001101",
  58277=>"000001101",
  58278=>"011001111",
  58279=>"110010000",
  58280=>"000000000",
  58281=>"000000000",
  58282=>"100110111",
  58283=>"000000000",
  58284=>"000000110",
  58285=>"110000100",
  58286=>"000000000",
  58287=>"001011101",
  58288=>"000000000",
  58289=>"111111111",
  58290=>"000000000",
  58291=>"110111111",
  58292=>"000100110",
  58293=>"101101111",
  58294=>"000001111",
  58295=>"000001001",
  58296=>"111101100",
  58297=>"000000000",
  58298=>"000000000",
  58299=>"000000100",
  58300=>"111111110",
  58301=>"000001101",
  58302=>"000111111",
  58303=>"101000101",
  58304=>"110111000",
  58305=>"011101101",
  58306=>"000000000",
  58307=>"111111111",
  58308=>"000000001",
  58309=>"111000100",
  58310=>"101001001",
  58311=>"000001111",
  58312=>"111101101",
  58313=>"111111111",
  58314=>"101001110",
  58315=>"111000000",
  58316=>"000000000",
  58317=>"010010001",
  58318=>"000000000",
  58319=>"000000000",
  58320=>"000000001",
  58321=>"110100000",
  58322=>"001101111",
  58323=>"011011000",
  58324=>"111111111",
  58325=>"111000000",
  58326=>"000001111",
  58327=>"000000000",
  58328=>"101101101",
  58329=>"111111111",
  58330=>"000110111",
  58331=>"111111010",
  58332=>"110111111",
  58333=>"000110111",
  58334=>"101001000",
  58335=>"100100001",
  58336=>"000001110",
  58337=>"001000000",
  58338=>"111111000",
  58339=>"111000000",
  58340=>"111110000",
  58341=>"000000111",
  58342=>"111110000",
  58343=>"000000000",
  58344=>"000000100",
  58345=>"001001001",
  58346=>"111000110",
  58347=>"001000001",
  58348=>"000000011",
  58349=>"001000100",
  58350=>"000000111",
  58351=>"000110110",
  58352=>"001001001",
  58353=>"000000110",
  58354=>"011111011",
  58355=>"111110000",
  58356=>"111111111",
  58357=>"000001000",
  58358=>"111111001",
  58359=>"000011011",
  58360=>"010111111",
  58361=>"000001000",
  58362=>"000001001",
  58363=>"101100100",
  58364=>"000000000",
  58365=>"001000000",
  58366=>"111111111",
  58367=>"011001101",
  58368=>"100000000",
  58369=>"110010000",
  58370=>"111110110",
  58371=>"010000000",
  58372=>"000110110",
  58373=>"001000000",
  58374=>"111001011",
  58375=>"111111111",
  58376=>"000011011",
  58377=>"000000000",
  58378=>"111111000",
  58379=>"111111111",
  58380=>"110110110",
  58381=>"111111001",
  58382=>"111000111",
  58383=>"000000011",
  58384=>"100000000",
  58385=>"010111110",
  58386=>"111010000",
  58387=>"000000000",
  58388=>"111111111",
  58389=>"110111111",
  58390=>"000000000",
  58391=>"111111110",
  58392=>"111111111",
  58393=>"001001011",
  58394=>"111111111",
  58395=>"111001000",
  58396=>"111111111",
  58397=>"111111111",
  58398=>"000000010",
  58399=>"000000100",
  58400=>"110110000",
  58401=>"001001001",
  58402=>"011011111",
  58403=>"110111011",
  58404=>"111111111",
  58405=>"001100000",
  58406=>"011000000",
  58407=>"111111011",
  58408=>"000000000",
  58409=>"110110100",
  58410=>"000000000",
  58411=>"000000000",
  58412=>"100111111",
  58413=>"000000000",
  58414=>"000000000",
  58415=>"111111110",
  58416=>"011011000",
  58417=>"111111111",
  58418=>"001111111",
  58419=>"000000000",
  58420=>"000111111",
  58421=>"000000011",
  58422=>"111001000",
  58423=>"000000000",
  58424=>"000000000",
  58425=>"100100100",
  58426=>"000000000",
  58427=>"110111110",
  58428=>"101000100",
  58429=>"111001000",
  58430=>"111111011",
  58431=>"111111111",
  58432=>"110010010",
  58433=>"111111111",
  58434=>"011111000",
  58435=>"001001001",
  58436=>"110110000",
  58437=>"000111110",
  58438=>"111011011",
  58439=>"000000000",
  58440=>"110110111",
  58441=>"111111111",
  58442=>"000000000",
  58443=>"100001011",
  58444=>"001000010",
  58445=>"111111000",
  58446=>"000000000",
  58447=>"000000000",
  58448=>"000000000",
  58449=>"111111000",
  58450=>"000000000",
  58451=>"100000000",
  58452=>"000000000",
  58453=>"000000000",
  58454=>"000000000",
  58455=>"000000010",
  58456=>"000000000",
  58457=>"100000000",
  58458=>"000000000",
  58459=>"000000011",
  58460=>"111101000",
  58461=>"000000000",
  58462=>"000000001",
  58463=>"111111111",
  58464=>"000000000",
  58465=>"001000000",
  58466=>"000110110",
  58467=>"000101111",
  58468=>"000000011",
  58469=>"010000000",
  58470=>"001001111",
  58471=>"110110100",
  58472=>"000110111",
  58473=>"100101111",
  58474=>"000000000",
  58475=>"111111111",
  58476=>"101100000",
  58477=>"111111111",
  58478=>"111000011",
  58479=>"000001001",
  58480=>"000000000",
  58481=>"111111111",
  58482=>"110110000",
  58483=>"000001000",
  58484=>"111000100",
  58485=>"000000000",
  58486=>"000100111",
  58487=>"110011001",
  58488=>"111111111",
  58489=>"111111100",
  58490=>"011010000",
  58491=>"111000000",
  58492=>"100110110",
  58493=>"111111010",
  58494=>"010000000",
  58495=>"000000000",
  58496=>"000111111",
  58497=>"111111011",
  58498=>"000000000",
  58499=>"000000000",
  58500=>"000000000",
  58501=>"111000000",
  58502=>"000000000",
  58503=>"000001001",
  58504=>"111000000",
  58505=>"111011111",
  58506=>"000001011",
  58507=>"110000000",
  58508=>"000110111",
  58509=>"111111111",
  58510=>"111111111",
  58511=>"111100001",
  58512=>"000000111",
  58513=>"100001001",
  58514=>"000000101",
  58515=>"100111111",
  58516=>"000100001",
  58517=>"011111000",
  58518=>"000000000",
  58519=>"000000000",
  58520=>"111100000",
  58521=>"111111110",
  58522=>"111110100",
  58523=>"000000111",
  58524=>"111111111",
  58525=>"000000101",
  58526=>"111111110",
  58527=>"000000000",
  58528=>"000000111",
  58529=>"110110010",
  58530=>"110111111",
  58531=>"000000010",
  58532=>"111111000",
  58533=>"001000000",
  58534=>"111101001",
  58535=>"000110010",
  58536=>"111000000",
  58537=>"111100111",
  58538=>"000000000",
  58539=>"011000000",
  58540=>"111110110",
  58541=>"000010111",
  58542=>"111100000",
  58543=>"110111111",
  58544=>"111111000",
  58545=>"000000011",
  58546=>"111111111",
  58547=>"000001111",
  58548=>"011011011",
  58549=>"000001000",
  58550=>"100111011",
  58551=>"100100111",
  58552=>"001001000",
  58553=>"111111111",
  58554=>"011011000",
  58555=>"111110111",
  58556=>"000000010",
  58557=>"000011001",
  58558=>"111111111",
  58559=>"111111111",
  58560=>"111111111",
  58561=>"000000000",
  58562=>"000000000",
  58563=>"000000011",
  58564=>"110111010",
  58565=>"000000111",
  58566=>"000000000",
  58567=>"000000000",
  58568=>"011011010",
  58569=>"111000000",
  58570=>"110100001",
  58571=>"111010000",
  58572=>"000011111",
  58573=>"000000000",
  58574=>"000000110",
  58575=>"000000000",
  58576=>"000000010",
  58577=>"000000000",
  58578=>"111111111",
  58579=>"000000000",
  58580=>"001001011",
  58581=>"111111111",
  58582=>"000000001",
  58583=>"000000000",
  58584=>"111111111",
  58585=>"000000000",
  58586=>"101111111",
  58587=>"010000000",
  58588=>"000000000",
  58589=>"111111011",
  58590=>"111111111",
  58591=>"110000000",
  58592=>"000000001",
  58593=>"000000000",
  58594=>"110110000",
  58595=>"011000000",
  58596=>"001000000",
  58597=>"011011111",
  58598=>"001011000",
  58599=>"000000000",
  58600=>"111111011",
  58601=>"000000000",
  58602=>"111000000",
  58603=>"000000000",
  58604=>"000000001",
  58605=>"000000000",
  58606=>"000000111",
  58607=>"010000010",
  58608=>"100100000",
  58609=>"000010000",
  58610=>"111111011",
  58611=>"111011000",
  58612=>"000000000",
  58613=>"110010001",
  58614=>"000000100",
  58615=>"111001101",
  58616=>"000000001",
  58617=>"111111111",
  58618=>"111000001",
  58619=>"000000000",
  58620=>"001011001",
  58621=>"111000001",
  58622=>"111111000",
  58623=>"000000000",
  58624=>"000000000",
  58625=>"000000001",
  58626=>"111111111",
  58627=>"010000000",
  58628=>"000000101",
  58629=>"000000000",
  58630=>"111111111",
  58631=>"110000000",
  58632=>"000000000",
  58633=>"000100100",
  58634=>"001001001",
  58635=>"001000000",
  58636=>"000001101",
  58637=>"000000000",
  58638=>"111111100",
  58639=>"000000000",
  58640=>"111111111",
  58641=>"111111111",
  58642=>"101000100",
  58643=>"100111111",
  58644=>"000000000",
  58645=>"100111000",
  58646=>"000000001",
  58647=>"111111111",
  58648=>"101001001",
  58649=>"011011011",
  58650=>"111111101",
  58651=>"100000000",
  58652=>"010110110",
  58653=>"000000000",
  58654=>"000000000",
  58655=>"111111111",
  58656=>"010010011",
  58657=>"011110111",
  58658=>"111111010",
  58659=>"111111111",
  58660=>"100100100",
  58661=>"111001000",
  58662=>"001001000",
  58663=>"100000100",
  58664=>"110100111",
  58665=>"000000000",
  58666=>"111000100",
  58667=>"111111111",
  58668=>"111111111",
  58669=>"011001000",
  58670=>"111000000",
  58671=>"000000000",
  58672=>"110011011",
  58673=>"000000000",
  58674=>"000000100",
  58675=>"110110110",
  58676=>"000000000",
  58677=>"000000000",
  58678=>"000000011",
  58679=>"000000000",
  58680=>"111111000",
  58681=>"111001100",
  58682=>"111111111",
  58683=>"000000000",
  58684=>"001000000",
  58685=>"111111111",
  58686=>"000111011",
  58687=>"111100111",
  58688=>"001000110",
  58689=>"101001001",
  58690=>"111111111",
  58691=>"111011100",
  58692=>"000000100",
  58693=>"011000001",
  58694=>"010010000",
  58695=>"000011111",
  58696=>"101100111",
  58697=>"110110111",
  58698=>"000000100",
  58699=>"000000001",
  58700=>"110000000",
  58701=>"011011111",
  58702=>"011000000",
  58703=>"000000000",
  58704=>"101111111",
  58705=>"010000110",
  58706=>"111100000",
  58707=>"000111111",
  58708=>"000010000",
  58709=>"011011011",
  58710=>"000000000",
  58711=>"100000111",
  58712=>"110111111",
  58713=>"111011111",
  58714=>"000000000",
  58715=>"000000000",
  58716=>"000100100",
  58717=>"111111111",
  58718=>"111111100",
  58719=>"010000000",
  58720=>"000000100",
  58721=>"111111111",
  58722=>"110110111",
  58723=>"101000001",
  58724=>"111111111",
  58725=>"111011001",
  58726=>"000001001",
  58727=>"111111111",
  58728=>"001000000",
  58729=>"000000000",
  58730=>"000000000",
  58731=>"001101110",
  58732=>"111011010",
  58733=>"011000000",
  58734=>"000000000",
  58735=>"000111111",
  58736=>"001111111",
  58737=>"000000000",
  58738=>"110110111",
  58739=>"111111011",
  58740=>"111110000",
  58741=>"000000000",
  58742=>"111111111",
  58743=>"000001000",
  58744=>"000000000",
  58745=>"111111011",
  58746=>"100100111",
  58747=>"000111111",
  58748=>"000100000",
  58749=>"111001101",
  58750=>"111111111",
  58751=>"111111111",
  58752=>"000000010",
  58753=>"111111111",
  58754=>"001011001",
  58755=>"111111000",
  58756=>"000000000",
  58757=>"111111110",
  58758=>"000100010",
  58759=>"100000000",
  58760=>"000000000",
  58761=>"111111110",
  58762=>"000000000",
  58763=>"000000000",
  58764=>"100111111",
  58765=>"011011011",
  58766=>"000000111",
  58767=>"000111111",
  58768=>"100000000",
  58769=>"111111111",
  58770=>"110100000",
  58771=>"000000000",
  58772=>"111111111",
  58773=>"010111110",
  58774=>"000000001",
  58775=>"011010000",
  58776=>"000000000",
  58777=>"110110001",
  58778=>"111000000",
  58779=>"000000000",
  58780=>"111000001",
  58781=>"000000000",
  58782=>"100100000",
  58783=>"000000000",
  58784=>"111111111",
  58785=>"111110110",
  58786=>"111111111",
  58787=>"111111000",
  58788=>"000000001",
  58789=>"111111000",
  58790=>"011111111",
  58791=>"111111111",
  58792=>"110100111",
  58793=>"111000000",
  58794=>"000000000",
  58795=>"111011011",
  58796=>"000000001",
  58797=>"000000000",
  58798=>"000000000",
  58799=>"110111111",
  58800=>"000000101",
  58801=>"111111111",
  58802=>"111111110",
  58803=>"000000111",
  58804=>"000000000",
  58805=>"111111000",
  58806=>"000110111",
  58807=>"000100111",
  58808=>"000111111",
  58809=>"011001000",
  58810=>"000000110",
  58811=>"111111111",
  58812=>"000100111",
  58813=>"111111110",
  58814=>"001101000",
  58815=>"010010000",
  58816=>"111000011",
  58817=>"111111111",
  58818=>"111111111",
  58819=>"111111111",
  58820=>"011001011",
  58821=>"001111110",
  58822=>"000000000",
  58823=>"001111111",
  58824=>"011010000",
  58825=>"111111111",
  58826=>"110000111",
  58827=>"110000000",
  58828=>"000000000",
  58829=>"000000000",
  58830=>"110100100",
  58831=>"000000100",
  58832=>"000000100",
  58833=>"000001111",
  58834=>"001101000",
  58835=>"111111101",
  58836=>"001000001",
  58837=>"000000000",
  58838=>"000000000",
  58839=>"001111110",
  58840=>"111000011",
  58841=>"111000000",
  58842=>"011001111",
  58843=>"000000000",
  58844=>"010111111",
  58845=>"111111111",
  58846=>"111110111",
  58847=>"111110000",
  58848=>"000000000",
  58849=>"111011000",
  58850=>"111011110",
  58851=>"111111011",
  58852=>"111011001",
  58853=>"011111111",
  58854=>"110100111",
  58855=>"000110111",
  58856=>"111111111",
  58857=>"000001001",
  58858=>"000100100",
  58859=>"011011000",
  58860=>"111111111",
  58861=>"010000000",
  58862=>"000000010",
  58863=>"111111111",
  58864=>"011011010",
  58865=>"000000111",
  58866=>"111111111",
  58867=>"000000100",
  58868=>"111111111",
  58869=>"011000000",
  58870=>"000000000",
  58871=>"000000111",
  58872=>"111110010",
  58873=>"111101001",
  58874=>"111111010",
  58875=>"000000000",
  58876=>"011000001",
  58877=>"100000000",
  58878=>"111111011",
  58879=>"111111111",
  58880=>"110000011",
  58881=>"111000001",
  58882=>"111111111",
  58883=>"000100101",
  58884=>"001001011",
  58885=>"100111111",
  58886=>"001000000",
  58887=>"101111111",
  58888=>"000000000",
  58889=>"111111111",
  58890=>"000000111",
  58891=>"011011111",
  58892=>"001011111",
  58893=>"000000000",
  58894=>"000100110",
  58895=>"111111001",
  58896=>"000000100",
  58897=>"011011111",
  58898=>"000000001",
  58899=>"010111111",
  58900=>"110110010",
  58901=>"111000000",
  58902=>"001000001",
  58903=>"111111011",
  58904=>"000000000",
  58905=>"100101111",
  58906=>"000010000",
  58907=>"101111111",
  58908=>"111111010",
  58909=>"111000000",
  58910=>"110110000",
  58911=>"010111110",
  58912=>"000000010",
  58913=>"110111111",
  58914=>"100111111",
  58915=>"011111111",
  58916=>"000100001",
  58917=>"111111000",
  58918=>"110110111",
  58919=>"111111111",
  58920=>"000000100",
  58921=>"000000000",
  58922=>"000111111",
  58923=>"000010000",
  58924=>"010000000",
  58925=>"001111111",
  58926=>"111111100",
  58927=>"100000010",
  58928=>"111100100",
  58929=>"000000000",
  58930=>"110000000",
  58931=>"010010000",
  58932=>"110111111",
  58933=>"111001011",
  58934=>"011111111",
  58935=>"001000100",
  58936=>"111000000",
  58937=>"110110100",
  58938=>"000001111",
  58939=>"110101000",
  58940=>"111111111",
  58941=>"000000010",
  58942=>"111111100",
  58943=>"000101111",
  58944=>"000100100",
  58945=>"001011000",
  58946=>"000001000",
  58947=>"000000100",
  58948=>"000000110",
  58949=>"011111111",
  58950=>"001111111",
  58951=>"000000000",
  58952=>"110111111",
  58953=>"111000100",
  58954=>"000000000",
  58955=>"110111100",
  58956=>"000111101",
  58957=>"111111111",
  58958=>"111111111",
  58959=>"000011111",
  58960=>"111111111",
  58961=>"000001001",
  58962=>"100100000",
  58963=>"000000001",
  58964=>"111111100",
  58965=>"011111100",
  58966=>"000000000",
  58967=>"110111111",
  58968=>"011111110",
  58969=>"000000101",
  58970=>"001000001",
  58971=>"111100100",
  58972=>"000000000",
  58973=>"111111111",
  58974=>"110110110",
  58975=>"100100100",
  58976=>"111111000",
  58977=>"000000000",
  58978=>"100111111",
  58979=>"000001000",
  58980=>"001001000",
  58981=>"000000000",
  58982=>"100111111",
  58983=>"000001011",
  58984=>"000000100",
  58985=>"110100100",
  58986=>"000000011",
  58987=>"111111111",
  58988=>"011111001",
  58989=>"010110111",
  58990=>"000000000",
  58991=>"000010110",
  58992=>"000000000",
  58993=>"000000000",
  58994=>"000010110",
  58995=>"110011011",
  58996=>"000111000",
  58997=>"000111000",
  58998=>"011111000",
  58999=>"000000000",
  59000=>"010011111",
  59001=>"110100110",
  59002=>"000001001",
  59003=>"111111000",
  59004=>"111111110",
  59005=>"000100100",
  59006=>"000110111",
  59007=>"110110000",
  59008=>"001010110",
  59009=>"110111101",
  59010=>"000000111",
  59011=>"110100110",
  59012=>"011001101",
  59013=>"110000000",
  59014=>"010110110",
  59015=>"111011111",
  59016=>"101000000",
  59017=>"111110000",
  59018=>"000000000",
  59019=>"001000000",
  59020=>"100000010",
  59021=>"000000000",
  59022=>"100000100",
  59023=>"000000000",
  59024=>"000000000",
  59025=>"111000000",
  59026=>"010000000",
  59027=>"000000000",
  59028=>"000000000",
  59029=>"111111111",
  59030=>"000000101",
  59031=>"111111111",
  59032=>"000000011",
  59033=>"000000000",
  59034=>"000001011",
  59035=>"001000000",
  59036=>"011000000",
  59037=>"000000000",
  59038=>"111111111",
  59039=>"000000000",
  59040=>"110110110",
  59041=>"101001000",
  59042=>"111000000",
  59043=>"111100110",
  59044=>"000000000",
  59045=>"110111110",
  59046=>"111111110",
  59047=>"010110111",
  59048=>"001101111",
  59049=>"000000000",
  59050=>"000100111",
  59051=>"110111000",
  59052=>"111011000",
  59053=>"100110111",
  59054=>"101101111",
  59055=>"111001000",
  59056=>"000100101",
  59057=>"111111111",
  59058=>"111111111",
  59059=>"000000000",
  59060=>"111011000",
  59061=>"001000111",
  59062=>"000000000",
  59063=>"110000000",
  59064=>"100100100",
  59065=>"111111111",
  59066=>"011000111",
  59067=>"001000001",
  59068=>"111111001",
  59069=>"011000000",
  59070=>"111111111",
  59071=>"011000000",
  59072=>"111111011",
  59073=>"111111100",
  59074=>"111100000",
  59075=>"001111111",
  59076=>"111111111",
  59077=>"000000110",
  59078=>"000001001",
  59079=>"111111111",
  59080=>"001000110",
  59081=>"100111011",
  59082=>"110111110",
  59083=>"111101111",
  59084=>"101111101",
  59085=>"111101100",
  59086=>"000000010",
  59087=>"101000000",
  59088=>"101111111",
  59089=>"111111110",
  59090=>"000110111",
  59091=>"111101111",
  59092=>"100100101",
  59093=>"000000000",
  59094=>"100111111",
  59095=>"010111111",
  59096=>"000000111",
  59097=>"111111000",
  59098=>"111000000",
  59099=>"011111100",
  59100=>"000000000",
  59101=>"111111100",
  59102=>"010010110",
  59103=>"100000000",
  59104=>"111111111",
  59105=>"000101111",
  59106=>"111111111",
  59107=>"000000000",
  59108=>"000000000",
  59109=>"000000000",
  59110=>"111100000",
  59111=>"011111111",
  59112=>"000000000",
  59113=>"000000000",
  59114=>"011011001",
  59115=>"111110111",
  59116=>"111111011",
  59117=>"111111111",
  59118=>"111101001",
  59119=>"001000000",
  59120=>"011111111",
  59121=>"000000000",
  59122=>"101000001",
  59123=>"001000000",
  59124=>"000011111",
  59125=>"001001001",
  59126=>"111110000",
  59127=>"111111100",
  59128=>"111111111",
  59129=>"010000010",
  59130=>"000011011",
  59131=>"000100111",
  59132=>"011011111",
  59133=>"110111000",
  59134=>"111111100",
  59135=>"100111111",
  59136=>"110110111",
  59137=>"111111110",
  59138=>"111111110",
  59139=>"010111111",
  59140=>"111111111",
  59141=>"110000000",
  59142=>"111111110",
  59143=>"100000000",
  59144=>"010011111",
  59145=>"000000000",
  59146=>"000000000",
  59147=>"000011111",
  59148=>"111111111",
  59149=>"111011111",
  59150=>"111111110",
  59151=>"000101111",
  59152=>"111100000",
  59153=>"100100100",
  59154=>"110110011",
  59155=>"000000000",
  59156=>"111111111",
  59157=>"111011111",
  59158=>"101001101",
  59159=>"000111111",
  59160=>"000011111",
  59161=>"001011111",
  59162=>"011010011",
  59163=>"111111000",
  59164=>"000000000",
  59165=>"100101111",
  59166=>"111111111",
  59167=>"000000000",
  59168=>"100001110",
  59169=>"011000011",
  59170=>"111110000",
  59171=>"101101111",
  59172=>"111001000",
  59173=>"000000001",
  59174=>"000100110",
  59175=>"001000110",
  59176=>"001001100",
  59177=>"000000000",
  59178=>"110110111",
  59179=>"110110010",
  59180=>"000000000",
  59181=>"111111111",
  59182=>"000000000",
  59183=>"000000111",
  59184=>"011111111",
  59185=>"000000000",
  59186=>"001110110",
  59187=>"111011111",
  59188=>"000000000",
  59189=>"111111110",
  59190=>"110000000",
  59191=>"001000000",
  59192=>"000101111",
  59193=>"111001000",
  59194=>"011010000",
  59195=>"011000000",
  59196=>"110000011",
  59197=>"111111000",
  59198=>"000000000",
  59199=>"111111001",
  59200=>"110111111",
  59201=>"111001001",
  59202=>"000000010",
  59203=>"101001000",
  59204=>"011111111",
  59205=>"000000000",
  59206=>"111111111",
  59207=>"111111111",
  59208=>"000000000",
  59209=>"011000000",
  59210=>"001001011",
  59211=>"011011011",
  59212=>"001000100",
  59213=>"000111111",
  59214=>"000001001",
  59215=>"111111000",
  59216=>"110011010",
  59217=>"001101101",
  59218=>"001001111",
  59219=>"000000010",
  59220=>"110100000",
  59221=>"000000000",
  59222=>"111100111",
  59223=>"000100110",
  59224=>"111000000",
  59225=>"111111111",
  59226=>"111111111",
  59227=>"111111111",
  59228=>"000000111",
  59229=>"111111011",
  59230=>"001000000",
  59231=>"110111111",
  59232=>"000000111",
  59233=>"000001111",
  59234=>"011011000",
  59235=>"100001001",
  59236=>"000011111",
  59237=>"111111111",
  59238=>"110111100",
  59239=>"100100100",
  59240=>"110111111",
  59241=>"110111000",
  59242=>"000000000",
  59243=>"000111111",
  59244=>"001001111",
  59245=>"011111111",
  59246=>"000000000",
  59247=>"111111101",
  59248=>"001111100",
  59249=>"011000000",
  59250=>"111111100",
  59251=>"000101111",
  59252=>"011010000",
  59253=>"111111111",
  59254=>"110100100",
  59255=>"011000111",
  59256=>"000000000",
  59257=>"111111111",
  59258=>"010011010",
  59259=>"000000000",
  59260=>"000111101",
  59261=>"111111111",
  59262=>"011001000",
  59263=>"000000001",
  59264=>"001011111",
  59265=>"000000000",
  59266=>"110110110",
  59267=>"001011011",
  59268=>"110111110",
  59269=>"111111011",
  59270=>"111011000",
  59271=>"001000000",
  59272=>"001000000",
  59273=>"001001000",
  59274=>"111100110",
  59275=>"101101101",
  59276=>"111111101",
  59277=>"111000000",
  59278=>"000000000",
  59279=>"111011001",
  59280=>"011110000",
  59281=>"000000111",
  59282=>"111110110",
  59283=>"101101110",
  59284=>"111111111",
  59285=>"000010011",
  59286=>"100110110",
  59287=>"001001001",
  59288=>"111111000",
  59289=>"000000000",
  59290=>"110110111",
  59291=>"000000000",
  59292=>"011000111",
  59293=>"011111111",
  59294=>"111001011",
  59295=>"000111111",
  59296=>"001000000",
  59297=>"000010011",
  59298=>"001010000",
  59299=>"000000100",
  59300=>"000000000",
  59301=>"111111111",
  59302=>"001000000",
  59303=>"111000000",
  59304=>"101000000",
  59305=>"100010110",
  59306=>"001000000",
  59307=>"111111111",
  59308=>"000010111",
  59309=>"111110110",
  59310=>"000000000",
  59311=>"000000000",
  59312=>"000000000",
  59313=>"000000000",
  59314=>"111111000",
  59315=>"111111111",
  59316=>"111111111",
  59317=>"000000000",
  59318=>"111110100",
  59319=>"111111111",
  59320=>"111110100",
  59321=>"111111111",
  59322=>"111011111",
  59323=>"000000000",
  59324=>"011111111",
  59325=>"000000000",
  59326=>"111101111",
  59327=>"110000100",
  59328=>"000001000",
  59329=>"110010010",
  59330=>"001000000",
  59331=>"000010110",
  59332=>"111001000",
  59333=>"111110100",
  59334=>"110110000",
  59335=>"111111111",
  59336=>"000111011",
  59337=>"000000000",
  59338=>"000000100",
  59339=>"111111111",
  59340=>"111100000",
  59341=>"000010000",
  59342=>"000010011",
  59343=>"000100000",
  59344=>"000000001",
  59345=>"001001111",
  59346=>"111111110",
  59347=>"111111111",
  59348=>"001111111",
  59349=>"111111001",
  59350=>"110110110",
  59351=>"111011001",
  59352=>"001001111",
  59353=>"111111100",
  59354=>"011111011",
  59355=>"001000000",
  59356=>"000000000",
  59357=>"000001111",
  59358=>"111110000",
  59359=>"011001000",
  59360=>"110000010",
  59361=>"001000000",
  59362=>"110111111",
  59363=>"000111111",
  59364=>"111011111",
  59365=>"000000110",
  59366=>"101001011",
  59367=>"000000111",
  59368=>"111111111",
  59369=>"111111111",
  59370=>"110111111",
  59371=>"111111111",
  59372=>"100110111",
  59373=>"000000000",
  59374=>"111111111",
  59375=>"111011001",
  59376=>"001000000",
  59377=>"111111111",
  59378=>"000000000",
  59379=>"000001111",
  59380=>"000001001",
  59381=>"111111101",
  59382=>"100000000",
  59383=>"100100000",
  59384=>"111111110",
  59385=>"001000000",
  59386=>"011111111",
  59387=>"111111011",
  59388=>"111110101",
  59389=>"000001000",
  59390=>"111110110",
  59391=>"111111111",
  59392=>"000000000",
  59393=>"000110000",
  59394=>"100100100",
  59395=>"011111111",
  59396=>"001000000",
  59397=>"001011111",
  59398=>"000000000",
  59399=>"111111111",
  59400=>"111000110",
  59401=>"111111000",
  59402=>"111101101",
  59403=>"100000000",
  59404=>"000010111",
  59405=>"000000100",
  59406=>"000100001",
  59407=>"111111101",
  59408=>"000000001",
  59409=>"000000011",
  59410=>"000000101",
  59411=>"111111111",
  59412=>"111100000",
  59413=>"010000000",
  59414=>"111111111",
  59415=>"111111110",
  59416=>"100100000",
  59417=>"011011011",
  59418=>"010000000",
  59419=>"111111010",
  59420=>"111111111",
  59421=>"000101111",
  59422=>"111111111",
  59423=>"000000000",
  59424=>"001111111",
  59425=>"000100100",
  59426=>"111000000",
  59427=>"100000001",
  59428=>"111011111",
  59429=>"111111011",
  59430=>"011011000",
  59431=>"111001000",
  59432=>"000000000",
  59433=>"000000000",
  59434=>"111111101",
  59435=>"111111111",
  59436=>"111001111",
  59437=>"111111111",
  59438=>"111111110",
  59439=>"111110110",
  59440=>"111011110",
  59441=>"000001001",
  59442=>"111111111",
  59443=>"110110000",
  59444=>"111000000",
  59445=>"000000111",
  59446=>"111111111",
  59447=>"100100000",
  59448=>"110110100",
  59449=>"001011001",
  59450=>"000000000",
  59451=>"111111111",
  59452=>"011000011",
  59453=>"011111111",
  59454=>"000000000",
  59455=>"100100100",
  59456=>"001000000",
  59457=>"111111100",
  59458=>"000000000",
  59459=>"111111111",
  59460=>"000001101",
  59461=>"111010000",
  59462=>"100111000",
  59463=>"111111111",
  59464=>"111011001",
  59465=>"111001101",
  59466=>"000000000",
  59467=>"001011110",
  59468=>"000110000",
  59469=>"100000111",
  59470=>"101000000",
  59471=>"000000000",
  59472=>"000000000",
  59473=>"000000001",
  59474=>"100000000",
  59475=>"000100110",
  59476=>"000000000",
  59477=>"000010001",
  59478=>"000000000",
  59479=>"000000111",
  59480=>"000001111",
  59481=>"000000100",
  59482=>"100001111",
  59483=>"000101111",
  59484=>"000110000",
  59485=>"111111111",
  59486=>"111111000",
  59487=>"111111100",
  59488=>"001111111",
  59489=>"110011111",
  59490=>"111111110",
  59491=>"011111111",
  59492=>"001101110",
  59493=>"000000000",
  59494=>"111000000",
  59495=>"111110100",
  59496=>"010110110",
  59497=>"011110011",
  59498=>"100001000",
  59499=>"000000111",
  59500=>"001001000",
  59501=>"000000111",
  59502=>"111111111",
  59503=>"000000000",
  59504=>"111111000",
  59505=>"001111111",
  59506=>"011000001",
  59507=>"111011000",
  59508=>"110111000",
  59509=>"111111111",
  59510=>"111111111",
  59511=>"000000000",
  59512=>"000000001",
  59513=>"010001111",
  59514=>"000000011",
  59515=>"000000111",
  59516=>"110110100",
  59517=>"101111110",
  59518=>"111111111",
  59519=>"010111111",
  59520=>"100100111",
  59521=>"011000000",
  59522=>"000000000",
  59523=>"001011011",
  59524=>"110010000",
  59525=>"111111101",
  59526=>"001000000",
  59527=>"000000000",
  59528=>"000000000",
  59529=>"111000000",
  59530=>"000000000",
  59531=>"000001111",
  59532=>"111111011",
  59533=>"000000000",
  59534=>"101111011",
  59535=>"111111001",
  59536=>"000000001",
  59537=>"010010011",
  59538=>"011001000",
  59539=>"111011000",
  59540=>"001011000",
  59541=>"000001000",
  59542=>"111111000",
  59543=>"000000101",
  59544=>"100100100",
  59545=>"111010010",
  59546=>"010100110",
  59547=>"001001000",
  59548=>"111111111",
  59549=>"111111001",
  59550=>"001010111",
  59551=>"000000001",
  59552=>"100110110",
  59553=>"011011000",
  59554=>"111111111",
  59555=>"111111111",
  59556=>"001001011",
  59557=>"000111111",
  59558=>"111111111",
  59559=>"001001001",
  59560=>"100000000",
  59561=>"011111011",
  59562=>"111111111",
  59563=>"000000000",
  59564=>"011000000",
  59565=>"110110111",
  59566=>"111111111",
  59567=>"000100000",
  59568=>"000000000",
  59569=>"111111101",
  59570=>"111000000",
  59571=>"111111111",
  59572=>"011000000",
  59573=>"111111111",
  59574=>"000000111",
  59575=>"001001111",
  59576=>"011111111",
  59577=>"111001000",
  59578=>"000000000",
  59579=>"000000010",
  59580=>"110110110",
  59581=>"000000000",
  59582=>"111110111",
  59583=>"111111000",
  59584=>"111000000",
  59585=>"000001011",
  59586=>"000000000",
  59587=>"111101000",
  59588=>"001000000",
  59589=>"110100111",
  59590=>"011011110",
  59591=>"000010000",
  59592=>"111001000",
  59593=>"011111111",
  59594=>"011111100",
  59595=>"000000000",
  59596=>"111111111",
  59597=>"111111000",
  59598=>"001001101",
  59599=>"000000001",
  59600=>"111100100",
  59601=>"111101000",
  59602=>"011111111",
  59603=>"000010111",
  59604=>"011110111",
  59605=>"111111110",
  59606=>"000001000",
  59607=>"111000000",
  59608=>"111111111",
  59609=>"100000111",
  59610=>"111111111",
  59611=>"111111111",
  59612=>"000000001",
  59613=>"100110111",
  59614=>"000000000",
  59615=>"111100001",
  59616=>"000000000",
  59617=>"111110111",
  59618=>"111111111",
  59619=>"111111101",
  59620=>"111111111",
  59621=>"001001111",
  59622=>"000000000",
  59623=>"111111101",
  59624=>"111011011",
  59625=>"000111000",
  59626=>"111111001",
  59627=>"000000110",
  59628=>"111111000",
  59629=>"000000000",
  59630=>"000000000",
  59631=>"111111001",
  59632=>"111000000",
  59633=>"000000000",
  59634=>"111111111",
  59635=>"001111111",
  59636=>"111111111",
  59637=>"000000100",
  59638=>"111111110",
  59639=>"000000000",
  59640=>"111000000",
  59641=>"111110100",
  59642=>"000101111",
  59643=>"011000000",
  59644=>"111110111",
  59645=>"111111101",
  59646=>"100001000",
  59647=>"111000000",
  59648=>"111101101",
  59649=>"011011011",
  59650=>"010000001",
  59651=>"111111111",
  59652=>"100000000",
  59653=>"111111111",
  59654=>"110110011",
  59655=>"101001000",
  59656=>"000000000",
  59657=>"111000000",
  59658=>"110110100",
  59659=>"000000000",
  59660=>"111100100",
  59661=>"000000000",
  59662=>"111111111",
  59663=>"111110000",
  59664=>"000100000",
  59665=>"010000000",
  59666=>"111111111",
  59667=>"111110111",
  59668=>"111111111",
  59669=>"000000000",
  59670=>"111100100",
  59671=>"000000000",
  59672=>"111111110",
  59673=>"000001001",
  59674=>"000000000",
  59675=>"111100001",
  59676=>"111111111",
  59677=>"111111111",
  59678=>"110111111",
  59679=>"111111111",
  59680=>"110111000",
  59681=>"000100000",
  59682=>"011110110",
  59683=>"000000100",
  59684=>"111111111",
  59685=>"000000100",
  59686=>"111011011",
  59687=>"001001001",
  59688=>"000111111",
  59689=>"111111100",
  59690=>"111110110",
  59691=>"000000100",
  59692=>"000000001",
  59693=>"011010011",
  59694=>"000000011",
  59695=>"100100001",
  59696=>"001000000",
  59697=>"000100000",
  59698=>"011111111",
  59699=>"110010000",
  59700=>"100000001",
  59701=>"000000000",
  59702=>"000000111",
  59703=>"111111111",
  59704=>"111011000",
  59705=>"100100111",
  59706=>"100111111",
  59707=>"111111111",
  59708=>"000000000",
  59709=>"110110110",
  59710=>"001011111",
  59711=>"101001001",
  59712=>"000000000",
  59713=>"111111111",
  59714=>"111111111",
  59715=>"101111111",
  59716=>"000000000",
  59717=>"111001000",
  59718=>"000000000",
  59719=>"000000010",
  59720=>"000000000",
  59721=>"000111111",
  59722=>"000100100",
  59723=>"111101100",
  59724=>"111000100",
  59725=>"110011000",
  59726=>"000100111",
  59727=>"111111100",
  59728=>"100110110",
  59729=>"000000011",
  59730=>"111110000",
  59731=>"111111111",
  59732=>"111111111",
  59733=>"000010111",
  59734=>"111111000",
  59735=>"000000000",
  59736=>"111111001",
  59737=>"000000000",
  59738=>"111111000",
  59739=>"000000000",
  59740=>"111111111",
  59741=>"111111111",
  59742=>"001000000",
  59743=>"001000000",
  59744=>"000110010",
  59745=>"001101000",
  59746=>"010101111",
  59747=>"000000000",
  59748=>"111111111",
  59749=>"011111111",
  59750=>"100111000",
  59751=>"000100100",
  59752=>"111001001",
  59753=>"000011000",
  59754=>"111111111",
  59755=>"001111110",
  59756=>"000001001",
  59757=>"011011001",
  59758=>"000000000",
  59759=>"010111101",
  59760=>"000000101",
  59761=>"000000000",
  59762=>"110111000",
  59763=>"111111111",
  59764=>"111000000",
  59765=>"000101111",
  59766=>"011000000",
  59767=>"001001001",
  59768=>"000000000",
  59769=>"011111000",
  59770=>"010000000",
  59771=>"111111111",
  59772=>"111111000",
  59773=>"010110110",
  59774=>"111000000",
  59775=>"000111111",
  59776=>"001001001",
  59777=>"110110000",
  59778=>"101001011",
  59779=>"000000000",
  59780=>"000000000",
  59781=>"000000000",
  59782=>"111111000",
  59783=>"000000000",
  59784=>"011111101",
  59785=>"011011111",
  59786=>"000111111",
  59787=>"000000001",
  59788=>"000000000",
  59789=>"000000111",
  59790=>"100111111",
  59791=>"111111110",
  59792=>"000111111",
  59793=>"111111111",
  59794=>"011111111",
  59795=>"000100010",
  59796=>"000000000",
  59797=>"000000111",
  59798=>"010000100",
  59799=>"000000110",
  59800=>"000000000",
  59801=>"100000000",
  59802=>"111111110",
  59803=>"100100111",
  59804=>"100110111",
  59805=>"111111111",
  59806=>"101001001",
  59807=>"000000000",
  59808=>"000000000",
  59809=>"000000000",
  59810=>"000000111",
  59811=>"111111111",
  59812=>"101100110",
  59813=>"101101111",
  59814=>"100000000",
  59815=>"000011000",
  59816=>"000000000",
  59817=>"011111111",
  59818=>"111111110",
  59819=>"000000011",
  59820=>"111111000",
  59821=>"000000000",
  59822=>"000001001",
  59823=>"000000000",
  59824=>"000000111",
  59825=>"111111111",
  59826=>"111011101",
  59827=>"001111111",
  59828=>"001000000",
  59829=>"100111111",
  59830=>"000000000",
  59831=>"111110000",
  59832=>"110111000",
  59833=>"000000000",
  59834=>"111001001",
  59835=>"110111111",
  59836=>"110110111",
  59837=>"101000000",
  59838=>"111110110",
  59839=>"100000111",
  59840=>"000000000",
  59841=>"111110000",
  59842=>"111111111",
  59843=>"000000000",
  59844=>"111110110",
  59845=>"000000000",
  59846=>"000111111",
  59847=>"000111111",
  59848=>"111111111",
  59849=>"000100110",
  59850=>"000000001",
  59851=>"010111111",
  59852=>"111000111",
  59853=>"111111000",
  59854=>"111111100",
  59855=>"000100101",
  59856=>"111111011",
  59857=>"000000011",
  59858=>"000000011",
  59859=>"111111111",
  59860=>"111111111",
  59861=>"100100100",
  59862=>"011111111",
  59863=>"000001101",
  59864=>"111111111",
  59865=>"000001000",
  59866=>"011110000",
  59867=>"001000111",
  59868=>"000000000",
  59869=>"101111101",
  59870=>"111111111",
  59871=>"011111001",
  59872=>"000001000",
  59873=>"000000000",
  59874=>"000000000",
  59875=>"000110111",
  59876=>"101000110",
  59877=>"111111111",
  59878=>"111100000",
  59879=>"100000000",
  59880=>"111110110",
  59881=>"111111111",
  59882=>"000000000",
  59883=>"000000001",
  59884=>"100101100",
  59885=>"011001001",
  59886=>"000000000",
  59887=>"001110000",
  59888=>"000000000",
  59889=>"111111010",
  59890=>"000110110",
  59891=>"001001000",
  59892=>"100111111",
  59893=>"110000001",
  59894=>"001000111",
  59895=>"001001101",
  59896=>"000000100",
  59897=>"010011111",
  59898=>"111011100",
  59899=>"110100000",
  59900=>"111110111",
  59901=>"100101110",
  59902=>"001111111",
  59903=>"000000000",
  59904=>"101101100",
  59905=>"000110111",
  59906=>"111111111",
  59907=>"000000001",
  59908=>"000000000",
  59909=>"000000001",
  59910=>"101111111",
  59911=>"001001111",
  59912=>"000000111",
  59913=>"010010000",
  59914=>"000000000",
  59915=>"100000000",
  59916=>"010000000",
  59917=>"100111101",
  59918=>"111111001",
  59919=>"110100110",
  59920=>"110110110",
  59921=>"000110111",
  59922=>"100100000",
  59923=>"011111111",
  59924=>"101000000",
  59925=>"111000000",
  59926=>"000000110",
  59927=>"111001000",
  59928=>"110101111",
  59929=>"000000100",
  59930=>"000000000",
  59931=>"100001001",
  59932=>"001000000",
  59933=>"011000000",
  59934=>"000100011",
  59935=>"000000000",
  59936=>"111111101",
  59937=>"000111111",
  59938=>"111111001",
  59939=>"000000000",
  59940=>"000000111",
  59941=>"110111111",
  59942=>"001011001",
  59943=>"110111010",
  59944=>"111111000",
  59945=>"110100100",
  59946=>"001001000",
  59947=>"111110100",
  59948=>"000000000",
  59949=>"010100100",
  59950=>"000000100",
  59951=>"000101001",
  59952=>"110111000",
  59953=>"011111010",
  59954=>"000000000",
  59955=>"000100111",
  59956=>"001010010",
  59957=>"100101100",
  59958=>"000100000",
  59959=>"101100000",
  59960=>"000001111",
  59961=>"000111111",
  59962=>"111111111",
  59963=>"010011111",
  59964=>"000000000",
  59965=>"000110000",
  59966=>"011000000",
  59967=>"110110111",
  59968=>"100110111",
  59969=>"000011001",
  59970=>"001111111",
  59971=>"000111111",
  59972=>"101100101",
  59973=>"000000000",
  59974=>"000000000",
  59975=>"000000000",
  59976=>"111111111",
  59977=>"111001001",
  59978=>"011000001",
  59979=>"101001011",
  59980=>"001000001",
  59981=>"110110000",
  59982=>"111110000",
  59983=>"001000000",
  59984=>"001000001",
  59985=>"001000001",
  59986=>"000000111",
  59987=>"111111110",
  59988=>"110110110",
  59989=>"111000000",
  59990=>"111000000",
  59991=>"111001000",
  59992=>"011011010",
  59993=>"111001111",
  59994=>"011011000",
  59995=>"000110011",
  59996=>"111000011",
  59997=>"111111111",
  59998=>"001001001",
  59999=>"000111110",
  60000=>"111111111",
  60001=>"111111011",
  60002=>"001000001",
  60003=>"010010010",
  60004=>"000000000",
  60005=>"110111111",
  60006=>"000110111",
  60007=>"111111100",
  60008=>"000111111",
  60009=>"111111111",
  60010=>"100100111",
  60011=>"100011000",
  60012=>"000000000",
  60013=>"111111111",
  60014=>"000101111",
  60015=>"011111000",
  60016=>"011001111",
  60017=>"110011001",
  60018=>"011111010",
  60019=>"011011111",
  60020=>"111000000",
  60021=>"111100101",
  60022=>"111111111",
  60023=>"000000001",
  60024=>"000000000",
  60025=>"111000000",
  60026=>"011001000",
  60027=>"111111001",
  60028=>"100110100",
  60029=>"110111011",
  60030=>"001000000",
  60031=>"011010110",
  60032=>"011011111",
  60033=>"111000010",
  60034=>"111111111",
  60035=>"111110111",
  60036=>"000111111",
  60037=>"101001000",
  60038=>"001101111",
  60039=>"111111111",
  60040=>"000000011",
  60041=>"100000000",
  60042=>"000000111",
  60043=>"010110111",
  60044=>"111011011",
  60045=>"100000000",
  60046=>"111111011",
  60047=>"111111000",
  60048=>"001001011",
  60049=>"000000000",
  60050=>"100110110",
  60051=>"000111111",
  60052=>"111111111",
  60053=>"000100111",
  60054=>"011111111",
  60055=>"011000000",
  60056=>"000000000",
  60057=>"111111111",
  60058=>"100000000",
  60059=>"000000000",
  60060=>"111000000",
  60061=>"110001101",
  60062=>"000000000",
  60063=>"001101000",
  60064=>"111111111",
  60065=>"110110111",
  60066=>"010110110",
  60067=>"001001000",
  60068=>"110100100",
  60069=>"110110110",
  60070=>"111111111",
  60071=>"000011000",
  60072=>"101000000",
  60073=>"010010111",
  60074=>"011011000",
  60075=>"111111111",
  60076=>"000100000",
  60077=>"000000000",
  60078=>"110000000",
  60079=>"000000010",
  60080=>"111111000",
  60081=>"110010000",
  60082=>"000010010",
  60083=>"001001000",
  60084=>"100100011",
  60085=>"000110110",
  60086=>"000000011",
  60087=>"111110100",
  60088=>"000000000",
  60089=>"011000111",
  60090=>"011000000",
  60091=>"000000000",
  60092=>"111000001",
  60093=>"000001111",
  60094=>"110000000",
  60095=>"101111111",
  60096=>"111000000",
  60097=>"110111111",
  60098=>"000000001",
  60099=>"111111000",
  60100=>"111111111",
  60101=>"000111111",
  60102=>"011111001",
  60103=>"001000000",
  60104=>"000000111",
  60105=>"000000111",
  60106=>"111011001",
  60107=>"011011111",
  60108=>"110010000",
  60109=>"100100000",
  60110=>"110110010",
  60111=>"001001000",
  60112=>"111110110",
  60113=>"001001111",
  60114=>"010110111",
  60115=>"001111111",
  60116=>"000000000",
  60117=>"100100110",
  60118=>"001001001",
  60119=>"111000000",
  60120=>"110000000",
  60121=>"000001001",
  60122=>"111000000",
  60123=>"000000000",
  60124=>"000000000",
  60125=>"000000000",
  60126=>"000000001",
  60127=>"000000000",
  60128=>"010000010",
  60129=>"000000000",
  60130=>"111000000",
  60131=>"000100000",
  60132=>"011111100",
  60133=>"100110111",
  60134=>"111111011",
  60135=>"111111111",
  60136=>"000000011",
  60137=>"110011000",
  60138=>"100000000",
  60139=>"100010111",
  60140=>"111111100",
  60141=>"111101000",
  60142=>"000000001",
  60143=>"110000110",
  60144=>"111111000",
  60145=>"001000000",
  60146=>"000000011",
  60147=>"110110110",
  60148=>"111111111",
  60149=>"110111111",
  60150=>"111011011",
  60151=>"111111000",
  60152=>"111111001",
  60153=>"111111011",
  60154=>"000110110",
  60155=>"000000000",
  60156=>"111110110",
  60157=>"001001111",
  60158=>"110111000",
  60159=>"111111111",
  60160=>"111111111",
  60161=>"001001001",
  60162=>"000100111",
  60163=>"000000000",
  60164=>"000110100",
  60165=>"010000100",
  60166=>"001111001",
  60167=>"111111111",
  60168=>"000000000",
  60169=>"011011011",
  60170=>"101111011",
  60171=>"110111111",
  60172=>"110000100",
  60173=>"111100000",
  60174=>"111111111",
  60175=>"010111111",
  60176=>"111111110",
  60177=>"000010111",
  60178=>"111001111",
  60179=>"010000001",
  60180=>"111100100",
  60181=>"110000100",
  60182=>"000100111",
  60183=>"000000000",
  60184=>"110010000",
  60185=>"111011000",
  60186=>"111111000",
  60187=>"111100001",
  60188=>"001000000",
  60189=>"000000000",
  60190=>"111001001",
  60191=>"111110110",
  60192=>"111111011",
  60193=>"001000011",
  60194=>"111111111",
  60195=>"111111111",
  60196=>"001001000",
  60197=>"000000001",
  60198=>"111100000",
  60199=>"000000100",
  60200=>"000011001",
  60201=>"000000000",
  60202=>"000010000",
  60203=>"001000000",
  60204=>"000000000",
  60205=>"100001000",
  60206=>"101111111",
  60207=>"110110010",
  60208=>"110110110",
  60209=>"100100000",
  60210=>"111111101",
  60211=>"011111111",
  60212=>"000100110",
  60213=>"100110110",
  60214=>"000000000",
  60215=>"000000011",
  60216=>"000000000",
  60217=>"001111111",
  60218=>"001011000",
  60219=>"000000011",
  60220=>"000000001",
  60221=>"110111110",
  60222=>"011101110",
  60223=>"000110111",
  60224=>"001001001",
  60225=>"111111110",
  60226=>"111111011",
  60227=>"000000001",
  60228=>"111111111",
  60229=>"100100000",
  60230=>"110100000",
  60231=>"000000111",
  60232=>"000000000",
  60233=>"000000001",
  60234=>"111010000",
  60235=>"000111111",
  60236=>"111100110",
  60237=>"111111110",
  60238=>"100100111",
  60239=>"001111111",
  60240=>"000110110",
  60241=>"000000000",
  60242=>"000000000",
  60243=>"111111111",
  60244=>"111111111",
  60245=>"001011001",
  60246=>"111111110",
  60247=>"111111100",
  60248=>"100101111",
  60249=>"011010000",
  60250=>"000000000",
  60251=>"001000001",
  60252=>"000000000",
  60253=>"111111111",
  60254=>"100100100",
  60255=>"111111011",
  60256=>"111000000",
  60257=>"111101000",
  60258=>"000000000",
  60259=>"000000011",
  60260=>"000001111",
  60261=>"000000000",
  60262=>"000000000",
  60263=>"111111111",
  60264=>"100111011",
  60265=>"111111111",
  60266=>"111011010",
  60267=>"000000000",
  60268=>"110110110",
  60269=>"011000100",
  60270=>"111000001",
  60271=>"000010000",
  60272=>"000000111",
  60273=>"110010000",
  60274=>"111111001",
  60275=>"001111111",
  60276=>"000000000",
  60277=>"000111111",
  60278=>"111011011",
  60279=>"000000000",
  60280=>"000000000",
  60281=>"000011111",
  60282=>"111001001",
  60283=>"011000000",
  60284=>"110110110",
  60285=>"111000000",
  60286=>"111100110",
  60287=>"101000000",
  60288=>"110101100",
  60289=>"111011100",
  60290=>"000100101",
  60291=>"000000000",
  60292=>"000000000",
  60293=>"011111000",
  60294=>"100100000",
  60295=>"111000000",
  60296=>"111111111",
  60297=>"000100111",
  60298=>"000000000",
  60299=>"111011111",
  60300=>"000011011",
  60301=>"111111110",
  60302=>"111111111",
  60303=>"001011111",
  60304=>"000000000",
  60305=>"000000000",
  60306=>"110110110",
  60307=>"000000000",
  60308=>"100000000",
  60309=>"000000000",
  60310=>"111001001",
  60311=>"000000011",
  60312=>"111111111",
  60313=>"010110110",
  60314=>"000000000",
  60315=>"000001010",
  60316=>"000000010",
  60317=>"111111111",
  60318=>"000111001",
  60319=>"111110000",
  60320=>"000110110",
  60321=>"111011011",
  60322=>"111111011",
  60323=>"111001001",
  60324=>"111111110",
  60325=>"000000000",
  60326=>"000000111",
  60327=>"100000000",
  60328=>"111011111",
  60329=>"000000000",
  60330=>"000000000",
  60331=>"110110110",
  60332=>"000000000",
  60333=>"100010011",
  60334=>"000111111",
  60335=>"111111111",
  60336=>"110111111",
  60337=>"000000000",
  60338=>"001000001",
  60339=>"000000000",
  60340=>"111111111",
  60341=>"010000000",
  60342=>"000100100",
  60343=>"001001111",
  60344=>"000000010",
  60345=>"011011000",
  60346=>"000010000",
  60347=>"110111111",
  60348=>"000000110",
  60349=>"101000000",
  60350=>"100000110",
  60351=>"000100101",
  60352=>"100000111",
  60353=>"111111111",
  60354=>"011000111",
  60355=>"010000000",
  60356=>"000100100",
  60357=>"100100100",
  60358=>"000000010",
  60359=>"000111110",
  60360=>"100100111",
  60361=>"000111011",
  60362=>"011000011",
  60363=>"000001111",
  60364=>"000000100",
  60365=>"111001000",
  60366=>"111111100",
  60367=>"111111111",
  60368=>"000110110",
  60369=>"110111111",
  60370=>"111001000",
  60371=>"000000000",
  60372=>"111111000",
  60373=>"000000100",
  60374=>"000000000",
  60375=>"110100111",
  60376=>"001000111",
  60377=>"110111010",
  60378=>"110110111",
  60379=>"011111111",
  60380=>"001011111",
  60381=>"110111010",
  60382=>"111110111",
  60383=>"100000101",
  60384=>"100110110",
  60385=>"010000001",
  60386=>"000001000",
  60387=>"000000100",
  60388=>"000001111",
  60389=>"001101101",
  60390=>"000000001",
  60391=>"000000000",
  60392=>"000000001",
  60393=>"111111011",
  60394=>"100111111",
  60395=>"000000001",
  60396=>"001000011",
  60397=>"000000000",
  60398=>"111000011",
  60399=>"111011000",
  60400=>"000000000",
  60401=>"100100000",
  60402=>"110111111",
  60403=>"000000000",
  60404=>"001000100",
  60405=>"010000000",
  60406=>"110000000",
  60407=>"101101000",
  60408=>"111111110",
  60409=>"000010010",
  60410=>"000000000",
  60411=>"010000000",
  60412=>"000000010",
  60413=>"101111111",
  60414=>"000110111",
  60415=>"000000111",
  60416=>"111110111",
  60417=>"000010000",
  60418=>"111111000",
  60419=>"000000000",
  60420=>"110111011",
  60421=>"000000000",
  60422=>"000000000",
  60423=>"111111101",
  60424=>"111111110",
  60425=>"111011000",
  60426=>"010111111",
  60427=>"100010000",
  60428=>"100110110",
  60429=>"100100000",
  60430=>"001000000",
  60431=>"000001011",
  60432=>"000000000",
  60433=>"001000101",
  60434=>"000000000",
  60435=>"111010000",
  60436=>"110111000",
  60437=>"000000000",
  60438=>"000111111",
  60439=>"000001011",
  60440=>"111111111",
  60441=>"000100110",
  60442=>"100111111",
  60443=>"111011001",
  60444=>"000001001",
  60445=>"000000000",
  60446=>"001000000",
  60447=>"000000000",
  60448=>"011001001",
  60449=>"011001111",
  60450=>"000000000",
  60451=>"001001000",
  60452=>"111111111",
  60453=>"111001111",
  60454=>"111111111",
  60455=>"001000000",
  60456=>"111111111",
  60457=>"000110110",
  60458=>"100100111",
  60459=>"100110111",
  60460=>"010111111",
  60461=>"000000000",
  60462=>"001000101",
  60463=>"000000000",
  60464=>"111001001",
  60465=>"111111110",
  60466=>"111111110",
  60467=>"111001111",
  60468=>"111111111",
  60469=>"111111110",
  60470=>"001000000",
  60471=>"000000000",
  60472=>"000000000",
  60473=>"000000101",
  60474=>"000000111",
  60475=>"000111111",
  60476=>"000000011",
  60477=>"000100110",
  60478=>"000111111",
  60479=>"101000111",
  60480=>"000001011",
  60481=>"100100000",
  60482=>"001001001",
  60483=>"000101111",
  60484=>"110001001",
  60485=>"111000000",
  60486=>"111000001",
  60487=>"000000000",
  60488=>"111111011",
  60489=>"110010000",
  60490=>"111001000",
  60491=>"111111111",
  60492=>"011111000",
  60493=>"000100110",
  60494=>"111101101",
  60495=>"111111111",
  60496=>"000000000",
  60497=>"001100110",
  60498=>"111011000",
  60499=>"110111111",
  60500=>"000000000",
  60501=>"100110111",
  60502=>"111111100",
  60503=>"111111111",
  60504=>"100100111",
  60505=>"111111111",
  60506=>"000000000",
  60507=>"110100100",
  60508=>"111111111",
  60509=>"000000000",
  60510=>"010000100",
  60511=>"000000000",
  60512=>"000000000",
  60513=>"110100100",
  60514=>"111111111",
  60515=>"000000001",
  60516=>"111111111",
  60517=>"000000110",
  60518=>"000000000",
  60519=>"111111101",
  60520=>"111111111",
  60521=>"000000000",
  60522=>"100111111",
  60523=>"111111111",
  60524=>"111100100",
  60525=>"000000000",
  60526=>"000000000",
  60527=>"000010111",
  60528=>"000100000",
  60529=>"000001100",
  60530=>"000010000",
  60531=>"011010110",
  60532=>"000000000",
  60533=>"011111010",
  60534=>"000001000",
  60535=>"000111111",
  60536=>"011011010",
  60537=>"101111111",
  60538=>"111111011",
  60539=>"111000000",
  60540=>"001011111",
  60541=>"111111110",
  60542=>"101000000",
  60543=>"110110000",
  60544=>"110111111",
  60545=>"000000000",
  60546=>"111111111",
  60547=>"011000000",
  60548=>"111101100",
  60549=>"000000111",
  60550=>"000001000",
  60551=>"110111000",
  60552=>"100000000",
  60553=>"111000000",
  60554=>"000000000",
  60555=>"111111110",
  60556=>"000100110",
  60557=>"111111111",
  60558=>"111001101",
  60559=>"100001011",
  60560=>"001011001",
  60561=>"000000000",
  60562=>"000000000",
  60563=>"000111100",
  60564=>"000100111",
  60565=>"100000000",
  60566=>"111111111",
  60567=>"111000000",
  60568=>"000000000",
  60569=>"011100111",
  60570=>"111111000",
  60571=>"010010010",
  60572=>"000000111",
  60573=>"111111000",
  60574=>"010110111",
  60575=>"000001011",
  60576=>"110110110",
  60577=>"111111111",
  60578=>"111111111",
  60579=>"000000000",
  60580=>"011001011",
  60581=>"010100111",
  60582=>"000000000",
  60583=>"111111111",
  60584=>"111111000",
  60585=>"111000000",
  60586=>"111000000",
  60587=>"010000001",
  60588=>"111111011",
  60589=>"111111111",
  60590=>"111101111",
  60591=>"000111111",
  60592=>"000110111",
  60593=>"000001100",
  60594=>"000000010",
  60595=>"010011000",
  60596=>"001000000",
  60597=>"111011111",
  60598=>"000001101",
  60599=>"011111111",
  60600=>"111111111",
  60601=>"000000000",
  60602=>"000001011",
  60603=>"010010111",
  60604=>"111001111",
  60605=>"110111000",
  60606=>"010000101",
  60607=>"100110110",
  60608=>"000000000",
  60609=>"001000000",
  60610=>"011111111",
  60611=>"000000001",
  60612=>"010111011",
  60613=>"111001011",
  60614=>"100111111",
  60615=>"111111111",
  60616=>"111011111",
  60617=>"111000000",
  60618=>"000000000",
  60619=>"111111111",
  60620=>"000000101",
  60621=>"000000000",
  60622=>"111101111",
  60623=>"000000000",
  60624=>"111110111",
  60625=>"111111111",
  60626=>"111111111",
  60627=>"111111111",
  60628=>"000101111",
  60629=>"001001101",
  60630=>"000001000",
  60631=>"000000000",
  60632=>"111111111",
  60633=>"000000011",
  60634=>"010010011",
  60635=>"000011001",
  60636=>"111111111",
  60637=>"000000000",
  60638=>"111011011",
  60639=>"000001111",
  60640=>"000000000",
  60641=>"100000000",
  60642=>"111111111",
  60643=>"000000000",
  60644=>"000100000",
  60645=>"011001001",
  60646=>"111111111",
  60647=>"000000111",
  60648=>"000000000",
  60649=>"111111001",
  60650=>"000001000",
  60651=>"110110101",
  60652=>"111111111",
  60653=>"000000000",
  60654=>"001011111",
  60655=>"011001011",
  60656=>"100011001",
  60657=>"100000100",
  60658=>"000111001",
  60659=>"000000110",
  60660=>"111001111",
  60661=>"000001000",
  60662=>"111011111",
  60663=>"111111111",
  60664=>"001101111",
  60665=>"111111111",
  60666=>"000000000",
  60667=>"111111111",
  60668=>"111110110",
  60669=>"000000000",
  60670=>"000001011",
  60671=>"001001111",
  60672=>"111011000",
  60673=>"001001001",
  60674=>"000000000",
  60675=>"000000000",
  60676=>"111101100",
  60677=>"100110111",
  60678=>"001001101",
  60679=>"111000000",
  60680=>"111111111",
  60681=>"111111100",
  60682=>"111111111",
  60683=>"011101110",
  60684=>"000000001",
  60685=>"110100101",
  60686=>"111000011",
  60687=>"111111010",
  60688=>"110110000",
  60689=>"000011111",
  60690=>"111111000",
  60691=>"010110000",
  60692=>"110000000",
  60693=>"000000000",
  60694=>"110110111",
  60695=>"011010110",
  60696=>"111111111",
  60697=>"111111111",
  60698=>"001001001",
  60699=>"000000111",
  60700=>"001000011",
  60701=>"000000000",
  60702=>"110111111",
  60703=>"010010101",
  60704=>"001110111",
  60705=>"000000000",
  60706=>"001111111",
  60707=>"000000000",
  60708=>"000000001",
  60709=>"000000000",
  60710=>"111111111",
  60711=>"111111111",
  60712=>"000000000",
  60713=>"111111111",
  60714=>"111101111",
  60715=>"000100111",
  60716=>"100111111",
  60717=>"000001001",
  60718=>"000000000",
  60719=>"001001111",
  60720=>"010000110",
  60721=>"000000000",
  60722=>"000000000",
  60723=>"111111000",
  60724=>"001111111",
  60725=>"111111111",
  60726=>"111111111",
  60727=>"000011001",
  60728=>"111110100",
  60729=>"000000000",
  60730=>"011000011",
  60731=>"111111111",
  60732=>"111111111",
  60733=>"000000000",
  60734=>"000000000",
  60735=>"000000010",
  60736=>"000001111",
  60737=>"111011000",
  60738=>"010000000",
  60739=>"111000000",
  60740=>"000000000",
  60741=>"111111111",
  60742=>"101100100",
  60743=>"111111111",
  60744=>"111111111",
  60745=>"111111111",
  60746=>"000000001",
  60747=>"000000111",
  60748=>"000001001",
  60749=>"000000000",
  60750=>"011001001",
  60751=>"100000111",
  60752=>"000000100",
  60753=>"110101101",
  60754=>"111111111",
  60755=>"011111001",
  60756=>"111000000",
  60757=>"000000010",
  60758=>"111000000",
  60759=>"001011111",
  60760=>"111001111",
  60761=>"111111000",
  60762=>"111111111",
  60763=>"111010010",
  60764=>"000000000",
  60765=>"000000011",
  60766=>"001101111",
  60767=>"011011011",
  60768=>"110010000",
  60769=>"111000000",
  60770=>"011100110",
  60771=>"000000000",
  60772=>"111111111",
  60773=>"001000001",
  60774=>"111001100",
  60775=>"000000000",
  60776=>"000001001",
  60777=>"000000000",
  60778=>"111111000",
  60779=>"000000000",
  60780=>"000000000",
  60781=>"111111011",
  60782=>"000000000",
  60783=>"011001000",
  60784=>"000000000",
  60785=>"000000000",
  60786=>"111010000",
  60787=>"111111111",
  60788=>"111110111",
  60789=>"111111011",
  60790=>"001001000",
  60791=>"000000000",
  60792=>"000111111",
  60793=>"111111000",
  60794=>"000000111",
  60795=>"111111111",
  60796=>"000000000",
  60797=>"010010000",
  60798=>"011011011",
  60799=>"111111111",
  60800=>"001011011",
  60801=>"011001000",
  60802=>"000111111",
  60803=>"000000000",
  60804=>"000000110",
  60805=>"110010000",
  60806=>"110000001",
  60807=>"001000000",
  60808=>"000000000",
  60809=>"010010011",
  60810=>"011011111",
  60811=>"111111111",
  60812=>"111111111",
  60813=>"000000111",
  60814=>"110010111",
  60815=>"111111111",
  60816=>"001001000",
  60817=>"000111111",
  60818=>"000000100",
  60819=>"001001001",
  60820=>"000000000",
  60821=>"000000000",
  60822=>"111111001",
  60823=>"000000110",
  60824=>"000000000",
  60825=>"000000000",
  60826=>"000000000",
  60827=>"000100000",
  60828=>"111111100",
  60829=>"000000001",
  60830=>"011011011",
  60831=>"111100100",
  60832=>"000000000",
  60833=>"111111100",
  60834=>"111000000",
  60835=>"011000010",
  60836=>"000000000",
  60837=>"111111111",
  60838=>"001000000",
  60839=>"000000000",
  60840=>"111111000",
  60841=>"110000000",
  60842=>"000010000",
  60843=>"110100111",
  60844=>"000010000",
  60845=>"011010011",
  60846=>"111000100",
  60847=>"000000000",
  60848=>"000011111",
  60849=>"000000000",
  60850=>"111011111",
  60851=>"111111111",
  60852=>"000001100",
  60853=>"000000000",
  60854=>"011111111",
  60855=>"111111111",
  60856=>"000011111",
  60857=>"000100000",
  60858=>"000100000",
  60859=>"100100000",
  60860=>"000000001",
  60861=>"100111111",
  60862=>"111111111",
  60863=>"001001000",
  60864=>"111111110",
  60865=>"111111111",
  60866=>"000011011",
  60867=>"111111111",
  60868=>"000000000",
  60869=>"111101000",
  60870=>"011100100",
  60871=>"000000000",
  60872=>"000000000",
  60873=>"001000000",
  60874=>"001000000",
  60875=>"010000000",
  60876=>"000111111",
  60877=>"111000000",
  60878=>"110110100",
  60879=>"000000000",
  60880=>"111001001",
  60881=>"011001001",
  60882=>"000000000",
  60883=>"000000011",
  60884=>"111111110",
  60885=>"101100001",
  60886=>"001000000",
  60887=>"101110100",
  60888=>"000000000",
  60889=>"000000011",
  60890=>"000000000",
  60891=>"001101111",
  60892=>"000000000",
  60893=>"000000100",
  60894=>"111111100",
  60895=>"001001011",
  60896=>"000000000",
  60897=>"000011011",
  60898=>"000000000",
  60899=>"111111000",
  60900=>"000001011",
  60901=>"110100100",
  60902=>"000101001",
  60903=>"000000000",
  60904=>"010000001",
  60905=>"000101101",
  60906=>"011100110",
  60907=>"111111011",
  60908=>"110111111",
  60909=>"111111111",
  60910=>"000001000",
  60911=>"000000111",
  60912=>"011011111",
  60913=>"000000000",
  60914=>"111000000",
  60915=>"000111011",
  60916=>"111111111",
  60917=>"100100000",
  60918=>"001000110",
  60919=>"110000011",
  60920=>"000000000",
  60921=>"001001001",
  60922=>"111100110",
  60923=>"111000000",
  60924=>"000001001",
  60925=>"111111111",
  60926=>"000000000",
  60927=>"000100110",
  60928=>"000000000",
  60929=>"111000111",
  60930=>"110000000",
  60931=>"111111000",
  60932=>"111111010",
  60933=>"111110110",
  60934=>"111111111",
  60935=>"111101111",
  60936=>"110110010",
  60937=>"110111111",
  60938=>"111110010",
  60939=>"111000010",
  60940=>"100110100",
  60941=>"111100100",
  60942=>"111111111",
  60943=>"000110110",
  60944=>"111111110",
  60945=>"100110110",
  60946=>"010111110",
  60947=>"011000000",
  60948=>"000000000",
  60949=>"111011111",
  60950=>"000000000",
  60951=>"001011111",
  60952=>"111100101",
  60953=>"110110110",
  60954=>"011010010",
  60955=>"100100100",
  60956=>"101000001",
  60957=>"000000011",
  60958=>"111111111",
  60959=>"000011011",
  60960=>"111111111",
  60961=>"000000101",
  60962=>"110110110",
  60963=>"010000000",
  60964=>"101111111",
  60965=>"111111111",
  60966=>"111010001",
  60967=>"111110010",
  60968=>"001000100",
  60969=>"000000000",
  60970=>"010000000",
  60971=>"001000111",
  60972=>"000000000",
  60973=>"111111010",
  60974=>"111111110",
  60975=>"001000001",
  60976=>"110000000",
  60977=>"010010000",
  60978=>"111111110",
  60979=>"111000000",
  60980=>"110110110",
  60981=>"100111111",
  60982=>"110000000",
  60983=>"001110110",
  60984=>"100110110",
  60985=>"000000101",
  60986=>"000110111",
  60987=>"111111111",
  60988=>"100100100",
  60989=>"100110111",
  60990=>"011000100",
  60991=>"000000000",
  60992=>"110110110",
  60993=>"000011000",
  60994=>"000000010",
  60995=>"010010111",
  60996=>"110110100",
  60997=>"001000100",
  60998=>"111111000",
  60999=>"101001000",
  61000=>"111111001",
  61001=>"000001111",
  61002=>"011111111",
  61003=>"001001111",
  61004=>"000000110",
  61005=>"000000110",
  61006=>"011000101",
  61007=>"111111111",
  61008=>"111111110",
  61009=>"111111111",
  61010=>"011111111",
  61011=>"001100100",
  61012=>"100000000",
  61013=>"111110000",
  61014=>"000000100",
  61015=>"101001001",
  61016=>"000100000",
  61017=>"101101101",
  61018=>"000000110",
  61019=>"110010000",
  61020=>"111000000",
  61021=>"111001101",
  61022=>"011011001",
  61023=>"001001000",
  61024=>"000000100",
  61025=>"000010010",
  61026=>"000000000",
  61027=>"110111000",
  61028=>"100100111",
  61029=>"111110000",
  61030=>"110111011",
  61031=>"111111111",
  61032=>"010000011",
  61033=>"111000111",
  61034=>"111110000",
  61035=>"000011011",
  61036=>"001101100",
  61037=>"110111111",
  61038=>"111111001",
  61039=>"000011011",
  61040=>"010111110",
  61041=>"110100110",
  61042=>"001010000",
  61043=>"001101100",
  61044=>"001001000",
  61045=>"000110100",
  61046=>"000000111",
  61047=>"010111110",
  61048=>"110010011",
  61049=>"111111111",
  61050=>"001000000",
  61051=>"000000001",
  61052=>"101101101",
  61053=>"111111000",
  61054=>"000100100",
  61055=>"010000000",
  61056=>"111000000",
  61057=>"000001111",
  61058=>"000001111",
  61059=>"111111000",
  61060=>"111111111",
  61061=>"111101111",
  61062=>"101101110",
  61063=>"000000000",
  61064=>"010000000",
  61065=>"000101011",
  61066=>"111111111",
  61067=>"111110000",
  61068=>"110111110",
  61069=>"000000000",
  61070=>"001000111",
  61071=>"000110110",
  61072=>"101000101",
  61073=>"111000000",
  61074=>"000000000",
  61075=>"111100100",
  61076=>"010010011",
  61077=>"101101111",
  61078=>"001000101",
  61079=>"000000100",
  61080=>"111001101",
  61081=>"000000101",
  61082=>"010000000",
  61083=>"000000000",
  61084=>"001101111",
  61085=>"111101111",
  61086=>"111111001",
  61087=>"000000011",
  61088=>"011111111",
  61089=>"011110111",
  61090=>"111110100",
  61091=>"111111111",
  61092=>"100100000",
  61093=>"000101001",
  61094=>"011000000",
  61095=>"111111101",
  61096=>"110000001",
  61097=>"000000001",
  61098=>"000001101",
  61099=>"101100101",
  61100=>"000000000",
  61101=>"000001101",
  61102=>"000000000",
  61103=>"111111111",
  61104=>"010000000",
  61105=>"000000001",
  61106=>"111111010",
  61107=>"111101111",
  61108=>"111011000",
  61109=>"111011111",
  61110=>"000000100",
  61111=>"110110000",
  61112=>"000000101",
  61113=>"111111010",
  61114=>"111101101",
  61115=>"010011000",
  61116=>"111111011",
  61117=>"110110110",
  61118=>"010000000",
  61119=>"001000101",
  61120=>"011111011",
  61121=>"111111111",
  61122=>"010110111",
  61123=>"000011011",
  61124=>"111101001",
  61125=>"010000000",
  61126=>"110010000",
  61127=>"111111110",
  61128=>"000000011",
  61129=>"001000101",
  61130=>"000100111",
  61131=>"111111111",
  61132=>"001110110",
  61133=>"000100111",
  61134=>"000000111",
  61135=>"011111111",
  61136=>"111111111",
  61137=>"111111111",
  61138=>"100111111",
  61139=>"101000001",
  61140=>"000110010",
  61141=>"001101110",
  61142=>"111111111",
  61143=>"111011011",
  61144=>"010000111",
  61145=>"110111110",
  61146=>"010010010",
  61147=>"010010111",
  61148=>"000000000",
  61149=>"001010010",
  61150=>"110100000",
  61151=>"000101111",
  61152=>"000100010",
  61153=>"110110010",
  61154=>"111111111",
  61155=>"000000101",
  61156=>"001000101",
  61157=>"111110011",
  61158=>"011011001",
  61159=>"000000101",
  61160=>"000000001",
  61161=>"000000000",
  61162=>"110110110",
  61163=>"111111111",
  61164=>"100111110",
  61165=>"111111011",
  61166=>"000000101",
  61167=>"111111000",
  61168=>"001111111",
  61169=>"011001101",
  61170=>"001000000",
  61171=>"111100110",
  61172=>"000110111",
  61173=>"111111011",
  61174=>"000111111",
  61175=>"111111111",
  61176=>"110110010",
  61177=>"100010000",
  61178=>"000000101",
  61179=>"111110110",
  61180=>"000011010",
  61181=>"111111111",
  61182=>"111011010",
  61183=>"000000101",
  61184=>"111110000",
  61185=>"111101100",
  61186=>"111111001",
  61187=>"111111100",
  61188=>"111111000",
  61189=>"000100101",
  61190=>"011000000",
  61191=>"001000111",
  61192=>"001000100",
  61193=>"000000000",
  61194=>"000000011",
  61195=>"110110110",
  61196=>"100000000",
  61197=>"111001000",
  61198=>"000000000",
  61199=>"111111111",
  61200=>"001001001",
  61201=>"000010111",
  61202=>"111111111",
  61203=>"110100111",
  61204=>"000000001",
  61205=>"000111111",
  61206=>"011111110",
  61207=>"101000000",
  61208=>"000000001",
  61209=>"111111101",
  61210=>"101101111",
  61211=>"000000000",
  61212=>"110110110",
  61213=>"100000000",
  61214=>"000000111",
  61215=>"111010100",
  61216=>"001000111",
  61217=>"110000000",
  61218=>"000000111",
  61219=>"111111110",
  61220=>"100111110",
  61221=>"010101110",
  61222=>"000111000",
  61223=>"000000011",
  61224=>"010010111",
  61225=>"000000000",
  61226=>"011110110",
  61227=>"000000000",
  61228=>"000001111",
  61229=>"000000000",
  61230=>"101000000",
  61231=>"000000000",
  61232=>"001001101",
  61233=>"100000000",
  61234=>"000001101",
  61235=>"111111011",
  61236=>"000110100",
  61237=>"110010000",
  61238=>"111111001",
  61239=>"100000100",
  61240=>"111111111",
  61241=>"111000000",
  61242=>"101000001",
  61243=>"111011000",
  61244=>"001100101",
  61245=>"001100111",
  61246=>"001001001",
  61247=>"110100100",
  61248=>"000100000",
  61249=>"111000000",
  61250=>"101001101",
  61251=>"001001111",
  61252=>"110110010",
  61253=>"111100011",
  61254=>"000001001",
  61255=>"001011111",
  61256=>"111001111",
  61257=>"110111011",
  61258=>"011000111",
  61259=>"100000101",
  61260=>"010111111",
  61261=>"000100000",
  61262=>"110000110",
  61263=>"000000001",
  61264=>"000000001",
  61265=>"011011011",
  61266=>"000000000",
  61267=>"111011010",
  61268=>"111011000",
  61269=>"001011001",
  61270=>"101001111",
  61271=>"100110111",
  61272=>"111111111",
  61273=>"001001000",
  61274=>"000100000",
  61275=>"111101001",
  61276=>"000000000",
  61277=>"100111111",
  61278=>"111111111",
  61279=>"111010001",
  61280=>"011111111",
  61281=>"111110000",
  61282=>"100001001",
  61283=>"101111011",
  61284=>"000001001",
  61285=>"101000000",
  61286=>"011111111",
  61287=>"000000101",
  61288=>"111011001",
  61289=>"011011111",
  61290=>"111000000",
  61291=>"110110110",
  61292=>"111111111",
  61293=>"111111000",
  61294=>"000010010",
  61295=>"000000000",
  61296=>"101000000",
  61297=>"111011101",
  61298=>"100000001",
  61299=>"011111001",
  61300=>"000000111",
  61301=>"111111111",
  61302=>"000000100",
  61303=>"111111010",
  61304=>"000001101",
  61305=>"000000010",
  61306=>"101011111",
  61307=>"000000101",
  61308=>"001101100",
  61309=>"001011111",
  61310=>"111011111",
  61311=>"010001000",
  61312=>"110110100",
  61313=>"000100110",
  61314=>"000000000",
  61315=>"111000000",
  61316=>"111000000",
  61317=>"000000010",
  61318=>"011101011",
  61319=>"010010110",
  61320=>"100110110",
  61321=>"011011011",
  61322=>"000000000",
  61323=>"111011011",
  61324=>"000001000",
  61325=>"101110111",
  61326=>"111111110",
  61327=>"000000000",
  61328=>"100110110",
  61329=>"000001000",
  61330=>"010110111",
  61331=>"000000000",
  61332=>"000000110",
  61333=>"000010011",
  61334=>"001000100",
  61335=>"000001111",
  61336=>"000000110",
  61337=>"000000000",
  61338=>"110110000",
  61339=>"000000010",
  61340=>"011111111",
  61341=>"000000000",
  61342=>"111011001",
  61343=>"010000000",
  61344=>"000000101",
  61345=>"010000101",
  61346=>"011011111",
  61347=>"000000001",
  61348=>"111111111",
  61349=>"000010010",
  61350=>"000000000",
  61351=>"111000000",
  61352=>"110111101",
  61353=>"000000001",
  61354=>"111111000",
  61355=>"111000000",
  61356=>"000000000",
  61357=>"111111111",
  61358=>"001000000",
  61359=>"111001101",
  61360=>"000000000",
  61361=>"101000000",
  61362=>"111110111",
  61363=>"001000000",
  61364=>"111111111",
  61365=>"011111111",
  61366=>"111100100",
  61367=>"100000001",
  61368=>"000000000",
  61369=>"111001000",
  61370=>"000100000",
  61371=>"100100100",
  61372=>"111111110",
  61373=>"010000000",
  61374=>"110110110",
  61375=>"100101101",
  61376=>"010010000",
  61377=>"111011110",
  61378=>"000111111",
  61379=>"011011111",
  61380=>"000000000",
  61381=>"000000111",
  61382=>"000000010",
  61383=>"100110110",
  61384=>"111000000",
  61385=>"000111011",
  61386=>"111101111",
  61387=>"010010111",
  61388=>"110110111",
  61389=>"011011111",
  61390=>"110100110",
  61391=>"001001111",
  61392=>"010110100",
  61393=>"000000000",
  61394=>"010000000",
  61395=>"110010000",
  61396=>"111011001",
  61397=>"000000111",
  61398=>"010000000",
  61399=>"011111110",
  61400=>"011101001",
  61401=>"001000000",
  61402=>"111111000",
  61403=>"111111010",
  61404=>"000111111",
  61405=>"111111101",
  61406=>"111011001",
  61407=>"110000000",
  61408=>"000011111",
  61409=>"001000101",
  61410=>"010000000",
  61411=>"001001101",
  61412=>"111011001",
  61413=>"110010111",
  61414=>"000000100",
  61415=>"001000001",
  61416=>"100100100",
  61417=>"111111010",
  61418=>"000000000",
  61419=>"111110110",
  61420=>"000000111",
  61421=>"001000000",
  61422=>"111110111",
  61423=>"110000000",
  61424=>"111111101",
  61425=>"000000000",
  61426=>"111000000",
  61427=>"111000000",
  61428=>"111001000",
  61429=>"111001001",
  61430=>"001000000",
  61431=>"000000001",
  61432=>"010000000",
  61433=>"000100100",
  61434=>"000000000",
  61435=>"001001101",
  61436=>"110110111",
  61437=>"110000000",
  61438=>"011010000",
  61439=>"000000000",
  61440=>"111111011",
  61441=>"000100000",
  61442=>"101000001",
  61443=>"111111111",
  61444=>"000000001",
  61445=>"111111100",
  61446=>"011111010",
  61447=>"001000000",
  61448=>"110010111",
  61449=>"110110110",
  61450=>"110111111",
  61451=>"100100100",
  61452=>"110110110",
  61453=>"011101111",
  61454=>"110100110",
  61455=>"001001001",
  61456=>"000000000",
  61457=>"000000101",
  61458=>"111111111",
  61459=>"000000000",
  61460=>"111111001",
  61461=>"001001101",
  61462=>"111101101",
  61463=>"011001000",
  61464=>"100100100",
  61465=>"111101101",
  61466=>"110000111",
  61467=>"100100100",
  61468=>"111101001",
  61469=>"000000000",
  61470=>"011011110",
  61471=>"101101000",
  61472=>"001000000",
  61473=>"011000000",
  61474=>"111111110",
  61475=>"000010010",
  61476=>"111111001",
  61477=>"000001001",
  61478=>"000000001",
  61479=>"010000101",
  61480=>"000000000",
  61481=>"100100000",
  61482=>"111100000",
  61483=>"110010010",
  61484=>"111111111",
  61485=>"111111010",
  61486=>"000000100",
  61487=>"000000000",
  61488=>"000000100",
  61489=>"101001101",
  61490=>"000010011",
  61491=>"000000000",
  61492=>"000001011",
  61493=>"100000100",
  61494=>"000000001",
  61495=>"000110110",
  61496=>"000000000",
  61497=>"100000111",
  61498=>"000010011",
  61499=>"000010001",
  61500=>"001001001",
  61501=>"000110000",
  61502=>"100100000",
  61503=>"111100000",
  61504=>"010111111",
  61505=>"111111110",
  61506=>"110111111",
  61507=>"000000000",
  61508=>"000000001",
  61509=>"001000000",
  61510=>"110010000",
  61511=>"000000000",
  61512=>"111111011",
  61513=>"000111111",
  61514=>"000010110",
  61515=>"000100001",
  61516=>"111110000",
  61517=>"000000000",
  61518=>"000000000",
  61519=>"110110110",
  61520=>"110111100",
  61521=>"000011000",
  61522=>"000000101",
  61523=>"110110100",
  61524=>"001000000",
  61525=>"000000100",
  61526=>"100000000",
  61527=>"110000000",
  61528=>"111111011",
  61529=>"111101111",
  61530=>"000000110",
  61531=>"100100100",
  61532=>"110100101",
  61533=>"000000001",
  61534=>"000000000",
  61535=>"111111000",
  61536=>"001000000",
  61537=>"000000000",
  61538=>"100100101",
  61539=>"110100000",
  61540=>"111111110",
  61541=>"101000000",
  61542=>"111010000",
  61543=>"000111011",
  61544=>"011111000",
  61545=>"000001101",
  61546=>"000000111",
  61547=>"000000000",
  61548=>"011010000",
  61549=>"000000000",
  61550=>"000000001",
  61551=>"010110110",
  61552=>"000000110",
  61553=>"111110110",
  61554=>"100110111",
  61555=>"011111000",
  61556=>"000000000",
  61557=>"000100111",
  61558=>"000010111",
  61559=>"111101111",
  61560=>"001101111",
  61561=>"110011001",
  61562=>"111010000",
  61563=>"001000000",
  61564=>"110111100",
  61565=>"111111110",
  61566=>"111111110",
  61567=>"000001001",
  61568=>"000000101",
  61569=>"000000000",
  61570=>"010110000",
  61571=>"001001001",
  61572=>"000100101",
  61573=>"001001001",
  61574=>"110100000",
  61575=>"110100000",
  61576=>"000010110",
  61577=>"110111111",
  61578=>"111111000",
  61579=>"000000000",
  61580=>"000000000",
  61581=>"010010010",
  61582=>"000000111",
  61583=>"111111111",
  61584=>"000000000",
  61585=>"100000000",
  61586=>"000000000",
  61587=>"111111110",
  61588=>"001011000",
  61589=>"100111111",
  61590=>"000010010",
  61591=>"011011011",
  61592=>"001000000",
  61593=>"010011011",
  61594=>"111111111",
  61595=>"100000000",
  61596=>"100100001",
  61597=>"001001001",
  61598=>"001000100",
  61599=>"010111111",
  61600=>"011011001",
  61601=>"000111111",
  61602=>"010011010",
  61603=>"111111111",
  61604=>"111001000",
  61605=>"011011011",
  61606=>"111101111",
  61607=>"000100111",
  61608=>"111111110",
  61609=>"101101101",
  61610=>"111000000",
  61611=>"011000000",
  61612=>"111111101",
  61613=>"111111001",
  61614=>"000000000",
  61615=>"111111110",
  61616=>"111011001",
  61617=>"010110111",
  61618=>"001001011",
  61619=>"010000000",
  61620=>"101110110",
  61621=>"100000000",
  61622=>"111101101",
  61623=>"110110110",
  61624=>"000000000",
  61625=>"000000001",
  61626=>"100000000",
  61627=>"110110010",
  61628=>"111111010",
  61629=>"000110010",
  61630=>"011010000",
  61631=>"000000000",
  61632=>"000000001",
  61633=>"001000000",
  61634=>"000000001",
  61635=>"110110110",
  61636=>"111111010",
  61637=>"000000011",
  61638=>"001000000",
  61639=>"100001001",
  61640=>"001011111",
  61641=>"000000000",
  61642=>"100110100",
  61643=>"000000000",
  61644=>"110111111",
  61645=>"011011011",
  61646=>"000000001",
  61647=>"111011001",
  61648=>"010111111",
  61649=>"001001000",
  61650=>"110100000",
  61651=>"111111011",
  61652=>"110100001",
  61653=>"000000111",
  61654=>"101000000",
  61655=>"111111111",
  61656=>"000000001",
  61657=>"000000000",
  61658=>"000000000",
  61659=>"101111111",
  61660=>"111111111",
  61661=>"111111111",
  61662=>"000000000",
  61663=>"111000000",
  61664=>"000000000",
  61665=>"000010010",
  61666=>"010110110",
  61667=>"111011000",
  61668=>"010111111",
  61669=>"001000000",
  61670=>"000000000",
  61671=>"000000000",
  61672=>"111111010",
  61673=>"011001000",
  61674=>"000000000",
  61675=>"000000000",
  61676=>"001001001",
  61677=>"111110010",
  61678=>"111111111",
  61679=>"001111111",
  61680=>"000100111",
  61681=>"111111111",
  61682=>"110111111",
  61683=>"000101001",
  61684=>"000100000",
  61685=>"011001000",
  61686=>"000100000",
  61687=>"000000010",
  61688=>"010110110",
  61689=>"001001001",
  61690=>"001000001",
  61691=>"000000000",
  61692=>"001000000",
  61693=>"110110110",
  61694=>"111111000",
  61695=>"000011111",
  61696=>"110000000",
  61697=>"111111101",
  61698=>"000001011",
  61699=>"111111110",
  61700=>"000010111",
  61701=>"000000110",
  61702=>"000000000",
  61703=>"110000111",
  61704=>"000000000",
  61705=>"000000111",
  61706=>"000100000",
  61707=>"000111111",
  61708=>"000000001",
  61709=>"001111000",
  61710=>"011011011",
  61711=>"000000000",
  61712=>"000000000",
  61713=>"000001001",
  61714=>"111111111",
  61715=>"000111111",
  61716=>"100000000",
  61717=>"100100100",
  61718=>"110110110",
  61719=>"000000001",
  61720=>"011001001",
  61721=>"001000111",
  61722=>"111111010",
  61723=>"011000001",
  61724=>"110110110",
  61725=>"101000100",
  61726=>"110111111",
  61727=>"000001000",
  61728=>"111111000",
  61729=>"000000000",
  61730=>"000000000",
  61731=>"001000000",
  61732=>"111100110",
  61733=>"110110000",
  61734=>"110111011",
  61735=>"110100000",
  61736=>"000000000",
  61737=>"001000000",
  61738=>"000001000",
  61739=>"000000000",
  61740=>"010110000",
  61741=>"000000000",
  61742=>"100011000",
  61743=>"000000101",
  61744=>"000000001",
  61745=>"000000000",
  61746=>"000000001",
  61747=>"000000000",
  61748=>"111111111",
  61749=>"111111111",
  61750=>"000000011",
  61751=>"000000000",
  61752=>"000001011",
  61753=>"100000111",
  61754=>"111111111",
  61755=>"110110111",
  61756=>"100110100",
  61757=>"111111001",
  61758=>"100111011",
  61759=>"000100100",
  61760=>"111111111",
  61761=>"000000000",
  61762=>"111000000",
  61763=>"001011011",
  61764=>"000000000",
  61765=>"111111000",
  61766=>"111001011",
  61767=>"000100111",
  61768=>"111111110",
  61769=>"110110000",
  61770=>"001111001",
  61771=>"111111100",
  61772=>"100101001",
  61773=>"010110110",
  61774=>"000000000",
  61775=>"000101101",
  61776=>"101100100",
  61777=>"000000000",
  61778=>"100001000",
  61779=>"000000001",
  61780=>"001111011",
  61781=>"011011011",
  61782=>"111111000",
  61783=>"111111111",
  61784=>"111101111",
  61785=>"100010010",
  61786=>"001101111",
  61787=>"000000000",
  61788=>"110110110",
  61789=>"111111110",
  61790=>"001001000",
  61791=>"111110000",
  61792=>"110111101",
  61793=>"111111111",
  61794=>"100110000",
  61795=>"001000000",
  61796=>"111111111",
  61797=>"000111111",
  61798=>"000111111",
  61799=>"010010000",
  61800=>"111111111",
  61801=>"010111111",
  61802=>"011011001",
  61803=>"111110110",
  61804=>"001001001",
  61805=>"110100111",
  61806=>"000000000",
  61807=>"000011011",
  61808=>"000000000",
  61809=>"000000000",
  61810=>"101000000",
  61811=>"101101101",
  61812=>"111111111",
  61813=>"000000100",
  61814=>"000100111",
  61815=>"000000000",
  61816=>"011011011",
  61817=>"000111111",
  61818=>"111111111",
  61819=>"111111111",
  61820=>"111100000",
  61821=>"000000000",
  61822=>"000000011",
  61823=>"000000000",
  61824=>"111111111",
  61825=>"000001011",
  61826=>"000000000",
  61827=>"111111000",
  61828=>"111111111",
  61829=>"010010010",
  61830=>"000011111",
  61831=>"100001111",
  61832=>"011011111",
  61833=>"111110110",
  61834=>"000000000",
  61835=>"000000000",
  61836=>"110101001",
  61837=>"100100101",
  61838=>"010010000",
  61839=>"000000000",
  61840=>"110111111",
  61841=>"111111111",
  61842=>"111111111",
  61843=>"100100100",
  61844=>"111011111",
  61845=>"000011011",
  61846=>"000000000",
  61847=>"000010000",
  61848=>"000000000",
  61849=>"000111111",
  61850=>"000000001",
  61851=>"001001001",
  61852=>"000001001",
  61853=>"110111011",
  61854=>"101000011",
  61855=>"000100000",
  61856=>"001000001",
  61857=>"000010010",
  61858=>"111111000",
  61859=>"000110111",
  61860=>"111111000",
  61861=>"111111111",
  61862=>"000000001",
  61863=>"000111010",
  61864=>"110111110",
  61865=>"000000100",
  61866=>"111100100",
  61867=>"111001001",
  61868=>"101111101",
  61869=>"101000000",
  61870=>"011010001",
  61871=>"100000100",
  61872=>"000000111",
  61873=>"000000001",
  61874=>"001000001",
  61875=>"001111101",
  61876=>"000101111",
  61877=>"111111110",
  61878=>"111111110",
  61879=>"110110010",
  61880=>"110110111",
  61881=>"000000000",
  61882=>"011000000",
  61883=>"101111000",
  61884=>"110110110",
  61885=>"000011001",
  61886=>"001111000",
  61887=>"100001000",
  61888=>"111111010",
  61889=>"001000111",
  61890=>"000010000",
  61891=>"111111111",
  61892=>"110100010",
  61893=>"111111111",
  61894=>"000000000",
  61895=>"010110111",
  61896=>"100000000",
  61897=>"000100101",
  61898=>"001001000",
  61899=>"001001000",
  61900=>"000000000",
  61901=>"000000001",
  61902=>"000000001",
  61903=>"000000000",
  61904=>"001111000",
  61905=>"100000000",
  61906=>"000000000",
  61907=>"000100111",
  61908=>"111111100",
  61909=>"001111111",
  61910=>"111111011",
  61911=>"011011001",
  61912=>"000000000",
  61913=>"001001000",
  61914=>"110111000",
  61915=>"000110111",
  61916=>"110111111",
  61917=>"110000000",
  61918=>"100000000",
  61919=>"110101001",
  61920=>"011011111",
  61921=>"110111111",
  61922=>"111010111",
  61923=>"000000001",
  61924=>"000000000",
  61925=>"001001111",
  61926=>"110110010",
  61927=>"100111111",
  61928=>"110110111",
  61929=>"001101110",
  61930=>"000000000",
  61931=>"111111111",
  61932=>"010110010",
  61933=>"110111000",
  61934=>"111111111",
  61935=>"111000000",
  61936=>"101001111",
  61937=>"011010000",
  61938=>"111111111",
  61939=>"001011011",
  61940=>"001001111",
  61941=>"111110111",
  61942=>"000001001",
  61943=>"011010110",
  61944=>"111111111",
  61945=>"001011001",
  61946=>"000000000",
  61947=>"000000000",
  61948=>"111110000",
  61949=>"001001001",
  61950=>"000000001",
  61951=>"111110110",
  61952=>"011010100",
  61953=>"000011011",
  61954=>"001000000",
  61955=>"110111111",
  61956=>"000000000",
  61957=>"110110100",
  61958=>"110100000",
  61959=>"111101001",
  61960=>"000100000",
  61961=>"111111000",
  61962=>"000000000",
  61963=>"000110111",
  61964=>"000000000",
  61965=>"111111111",
  61966=>"100100000",
  61967=>"010000111",
  61968=>"100000011",
  61969=>"111111111",
  61970=>"000001001",
  61971=>"111000000",
  61972=>"000000000",
  61973=>"000000000",
  61974=>"100000000",
  61975=>"000001001",
  61976=>"111111111",
  61977=>"000001111",
  61978=>"111111111",
  61979=>"111111000",
  61980=>"001000000",
  61981=>"111111110",
  61982=>"111000000",
  61983=>"100111111",
  61984=>"000000000",
  61985=>"001000111",
  61986=>"001000000",
  61987=>"101101111",
  61988=>"000000000",
  61989=>"000000100",
  61990=>"010110110",
  61991=>"000000000",
  61992=>"000000000",
  61993=>"000110100",
  61994=>"011011111",
  61995=>"111111000",
  61996=>"000000000",
  61997=>"111111110",
  61998=>"111110100",
  61999=>"000001111",
  62000=>"111111110",
  62001=>"000000000",
  62002=>"000000011",
  62003=>"100111111",
  62004=>"001011111",
  62005=>"100011001",
  62006=>"011001001",
  62007=>"000000000",
  62008=>"000100000",
  62009=>"000000110",
  62010=>"000001111",
  62011=>"111111110",
  62012=>"110000111",
  62013=>"111001000",
  62014=>"111111011",
  62015=>"001111111",
  62016=>"100101011",
  62017=>"000000101",
  62018=>"011111111",
  62019=>"000000010",
  62020=>"001000100",
  62021=>"000000000",
  62022=>"000111110",
  62023=>"111111110",
  62024=>"000001001",
  62025=>"000000001",
  62026=>"111111110",
  62027=>"111111111",
  62028=>"101111010",
  62029=>"110111111",
  62030=>"010011100",
  62031=>"101000000",
  62032=>"111000000",
  62033=>"100000000",
  62034=>"000000000",
  62035=>"000001000",
  62036=>"000000000",
  62037=>"111100000",
  62038=>"101111111",
  62039=>"000000000",
  62040=>"000000000",
  62041=>"101101111",
  62042=>"111100100",
  62043=>"010111111",
  62044=>"011011010",
  62045=>"110110111",
  62046=>"101111111",
  62047=>"100100000",
  62048=>"101111111",
  62049=>"100100111",
  62050=>"101000000",
  62051=>"010001000",
  62052=>"000000000",
  62053=>"011111111",
  62054=>"111101000",
  62055=>"011100100",
  62056=>"111111111",
  62057=>"111111010",
  62058=>"000000000",
  62059=>"100000000",
  62060=>"111011000",
  62061=>"111111110",
  62062=>"111000000",
  62063=>"111111111",
  62064=>"000011000",
  62065=>"011000000",
  62066=>"111111100",
  62067=>"101000011",
  62068=>"100111000",
  62069=>"110100000",
  62070=>"000000000",
  62071=>"100111010",
  62072=>"000000111",
  62073=>"111101111",
  62074=>"000000000",
  62075=>"111001000",
  62076=>"001001111",
  62077=>"000000000",
  62078=>"000000000",
  62079=>"000000000",
  62080=>"011000010",
  62081=>"000000000",
  62082=>"000001111",
  62083=>"000000000",
  62084=>"101100111",
  62085=>"011000000",
  62086=>"111111000",
  62087=>"000000000",
  62088=>"000110000",
  62089=>"001011011",
  62090=>"000000000",
  62091=>"111101000",
  62092=>"100100000",
  62093=>"000000000",
  62094=>"101000111",
  62095=>"111000111",
  62096=>"000000001",
  62097=>"110110100",
  62098=>"000000011",
  62099=>"000000110",
  62100=>"000111111",
  62101=>"000000000",
  62102=>"000001011",
  62103=>"111001001",
  62104=>"100000000",
  62105=>"000000000",
  62106=>"110000000",
  62107=>"111001111",
  62108=>"000111000",
  62109=>"111111111",
  62110=>"001100000",
  62111=>"000000000",
  62112=>"000000000",
  62113=>"000010001",
  62114=>"000000111",
  62115=>"111111111",
  62116=>"000000000",
  62117=>"100100111",
  62118=>"111111111",
  62119=>"000100111",
  62120=>"000000111",
  62121=>"000000000",
  62122=>"111001000",
  62123=>"100111100",
  62124=>"100100111",
  62125=>"001001000",
  62126=>"101101001",
  62127=>"000111111",
  62128=>"000000000",
  62129=>"000110111",
  62130=>"011111111",
  62131=>"111011111",
  62132=>"101000010",
  62133=>"000001011",
  62134=>"000000000",
  62135=>"111000000",
  62136=>"000001111",
  62137=>"000000000",
  62138=>"000101101",
  62139=>"101000000",
  62140=>"000000000",
  62141=>"000000000",
  62142=>"000000000",
  62143=>"000000000",
  62144=>"000000000",
  62145=>"011011011",
  62146=>"111000000",
  62147=>"000000000",
  62148=>"011111111",
  62149=>"111111000",
  62150=>"000000000",
  62151=>"111101100",
  62152=>"111111111",
  62153=>"101101111",
  62154=>"000111111",
  62155=>"000010111",
  62156=>"000100111",
  62157=>"111111110",
  62158=>"000101111",
  62159=>"100000000",
  62160=>"111111111",
  62161=>"011010000",
  62162=>"000000101",
  62163=>"000000000",
  62164=>"000001111",
  62165=>"100111111",
  62166=>"111111011",
  62167=>"111000101",
  62168=>"111111110",
  62169=>"011000101",
  62170=>"011000011",
  62171=>"000101101",
  62172=>"000001000",
  62173=>"000000111",
  62174=>"000110000",
  62175=>"111101111",
  62176=>"000011011",
  62177=>"111111111",
  62178=>"000100110",
  62179=>"111000000",
  62180=>"110111111",
  62181=>"001110110",
  62182=>"000000000",
  62183=>"000000000",
  62184=>"111111100",
  62185=>"000110111",
  62186=>"001001111",
  62187=>"110110100",
  62188=>"000000001",
  62189=>"110000000",
  62190=>"101001000",
  62191=>"000010000",
  62192=>"111111000",
  62193=>"111111111",
  62194=>"111001000",
  62195=>"100100110",
  62196=>"011000000",
  62197=>"011011010",
  62198=>"110111111",
  62199=>"100100000",
  62200=>"100000111",
  62201=>"111111111",
  62202=>"000000111",
  62203=>"111110111",
  62204=>"110110110",
  62205=>"101011000",
  62206=>"100000100",
  62207=>"100100000",
  62208=>"000000000",
  62209=>"000100101",
  62210=>"000000001",
  62211=>"101101000",
  62212=>"100100100",
  62213=>"011111111",
  62214=>"111111111",
  62215=>"001111111",
  62216=>"111111111",
  62217=>"001000000",
  62218=>"100000000",
  62219=>"111111111",
  62220=>"110111111",
  62221=>"100111110",
  62222=>"001001000",
  62223=>"111111011",
  62224=>"011011111",
  62225=>"000001111",
  62226=>"000000111",
  62227=>"000001111",
  62228=>"111011000",
  62229=>"111111011",
  62230=>"111011000",
  62231=>"111111111",
  62232=>"011001001",
  62233=>"111111111",
  62234=>"001001001",
  62235=>"000000000",
  62236=>"000100111",
  62237=>"000000000",
  62238=>"000010111",
  62239=>"000011011",
  62240=>"000100000",
  62241=>"001011000",
  62242=>"110111110",
  62243=>"100000000",
  62244=>"001111111",
  62245=>"111111001",
  62246=>"111101000",
  62247=>"111111000",
  62248=>"011010100",
  62249=>"011000010",
  62250=>"001000100",
  62251=>"001011000",
  62252=>"000000111",
  62253=>"111101000",
  62254=>"001111101",
  62255=>"100100111",
  62256=>"001000000",
  62257=>"000000110",
  62258=>"011001111",
  62259=>"000000000",
  62260=>"000000010",
  62261=>"001011111",
  62262=>"100100000",
  62263=>"001001001",
  62264=>"111110100",
  62265=>"111000000",
  62266=>"000000000",
  62267=>"111111000",
  62268=>"001101111",
  62269=>"000001101",
  62270=>"111111000",
  62271=>"001100101",
  62272=>"111111010",
  62273=>"000101111",
  62274=>"000111111",
  62275=>"101000000",
  62276=>"001011001",
  62277=>"000100111",
  62278=>"000000000",
  62279=>"111111111",
  62280=>"000111110",
  62281=>"000000000",
  62282=>"000000000",
  62283=>"111011111",
  62284=>"111101000",
  62285=>"110110111",
  62286=>"110111110",
  62287=>"111111100",
  62288=>"010001001",
  62289=>"111111111",
  62290=>"011000001",
  62291=>"000100111",
  62292=>"101111111",
  62293=>"100111111",
  62294=>"111111111",
  62295=>"000001000",
  62296=>"000000000",
  62297=>"000000110",
  62298=>"101011011",
  62299=>"000001001",
  62300=>"111111111",
  62301=>"000000100",
  62302=>"111111111",
  62303=>"111111111",
  62304=>"000000100",
  62305=>"111111110",
  62306=>"100000000",
  62307=>"000000000",
  62308=>"110100000",
  62309=>"111111100",
  62310=>"111111000",
  62311=>"111111110",
  62312=>"101000011",
  62313=>"000011111",
  62314=>"001011111",
  62315=>"000000000",
  62316=>"011111110",
  62317=>"000000000",
  62318=>"000000000",
  62319=>"000000110",
  62320=>"100000111",
  62321=>"000000000",
  62322=>"111111111",
  62323=>"000111011",
  62324=>"111111111",
  62325=>"111111111",
  62326=>"111111111",
  62327=>"111111111",
  62328=>"000000000",
  62329=>"000111000",
  62330=>"000101111",
  62331=>"111000000",
  62332=>"011011000",
  62333=>"011011011",
  62334=>"111011000",
  62335=>"000000000",
  62336=>"001000111",
  62337=>"101100101",
  62338=>"000101001",
  62339=>"000010010",
  62340=>"000100111",
  62341=>"011001001",
  62342=>"000000000",
  62343=>"001011000",
  62344=>"010111111",
  62345=>"001000000",
  62346=>"111111110",
  62347=>"000000000",
  62348=>"000000111",
  62349=>"111110111",
  62350=>"111110110",
  62351=>"011011111",
  62352=>"110110110",
  62353=>"111011111",
  62354=>"111111111",
  62355=>"100000111",
  62356=>"000100110",
  62357=>"000010000",
  62358=>"111111111",
  62359=>"011011001",
  62360=>"000000000",
  62361=>"111111111",
  62362=>"100100110",
  62363=>"000000100",
  62364=>"001100100",
  62365=>"011111111",
  62366=>"111101101",
  62367=>"111000000",
  62368=>"100100000",
  62369=>"111111100",
  62370=>"001000100",
  62371=>"000000111",
  62372=>"100100111",
  62373=>"111111111",
  62374=>"011111111",
  62375=>"011111111",
  62376=>"000111100",
  62377=>"110110110",
  62378=>"111000011",
  62379=>"111111000",
  62380=>"111000010",
  62381=>"011001011",
  62382=>"111111110",
  62383=>"000000000",
  62384=>"000000011",
  62385=>"000000000",
  62386=>"011000000",
  62387=>"000000100",
  62388=>"111000000",
  62389=>"011111000",
  62390=>"000000111",
  62391=>"000000101",
  62392=>"100000000",
  62393=>"000111111",
  62394=>"111011011",
  62395=>"011000000",
  62396=>"001001000",
  62397=>"001101111",
  62398=>"111010000",
  62399=>"111100001",
  62400=>"000111110",
  62401=>"000111111",
  62402=>"001011011",
  62403=>"110100111",
  62404=>"001111111",
  62405=>"111111011",
  62406=>"111100000",
  62407=>"100100000",
  62408=>"100101101",
  62409=>"111000000",
  62410=>"000000000",
  62411=>"110110110",
  62412=>"000000111",
  62413=>"011111110",
  62414=>"000000100",
  62415=>"000111111",
  62416=>"111111111",
  62417=>"111111110",
  62418=>"111001000",
  62419=>"000000111",
  62420=>"101111111",
  62421=>"101111101",
  62422=>"111111111",
  62423=>"000000000",
  62424=>"000111111",
  62425=>"111000000",
  62426=>"011111101",
  62427=>"001000001",
  62428=>"111110010",
  62429=>"000000000",
  62430=>"111111111",
  62431=>"000000100",
  62432=>"000011011",
  62433=>"111010000",
  62434=>"000011111",
  62435=>"011011111",
  62436=>"001111111",
  62437=>"011111111",
  62438=>"001011111",
  62439=>"100000110",
  62440=>"001011000",
  62441=>"111000000",
  62442=>"011001000",
  62443=>"000000111",
  62444=>"111111001",
  62445=>"110100110",
  62446=>"111111010",
  62447=>"011001000",
  62448=>"000000000",
  62449=>"001101100",
  62450=>"110100101",
  62451=>"000011111",
  62452=>"000001011",
  62453=>"000000100",
  62454=>"111111000",
  62455=>"001001110",
  62456=>"111001000",
  62457=>"001000100",
  62458=>"110110100",
  62459=>"000111000",
  62460=>"000000100",
  62461=>"111001000",
  62462=>"111111111",
  62463=>"000011111",
  62464=>"011011110",
  62465=>"110100100",
  62466=>"111111111",
  62467=>"000100111",
  62468=>"000100000",
  62469=>"001000001",
  62470=>"100000101",
  62471=>"000000010",
  62472=>"111110111",
  62473=>"000100111",
  62474=>"111110111",
  62475=>"000100001",
  62476=>"100110110",
  62477=>"000000000",
  62478=>"100001111",
  62479=>"100111111",
  62480=>"100111111",
  62481=>"000000000",
  62482=>"111111111",
  62483=>"000000000",
  62484=>"010000000",
  62485=>"000000111",
  62486=>"100000100",
  62487=>"111111111",
  62488=>"000001111",
  62489=>"000010000",
  62490=>"000000000",
  62491=>"111111111",
  62492=>"000000000",
  62493=>"000001111",
  62494=>"001000000",
  62495=>"000110111",
  62496=>"001000110",
  62497=>"110010011",
  62498=>"111110000",
  62499=>"000000000",
  62500=>"000000000",
  62501=>"000000000",
  62502=>"111111111",
  62503=>"000011010",
  62504=>"111001111",
  62505=>"000000000",
  62506=>"001000111",
  62507=>"011000000",
  62508=>"000000000",
  62509=>"001011111",
  62510=>"111111010",
  62511=>"000110111",
  62512=>"110111111",
  62513=>"000000011",
  62514=>"000000011",
  62515=>"000000000",
  62516=>"011000000",
  62517=>"000000000",
  62518=>"000000001",
  62519=>"000000111",
  62520=>"110110100",
  62521=>"010010000",
  62522=>"001001011",
  62523=>"111111111",
  62524=>"001111101",
  62525=>"011111000",
  62526=>"000000101",
  62527=>"000000001",
  62528=>"001000000",
  62529=>"000000000",
  62530=>"110111111",
  62531=>"100000000",
  62532=>"000000001",
  62533=>"001000000",
  62534=>"001001000",
  62535=>"000000000",
  62536=>"001001001",
  62537=>"111111111",
  62538=>"111111110",
  62539=>"000000000",
  62540=>"111111011",
  62541=>"110110000",
  62542=>"111111000",
  62543=>"111111010",
  62544=>"111100111",
  62545=>"000000000",
  62546=>"000000000",
  62547=>"010000000",
  62548=>"000110000",
  62549=>"100010000",
  62550=>"000000111",
  62551=>"000000000",
  62552=>"001001110",
  62553=>"001000000",
  62554=>"000111100",
  62555=>"000000001",
  62556=>"111111010",
  62557=>"111001000",
  62558=>"000000000",
  62559=>"010111100",
  62560=>"011111110",
  62561=>"000000000",
  62562=>"000000001",
  62563=>"000000000",
  62564=>"000110010",
  62565=>"000010111",
  62566=>"110110111",
  62567=>"111000111",
  62568=>"111000000",
  62569=>"000000000",
  62570=>"111111111",
  62571=>"000000100",
  62572=>"000000011",
  62573=>"111011011",
  62574=>"111111100",
  62575=>"111110110",
  62576=>"000010000",
  62577=>"110110001",
  62578=>"000001001",
  62579=>"000000110",
  62580=>"000000000",
  62581=>"111110010",
  62582=>"111111111",
  62583=>"000000001",
  62584=>"010111101",
  62585=>"001011000",
  62586=>"000000000",
  62587=>"001001001",
  62588=>"000010000",
  62589=>"111001111",
  62590=>"111000000",
  62591=>"000000001",
  62592=>"000000000",
  62593=>"000000111",
  62594=>"111110110",
  62595=>"001111111",
  62596=>"100000000",
  62597=>"010011011",
  62598=>"111111111",
  62599=>"000000000",
  62600=>"110111111",
  62601=>"011011011",
  62602=>"000000000",
  62603=>"111111111",
  62604=>"111101001",
  62605=>"111111111",
  62606=>"001001001",
  62607=>"111111111",
  62608=>"000000000",
  62609=>"110111111",
  62610=>"011111110",
  62611=>"011111111",
  62612=>"000111111",
  62613=>"111111111",
  62614=>"110100100",
  62615=>"011001000",
  62616=>"111000001",
  62617=>"001001011",
  62618=>"100000000",
  62619=>"000000100",
  62620=>"110110111",
  62621=>"011010111",
  62622=>"011111001",
  62623=>"011001001",
  62624=>"111111111",
  62625=>"100000000",
  62626=>"000000111",
  62627=>"010011111",
  62628=>"000000000",
  62629=>"111111111",
  62630=>"000111000",
  62631=>"101100001",
  62632=>"100111111",
  62633=>"000100101",
  62634=>"100111111",
  62635=>"000000010",
  62636=>"111111010",
  62637=>"000000000",
  62638=>"000000000",
  62639=>"110000001",
  62640=>"000111001",
  62641=>"011111001",
  62642=>"000011011",
  62643=>"111011010",
  62644=>"111111111",
  62645=>"000111110",
  62646=>"000000001",
  62647=>"001011111",
  62648=>"111001001",
  62649=>"111111000",
  62650=>"000000000",
  62651=>"010001111",
  62652=>"111111110",
  62653=>"111001000",
  62654=>"010111110",
  62655=>"110111111",
  62656=>"000000000",
  62657=>"111011011",
  62658=>"001001000",
  62659=>"111111000",
  62660=>"111111011",
  62661=>"001000100",
  62662=>"011111010",
  62663=>"000000111",
  62664=>"111111101",
  62665=>"100111001",
  62666=>"010000011",
  62667=>"110110110",
  62668=>"111011001",
  62669=>"100111101",
  62670=>"000011111",
  62671=>"000000000",
  62672=>"000100110",
  62673=>"111010011",
  62674=>"000000111",
  62675=>"000000000",
  62676=>"011111011",
  62677=>"000000001",
  62678=>"111111110",
  62679=>"111111011",
  62680=>"000000100",
  62681=>"000000000",
  62682=>"001000000",
  62683=>"111111111",
  62684=>"111110110",
  62685=>"100111111",
  62686=>"011111000",
  62687=>"000000000",
  62688=>"111111110",
  62689=>"000000100",
  62690=>"000111111",
  62691=>"111111100",
  62692=>"000111000",
  62693=>"011000001",
  62694=>"000000110",
  62695=>"000000111",
  62696=>"011111110",
  62697=>"000000000",
  62698=>"010010111",
  62699=>"111111111",
  62700=>"000000111",
  62701=>"110110110",
  62702=>"011011011",
  62703=>"000000000",
  62704=>"100010001",
  62705=>"000000000",
  62706=>"111111111",
  62707=>"000000000",
  62708=>"111000000",
  62709=>"111110100",
  62710=>"111111100",
  62711=>"111110100",
  62712=>"111000010",
  62713=>"111111000",
  62714=>"000000000",
  62715=>"001111111",
  62716=>"111111001",
  62717=>"111110001",
  62718=>"110000000",
  62719=>"111111111",
  62720=>"000000000",
  62721=>"001000000",
  62722=>"111111111",
  62723=>"100110001",
  62724=>"000000101",
  62725=>"000000000",
  62726=>"111011011",
  62727=>"000111111",
  62728=>"111111110",
  62729=>"000110100",
  62730=>"000000001",
  62731=>"000110111",
  62732=>"001001001",
  62733=>"000000111",
  62734=>"100000000",
  62735=>"111111111",
  62736=>"110110110",
  62737=>"000000100",
  62738=>"000001111",
  62739=>"001100100",
  62740=>"000000000",
  62741=>"111111000",
  62742=>"100000000",
  62743=>"000110101",
  62744=>"100111000",
  62745=>"010000000",
  62746=>"111111111",
  62747=>"100110110",
  62748=>"011001000",
  62749=>"000101111",
  62750=>"111111111",
  62751=>"111111000",
  62752=>"011011000",
  62753=>"000100111",
  62754=>"000101001",
  62755=>"000000101",
  62756=>"011110110",
  62757=>"000000001",
  62758=>"111111111",
  62759=>"111010000",
  62760=>"000111111",
  62761=>"101101100",
  62762=>"110000000",
  62763=>"011000000",
  62764=>"011011001",
  62765=>"000000100",
  62766=>"111111111",
  62767=>"100111111",
  62768=>"000111010",
  62769=>"000000000",
  62770=>"000000000",
  62771=>"111111000",
  62772=>"111101000",
  62773=>"111111111",
  62774=>"110000111",
  62775=>"111011001",
  62776=>"001001011",
  62777=>"000000000",
  62778=>"111000110",
  62779=>"000000000",
  62780=>"000000000",
  62781=>"000001111",
  62782=>"010000000",
  62783=>"010111111",
  62784=>"000000000",
  62785=>"000111111",
  62786=>"110000000",
  62787=>"000000001",
  62788=>"000001011",
  62789=>"100110100",
  62790=>"100100110",
  62791=>"111111111",
  62792=>"111000000",
  62793=>"000111111",
  62794=>"000000100",
  62795=>"011011011",
  62796=>"111010100",
  62797=>"100000000",
  62798=>"010000000",
  62799=>"001001000",
  62800=>"111100110",
  62801=>"111111100",
  62802=>"001111000",
  62803=>"111000000",
  62804=>"111111111",
  62805=>"000010000",
  62806=>"111011111",
  62807=>"110111111",
  62808=>"110111111",
  62809=>"001001000",
  62810=>"010000000",
  62811=>"111111010",
  62812=>"101000000",
  62813=>"000000000",
  62814=>"010000011",
  62815=>"100110010",
  62816=>"111110100",
  62817=>"000000000",
  62818=>"001001101",
  62819=>"011111111",
  62820=>"000000000",
  62821=>"001000101",
  62822=>"000000100",
  62823=>"100110000",
  62824=>"000000000",
  62825=>"011011000",
  62826=>"001000000",
  62827=>"111111111",
  62828=>"000110000",
  62829=>"010111111",
  62830=>"111111111",
  62831=>"000000000",
  62832=>"100000000",
  62833=>"100010000",
  62834=>"011010000",
  62835=>"001001001",
  62836=>"111111110",
  62837=>"000000111",
  62838=>"000000011",
  62839=>"000000111",
  62840=>"000000000",
  62841=>"000000011",
  62842=>"001001000",
  62843=>"010011111",
  62844=>"000000010",
  62845=>"111111111",
  62846=>"111111011",
  62847=>"111101000",
  62848=>"000000011",
  62849=>"100000000",
  62850=>"100100100",
  62851=>"010111110",
  62852=>"111111111",
  62853=>"001000001",
  62854=>"011000000",
  62855=>"000011011",
  62856=>"000001001",
  62857=>"111101100",
  62858=>"110011011",
  62859=>"011001001",
  62860=>"011000111",
  62861=>"000001011",
  62862=>"111111000",
  62863=>"000110111",
  62864=>"110111100",
  62865=>"110110000",
  62866=>"111110111",
  62867=>"000000000",
  62868=>"000000010",
  62869=>"000010000",
  62870=>"001000001",
  62871=>"001111111",
  62872=>"111111011",
  62873=>"000000000",
  62874=>"000000000",
  62875=>"101000000",
  62876=>"100100111",
  62877=>"000000000",
  62878=>"100100100",
  62879=>"111000000",
  62880=>"111111111",
  62881=>"001111000",
  62882=>"001011111",
  62883=>"111110111",
  62884=>"111111110",
  62885=>"000000000",
  62886=>"111111000",
  62887=>"000000000",
  62888=>"000001000",
  62889=>"101111111",
  62890=>"111110000",
  62891=>"000100110",
  62892=>"100110111",
  62893=>"000000001",
  62894=>"110000000",
  62895=>"111111111",
  62896=>"000000011",
  62897=>"011000011",
  62898=>"001001111",
  62899=>"000100100",
  62900=>"111100000",
  62901=>"000000100",
  62902=>"011011111",
  62903=>"011000001",
  62904=>"110110011",
  62905=>"011111100",
  62906=>"111111010",
  62907=>"111111111",
  62908=>"001111111",
  62909=>"111101011",
  62910=>"011011111",
  62911=>"000000000",
  62912=>"011011111",
  62913=>"111000000",
  62914=>"111111111",
  62915=>"000000000",
  62916=>"000000000",
  62917=>"111100100",
  62918=>"000000000",
  62919=>"111111001",
  62920=>"111110100",
  62921=>"111111000",
  62922=>"000000001",
  62923=>"111011100",
  62924=>"100001011",
  62925=>"011000111",
  62926=>"100100001",
  62927=>"110110111",
  62928=>"011010111",
  62929=>"111111101",
  62930=>"111111111",
  62931=>"000000110",
  62932=>"111111111",
  62933=>"000111111",
  62934=>"000011111",
  62935=>"010011001",
  62936=>"000001011",
  62937=>"110010000",
  62938=>"111111111",
  62939=>"111000001",
  62940=>"000000000",
  62941=>"000000111",
  62942=>"000110111",
  62943=>"101001000",
  62944=>"011001000",
  62945=>"011111111",
  62946=>"000000000",
  62947=>"011001100",
  62948=>"111111100",
  62949=>"111111111",
  62950=>"101100111",
  62951=>"100000100",
  62952=>"001100000",
  62953=>"111111111",
  62954=>"010011011",
  62955=>"000100111",
  62956=>"000000111",
  62957=>"111111011",
  62958=>"011000000",
  62959=>"011001000",
  62960=>"000000000",
  62961=>"001111000",
  62962=>"111011011",
  62963=>"000000001",
  62964=>"111111111",
  62965=>"100111111",
  62966=>"000000110",
  62967=>"011001001",
  62968=>"000111111",
  62969=>"111111101",
  62970=>"110000000",
  62971=>"011001111",
  62972=>"010000111",
  62973=>"111111111",
  62974=>"011001001",
  62975=>"000000000",
  62976=>"110110110",
  62977=>"111011000",
  62978=>"111000101",
  62979=>"011111010",
  62980=>"000000110",
  62981=>"100000000",
  62982=>"101101111",
  62983=>"000000000",
  62984=>"100000110",
  62985=>"001001011",
  62986=>"111111111",
  62987=>"111111110",
  62988=>"011010111",
  62989=>"000000000",
  62990=>"000000111",
  62991=>"000100111",
  62992=>"110110010",
  62993=>"110111101",
  62994=>"111111111",
  62995=>"011001000",
  62996=>"100000000",
  62997=>"100100000",
  62998=>"111100000",
  62999=>"000001000",
  63000=>"010000000",
  63001=>"111111111",
  63002=>"000000000",
  63003=>"000000000",
  63004=>"111111111",
  63005=>"011111111",
  63006=>"000011000",
  63007=>"111111111",
  63008=>"111111111",
  63009=>"110110111",
  63010=>"001000111",
  63011=>"111110110",
  63012=>"000000000",
  63013=>"001000100",
  63014=>"111100100",
  63015=>"000000101",
  63016=>"000000110",
  63017=>"010000000",
  63018=>"000000111",
  63019=>"111111001",
  63020=>"000000110",
  63021=>"111000111",
  63022=>"000000001",
  63023=>"110110100",
  63024=>"000000000",
  63025=>"101001111",
  63026=>"001100100",
  63027=>"000001001",
  63028=>"000001000",
  63029=>"000000000",
  63030=>"100000000",
  63031=>"011000110",
  63032=>"000000000",
  63033=>"101001111",
  63034=>"000000001",
  63035=>"010100000",
  63036=>"111100000",
  63037=>"000110111",
  63038=>"101111111",
  63039=>"000000111",
  63040=>"111111111",
  63041=>"111111111",
  63042=>"000000000",
  63043=>"110110111",
  63044=>"000000000",
  63045=>"000000000",
  63046=>"000000011",
  63047=>"111111111",
  63048=>"001001011",
  63049=>"000000000",
  63050=>"111111001",
  63051=>"111111110",
  63052=>"000000000",
  63053=>"111011111",
  63054=>"011000000",
  63055=>"111101101",
  63056=>"010111111",
  63057=>"111110000",
  63058=>"111111111",
  63059=>"011011011",
  63060=>"000000000",
  63061=>"000000111",
  63062=>"110000111",
  63063=>"000000000",
  63064=>"111000000",
  63065=>"100000000",
  63066=>"000110000",
  63067=>"110110110",
  63068=>"000000111",
  63069=>"000000000",
  63070=>"000111111",
  63071=>"110111111",
  63072=>"111100000",
  63073=>"000000100",
  63074=>"100000111",
  63075=>"101001000",
  63076=>"000000000",
  63077=>"110111000",
  63078=>"010010010",
  63079=>"000111111",
  63080=>"000111111",
  63081=>"001001001",
  63082=>"111010000",
  63083=>"110100000",
  63084=>"110110100",
  63085=>"111111111",
  63086=>"000000111",
  63087=>"110111011",
  63088=>"000000100",
  63089=>"000000001",
  63090=>"100111111",
  63091=>"111001011",
  63092=>"100000000",
  63093=>"100100000",
  63094=>"000000000",
  63095=>"000000000",
  63096=>"010000000",
  63097=>"111111111",
  63098=>"111000000",
  63099=>"001000111",
  63100=>"110110110",
  63101=>"000000000",
  63102=>"000000000",
  63103=>"000000000",
  63104=>"111111100",
  63105=>"000000000",
  63106=>"000000000",
  63107=>"000000000",
  63108=>"000000100",
  63109=>"111100111",
  63110=>"110110110",
  63111=>"110111110",
  63112=>"111101000",
  63113=>"000000000",
  63114=>"000000101",
  63115=>"000000000",
  63116=>"110000000",
  63117=>"111111111",
  63118=>"010111111",
  63119=>"000001001",
  63120=>"111100101",
  63121=>"000000000",
  63122=>"111111111",
  63123=>"000000000",
  63124=>"000000000",
  63125=>"010000000",
  63126=>"100000000",
  63127=>"100000101",
  63128=>"000000000",
  63129=>"000000011",
  63130=>"000000000",
  63131=>"001001111",
  63132=>"110110111",
  63133=>"001111111",
  63134=>"100000000",
  63135=>"111011001",
  63136=>"111111111",
  63137=>"000000000",
  63138=>"101001001",
  63139=>"110111111",
  63140=>"000000000",
  63141=>"001111111",
  63142=>"111111111",
  63143=>"111110010",
  63144=>"000000111",
  63145=>"111111111",
  63146=>"111111111",
  63147=>"011001000",
  63148=>"000101111",
  63149=>"011011111",
  63150=>"010111111",
  63151=>"000011111",
  63152=>"111011001",
  63153=>"100000011",
  63154=>"111111111",
  63155=>"110100100",
  63156=>"111010000",
  63157=>"110111110",
  63158=>"111111111",
  63159=>"111111111",
  63160=>"111111111",
  63161=>"000000000",
  63162=>"001000000",
  63163=>"110010000",
  63164=>"111111111",
  63165=>"111000111",
  63166=>"111101111",
  63167=>"111111111",
  63168=>"010111111",
  63169=>"001111011",
  63170=>"111111111",
  63171=>"010111111",
  63172=>"110111111",
  63173=>"111111000",
  63174=>"111111111",
  63175=>"010000111",
  63176=>"000111010",
  63177=>"000000001",
  63178=>"001000000",
  63179=>"110110111",
  63180=>"100111111",
  63181=>"110111001",
  63182=>"000000000",
  63183=>"001000000",
  63184=>"111111101",
  63185=>"011000000",
  63186=>"111111111",
  63187=>"001001000",
  63188=>"001000000",
  63189=>"000001000",
  63190=>"000000000",
  63191=>"001000111",
  63192=>"111111111",
  63193=>"111111111",
  63194=>"000000000",
  63195=>"000010000",
  63196=>"111111111",
  63197=>"111101101",
  63198=>"000000000",
  63199=>"100001000",
  63200=>"001111111",
  63201=>"000000111",
  63202=>"110110110",
  63203=>"111111111",
  63204=>"100000000",
  63205=>"010011111",
  63206=>"111111111",
  63207=>"100111111",
  63208=>"111111111",
  63209=>"011111111",
  63210=>"000000000",
  63211=>"111000000",
  63212=>"000000000",
  63213=>"100000000",
  63214=>"111111111",
  63215=>"111111111",
  63216=>"000000000",
  63217=>"100000001",
  63218=>"000110110",
  63219=>"000000000",
  63220=>"111011001",
  63221=>"011011011",
  63222=>"111111000",
  63223=>"101101000",
  63224=>"101110110",
  63225=>"010110111",
  63226=>"011111111",
  63227=>"000000000",
  63228=>"011000000",
  63229=>"011001011",
  63230=>"000000000",
  63231=>"001111111",
  63232=>"110111111",
  63233=>"011011000",
  63234=>"000000111",
  63235=>"111111110",
  63236=>"000000101",
  63237=>"000000000",
  63238=>"111101000",
  63239=>"000000001",
  63240=>"100000000",
  63241=>"000000000",
  63242=>"000111111",
  63243=>"000000000",
  63244=>"000000000",
  63245=>"000000000",
  63246=>"000000001",
  63247=>"110000000",
  63248=>"000000100",
  63249=>"000000011",
  63250=>"000000001",
  63251=>"111000000",
  63252=>"111111111",
  63253=>"000000000",
  63254=>"011011001",
  63255=>"110000000",
  63256=>"000000000",
  63257=>"001000001",
  63258=>"000000000",
  63259=>"111101111",
  63260=>"000000001",
  63261=>"000000001",
  63262=>"000000000",
  63263=>"111111111",
  63264=>"101111010",
  63265=>"001000101",
  63266=>"100100000",
  63267=>"111111111",
  63268=>"000000001",
  63269=>"111111001",
  63270=>"100110100",
  63271=>"000000101",
  63272=>"000000000",
  63273=>"011111000",
  63274=>"101100101",
  63275=>"111111000",
  63276=>"000110110",
  63277=>"110110100",
  63278=>"111111111",
  63279=>"000000000",
  63280=>"110111011",
  63281=>"100111111",
  63282=>"000000000",
  63283=>"111111110",
  63284=>"111111000",
  63285=>"000000101",
  63286=>"000000000",
  63287=>"000000000",
  63288=>"000000000",
  63289=>"000000111",
  63290=>"000000100",
  63291=>"111111000",
  63292=>"111111111",
  63293=>"100000101",
  63294=>"000101111",
  63295=>"011000000",
  63296=>"111000000",
  63297=>"000000000",
  63298=>"010011111",
  63299=>"000100111",
  63300=>"111111111",
  63301=>"101111111",
  63302=>"111110111",
  63303=>"000111111",
  63304=>"000000111",
  63305=>"111100100",
  63306=>"111111111",
  63307=>"111110100",
  63308=>"101001111",
  63309=>"101000111",
  63310=>"000000000",
  63311=>"110110100",
  63312=>"100110101",
  63313=>"001011111",
  63314=>"000100100",
  63315=>"011000011",
  63316=>"000000000",
  63317=>"011011011",
  63318=>"011000000",
  63319=>"111111111",
  63320=>"000000000",
  63321=>"111110111",
  63322=>"111111000",
  63323=>"111001111",
  63324=>"000101111",
  63325=>"111111011",
  63326=>"111001001",
  63327=>"000111001",
  63328=>"111111111",
  63329=>"001000000",
  63330=>"110111000",
  63331=>"100111111",
  63332=>"111111110",
  63333=>"000000001",
  63334=>"000000110",
  63335=>"111101111",
  63336=>"011011001",
  63337=>"000010111",
  63338=>"000000000",
  63339=>"111110110",
  63340=>"100000000",
  63341=>"000000000",
  63342=>"001111111",
  63343=>"011001001",
  63344=>"000000000",
  63345=>"111111111",
  63346=>"011011111",
  63347=>"111000001",
  63348=>"000000000",
  63349=>"001001111",
  63350=>"101000111",
  63351=>"111000000",
  63352=>"000000111",
  63353=>"011000000",
  63354=>"000000111",
  63355=>"000111111",
  63356=>"000000000",
  63357=>"011111111",
  63358=>"011111111",
  63359=>"001111111",
  63360=>"000000000",
  63361=>"000011001",
  63362=>"000000000",
  63363=>"101000000",
  63364=>"000111111",
  63365=>"000000111",
  63366=>"000001111",
  63367=>"000000000",
  63368=>"000000000",
  63369=>"000100110",
  63370=>"010011111",
  63371=>"111110000",
  63372=>"101101111",
  63373=>"011110100",
  63374=>"111011001",
  63375=>"011001001",
  63376=>"000000000",
  63377=>"111111111",
  63378=>"101001100",
  63379=>"110110111",
  63380=>"010110010",
  63381=>"000000000",
  63382=>"111111111",
  63383=>"000001001",
  63384=>"000101111",
  63385=>"111101000",
  63386=>"000000010",
  63387=>"011000000",
  63388=>"100100010",
  63389=>"111111111",
  63390=>"000000000",
  63391=>"000000000",
  63392=>"100100000",
  63393=>"111111011",
  63394=>"001001111",
  63395=>"000000000",
  63396=>"111111111",
  63397=>"000000010",
  63398=>"000000000",
  63399=>"111101111",
  63400=>"000011111",
  63401=>"010000001",
  63402=>"000111100",
  63403=>"000000010",
  63404=>"000000000",
  63405=>"011011000",
  63406=>"001111001",
  63407=>"110111110",
  63408=>"000110000",
  63409=>"000100111",
  63410=>"001111110",
  63411=>"000000000",
  63412=>"111110110",
  63413=>"001111111",
  63414=>"111111111",
  63415=>"001010100",
  63416=>"000000111",
  63417=>"010111111",
  63418=>"011000000",
  63419=>"000100100",
  63420=>"000000000",
  63421=>"000001111",
  63422=>"000000000",
  63423=>"000000000",
  63424=>"000000000",
  63425=>"111100000",
  63426=>"000000000",
  63427=>"000000000",
  63428=>"000000000",
  63429=>"111001011",
  63430=>"000000010",
  63431=>"000000000",
  63432=>"000000000",
  63433=>"010001111",
  63434=>"111111111",
  63435=>"000000000",
  63436=>"011010000",
  63437=>"000000000",
  63438=>"111000000",
  63439=>"000000000",
  63440=>"000000000",
  63441=>"000000000",
  63442=>"111111001",
  63443=>"000000000",
  63444=>"111111111",
  63445=>"111111111",
  63446=>"000000000",
  63447=>"111110111",
  63448=>"000000000",
  63449=>"111101011",
  63450=>"000000000",
  63451=>"111111111",
  63452=>"000000110",
  63453=>"111000111",
  63454=>"111111111",
  63455=>"000000000",
  63456=>"100000000",
  63457=>"111111011",
  63458=>"111111111",
  63459=>"000000000",
  63460=>"111111111",
  63461=>"110110111",
  63462=>"111111000",
  63463=>"101000000",
  63464=>"010000111",
  63465=>"111110111",
  63466=>"011000000",
  63467=>"000000100",
  63468=>"000000000",
  63469=>"000100110",
  63470=>"111111111",
  63471=>"000000000",
  63472=>"100000001",
  63473=>"111111110",
  63474=>"000010111",
  63475=>"111111111",
  63476=>"111111111",
  63477=>"000000000",
  63478=>"000000000",
  63479=>"111111110",
  63480=>"010111110",
  63481=>"110000100",
  63482=>"101001111",
  63483=>"000000000",
  63484=>"111111010",
  63485=>"000000001",
  63486=>"010001000",
  63487=>"111111111",
  63488=>"111111000",
  63489=>"111000000",
  63490=>"000000000",
  63491=>"111111010",
  63492=>"011111111",
  63493=>"101000000",
  63494=>"111110000",
  63495=>"000000000",
  63496=>"111111000",
  63497=>"111111100",
  63498=>"000110100",
  63499=>"110100111",
  63500=>"111111110",
  63501=>"100000000",
  63502=>"000000111",
  63503=>"000000011",
  63504=>"110111111",
  63505=>"111111111",
  63506=>"111111111",
  63507=>"101000000",
  63508=>"000000000",
  63509=>"111011001",
  63510=>"111100100",
  63511=>"100100111",
  63512=>"110110110",
  63513=>"111111111",
  63514=>"000000111",
  63515=>"000000000",
  63516=>"110000111",
  63517=>"000000100",
  63518=>"011111111",
  63519=>"011110000",
  63520=>"000000101",
  63521=>"110111111",
  63522=>"010110000",
  63523=>"000000000",
  63524=>"111111111",
  63525=>"000000000",
  63526=>"000000000",
  63527=>"111111100",
  63528=>"000000100",
  63529=>"111111111",
  63530=>"111000101",
  63531=>"000000111",
  63532=>"000000111",
  63533=>"000001000",
  63534=>"111111111",
  63535=>"001111111",
  63536=>"000011111",
  63537=>"000000000",
  63538=>"000000010",
  63539=>"000100100",
  63540=>"111010111",
  63541=>"111111111",
  63542=>"000000010",
  63543=>"000000000",
  63544=>"100001001",
  63545=>"111111111",
  63546=>"000000000",
  63547=>"001001001",
  63548=>"000000111",
  63549=>"100111000",
  63550=>"011001001",
  63551=>"000101111",
  63552=>"000000000",
  63553=>"000000000",
  63554=>"111111111",
  63555=>"111001111",
  63556=>"110110110",
  63557=>"000000100",
  63558=>"000000000",
  63559=>"111111111",
  63560=>"111100000",
  63561=>"000000000",
  63562=>"111111111",
  63563=>"001000111",
  63564=>"000000000",
  63565=>"110000101",
  63566=>"001000000",
  63567=>"111111100",
  63568=>"000111000",
  63569=>"111111111",
  63570=>"110111111",
  63571=>"111111111",
  63572=>"000111010",
  63573=>"001001001",
  63574=>"101101000",
  63575=>"000000000",
  63576=>"000000000",
  63577=>"101100101",
  63578=>"000001111",
  63579=>"111110000",
  63580=>"000000011",
  63581=>"000000011",
  63582=>"001101001",
  63583=>"000100100",
  63584=>"000101111",
  63585=>"111111011",
  63586=>"000110111",
  63587=>"110010110",
  63588=>"000101001",
  63589=>"000011111",
  63590=>"000000000",
  63591=>"001010011",
  63592=>"010111111",
  63593=>"000000101",
  63594=>"110000000",
  63595=>"100111111",
  63596=>"101101111",
  63597=>"000011111",
  63598=>"100000111",
  63599=>"000000000",
  63600=>"010111111",
  63601=>"111011011",
  63602=>"000000000",
  63603=>"000000000",
  63604=>"001111000",
  63605=>"000001011",
  63606=>"111111111",
  63607=>"111111111",
  63608=>"000000000",
  63609=>"111111111",
  63610=>"111111111",
  63611=>"000000000",
  63612=>"100110111",
  63613=>"111100000",
  63614=>"111111111",
  63615=>"000011111",
  63616=>"111000000",
  63617=>"000000100",
  63618=>"111000000",
  63619=>"110111010",
  63620=>"000000000",
  63621=>"000001111",
  63622=>"100111100",
  63623=>"000001011",
  63624=>"000000010",
  63625=>"000100110",
  63626=>"000000000",
  63627=>"111000000",
  63628=>"011000101",
  63629=>"111111011",
  63630=>"000000000",
  63631=>"111111111",
  63632=>"000000111",
  63633=>"100000000",
  63634=>"101111111",
  63635=>"111110111",
  63636=>"000000001",
  63637=>"111101111",
  63638=>"000000111",
  63639=>"111001000",
  63640=>"000000111",
  63641=>"000000001",
  63642=>"111111111",
  63643=>"000000000",
  63644=>"000000000",
  63645=>"000000000",
  63646=>"100000000",
  63647=>"110000000",
  63648=>"010000000",
  63649=>"111110010",
  63650=>"000000000",
  63651=>"111000011",
  63652=>"111001001",
  63653=>"110101100",
  63654=>"000000110",
  63655=>"011011001",
  63656=>"010010010",
  63657=>"011111111",
  63658=>"000000000",
  63659=>"000000111",
  63660=>"000100000",
  63661=>"011111110",
  63662=>"111111001",
  63663=>"000001111",
  63664=>"000001000",
  63665=>"111001111",
  63666=>"111111111",
  63667=>"111000100",
  63668=>"110110111",
  63669=>"001000111",
  63670=>"110110000",
  63671=>"111111111",
  63672=>"110111111",
  63673=>"111111010",
  63674=>"000000000",
  63675=>"110100110",
  63676=>"101111001",
  63677=>"000111111",
  63678=>"000111001",
  63679=>"011000000",
  63680=>"011011000",
  63681=>"111111111",
  63682=>"111000000",
  63683=>"001111000",
  63684=>"111111111",
  63685=>"000000000",
  63686=>"111111000",
  63687=>"101001000",
  63688=>"000000001",
  63689=>"000000000",
  63690=>"000000000",
  63691=>"100101111",
  63692=>"111111111",
  63693=>"111111000",
  63694=>"000110111",
  63695=>"000000101",
  63696=>"111001001",
  63697=>"101000000",
  63698=>"000100000",
  63699=>"111111111",
  63700=>"111110111",
  63701=>"000000111",
  63702=>"000111111",
  63703=>"000111111",
  63704=>"011001111",
  63705=>"000101000",
  63706=>"110000000",
  63707=>"000000111",
  63708=>"100000000",
  63709=>"000001111",
  63710=>"000000111",
  63711=>"000000000",
  63712=>"111000001",
  63713=>"000000010",
  63714=>"111111000",
  63715=>"000000000",
  63716=>"111111000",
  63717=>"011001011",
  63718=>"000000101",
  63719=>"110111111",
  63720=>"000000000",
  63721=>"111111111",
  63722=>"110110001",
  63723=>"101111111",
  63724=>"110000000",
  63725=>"001011000",
  63726=>"110111011",
  63727=>"111111100",
  63728=>"111111111",
  63729=>"111111111",
  63730=>"000000000",
  63731=>"001000100",
  63732=>"111111001",
  63733=>"000000011",
  63734=>"000000000",
  63735=>"101000101",
  63736=>"111111111",
  63737=>"000011011",
  63738=>"000000000",
  63739=>"111111001",
  63740=>"111001000",
  63741=>"001001000",
  63742=>"111000000",
  63743=>"000000000",
  63744=>"000000000",
  63745=>"111000110",
  63746=>"111111111",
  63747=>"000000000",
  63748=>"011111110",
  63749=>"011000011",
  63750=>"000100000",
  63751=>"111101101",
  63752=>"111111111",
  63753=>"000100110",
  63754=>"000000000",
  63755=>"101000001",
  63756=>"001000111",
  63757=>"111111111",
  63758=>"100001000",
  63759=>"000111111",
  63760=>"100000111",
  63761=>"110000100",
  63762=>"000000110",
  63763=>"000000001",
  63764=>"011111000",
  63765=>"010010111",
  63766=>"011111111",
  63767=>"000111111",
  63768=>"001001011",
  63769=>"000000000",
  63770=>"000000000",
  63771=>"000001001",
  63772=>"100100000",
  63773=>"100100000",
  63774=>"000000000",
  63775=>"111000000",
  63776=>"100001111",
  63777=>"111011111",
  63778=>"111101111",
  63779=>"100000111",
  63780=>"000000001",
  63781=>"111111111",
  63782=>"111111101",
  63783=>"111111111",
  63784=>"111000000",
  63785=>"111111111",
  63786=>"000000001",
  63787=>"000000100",
  63788=>"110000100",
  63789=>"001000001",
  63790=>"111111000",
  63791=>"000000000",
  63792=>"000000000",
  63793=>"001000000",
  63794=>"001000000",
  63795=>"001111111",
  63796=>"000110100",
  63797=>"100111000",
  63798=>"000100100",
  63799=>"110111111",
  63800=>"000000111",
  63801=>"111111111",
  63802=>"000000111",
  63803=>"000000000",
  63804=>"000000000",
  63805=>"001011111",
  63806=>"110111111",
  63807=>"000000000",
  63808=>"000000001",
  63809=>"001001111",
  63810=>"110000000",
  63811=>"001000000",
  63812=>"000110000",
  63813=>"111111111",
  63814=>"110011000",
  63815=>"111111111",
  63816=>"000000111",
  63817=>"000000000",
  63818=>"001000001",
  63819=>"110110001",
  63820=>"111111111",
  63821=>"101000000",
  63822=>"111111000",
  63823=>"011011000",
  63824=>"111000001",
  63825=>"100000000",
  63826=>"111111111",
  63827=>"000000000",
  63828=>"000000001",
  63829=>"011011011",
  63830=>"111111111",
  63831=>"000110111",
  63832=>"000111111",
  63833=>"000000111",
  63834=>"000110110",
  63835=>"000000001",
  63836=>"101000000",
  63837=>"000000000",
  63838=>"111111110",
  63839=>"100111111",
  63840=>"100000000",
  63841=>"000000000",
  63842=>"000111111",
  63843=>"000000000",
  63844=>"110110110",
  63845=>"000000000",
  63846=>"111101111",
  63847=>"000100000",
  63848=>"000110010",
  63849=>"111111111",
  63850=>"100111101",
  63851=>"000000101",
  63852=>"011111111",
  63853=>"111111111",
  63854=>"000000000",
  63855=>"000011111",
  63856=>"111000000",
  63857=>"000000001",
  63858=>"111111011",
  63859=>"111111111",
  63860=>"101111111",
  63861=>"000000000",
  63862=>"111110000",
  63863=>"011011000",
  63864=>"111111111",
  63865=>"000001001",
  63866=>"111111111",
  63867=>"111111111",
  63868=>"000010111",
  63869=>"011011111",
  63870=>"000000000",
  63871=>"000110111",
  63872=>"011111011",
  63873=>"111111111",
  63874=>"000000000",
  63875=>"000000000",
  63876=>"111000001",
  63877=>"000000000",
  63878=>"000000000",
  63879=>"000100111",
  63880=>"000000000",
  63881=>"111000000",
  63882=>"000100110",
  63883=>"111000000",
  63884=>"101111111",
  63885=>"111111111",
  63886=>"011111111",
  63887=>"000011111",
  63888=>"000000111",
  63889=>"000000000",
  63890=>"111111111",
  63891=>"000000000",
  63892=>"000000111",
  63893=>"000000000",
  63894=>"000111100",
  63895=>"111110100",
  63896=>"111000111",
  63897=>"111000000",
  63898=>"111111010",
  63899=>"111111111",
  63900=>"111111111",
  63901=>"000000000",
  63902=>"000001111",
  63903=>"111111111",
  63904=>"111000000",
  63905=>"111111100",
  63906=>"000001111",
  63907=>"001000001",
  63908=>"100100000",
  63909=>"111111111",
  63910=>"111111111",
  63911=>"011011010",
  63912=>"011111000",
  63913=>"001111111",
  63914=>"110000000",
  63915=>"011111001",
  63916=>"000000000",
  63917=>"000000000",
  63918=>"000000000",
  63919=>"000111111",
  63920=>"000000111",
  63921=>"111001111",
  63922=>"111000000",
  63923=>"000000001",
  63924=>"111111100",
  63925=>"111111111",
  63926=>"000111111",
  63927=>"101011111",
  63928=>"111001111",
  63929=>"111111111",
  63930=>"100110110",
  63931=>"111100100",
  63932=>"111101111",
  63933=>"000000000",
  63934=>"111001000",
  63935=>"111101101",
  63936=>"111111000",
  63937=>"000000111",
  63938=>"111111111",
  63939=>"010111111",
  63940=>"110000000",
  63941=>"000000001",
  63942=>"001000111",
  63943=>"111101100",
  63944=>"111111110",
  63945=>"111111111",
  63946=>"000000000",
  63947=>"111011010",
  63948=>"000000000",
  63949=>"000011011",
  63950=>"001111110",
  63951=>"111111010",
  63952=>"001001000",
  63953=>"000000111",
  63954=>"000000000",
  63955=>"111111111",
  63956=>"100000000",
  63957=>"100110100",
  63958=>"000000111",
  63959=>"110010000",
  63960=>"101101100",
  63961=>"100110000",
  63962=>"000111111",
  63963=>"111110000",
  63964=>"000000000",
  63965=>"111111001",
  63966=>"000011001",
  63967=>"100000000",
  63968=>"001001111",
  63969=>"111111011",
  63970=>"000000111",
  63971=>"100110011",
  63972=>"001000101",
  63973=>"000011111",
  63974=>"000000000",
  63975=>"111111111",
  63976=>"000100001",
  63977=>"111111111",
  63978=>"000000000",
  63979=>"110101111",
  63980=>"000000000",
  63981=>"100100100",
  63982=>"001000000",
  63983=>"100000000",
  63984=>"000000111",
  63985=>"011111111",
  63986=>"111111110",
  63987=>"110001001",
  63988=>"111111111",
  63989=>"000010000",
  63990=>"000000000",
  63991=>"001100001",
  63992=>"000000000",
  63993=>"111000001",
  63994=>"000111111",
  63995=>"001001101",
  63996=>"111111111",
  63997=>"111000000",
  63998=>"011011111",
  63999=>"011011001",
  64000=>"001101101",
  64001=>"000000000",
  64002=>"111111111",
  64003=>"111111111",
  64004=>"000000000",
  64005=>"111000001",
  64006=>"000000000",
  64007=>"001000001",
  64008=>"011000000",
  64009=>"110100000",
  64010=>"110111111",
  64011=>"100111111",
  64012=>"000100110",
  64013=>"111000100",
  64014=>"011011111",
  64015=>"000111111",
  64016=>"011001111",
  64017=>"100000011",
  64018=>"101110111",
  64019=>"111111111",
  64020=>"000000000",
  64021=>"000000010",
  64022=>"000110000",
  64023=>"111101111",
  64024=>"111111111",
  64025=>"000000000",
  64026=>"000010111",
  64027=>"111111011",
  64028=>"111111111",
  64029=>"111110100",
  64030=>"000000000",
  64031=>"000000000",
  64032=>"111111000",
  64033=>"000000000",
  64034=>"111111111",
  64035=>"000000000",
  64036=>"001000000",
  64037=>"000110111",
  64038=>"111000000",
  64039=>"010000000",
  64040=>"001001001",
  64041=>"111111000",
  64042=>"111111111",
  64043=>"000000000",
  64044=>"111110111",
  64045=>"101101111",
  64046=>"111111111",
  64047=>"011000111",
  64048=>"111111111",
  64049=>"000000000",
  64050=>"000000100",
  64051=>"010000110",
  64052=>"000000000",
  64053=>"010100000",
  64054=>"111000000",
  64055=>"000000000",
  64056=>"111111111",
  64057=>"011010000",
  64058=>"111111111",
  64059=>"000000000",
  64060=>"000000000",
  64061=>"111111001",
  64062=>"111011001",
  64063=>"000000101",
  64064=>"111111000",
  64065=>"000100111",
  64066=>"111111111",
  64067=>"011000000",
  64068=>"111001000",
  64069=>"000000000",
  64070=>"000000110",
  64071=>"111111111",
  64072=>"111111111",
  64073=>"111111111",
  64074=>"011111000",
  64075=>"100000111",
  64076=>"000000000",
  64077=>"000000000",
  64078=>"110111111",
  64079=>"111111111",
  64080=>"000011000",
  64081=>"000110000",
  64082=>"000000000",
  64083=>"000000110",
  64084=>"111111111",
  64085=>"110110110",
  64086=>"111111111",
  64087=>"000001011",
  64088=>"111111111",
  64089=>"001000001",
  64090=>"010111011",
  64091=>"000000000",
  64092=>"000000010",
  64093=>"000000000",
  64094=>"111111111",
  64095=>"011001001",
  64096=>"111111111",
  64097=>"000000000",
  64098=>"000100111",
  64099=>"000000000",
  64100=>"001000111",
  64101=>"111111111",
  64102=>"111101111",
  64103=>"000000000",
  64104=>"000000000",
  64105=>"000000000",
  64106=>"000100110",
  64107=>"000000000",
  64108=>"001001001",
  64109=>"000000001",
  64110=>"000100000",
  64111=>"000000110",
  64112=>"100001100",
  64113=>"000000000",
  64114=>"101111111",
  64115=>"111111111",
  64116=>"111111000",
  64117=>"111010111",
  64118=>"000000000",
  64119=>"111111000",
  64120=>"111111111",
  64121=>"000000000",
  64122=>"101101111",
  64123=>"000001111",
  64124=>"110110100",
  64125=>"000101111",
  64126=>"000000000",
  64127=>"000000000",
  64128=>"000010111",
  64129=>"111110100",
  64130=>"001000000",
  64131=>"000100100",
  64132=>"000000001",
  64133=>"111111111",
  64134=>"000110110",
  64135=>"010000100",
  64136=>"111111111",
  64137=>"000000000",
  64138=>"000000000",
  64139=>"000000100",
  64140=>"100111111",
  64141=>"111111110",
  64142=>"000000000",
  64143=>"000000000",
  64144=>"111111111",
  64145=>"111010000",
  64146=>"001111001",
  64147=>"111111001",
  64148=>"111111111",
  64149=>"111111111",
  64150=>"111111000",
  64151=>"111000000",
  64152=>"111111001",
  64153=>"111111111",
  64154=>"000000100",
  64155=>"000000000",
  64156=>"100000000",
  64157=>"111110000",
  64158=>"000101111",
  64159=>"000000001",
  64160=>"100100000",
  64161=>"001001000",
  64162=>"111111111",
  64163=>"111011000",
  64164=>"000000000",
  64165=>"010010111",
  64166=>"111111111",
  64167=>"111111011",
  64168=>"100100100",
  64169=>"000000000",
  64170=>"100000000",
  64171=>"000000000",
  64172=>"001011111",
  64173=>"100100000",
  64174=>"000000100",
  64175=>"000000000",
  64176=>"111111111",
  64177=>"001001001",
  64178=>"000110010",
  64179=>"111111000",
  64180=>"000100101",
  64181=>"110111111",
  64182=>"111110100",
  64183=>"001000000",
  64184=>"111101001",
  64185=>"111001011",
  64186=>"101001001",
  64187=>"000000000",
  64188=>"000100111",
  64189=>"000100111",
  64190=>"000000000",
  64191=>"000110000",
  64192=>"000000100",
  64193=>"010110000",
  64194=>"111111111",
  64195=>"000100000",
  64196=>"001000000",
  64197=>"000000000",
  64198=>"000000000",
  64199=>"111000000",
  64200=>"000100110",
  64201=>"111000000",
  64202=>"100000001",
  64203=>"000110111",
  64204=>"101101111",
  64205=>"000111111",
  64206=>"000000000",
  64207=>"111111000",
  64208=>"111101101",
  64209=>"010100111",
  64210=>"111111111",
  64211=>"011011001",
  64212=>"111111111",
  64213=>"000000000",
  64214=>"000101111",
  64215=>"000000001",
  64216=>"111010111",
  64217=>"111110111",
  64218=>"000000000",
  64219=>"011011111",
  64220=>"111111111",
  64221=>"111111111",
  64222=>"110111111",
  64223=>"111000000",
  64224=>"000000000",
  64225=>"011010000",
  64226=>"111111011",
  64227=>"000000000",
  64228=>"000000000",
  64229=>"000000000",
  64230=>"000000000",
  64231=>"111111111",
  64232=>"000000000",
  64233=>"000110111",
  64234=>"001000111",
  64235=>"000000000",
  64236=>"111111111",
  64237=>"000000000",
  64238=>"111111111",
  64239=>"000111111",
  64240=>"100000000",
  64241=>"000000000",
  64242=>"111111001",
  64243=>"000000000",
  64244=>"111111111",
  64245=>"110011000",
  64246=>"011011111",
  64247=>"111111111",
  64248=>"111111111",
  64249=>"000000000",
  64250=>"101111000",
  64251=>"110111110",
  64252=>"111111111",
  64253=>"100111010",
  64254=>"001011011",
  64255=>"100110111",
  64256=>"111000111",
  64257=>"010010010",
  64258=>"110111000",
  64259=>"001001011",
  64260=>"001000000",
  64261=>"000000000",
  64262=>"111111111",
  64263=>"111111111",
  64264=>"111100110",
  64265=>"000000000",
  64266=>"000000000",
  64267=>"010000000",
  64268=>"000000000",
  64269=>"111000000",
  64270=>"000000000",
  64271=>"000000000",
  64272=>"111111111",
  64273=>"111111111",
  64274=>"100101111",
  64275=>"100110000",
  64276=>"111111111",
  64277=>"000000111",
  64278=>"111110110",
  64279=>"011011000",
  64280=>"001001010",
  64281=>"000000100",
  64282=>"101001001",
  64283=>"100111111",
  64284=>"111011010",
  64285=>"001110000",
  64286=>"000000000",
  64287=>"011000000",
  64288=>"110000000",
  64289=>"000000000",
  64290=>"101110000",
  64291=>"000000001",
  64292=>"000000000",
  64293=>"111101111",
  64294=>"111111111",
  64295=>"000000001",
  64296=>"001001111",
  64297=>"011111111",
  64298=>"111000000",
  64299=>"111111000",
  64300=>"111001000",
  64301=>"111011001",
  64302=>"000000111",
  64303=>"111111111",
  64304=>"111000000",
  64305=>"000000000",
  64306=>"111111111",
  64307=>"000000111",
  64308=>"111111111",
  64309=>"111000010",
  64310=>"000000000",
  64311=>"111111111",
  64312=>"000000000",
  64313=>"101000000",
  64314=>"111111111",
  64315=>"100111111",
  64316=>"000000100",
  64317=>"111111111",
  64318=>"000000000",
  64319=>"111111111",
  64320=>"000000000",
  64321=>"100100000",
  64322=>"011000000",
  64323=>"111111111",
  64324=>"111111011",
  64325=>"011001000",
  64326=>"000000000",
  64327=>"000000000",
  64328=>"000100000",
  64329=>"000011111",
  64330=>"000100111",
  64331=>"100000000",
  64332=>"000001001",
  64333=>"000000000",
  64334=>"111111001",
  64335=>"111111100",
  64336=>"001001000",
  64337=>"100000000",
  64338=>"111100100",
  64339=>"000000000",
  64340=>"000000111",
  64341=>"011001011",
  64342=>"110111000",
  64343=>"111111100",
  64344=>"110111110",
  64345=>"111111111",
  64346=>"111111001",
  64347=>"101000000",
  64348=>"000000000",
  64349=>"000000000",
  64350=>"000000000",
  64351=>"000000000",
  64352=>"111000010",
  64353=>"000000000",
  64354=>"000000000",
  64355=>"000001001",
  64356=>"110111111",
  64357=>"000000000",
  64358=>"111101111",
  64359=>"111000000",
  64360=>"001001111",
  64361=>"000000110",
  64362=>"000010111",
  64363=>"000000010",
  64364=>"100100110",
  64365=>"100110000",
  64366=>"110111111",
  64367=>"000000000",
  64368=>"000100111",
  64369=>"000000000",
  64370=>"000011011",
  64371=>"111111111",
  64372=>"000000000",
  64373=>"011111111",
  64374=>"000000000",
  64375=>"111001000",
  64376=>"111111101",
  64377=>"111111111",
  64378=>"110000001",
  64379=>"000001011",
  64380=>"000000001",
  64381=>"001000100",
  64382=>"000101111",
  64383=>"000000000",
  64384=>"010000000",
  64385=>"010000000",
  64386=>"000000000",
  64387=>"110111111",
  64388=>"111111111",
  64389=>"011000000",
  64390=>"111000001",
  64391=>"110001000",
  64392=>"000000000",
  64393=>"000001111",
  64394=>"111111111",
  64395=>"111111111",
  64396=>"011001001",
  64397=>"011111111",
  64398=>"000000111",
  64399=>"000000000",
  64400=>"000000000",
  64401=>"111111111",
  64402=>"101110110",
  64403=>"000000001",
  64404=>"011001000",
  64405=>"000000000",
  64406=>"001000000",
  64407=>"001000000",
  64408=>"000000110",
  64409=>"000110100",
  64410=>"111101111",
  64411=>"111000000",
  64412=>"111011011",
  64413=>"000000000",
  64414=>"000000000",
  64415=>"000000000",
  64416=>"000000000",
  64417=>"011001001",
  64418=>"000000001",
  64419=>"001001000",
  64420=>"111111111",
  64421=>"111111111",
  64422=>"111111111",
  64423=>"000000111",
  64424=>"000000000",
  64425=>"111111111",
  64426=>"111111111",
  64427=>"011000000",
  64428=>"001011000",
  64429=>"001000000",
  64430=>"000000000",
  64431=>"000000011",
  64432=>"100111111",
  64433=>"111111111",
  64434=>"111111000",
  64435=>"000000100",
  64436=>"111111111",
  64437=>"000000001",
  64438=>"000000111",
  64439=>"000011111",
  64440=>"111111000",
  64441=>"000110111",
  64442=>"111111111",
  64443=>"111101101",
  64444=>"000001111",
  64445=>"111111111",
  64446=>"110111111",
  64447=>"011110111",
  64448=>"010000000",
  64449=>"000000000",
  64450=>"000000000",
  64451=>"000000000",
  64452=>"001000000",
  64453=>"001001110",
  64454=>"000000000",
  64455=>"000000111",
  64456=>"000000000",
  64457=>"010010000",
  64458=>"000000000",
  64459=>"110111111",
  64460=>"000000000",
  64461=>"111111000",
  64462=>"111111111",
  64463=>"000000001",
  64464=>"100111111",
  64465=>"000000000",
  64466=>"000000000",
  64467=>"000000000",
  64468=>"111111111",
  64469=>"000001001",
  64470=>"111001001",
  64471=>"000010110",
  64472=>"000000000",
  64473=>"100000000",
  64474=>"111111111",
  64475=>"111101111",
  64476=>"000000001",
  64477=>"000000000",
  64478=>"000000010",
  64479=>"000000011",
  64480=>"000100111",
  64481=>"111111000",
  64482=>"111111111",
  64483=>"111111000",
  64484=>"100100001",
  64485=>"000000000",
  64486=>"101000000",
  64487=>"000001000",
  64488=>"000000000",
  64489=>"000001001",
  64490=>"110111111",
  64491=>"000000000",
  64492=>"000000001",
  64493=>"111011000",
  64494=>"000000110",
  64495=>"111100111",
  64496=>"000000000",
  64497=>"111111111",
  64498=>"000000000",
  64499=>"100000110",
  64500=>"111111111",
  64501=>"111111111",
  64502=>"000011111",
  64503=>"110100100",
  64504=>"010011000",
  64505=>"101101101",
  64506=>"001001000",
  64507=>"111111111",
  64508=>"000000010",
  64509=>"111100000",
  64510=>"011111111",
  64511=>"000100111",
  64512=>"000000101",
  64513=>"111010000",
  64514=>"111110000",
  64515=>"100000000",
  64516=>"110110000",
  64517=>"000000000",
  64518=>"111110111",
  64519=>"101111111",
  64520=>"101100000",
  64521=>"000000000",
  64522=>"100000000",
  64523=>"011000000",
  64524=>"011111011",
  64525=>"001101111",
  64526=>"000101111",
  64527=>"100110100",
  64528=>"001001001",
  64529=>"110110010",
  64530=>"000000110",
  64531=>"111111100",
  64532=>"000000000",
  64533=>"111000100",
  64534=>"001001000",
  64535=>"000011111",
  64536=>"111110000",
  64537=>"100100110",
  64538=>"001000000",
  64539=>"100001111",
  64540=>"100110111",
  64541=>"010011111",
  64542=>"001001001",
  64543=>"001100111",
  64544=>"000000111",
  64545=>"110110110",
  64546=>"001001001",
  64547=>"000000001",
  64548=>"000110000",
  64549=>"111110111",
  64550=>"111111100",
  64551=>"111110000",
  64552=>"110111111",
  64553=>"000000001",
  64554=>"000001001",
  64555=>"101110000",
  64556=>"000000000",
  64557=>"000000000",
  64558=>"001001111",
  64559=>"011111100",
  64560=>"110011111",
  64561=>"000000000",
  64562=>"110111000",
  64563=>"010010011",
  64564=>"000100110",
  64565=>"111111111",
  64566=>"110010010",
  64567=>"001001101",
  64568=>"101001001",
  64569=>"000010111",
  64570=>"111111111",
  64571=>"000000000",
  64572=>"000000101",
  64573=>"111111110",
  64574=>"111111111",
  64575=>"100100100",
  64576=>"111000110",
  64577=>"000000001",
  64578=>"000000000",
  64579=>"110110001",
  64580=>"111110111",
  64581=>"001001000",
  64582=>"101000000",
  64583=>"000000000",
  64584=>"111111100",
  64585=>"111001111",
  64586=>"101001111",
  64587=>"110110000",
  64588=>"101110111",
  64589=>"000001001",
  64590=>"001001000",
  64591=>"100111111",
  64592=>"000000000",
  64593=>"110111100",
  64594=>"111111000",
  64595=>"000101100",
  64596=>"010110000",
  64597=>"000000001",
  64598=>"000000000",
  64599=>"001111111",
  64600=>"110110110",
  64601=>"111101001",
  64602=>"000000000",
  64603=>"010000000",
  64604=>"000110111",
  64605=>"001001000",
  64606=>"111110000",
  64607=>"011111110",
  64608=>"011011011",
  64609=>"000000100",
  64610=>"111111010",
  64611=>"111111111",
  64612=>"110110000",
  64613=>"101000001",
  64614=>"000000111",
  64615=>"001000001",
  64616=>"001001001",
  64617=>"010000110",
  64618=>"100100000",
  64619=>"010000000",
  64620=>"101111111",
  64621=>"111111010",
  64622=>"000001000",
  64623=>"111111000",
  64624=>"000000000",
  64625=>"000001000",
  64626=>"000000001",
  64627=>"100010011",
  64628=>"000000000",
  64629=>"111111011",
  64630=>"000110000",
  64631=>"100100111",
  64632=>"110000000",
  64633=>"001111111",
  64634=>"011001101",
  64635=>"000000000",
  64636=>"110110111",
  64637=>"001111111",
  64638=>"010011000",
  64639=>"001000000",
  64640=>"101101000",
  64641=>"111110000",
  64642=>"000000000",
  64643=>"010010110",
  64644=>"111111111",
  64645=>"000001101",
  64646=>"111100000",
  64647=>"000000001",
  64648=>"000000110",
  64649=>"001001000",
  64650=>"111111111",
  64651=>"000000110",
  64652=>"000000000",
  64653=>"000000100",
  64654=>"010111111",
  64655=>"000000000",
  64656=>"001001101",
  64657=>"001000001",
  64658=>"000010000",
  64659=>"111100000",
  64660=>"000110110",
  64661=>"110111111",
  64662=>"111001100",
  64663=>"001000001",
  64664=>"000001001",
  64665=>"001000101",
  64666=>"001001101",
  64667=>"000100100",
  64668=>"001001001",
  64669=>"000011001",
  64670=>"111110000",
  64671=>"110110110",
  64672=>"101111111",
  64673=>"110000000",
  64674=>"110111001",
  64675=>"001001111",
  64676=>"000000100",
  64677=>"110110110",
  64678=>"111100100",
  64679=>"001011111",
  64680=>"110110001",
  64681=>"111111111",
  64682=>"001001001",
  64683=>"001011001",
  64684=>"111110100",
  64685=>"000100111",
  64686=>"111100000",
  64687=>"111111000",
  64688=>"111111111",
  64689=>"111111111",
  64690=>"010110000",
  64691=>"111101000",
  64692=>"101001001",
  64693=>"001001100",
  64694=>"000000000",
  64695=>"111100100",
  64696=>"001001011",
  64697=>"000010111",
  64698=>"111001001",
  64699=>"000000000",
  64700=>"001000111",
  64701=>"110110000",
  64702=>"000000110",
  64703=>"001001001",
  64704=>"111111010",
  64705=>"111001111",
  64706=>"000001001",
  64707=>"110111000",
  64708=>"111111111",
  64709=>"000000000",
  64710=>"111101100",
  64711=>"111010000",
  64712=>"111001001",
  64713=>"110101111",
  64714=>"000000001",
  64715=>"111001000",
  64716=>"000011010",
  64717=>"000010111",
  64718=>"111111111",
  64719=>"000000000",
  64720=>"011111111",
  64721=>"011000111",
  64722=>"000000111",
  64723=>"000000000",
  64724=>"000110110",
  64725=>"111110100",
  64726=>"000000000",
  64727=>"111111100",
  64728=>"000001000",
  64729=>"110010000",
  64730=>"110111111",
  64731=>"000110111",
  64732=>"011001001",
  64733=>"000000111",
  64734=>"110110000",
  64735=>"111001000",
  64736=>"000001101",
  64737=>"000000000",
  64738=>"000011111",
  64739=>"100100100",
  64740=>"000000000",
  64741=>"111000000",
  64742=>"000000000",
  64743=>"001001001",
  64744=>"001001000",
  64745=>"111111111",
  64746=>"100100100",
  64747=>"111001111",
  64748=>"111101111",
  64749=>"110000000",
  64750=>"001000001",
  64751=>"111111101",
  64752=>"100000110",
  64753=>"111110111",
  64754=>"001000100",
  64755=>"001000011",
  64756=>"111111111",
  64757=>"100111011",
  64758=>"011111001",
  64759=>"111001001",
  64760=>"111100000",
  64761=>"001010111",
  64762=>"100111111",
  64763=>"001001111",
  64764=>"011111011",
  64765=>"001111111",
  64766=>"000000000",
  64767=>"000001110",
  64768=>"000000111",
  64769=>"000000001",
  64770=>"000000011",
  64771=>"111111111",
  64772=>"001101111",
  64773=>"000000000",
  64774=>"111111001",
  64775=>"110000000",
  64776=>"111110000",
  64777=>"111011000",
  64778=>"100110110",
  64779=>"000000011",
  64780=>"110000000",
  64781=>"010111001",
  64782=>"110110001",
  64783=>"111000001",
  64784=>"100100000",
  64785=>"000000000",
  64786=>"001001001",
  64787=>"000000000",
  64788=>"100000101",
  64789=>"110111000",
  64790=>"111111111",
  64791=>"000000000",
  64792=>"110010000",
  64793=>"001001001",
  64794=>"101100100",
  64795=>"000001111",
  64796=>"000000011",
  64797=>"000000010",
  64798=>"001001101",
  64799=>"111010000",
  64800=>"111110000",
  64801=>"001000000",
  64802=>"000000000",
  64803=>"111111110",
  64804=>"110100101",
  64805=>"110100000",
  64806=>"001001111",
  64807=>"000000000",
  64808=>"111111111",
  64809=>"000000111",
  64810=>"110110000",
  64811=>"000000000",
  64812=>"101111001",
  64813=>"000000000",
  64814=>"000011000",
  64815=>"000000100",
  64816=>"010010000",
  64817=>"000000000",
  64818=>"001111111",
  64819=>"100000000",
  64820=>"110110111",
  64821=>"000000000",
  64822=>"000000000",
  64823=>"000000000",
  64824=>"000010000",
  64825=>"111101111",
  64826=>"000001111",
  64827=>"001000111",
  64828=>"000000000",
  64829=>"110010000",
  64830=>"100100100",
  64831=>"000000110",
  64832=>"001001000",
  64833=>"010000000",
  64834=>"001000101",
  64835=>"011011011",
  64836=>"000001011",
  64837=>"000000111",
  64838=>"000000111",
  64839=>"000000100",
  64840=>"111111001",
  64841=>"000000011",
  64842=>"100110001",
  64843=>"110110000",
  64844=>"001000100",
  64845=>"111111011",
  64846=>"000000000",
  64847=>"000111111",
  64848=>"001000100",
  64849=>"000000111",
  64850=>"111111111",
  64851=>"001001111",
  64852=>"101111000",
  64853=>"011001001",
  64854=>"001101111",
  64855=>"111111111",
  64856=>"000000111",
  64857=>"000100100",
  64858=>"010001001",
  64859=>"111111110",
  64860=>"010100100",
  64861=>"001001011",
  64862=>"000000000",
  64863=>"000000100",
  64864=>"000000000",
  64865=>"001000000",
  64866=>"000001011",
  64867=>"000000111",
  64868=>"111111011",
  64869=>"000000101",
  64870=>"000000000",
  64871=>"001000001",
  64872=>"101000100",
  64873=>"011000000",
  64874=>"010010011",
  64875=>"110000001",
  64876=>"110110100",
  64877=>"101100111",
  64878=>"111111111",
  64879=>"101001001",
  64880=>"111000000",
  64881=>"101000111",
  64882=>"110110110",
  64883=>"111111110",
  64884=>"111011001",
  64885=>"001001001",
  64886=>"000111111",
  64887=>"000000000",
  64888=>"100000000",
  64889=>"000000110",
  64890=>"000000101",
  64891=>"000001111",
  64892=>"110110111",
  64893=>"000000000",
  64894=>"011010001",
  64895=>"000000000",
  64896=>"110110000",
  64897=>"111111010",
  64898=>"100100100",
  64899=>"001001101",
  64900=>"111001000",
  64901=>"111001111",
  64902=>"000000000",
  64903=>"111111111",
  64904=>"100100001",
  64905=>"010000000",
  64906=>"000001111",
  64907=>"000011011",
  64908=>"111111111",
  64909=>"010011011",
  64910=>"110110000",
  64911=>"111111000",
  64912=>"000000000",
  64913=>"001001011",
  64914=>"110111001",
  64915=>"000001001",
  64916=>"000110111",
  64917=>"000000010",
  64918=>"011111001",
  64919=>"111001001",
  64920=>"111011111",
  64921=>"111110000",
  64922=>"111111111",
  64923=>"010010000",
  64924=>"000000010",
  64925=>"111111111",
  64926=>"011001001",
  64927=>"111111000",
  64928=>"000111101",
  64929=>"001011011",
  64930=>"110110011",
  64931=>"111111101",
  64932=>"111111101",
  64933=>"111111111",
  64934=>"111111111",
  64935=>"000111111",
  64936=>"000111111",
  64937=>"111111111",
  64938=>"110110010",
  64939=>"111011001",
  64940=>"000000110",
  64941=>"110100111",
  64942=>"110100000",
  64943=>"000000100",
  64944=>"110000000",
  64945=>"111111000",
  64946=>"000000111",
  64947=>"110110010",
  64948=>"000000011",
  64949=>"011000000",
  64950=>"001001101",
  64951=>"001001000",
  64952=>"011111111",
  64953=>"110110111",
  64954=>"110110111",
  64955=>"001111111",
  64956=>"000000000",
  64957=>"000001111",
  64958=>"001000000",
  64959=>"000000000",
  64960=>"000000000",
  64961=>"101110000",
  64962=>"000110111",
  64963=>"000000011",
  64964=>"000000000",
  64965=>"100010111",
  64966=>"000000001",
  64967=>"000010000",
  64968=>"000000011",
  64969=>"111110000",
  64970=>"001001100",
  64971=>"000010000",
  64972=>"011000000",
  64973=>"000000000",
  64974=>"110110100",
  64975=>"000000011",
  64976=>"111011000",
  64977=>"011111110",
  64978=>"101101111",
  64979=>"001000001",
  64980=>"111111111",
  64981=>"000000010",
  64982=>"000010010",
  64983=>"110110110",
  64984=>"000001001",
  64985=>"001001000",
  64986=>"011111111",
  64987=>"011000000",
  64988=>"001011110",
  64989=>"111001000",
  64990=>"001000001",
  64991=>"101111101",
  64992=>"001100111",
  64993=>"000000000",
  64994=>"001000000",
  64995=>"010100111",
  64996=>"001000100",
  64997=>"000111100",
  64998=>"110110010",
  64999=>"000000000",
  65000=>"111000001",
  65001=>"000000110",
  65002=>"111000000",
  65003=>"010100000",
  65004=>"111111111",
  65005=>"000000000",
  65006=>"001000000",
  65007=>"000000000",
  65008=>"101100101",
  65009=>"000000010",
  65010=>"111111110",
  65011=>"001000110",
  65012=>"111111101",
  65013=>"000001111",
  65014=>"001101101",
  65015=>"100000000",
  65016=>"000000000",
  65017=>"100110110",
  65018=>"111111110",
  65019=>"000000000",
  65020=>"110000000",
  65021=>"000001111",
  65022=>"010001001",
  65023=>"001111111",
  65024=>"111000000",
  65025=>"101000000",
  65026=>"000101111",
  65027=>"001111111",
  65028=>"001001000",
  65029=>"100000000",
  65030=>"110111110",
  65031=>"111111111",
  65032=>"111100000",
  65033=>"100000001",
  65034=>"111111111",
  65035=>"000000100",
  65036=>"011001000",
  65037=>"110001000",
  65038=>"000001011",
  65039=>"000000001",
  65040=>"111111111",
  65041=>"111101000",
  65042=>"111001001",
  65043=>"110100101",
  65044=>"000000111",
  65045=>"011000000",
  65046=>"000000000",
  65047=>"011000000",
  65048=>"000000100",
  65049=>"000111111",
  65050=>"000100000",
  65051=>"111110000",
  65052=>"111111100",
  65053=>"111111001",
  65054=>"111011000",
  65055=>"000000000",
  65056=>"101100000",
  65057=>"111111100",
  65058=>"111100111",
  65059=>"000111100",
  65060=>"000000000",
  65061=>"001000000",
  65062=>"111110100",
  65063=>"000111110",
  65064=>"110100001",
  65065=>"111000000",
  65066=>"011011111",
  65067=>"001001111",
  65068=>"111111000",
  65069=>"111000000",
  65070=>"000111111",
  65071=>"011000000",
  65072=>"011000111",
  65073=>"000000000",
  65074=>"101100000",
  65075=>"111111110",
  65076=>"011000000",
  65077=>"000000010",
  65078=>"001001001",
  65079=>"000000000",
  65080=>"000000000",
  65081=>"000000000",
  65082=>"000000111",
  65083=>"000001111",
  65084=>"111111000",
  65085=>"111101000",
  65086=>"111111011",
  65087=>"000000110",
  65088=>"111011001",
  65089=>"111000000",
  65090=>"111001111",
  65091=>"000000100",
  65092=>"011001110",
  65093=>"000000111",
  65094=>"110110000",
  65095=>"111101001",
  65096=>"111100000",
  65097=>"000100000",
  65098=>"111111100",
  65099=>"001001001",
  65100=>"000110111",
  65101=>"101100000",
  65102=>"100110111",
  65103=>"111110110",
  65104=>"100000000",
  65105=>"111111111",
  65106=>"111000000",
  65107=>"000000000",
  65108=>"000011111",
  65109=>"111111000",
  65110=>"111001111",
  65111=>"111000000",
  65112=>"000001001",
  65113=>"000001000",
  65114=>"111101100",
  65115=>"111001000",
  65116=>"000000011",
  65117=>"111101111",
  65118=>"000001100",
  65119=>"000000101",
  65120=>"111011000",
  65121=>"111111111",
  65122=>"000110111",
  65123=>"101110110",
  65124=>"001111111",
  65125=>"000111111",
  65126=>"001001111",
  65127=>"111001000",
  65128=>"000111111",
  65129=>"011001011",
  65130=>"000001111",
  65131=>"111110110",
  65132=>"110110000",
  65133=>"000001000",
  65134=>"111111111",
  65135=>"100110100",
  65136=>"000000000",
  65137=>"111000000",
  65138=>"001011111",
  65139=>"111001000",
  65140=>"000000000",
  65141=>"001000000",
  65142=>"000000000",
  65143=>"001001111",
  65144=>"100000000",
  65145=>"000000000",
  65146=>"000000000",
  65147=>"000000000",
  65148=>"001001000",
  65149=>"100000000",
  65150=>"000000100",
  65151=>"111100111",
  65152=>"001001101",
  65153=>"011011000",
  65154=>"111111110",
  65155=>"000000011",
  65156=>"100000000",
  65157=>"010110100",
  65158=>"000100100",
  65159=>"111000000",
  65160=>"111111011",
  65161=>"111001000",
  65162=>"000000000",
  65163=>"101101010",
  65164=>"100000000",
  65165=>"010000000",
  65166=>"000011110",
  65167=>"111011001",
  65168=>"111110110",
  65169=>"111000000",
  65170=>"100101000",
  65171=>"101000110",
  65172=>"000000001",
  65173=>"000000111",
  65174=>"111000001",
  65175=>"000111111",
  65176=>"101000111",
  65177=>"111111111",
  65178=>"111000000",
  65179=>"000000111",
  65180=>"111000001",
  65181=>"100101111",
  65182=>"110000000",
  65183=>"111111111",
  65184=>"000011111",
  65185=>"101111111",
  65186=>"000000111",
  65187=>"111111111",
  65188=>"011000000",
  65189=>"001111100",
  65190=>"010111010",
  65191=>"001000000",
  65192=>"000100000",
  65193=>"001001111",
  65194=>"011111111",
  65195=>"111000000",
  65196=>"111111000",
  65197=>"000000011",
  65198=>"001101111",
  65199=>"100000111",
  65200=>"000000111",
  65201=>"001111011",
  65202=>"010010111",
  65203=>"000000111",
  65204=>"111111001",
  65205=>"001111111",
  65206=>"000111111",
  65207=>"110000110",
  65208=>"101000111",
  65209=>"111000000",
  65210=>"011111100",
  65211=>"001000110",
  65212=>"000011111",
  65213=>"111101101",
  65214=>"111111101",
  65215=>"001000101",
  65216=>"111111111",
  65217=>"111111100",
  65218=>"111100100",
  65219=>"000100110",
  65220=>"000111011",
  65221=>"000100111",
  65222=>"110111011",
  65223=>"000100111",
  65224=>"000000000",
  65225=>"111110000",
  65226=>"000000000",
  65227=>"111110110",
  65228=>"000000111",
  65229=>"001001111",
  65230=>"101000011",
  65231=>"011110000",
  65232=>"101100010",
  65233=>"000111111",
  65234=>"000111111",
  65235=>"000000000",
  65236=>"101001111",
  65237=>"110100110",
  65238=>"000001000",
  65239=>"100101001",
  65240=>"111000000",
  65241=>"001111111",
  65242=>"111111111",
  65243=>"111100100",
  65244=>"111111000",
  65245=>"110111111",
  65246=>"110111111",
  65247=>"111101111",
  65248=>"000000011",
  65249=>"110000000",
  65250=>"000111111",
  65251=>"001000000",
  65252=>"111111001",
  65253=>"111110100",
  65254=>"000110100",
  65255=>"111000000",
  65256=>"000001000",
  65257=>"111101001",
  65258=>"101100111",
  65259=>"000000000",
  65260=>"000000011",
  65261=>"111111100",
  65262=>"111001111",
  65263=>"111000000",
  65264=>"000001000",
  65265=>"000000111",
  65266=>"111111000",
  65267=>"000000110",
  65268=>"110100111",
  65269=>"011000001",
  65270=>"010001011",
  65271=>"001000000",
  65272=>"000011000",
  65273=>"111111111",
  65274=>"011001000",
  65275=>"111111111",
  65276=>"100101100",
  65277=>"111110010",
  65278=>"110000000",
  65279=>"000000111",
  65280=>"000100000",
  65281=>"011011000",
  65282=>"000000000",
  65283=>"000000000",
  65284=>"000000000",
  65285=>"001011111",
  65286=>"111111111",
  65287=>"000000100",
  65288=>"111111000",
  65289=>"000111111",
  65290=>"111100000",
  65291=>"111111111",
  65292=>"111111111",
  65293=>"000000111",
  65294=>"111111111",
  65295=>"000001000",
  65296=>"000000111",
  65297=>"101000101",
  65298=>"111111111",
  65299=>"100001000",
  65300=>"010010111",
  65301=>"111111010",
  65302=>"111010110",
  65303=>"000100000",
  65304=>"011011011",
  65305=>"000100000",
  65306=>"000000000",
  65307=>"111110110",
  65308=>"111101000",
  65309=>"000000000",
  65310=>"111111111",
  65311=>"111110111",
  65312=>"111110100",
  65313=>"001000111",
  65314=>"000000010",
  65315=>"000001011",
  65316=>"110010000",
  65317=>"001000000",
  65318=>"111100111",
  65319=>"000000000",
  65320=>"000011111",
  65321=>"111110110",
  65322=>"101000000",
  65323=>"111010000",
  65324=>"110000000",
  65325=>"100101000",
  65326=>"000011111",
  65327=>"000001110",
  65328=>"000000000",
  65329=>"111101100",
  65330=>"111001111",
  65331=>"111111111",
  65332=>"000000000",
  65333=>"111111111",
  65334=>"000000000",
  65335=>"111000000",
  65336=>"001000000",
  65337=>"000001000",
  65338=>"111111000",
  65339=>"111111011",
  65340=>"110110111",
  65341=>"000000110",
  65342=>"000111111",
  65343=>"000000011",
  65344=>"001000111",
  65345=>"111110000",
  65346=>"000001101",
  65347=>"000011001",
  65348=>"000011111",
  65349=>"000000000",
  65350=>"111111011",
  65351=>"000000101",
  65352=>"111000000",
  65353=>"111000000",
  65354=>"101111111",
  65355=>"111111101",
  65356=>"110100100",
  65357=>"000111111",
  65358=>"110000000",
  65359=>"111101000",
  65360=>"000100110",
  65361=>"111111000",
  65362=>"101101001",
  65363=>"011111111",
  65364=>"000000000",
  65365=>"111011001",
  65366=>"111001001",
  65367=>"011001111",
  65368=>"000111111",
  65369=>"101111010",
  65370=>"001000000",
  65371=>"100100111",
  65372=>"111100101",
  65373=>"000111111",
  65374=>"001011111",
  65375=>"000011110",
  65376=>"000000000",
  65377=>"000111111",
  65378=>"111100100",
  65379=>"100000000",
  65380=>"011111111",
  65381=>"111111000",
  65382=>"101111111",
  65383=>"111111110",
  65384=>"111111111",
  65385=>"111111111",
  65386=>"111000000",
  65387=>"111111101",
  65388=>"111111000",
  65389=>"110101000",
  65390=>"111000000",
  65391=>"000000000",
  65392=>"010101111",
  65393=>"101001000",
  65394=>"011001111",
  65395=>"000000011",
  65396=>"111011000",
  65397=>"001001100",
  65398=>"000101111",
  65399=>"001100000",
  65400=>"000101000",
  65401=>"111100110",
  65402=>"001111111",
  65403=>"111000000",
  65404=>"000000000",
  65405=>"111010110",
  65406=>"000001111",
  65407=>"111101101",
  65408=>"000001011",
  65409=>"000000000",
  65410=>"000000111",
  65411=>"001000000",
  65412=>"000000110",
  65413=>"101111110",
  65414=>"111110011",
  65415=>"111000000",
  65416=>"011011000",
  65417=>"111101100",
  65418=>"111000000",
  65419=>"000111111",
  65420=>"000100111",
  65421=>"111001111",
  65422=>"001000000",
  65423=>"000111111",
  65424=>"100000000",
  65425=>"000110111",
  65426=>"000000000",
  65427=>"111001111",
  65428=>"111101001",
  65429=>"011011000",
  65430=>"110111111",
  65431=>"011111111",
  65432=>"000011111",
  65433=>"000000000",
  65434=>"111111111",
  65435=>"000101111",
  65436=>"010000000",
  65437=>"111000000",
  65438=>"001011011",
  65439=>"000011111",
  65440=>"000001000",
  65441=>"100000001",
  65442=>"010110001",
  65443=>"000000000",
  65444=>"000111111",
  65445=>"101111010",
  65446=>"000000100",
  65447=>"111000111",
  65448=>"111000000",
  65449=>"000000000",
  65450=>"111100100",
  65451=>"000000111",
  65452=>"000000000",
  65453=>"110111111",
  65454=>"111100000",
  65455=>"111010000",
  65456=>"111111111",
  65457=>"001111101",
  65458=>"111111111",
  65459=>"111111000",
  65460=>"000000000",
  65461=>"111101111",
  65462=>"111111111",
  65463=>"111111001",
  65464=>"100000111",
  65465=>"111111110",
  65466=>"001001000",
  65467=>"111111111",
  65468=>"100000001",
  65469=>"001111000",
  65470=>"000000111",
  65471=>"101100100",
  65472=>"000000110",
  65473=>"011001000",
  65474=>"111111111",
  65475=>"111001000",
  65476=>"111111111",
  65477=>"111000000",
  65478=>"111000000",
  65479=>"001011111",
  65480=>"101100100",
  65481=>"111111000",
  65482=>"000000111",
  65483=>"000000000",
  65484=>"000000000",
  65485=>"010000000",
  65486=>"000000101",
  65487=>"111111001",
  65488=>"100110110",
  65489=>"000111011",
  65490=>"001000000",
  65491=>"001001111",
  65492=>"000000011",
  65493=>"100001000",
  65494=>"000100000",
  65495=>"001001011",
  65496=>"100111111",
  65497=>"011000000",
  65498=>"110000000",
  65499=>"111100101",
  65500=>"000010111",
  65501=>"011000111",
  65502=>"110100101",
  65503=>"011011010",
  65504=>"001001111",
  65505=>"111111111",
  65506=>"000111111",
  65507=>"100111111",
  65508=>"000110110",
  65509=>"111000000",
  65510=>"100110111",
  65511=>"111110111",
  65512=>"111001001",
  65513=>"100111101",
  65514=>"100100110",
  65515=>"000000111",
  65516=>"111111111",
  65517=>"110100100",
  65518=>"011111111",
  65519=>"111001001",
  65520=>"101000000",
  65521=>"011001011",
  65522=>"000000100",
  65523=>"000000111",
  65524=>"000000110",
  65525=>"000000000",
  65526=>"010111111",
  65527=>"001000111",
  65528=>"001100000",
  65529=>"111001001",
  65530=>"101000000",
  65531=>"000000000",
  65532=>"000000000",
  65533=>"111111110",
  65534=>"000011001",
  65535=>"111001000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;