LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L3_2_BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- Instruction bus
        address : IN unsigned(4 DOWNTO 0));
END L3_2_BNROM;

ARCHITECTURE RTL OF L3_2_BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 31) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"1111110000100000"&"0001010111111111",
    1=>"0000100101001101"&"0001010011110101",
    2=>"0000000011000111"&"0001100001101010",
    3=>"1101100100011110"&"0001111010111001",
    4=>"0000001100100011"&"0001101001011011",
    5=>"0000101001111111"&"0001010110001010",
    6=>"0000101100101101"&"0001011011010001",
    7=>"1111111010001010"&"0001010111010111",
    8=>"0000000111010011"&"0001100001111101",
    9=>"0000010011001101"&"0000110000101010",
    10=>"0000101111000111"&"0010001000111101",
    11=>"0000101101101111"&"0001011010010000",
    12=>"1111111111101000"&"0001100110000111",
    13=>"0000011001110110"&"0001101010000100",
    14=>"0000011110100000"&"0001100110110111",
    15=>"0000001001011010"&"0001110001011000",
    16=>"0001001010100010"&"0000111010100000",
    17=>"0000000110110010"&"0001001100010010",
    18=>"1111111111001101"&"0001011100011011",
    19=>"0000000010010000"&"0001110101101100",
    20=>"0001000100111100"&"0000110100111100",
    21=>"1111110000111111"&"0001101101011000",
    22=>"0000001001010001"&"0010000010010000",
    23=>"1111101111001000"&"0001010110111010",
    24=>"0000000101101101"&"0001101001101010",
    25=>"0001000101000000"&"0010001001100110",
    26=>"0000000110010100"&"0001100010111101",
    27=>"0000100010110111"&"0001101101000101",
    28=>"1111101001000100"&"0001010000110100",
    29=>"1110111001110111"&"0001101110110000",
    30=>"0000010111000101"&"0001011110010000",
    31=>"1111111011110001"&"0000111000010101");
    
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;