LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_3_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_3_BNROM;

ARCHITECTURE RTL OF L8_3_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0001110100011011"&"0010000011011011",
  1=>"0001110011011100"&"0010010110111000",
  2=>"0000101011100101"&"0010000111101111",
  3=>"0010000100000101"&"0010011100101001",
  4=>"0000111100110000"&"0010000101011000",
  5=>"0011110101010101"&"0010000100111001",
  6=>"0010010100110110"&"0001110110001011",
  7=>"0000100010000111"&"0010010011010011",
  8=>"0010110000001011"&"0010010011001000",
  9=>"0001011010010010"&"0010001000000001",
  10=>"0000010010101000"&"0010000110110101",
  11=>"0001100100000001"&"0010011101100100",
  12=>"0001001001111011"&"0010011101111001",
  13=>"0001010101111110"&"0001101000011101",
  14=>"0001001101011010"&"0010001111111101",
  15=>"1111110010001000"&"0010000101100000",
  16=>"1110010010011110"&"0001101110110100",
  17=>"0001011011001101"&"0010000011000000",
  18=>"0001110111000000"&"0001111011101100",
  19=>"0000001010001100"&"0010000011011001",
  20=>"0001101100111011"&"0010001111010100",
  21=>"0001111110111001"&"0010010101100000",
  22=>"0001101101011101"&"0010011100101010",
  23=>"0001110001110100"&"0010001001101111",
  24=>"0001111001101001"&"0010011010111011",
  25=>"0001110000100011"&"0010011011101001",
  26=>"0010000101011010"&"0010011000000101",
  27=>"0000110010100110"&"0010010111010000",
  28=>"0010000000101111"&"0001111001110001",
  29=>"0001100100111100"&"0010000110101111",
  30=>"0001011100010101"&"0001101100000011",
  31=>"0000110111010110"&"0010011010110000",
  32=>"0001010101111100"&"0010001111000000",
  33=>"0001010001101000"&"0010000110011100",
  34=>"0001000100110110"&"0010001100100111",
  35=>"0001100011100110"&"0010000001100010",
  36=>"0001111111001100"&"0001110111110011",
  37=>"0001000010000110"&"0010010110101010",
  38=>"0001001001101010"&"0010011010010111",
  39=>"0001010001101100"&"0010000111100111",
  40=>"0000110011101101"&"0010010100100011",
  41=>"1110101001101000"&"0001011010011111",
  42=>"0000110011111111"&"0010001000010010",
  43=>"0000011101011011"&"0010001111110100",
  44=>"0001101110000010"&"0010001000111111",
  45=>"0000101001101110"&"0010000110110101",
  46=>"0001111110110001"&"0010001001000011",
  47=>"0001001010101000"&"0010000110000010",
  48=>"0010000011001001"&"0010011110100000",
  49=>"0010001000001000"&"0010010010011100",
  50=>"0001110000011101"&"0010001100100101",
  51=>"0000001000101000"&"0010011000110011",
  52=>"0000110011111101"&"0010001111010110",
  53=>"0001110100011000"&"0010001111110000",
  54=>"0000100111000111"&"0010011010111011",
  55=>"0000100110001010"&"0010100001101001",
  56=>"0010110110111110"&"0010011110010000",
  57=>"0000101110100100"&"0001110101111110",
  58=>"0001000101000111"&"0010001010000111",
  59=>"0000100010011100"&"0010010011100101",
  60=>"1110110100000010"&"0001111110010101",
  61=>"0010000111001111"&"0001011110110110",
  62=>"1111110111101000"&"0010000111101111",
  63=>"0001010111000010"&"0010010010010001");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;